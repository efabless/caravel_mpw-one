VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2994.580 BY 3583.920 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 61.400 2957.480 62.000 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2407.400 2957.480 2408.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2642.000 2957.480 2642.600 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2876.600 2957.480 2877.200 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3111.200 2957.480 3111.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3345.800 2957.480 3346.400 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2916.710 3549.720 2916.990 3552.120 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2592.410 3549.720 2592.690 3552.120 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2268.110 3549.720 2268.390 3552.120 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1943.350 3549.720 1943.630 3552.120 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1619.050 3549.720 1619.330 3552.120 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 296.000 2957.480 296.600 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1294.750 3549.720 1295.030 3552.120 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 969.990 3549.720 970.270 3552.120 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 645.690 3549.720 645.970 3552.120 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 321.390 3549.720 321.670 3552.120 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 3515.120 39.880 3515.720 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 3227.480 39.880 3228.080 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2940.520 39.880 2941.120 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2652.880 39.880 2653.480 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2365.920 39.880 2366.520 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2078.280 39.880 2078.880 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 530.600 2957.480 531.200 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 1791.320 39.880 1791.920 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 765.200 2957.480 765.800 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 999.800 2957.480 1000.400 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1234.400 2957.480 1235.000 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1469.000 2957.480 1469.600 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1703.600 2957.480 1704.200 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1938.200 2957.480 1938.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2172.800 2957.480 2173.400 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 119.880 2957.480 120.480 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2465.880 2957.480 2466.480 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2701.160 2957.480 2701.760 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2935.760 2957.480 2936.360 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3170.360 2957.480 3170.960 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3404.960 2957.480 3405.560 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2835.750 3549.720 2836.030 3552.120 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2511.450 3549.720 2511.730 3552.120 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2186.690 3549.720 2186.970 3552.120 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1862.390 3549.720 1862.670 3552.120 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1538.090 3549.720 1538.370 3552.120 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 354.480 2957.480 355.080 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.330 3549.720 1213.610 3552.120 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 889.030 3549.720 889.310 3552.120 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.730 3549.720 565.010 3552.120 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.970 3549.720 240.250 3552.120 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 3443.040 39.880 3443.640 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 3156.080 39.880 3156.680 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2868.440 39.880 2869.040 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2581.480 39.880 2582.080 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2293.840 39.880 2294.440 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 2006.880 39.880 2007.480 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 589.080 2957.480 589.680 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 1719.240 39.880 1719.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 1503.680 39.880 1504.280 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 1288.120 39.880 1288.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 1072.560 39.880 1073.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 857.000 39.880 857.600 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 642.120 39.880 642.720 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 426.560 39.880 427.160 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 37.480 211.000 39.880 211.600 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 823.680 2957.480 824.280 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1058.280 2957.480 1058.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1292.880 2957.480 1293.480 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1527.480 2957.480 1528.080 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1762.080 2957.480 1762.680 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1996.680 2957.480 1997.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2231.280 2957.480 2231.880 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 236.840 2957.480 237.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2583.520 2957.480 2584.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2818.120 2957.480 2818.720 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3052.720 2957.480 3053.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3287.320 2957.480 3287.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3521.920 2957.480 3522.520 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2673.370 3549.720 2673.650 3552.120 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2349.070 3549.720 2349.350 3552.120 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2024.770 3549.720 2025.050 3552.120 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1700.010 3549.720 1700.290 3552.120 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.710 3549.720 1375.990 3552.120 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 471.440 2957.480 472.040 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1051.410 3549.720 1051.690 3552.120 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 726.650 3549.720 726.930 3552.120 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.350 3549.720 402.630 3552.120 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.050 3549.720 78.330 3552.120 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 3299.560 39.880 3300.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 3011.920 39.880 3012.520 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 2724.960 39.880 2725.560 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 2437.320 39.880 2437.920 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 2150.360 39.880 2150.960 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1862.720 39.880 1863.320 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 706.040 2957.480 706.640 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1575.760 39.880 1576.360 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1360.200 39.880 1360.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1144.640 39.880 1145.240 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 929.080 39.880 929.680 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 713.520 39.880 714.120 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 497.960 39.880 498.560 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 282.400 39.880 283.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 67.520 39.880 68.120 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 941.320 2957.480 941.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1175.920 2957.480 1176.520 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1410.520 2957.480 1411.120 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1645.120 2957.480 1645.720 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1879.720 2957.480 1880.320 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2114.320 2957.480 2114.920 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2348.920 2957.480 2349.520 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 178.360 2957.480 178.960 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2525.040 2957.480 2525.640 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2759.640 2957.480 2760.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2994.240 2957.480 2994.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3228.840 2957.480 3229.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 3463.440 2957.480 3464.040 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2754.790 3549.720 2755.070 3552.120 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2430.030 3549.720 2430.310 3552.120 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2105.730 3549.720 2106.010 3552.120 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1781.430 3549.720 1781.710 3552.120 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1456.670 3549.720 1456.950 3552.120 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 412.960 2957.480 413.560 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1132.370 3549.720 1132.650 3552.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 808.070 3549.720 808.350 3552.120 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.310 3549.720 483.590 3552.120 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.010 3549.720 159.290 3552.120 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 3371.640 39.880 3372.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 3084.000 39.880 3084.600 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 2797.040 39.880 2797.640 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 2509.400 39.880 2510.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 2221.760 39.880 2222.360 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1934.800 39.880 1935.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 647.560 2957.480 648.160 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1647.160 39.880 1647.760 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1432.280 39.880 1432.880 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1216.720 39.880 1217.320 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 1001.160 39.880 1001.760 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 785.600 39.880 786.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 570.040 39.880 570.640 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 354.480 39.880 355.080 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 37.480 138.920 39.880 139.520 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 882.160 2957.480 882.760 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1116.760 2957.480 1117.360 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1351.360 2957.480 1351.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1585.960 2957.480 1586.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 1821.240 2957.480 1821.840 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2055.840 2957.480 2056.440 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2955.080 2290.440 2957.480 2291.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.530 32.120 670.810 34.520 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2454.870 32.120 2455.150 34.520 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2472.350 32.120 2472.630 34.520 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2490.290 32.120 2490.570 34.520 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2508.230 32.120 2508.510 34.520 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2526.170 32.120 2526.450 34.520 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2543.650 32.120 2543.930 34.520 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2561.590 32.120 2561.870 34.520 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2579.530 32.120 2579.810 34.520 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2597.470 32.120 2597.750 34.520 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2615.410 32.120 2615.690 34.520 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 849.010 32.120 849.290 34.520 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2632.890 32.120 2633.170 34.520 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2650.830 32.120 2651.110 34.520 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2668.770 32.120 2669.050 34.520 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2686.710 32.120 2686.990 34.520 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2704.650 32.120 2704.930 34.520 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2722.130 32.120 2722.410 34.520 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2740.070 32.120 2740.350 34.520 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2758.010 32.120 2758.290 34.520 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2775.950 32.120 2776.230 34.520 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2793.430 32.120 2793.710 34.520 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.950 32.120 867.230 34.520 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2811.370 32.120 2811.650 34.520 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2829.310 32.120 2829.590 34.520 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2847.250 32.120 2847.530 34.520 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2865.190 32.120 2865.470 34.520 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2882.670 32.120 2882.950 34.520 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2900.610 32.120 2900.890 34.520 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2918.550 32.120 2918.830 34.520 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2936.490 32.120 2936.770 34.520 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.430 32.120 884.710 34.520 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.370 32.120 902.650 34.520 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.310 32.120 920.590 34.520 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.250 32.120 938.530 34.520 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.190 32.120 956.470 34.520 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.670 32.120 973.950 34.520 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.610 32.120 991.890 34.520 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.550 32.120 1009.830 34.520 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 688.470 32.120 688.750 34.520 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.490 32.120 1027.770 34.520 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.970 32.120 1045.250 34.520 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.910 32.120 1063.190 34.520 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.850 32.120 1081.130 34.520 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.790 32.120 1099.070 34.520 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.730 32.120 1117.010 34.520 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1134.210 32.120 1134.490 34.520 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.150 32.120 1152.430 34.520 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.090 32.120 1170.370 34.520 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1188.030 32.120 1188.310 34.520 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 706.410 32.120 706.690 34.520 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1205.970 32.120 1206.250 34.520 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1223.450 32.120 1223.730 34.520 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1241.390 32.120 1241.670 34.520 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.330 32.120 1259.610 34.520 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.270 32.120 1277.550 34.520 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.750 32.120 1295.030 34.520 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1312.690 32.120 1312.970 34.520 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1330.630 32.120 1330.910 34.520 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.570 32.120 1348.850 34.520 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1366.510 32.120 1366.790 34.520 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.890 32.120 724.170 34.520 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1383.990 32.120 1384.270 34.520 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1401.930 32.120 1402.210 34.520 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1419.870 32.120 1420.150 34.520 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1437.810 32.120 1438.090 34.520 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.750 32.120 1456.030 34.520 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1473.230 32.120 1473.510 34.520 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1491.170 32.120 1491.450 34.520 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1509.110 32.120 1509.390 34.520 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1527.050 32.120 1527.330 34.520 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1544.530 32.120 1544.810 34.520 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.830 32.120 742.110 34.520 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1562.470 32.120 1562.750 34.520 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1580.410 32.120 1580.690 34.520 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1598.350 32.120 1598.630 34.520 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1616.290 32.120 1616.570 34.520 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1633.770 32.120 1634.050 34.520 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1651.710 32.120 1651.990 34.520 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1669.650 32.120 1669.930 34.520 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1687.590 32.120 1687.870 34.520 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1705.530 32.120 1705.810 34.520 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1723.010 32.120 1723.290 34.520 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.770 32.120 760.050 34.520 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1740.950 32.120 1741.230 34.520 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1758.890 32.120 1759.170 34.520 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1776.830 32.120 1777.110 34.520 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1794.310 32.120 1794.590 34.520 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1812.250 32.120 1812.530 34.520 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1830.190 32.120 1830.470 34.520 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1848.130 32.120 1848.410 34.520 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1866.070 32.120 1866.350 34.520 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1883.550 32.120 1883.830 34.520 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1901.490 32.120 1901.770 34.520 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 777.710 32.120 777.990 34.520 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1919.430 32.120 1919.710 34.520 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1937.370 32.120 1937.650 34.520 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1955.310 32.120 1955.590 34.520 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1972.790 32.120 1973.070 34.520 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1990.730 32.120 1991.010 34.520 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2008.670 32.120 2008.950 34.520 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2026.610 32.120 2026.890 34.520 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2044.090 32.120 2044.370 34.520 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2062.030 32.120 2062.310 34.520 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2079.970 32.120 2080.250 34.520 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 795.190 32.120 795.470 34.520 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2097.910 32.120 2098.190 34.520 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2115.850 32.120 2116.130 34.520 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2133.330 32.120 2133.610 34.520 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2151.270 32.120 2151.550 34.520 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2169.210 32.120 2169.490 34.520 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2187.150 32.120 2187.430 34.520 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2205.090 32.120 2205.370 34.520 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2222.570 32.120 2222.850 34.520 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2240.510 32.120 2240.790 34.520 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2258.450 32.120 2258.730 34.520 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 813.130 32.120 813.410 34.520 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2276.390 32.120 2276.670 34.520 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2293.870 32.120 2294.150 34.520 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2311.810 32.120 2312.090 34.520 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2329.750 32.120 2330.030 34.520 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2347.690 32.120 2347.970 34.520 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2365.630 32.120 2365.910 34.520 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2383.110 32.120 2383.390 34.520 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2401.050 32.120 2401.330 34.520 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2418.990 32.120 2419.270 34.520 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2436.930 32.120 2437.210 34.520 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.070 32.120 831.350 34.520 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.510 32.120 676.790 34.520 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2460.390 32.120 2460.670 34.520 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2478.330 32.120 2478.610 34.520 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2496.270 32.120 2496.550 34.520 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2514.210 32.120 2514.490 34.520 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2532.150 32.120 2532.430 34.520 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2549.630 32.120 2549.910 34.520 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2567.570 32.120 2567.850 34.520 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2585.510 32.120 2585.790 34.520 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2603.450 32.120 2603.730 34.520 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2621.390 32.120 2621.670 34.520 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 854.990 32.120 855.270 34.520 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2638.870 32.120 2639.150 34.520 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2656.810 32.120 2657.090 34.520 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2674.750 32.120 2675.030 34.520 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2692.690 32.120 2692.970 34.520 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2710.170 32.120 2710.450 34.520 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2728.110 32.120 2728.390 34.520 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2746.050 32.120 2746.330 34.520 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2763.990 32.120 2764.270 34.520 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2781.930 32.120 2782.210 34.520 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2799.410 32.120 2799.690 34.520 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 872.930 32.120 873.210 34.520 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2817.350 32.120 2817.630 34.520 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2835.290 32.120 2835.570 34.520 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2853.230 32.120 2853.510 34.520 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2871.170 32.120 2871.450 34.520 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2888.650 32.120 2888.930 34.520 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2906.590 32.120 2906.870 34.520 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2924.530 32.120 2924.810 34.520 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2942.470 32.120 2942.750 34.520 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 890.410 32.120 890.690 34.520 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 908.350 32.120 908.630 34.520 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.290 32.120 926.570 34.520 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.230 32.120 944.510 34.520 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.710 32.120 961.990 34.520 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.650 32.120 979.930 34.520 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.590 32.120 997.870 34.520 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1015.530 32.120 1015.810 34.520 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.450 32.120 694.730 34.520 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1033.470 32.120 1033.750 34.520 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1050.950 32.120 1051.230 34.520 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.890 32.120 1069.170 34.520 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1086.830 32.120 1087.110 34.520 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1104.770 32.120 1105.050 34.520 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1122.710 32.120 1122.990 34.520 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1140.190 32.120 1140.470 34.520 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1158.130 32.120 1158.410 34.520 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1176.070 32.120 1176.350 34.520 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1194.010 32.120 1194.290 34.520 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 711.930 32.120 712.210 34.520 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1211.490 32.120 1211.770 34.520 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1229.430 32.120 1229.710 34.520 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1247.370 32.120 1247.650 34.520 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.310 32.120 1265.590 34.520 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.250 32.120 1283.530 34.520 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1300.730 32.120 1301.010 34.520 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1318.670 32.120 1318.950 34.520 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1336.610 32.120 1336.890 34.520 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1354.550 32.120 1354.830 34.520 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1372.490 32.120 1372.770 34.520 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 729.870 32.120 730.150 34.520 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1389.970 32.120 1390.250 34.520 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1407.910 32.120 1408.190 34.520 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1425.850 32.120 1426.130 34.520 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1443.790 32.120 1444.070 34.520 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1461.270 32.120 1461.550 34.520 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1479.210 32.120 1479.490 34.520 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1497.150 32.120 1497.430 34.520 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1515.090 32.120 1515.370 34.520 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1533.030 32.120 1533.310 34.520 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1550.510 32.120 1550.790 34.520 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 747.810 32.120 748.090 34.520 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1568.450 32.120 1568.730 34.520 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1586.390 32.120 1586.670 34.520 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1604.330 32.120 1604.610 34.520 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1622.270 32.120 1622.550 34.520 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1639.750 32.120 1640.030 34.520 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1657.690 32.120 1657.970 34.520 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1675.630 32.120 1675.910 34.520 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1693.570 32.120 1693.850 34.520 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1711.050 32.120 1711.330 34.520 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1728.990 32.120 1729.270 34.520 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.750 32.120 766.030 34.520 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1746.930 32.120 1747.210 34.520 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1764.870 32.120 1765.150 34.520 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1782.810 32.120 1783.090 34.520 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1800.290 32.120 1800.570 34.520 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1818.230 32.120 1818.510 34.520 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1836.170 32.120 1836.450 34.520 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1854.110 32.120 1854.390 34.520 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1872.050 32.120 1872.330 34.520 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1889.530 32.120 1889.810 34.520 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1907.470 32.120 1907.750 34.520 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.690 32.120 783.970 34.520 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1925.410 32.120 1925.690 34.520 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1943.350 32.120 1943.630 34.520 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1960.830 32.120 1961.110 34.520 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1978.770 32.120 1979.050 34.520 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1996.710 32.120 1996.990 34.520 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2014.650 32.120 2014.930 34.520 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2032.590 32.120 2032.870 34.520 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2050.070 32.120 2050.350 34.520 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.010 32.120 2068.290 34.520 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2085.950 32.120 2086.230 34.520 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 801.170 32.120 801.450 34.520 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2103.890 32.120 2104.170 34.520 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2121.830 32.120 2122.110 34.520 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2139.310 32.120 2139.590 34.520 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2157.250 32.120 2157.530 34.520 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2175.190 32.120 2175.470 34.520 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2193.130 32.120 2193.410 34.520 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2210.610 32.120 2210.890 34.520 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2228.550 32.120 2228.830 34.520 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2246.490 32.120 2246.770 34.520 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2264.430 32.120 2264.710 34.520 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.110 32.120 819.390 34.520 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2282.370 32.120 2282.650 34.520 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2299.850 32.120 2300.130 34.520 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2317.790 32.120 2318.070 34.520 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2335.730 32.120 2336.010 34.520 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2353.670 32.120 2353.950 34.520 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2371.610 32.120 2371.890 34.520 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2389.090 32.120 2389.370 34.520 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2407.030 32.120 2407.310 34.520 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2424.970 32.120 2425.250 34.520 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2442.910 32.120 2443.190 34.520 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 837.050 32.120 837.330 34.520 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 682.490 32.120 682.770 34.520 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2466.370 32.120 2466.650 34.520 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2484.310 32.120 2484.590 34.520 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2502.250 32.120 2502.530 34.520 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2520.190 32.120 2520.470 34.520 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2538.130 32.120 2538.410 34.520 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2555.610 32.120 2555.890 34.520 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2573.550 32.120 2573.830 34.520 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2591.490 32.120 2591.770 34.520 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2609.430 32.120 2609.710 34.520 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2626.910 32.120 2627.190 34.520 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 860.970 32.120 861.250 34.520 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2644.850 32.120 2645.130 34.520 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2662.790 32.120 2663.070 34.520 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2680.730 32.120 2681.010 34.520 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2698.670 32.120 2698.950 34.520 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2716.150 32.120 2716.430 34.520 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2734.090 32.120 2734.370 34.520 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2752.030 32.120 2752.310 34.520 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2769.970 32.120 2770.250 34.520 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2787.910 32.120 2788.190 34.520 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2805.390 32.120 2805.670 34.520 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 878.450 32.120 878.730 34.520 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2823.330 32.120 2823.610 34.520 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2841.270 32.120 2841.550 34.520 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2859.210 32.120 2859.490 34.520 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2876.690 32.120 2876.970 34.520 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2894.630 32.120 2894.910 34.520 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2912.570 32.120 2912.850 34.520 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2930.510 32.120 2930.790 34.520 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2948.450 32.120 2948.730 34.520 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.390 32.120 896.670 34.520 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 914.330 32.120 914.610 34.520 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.270 32.120 932.550 34.520 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.210 32.120 950.490 34.520 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.690 32.120 967.970 34.520 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.630 32.120 985.910 34.520 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.570 32.120 1003.850 34.520 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.510 32.120 1021.790 34.520 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.430 32.120 700.710 34.520 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.450 32.120 1039.730 34.520 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1056.930 32.120 1057.210 34.520 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1074.870 32.120 1075.150 34.520 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.810 32.120 1093.090 34.520 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.750 32.120 1111.030 34.520 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.230 32.120 1128.510 34.520 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1146.170 32.120 1146.450 34.520 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1164.110 32.120 1164.390 34.520 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1182.050 32.120 1182.330 34.520 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.990 32.120 1200.270 34.520 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 717.910 32.120 718.190 34.520 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1217.470 32.120 1217.750 34.520 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1235.410 32.120 1235.690 34.520 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1253.350 32.120 1253.630 34.520 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.290 32.120 1271.570 34.520 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1289.230 32.120 1289.510 34.520 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1306.710 32.120 1306.990 34.520 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1324.650 32.120 1324.930 34.520 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1342.590 32.120 1342.870 34.520 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.530 32.120 1360.810 34.520 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1378.010 32.120 1378.290 34.520 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 735.850 32.120 736.130 34.520 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1395.950 32.120 1396.230 34.520 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1413.890 32.120 1414.170 34.520 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1431.830 32.120 1432.110 34.520 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1449.770 32.120 1450.050 34.520 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1467.250 32.120 1467.530 34.520 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1485.190 32.120 1485.470 34.520 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1503.130 32.120 1503.410 34.520 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1521.070 32.120 1521.350 34.520 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1539.010 32.120 1539.290 34.520 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1556.490 32.120 1556.770 34.520 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.790 32.120 754.070 34.520 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1574.430 32.120 1574.710 34.520 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1592.370 32.120 1592.650 34.520 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1610.310 32.120 1610.590 34.520 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.790 32.120 1628.070 34.520 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1645.730 32.120 1646.010 34.520 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1663.670 32.120 1663.950 34.520 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1681.610 32.120 1681.890 34.520 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1699.550 32.120 1699.830 34.520 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1717.030 32.120 1717.310 34.520 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1734.970 32.120 1735.250 34.520 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.730 32.120 772.010 34.520 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1752.910 32.120 1753.190 34.520 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1770.850 32.120 1771.130 34.520 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1788.790 32.120 1789.070 34.520 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1806.270 32.120 1806.550 34.520 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.210 32.120 1824.490 34.520 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1842.150 32.120 1842.430 34.520 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1860.090 32.120 1860.370 34.520 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1877.570 32.120 1877.850 34.520 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1895.510 32.120 1895.790 34.520 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1913.450 32.120 1913.730 34.520 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.670 32.120 789.950 34.520 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1931.390 32.120 1931.670 34.520 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1949.330 32.120 1949.610 34.520 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1966.810 32.120 1967.090 34.520 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1984.750 32.120 1985.030 34.520 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2002.690 32.120 2002.970 34.520 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2020.630 32.120 2020.910 34.520 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2038.570 32.120 2038.850 34.520 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2056.050 32.120 2056.330 34.520 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2073.990 32.120 2074.270 34.520 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2091.930 32.120 2092.210 34.520 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.150 32.120 807.430 34.520 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2109.870 32.120 2110.150 34.520 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2127.350 32.120 2127.630 34.520 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2145.290 32.120 2145.570 34.520 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2163.230 32.120 2163.510 34.520 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2181.170 32.120 2181.450 34.520 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2199.110 32.120 2199.390 34.520 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2216.590 32.120 2216.870 34.520 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2234.530 32.120 2234.810 34.520 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2252.470 32.120 2252.750 34.520 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2270.410 32.120 2270.690 34.520 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.090 32.120 825.370 34.520 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2288.350 32.120 2288.630 34.520 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2305.830 32.120 2306.110 34.520 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2323.770 32.120 2324.050 34.520 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2341.710 32.120 2341.990 34.520 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2359.650 32.120 2359.930 34.520 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2377.130 32.120 2377.410 34.520 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2395.070 32.120 2395.350 34.520 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2413.010 32.120 2413.290 34.520 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2430.950 32.120 2431.230 34.520 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2448.890 32.120 2449.170 34.520 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 843.030 32.120 843.310 34.520 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2954.430 32.120 2954.710 34.520 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.330 32.120 40.610 34.520 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 91.830 44.445 93.490 44.645 ;
      LAYER L1M1_PR_C ;
        RECT 91.835 44.445 92.005 44.615 ;
      LAYER met1 ;
        RECT 45.760 48.000 46.080 48.060 ;
        RECT 77.960 48.000 78.280 48.060 ;
        RECT 45.760 47.860 78.280 48.000 ;
        RECT 45.760 47.800 46.080 47.860 ;
        RECT 77.960 47.800 78.280 47.860 ;
        RECT 91.775 44.415 92.065 44.645 ;
        RECT 77.960 43.920 78.280 43.980 ;
        RECT 91.850 43.920 91.990 44.415 ;
        RECT 77.960 43.780 91.990 43.920 ;
        RECT 77.960 43.720 78.280 43.780 ;
      LAYER via ;
        RECT 45.790 47.800 46.050 48.060 ;
        RECT 77.990 47.800 78.250 48.060 ;
        RECT 77.990 43.720 78.250 43.980 ;
      LAYER met2 ;
        RECT 45.790 47.770 46.050 48.090 ;
        RECT 77.990 47.770 78.250 48.090 ;
        RECT 45.850 34.520 45.990 47.770 ;
        RECT 78.050 44.010 78.190 47.770 ;
        RECT 77.990 43.690 78.250 44.010 ;
        RECT 45.780 32.120 46.130 34.520 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 51.740 51.740 52.060 51.800 ;
        RECT 77.040 51.740 77.360 51.800 ;
        RECT 51.740 51.600 77.360 51.740 ;
        RECT 51.740 51.540 52.060 51.600 ;
        RECT 77.040 51.540 77.360 51.600 ;
      LAYER via ;
        RECT 51.770 51.540 52.030 51.800 ;
        RECT 77.070 51.540 77.330 51.800 ;
      LAYER met2 ;
        RECT 77.130 51.830 77.270 54.000 ;
        RECT 51.770 51.510 52.030 51.830 ;
        RECT 77.070 51.510 77.330 51.830 ;
        RECT 51.830 34.520 51.970 51.510 ;
        RECT 51.760 32.120 52.110 34.520 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.750 32.120 76.030 34.520 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.150 32.120 278.430 34.520 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 281.280 38.820 281.600 38.880 ;
        RECT 295.540 38.820 295.860 38.880 ;
        RECT 281.280 38.680 295.860 38.820 ;
        RECT 281.280 38.620 281.600 38.680 ;
        RECT 295.540 38.620 295.860 38.680 ;
      LAYER via ;
        RECT 281.310 38.620 281.570 38.880 ;
        RECT 295.570 38.620 295.830 38.880 ;
      LAYER met2 ;
        RECT 281.370 38.910 281.510 54.000 ;
        RECT 281.310 38.590 281.570 38.910 ;
        RECT 295.570 38.590 295.830 38.910 ;
        RECT 295.630 34.520 295.770 38.590 ;
        RECT 295.560 32.120 295.910 34.520 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.570 32.120 313.850 34.520 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.510 32.120 331.790 34.520 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 342.000 45.280 342.320 45.340 ;
        RECT 349.360 45.280 349.680 45.340 ;
        RECT 342.000 45.140 349.680 45.280 ;
        RECT 342.000 45.080 342.320 45.140 ;
        RECT 349.360 45.080 349.680 45.140 ;
      LAYER via ;
        RECT 342.030 45.080 342.290 45.340 ;
        RECT 349.390 45.080 349.650 45.340 ;
      LAYER met2 ;
        RECT 342.090 45.370 342.230 54.000 ;
        RECT 342.030 45.050 342.290 45.370 ;
        RECT 349.390 45.050 349.650 45.370 ;
        RECT 349.450 34.520 349.590 45.050 ;
        RECT 349.380 32.120 349.730 34.520 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.390 32.120 367.670 34.520 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 395.605 46.635 396.125 48.185 ;
      LAYER L1M1_PR_C ;
        RECT 395.895 47.165 396.065 47.335 ;
      LAYER met1 ;
        RECT 384.780 47.320 385.100 47.380 ;
        RECT 395.835 47.320 396.125 47.365 ;
        RECT 384.780 47.180 396.125 47.320 ;
        RECT 384.780 47.120 385.100 47.180 ;
        RECT 395.835 47.135 396.125 47.180 ;
      LAYER via ;
        RECT 384.810 47.120 385.070 47.380 ;
      LAYER met2 ;
        RECT 384.810 47.090 385.070 47.410 ;
        RECT 384.870 34.520 385.010 47.090 ;
        RECT 384.800 32.120 385.150 34.520 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 402.810 32.120 403.090 34.520 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.750 32.120 421.030 34.520 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.620 32.120 438.970 34.520 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 148.355 50.430 148.690 50.855 ;
        RECT 149.210 50.430 149.545 50.855 ;
        RECT 148.355 50.260 150.025 50.430 ;
        RECT 149.780 49.695 150.025 50.260 ;
        RECT 148.355 49.525 150.025 49.695 ;
        RECT 148.355 48.765 148.690 49.525 ;
        RECT 149.210 48.765 149.540 49.525 ;
      LAYER L1M1_PR_C ;
        RECT 148.415 48.865 148.585 49.035 ;
      LAYER met1 ;
        RECT 148.340 49.020 148.660 49.080 ;
        RECT 148.145 48.880 148.660 49.020 ;
        RECT 148.340 48.820 148.660 48.880 ;
        RECT 99.580 48.000 99.900 48.060 ;
        RECT 146.960 48.000 147.280 48.060 ;
        RECT 148.340 48.000 148.660 48.060 ;
        RECT 99.580 47.860 106.710 48.000 ;
        RECT 99.580 47.800 99.900 47.860 ;
        RECT 106.570 47.660 106.710 47.860 ;
        RECT 146.960 47.860 148.660 48.000 ;
        RECT 146.960 47.800 147.280 47.860 ;
        RECT 148.340 47.800 148.660 47.860 ;
        RECT 113.380 47.660 113.700 47.720 ;
        RECT 106.570 47.520 113.700 47.660 ;
        RECT 113.380 47.460 113.700 47.520 ;
      LAYER via ;
        RECT 148.370 48.820 148.630 49.080 ;
        RECT 99.610 47.800 99.870 48.060 ;
        RECT 146.990 47.800 147.250 48.060 ;
        RECT 148.370 47.800 148.630 48.060 ;
        RECT 113.410 47.460 113.670 47.720 ;
      LAYER met2 ;
        RECT 138.310 48.285 138.450 54.000 ;
        RECT 148.370 48.790 148.630 49.110 ;
        RECT 99.610 47.770 99.870 48.090 ;
        RECT 113.400 47.915 113.680 48.285 ;
        RECT 138.240 47.915 138.520 48.285 ;
        RECT 146.980 47.915 147.260 48.285 ;
        RECT 148.430 48.090 148.570 48.790 ;
        RECT 99.670 34.520 99.810 47.770 ;
        RECT 113.470 47.750 113.610 47.915 ;
        RECT 146.990 47.770 147.250 47.915 ;
        RECT 148.370 47.770 148.630 48.090 ;
        RECT 113.410 47.430 113.670 47.750 ;
        RECT 99.600 32.120 99.950 34.520 ;
      LAYER via2 ;
        RECT 113.400 47.960 113.680 48.240 ;
        RECT 138.240 47.960 138.520 48.240 ;
        RECT 146.980 47.960 147.260 48.240 ;
      LAYER met3 ;
        RECT 113.375 48.250 113.705 48.265 ;
        RECT 138.215 48.250 138.545 48.265 ;
        RECT 146.955 48.250 147.285 48.265 ;
        RECT 113.375 47.950 147.285 48.250 ;
        RECT 113.375 47.935 113.705 47.950 ;
        RECT 138.215 47.935 138.545 47.950 ;
        RECT 146.955 47.935 147.285 47.950 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 456.630 32.120 456.910 34.520 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.110 32.120 474.390 34.520 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.050 32.120 492.330 34.520 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 512.905 46.635 513.425 48.185 ;
      LAYER L1M1_PR_C ;
        RECT 513.195 46.825 513.365 46.995 ;
      LAYER met1 ;
        RECT 509.900 46.980 510.220 47.040 ;
        RECT 513.135 46.980 513.425 47.025 ;
        RECT 509.900 46.840 513.425 46.980 ;
        RECT 509.900 46.780 510.220 46.840 ;
        RECT 513.135 46.795 513.425 46.840 ;
      LAYER via ;
        RECT 509.930 46.780 510.190 47.040 ;
      LAYER met2 ;
        RECT 509.930 46.750 510.190 47.070 ;
        RECT 509.990 34.520 510.130 46.750 ;
        RECT 509.920 32.120 510.270 34.520 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.930 32.120 528.210 34.520 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 545.340 32.120 545.690 34.520 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 563.350 32.120 563.630 34.520 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.290 32.120 581.570 34.520 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.160 32.120 599.510 34.520 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 617.170 32.120 617.450 34.520 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.590 32.120 123.870 34.520 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 622.845 43.255 623.365 44.805 ;
      LAYER L1M1_PR_C ;
        RECT 623.135 44.445 623.305 44.615 ;
      LAYER met1 ;
        RECT 623.060 46.300 623.380 46.360 ;
        RECT 634.560 46.300 634.880 46.360 ;
        RECT 623.060 46.160 634.880 46.300 ;
        RECT 623.060 46.100 623.380 46.160 ;
        RECT 634.560 46.100 634.880 46.160 ;
        RECT 623.060 44.600 623.380 44.660 ;
        RECT 622.865 44.460 623.380 44.600 ;
        RECT 623.060 44.400 623.380 44.460 ;
      LAYER via ;
        RECT 623.090 46.100 623.350 46.360 ;
        RECT 634.590 46.100 634.850 46.360 ;
        RECT 623.090 44.400 623.350 44.660 ;
      LAYER met2 ;
        RECT 623.090 46.070 623.350 46.390 ;
        RECT 634.590 46.070 634.850 46.390 ;
        RECT 623.150 44.690 623.290 46.070 ;
        RECT 623.090 44.370 623.350 44.690 ;
        RECT 634.650 34.520 634.790 46.070 ;
        RECT 634.580 32.120 634.930 34.520 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 652.590 32.120 652.870 34.520 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.050 32.120 147.330 34.520 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.900 32.120 171.250 34.520 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.840 32.120 189.190 34.520 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.850 32.120 207.130 34.520 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.330 32.120 224.610 34.520 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.270 32.120 242.550 34.520 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 338.850 50.330 339.105 50.905 ;
        RECT 338.935 49.600 339.105 50.330 ;
        RECT 338.850 48.695 339.105 49.600 ;
      LAYER L1M1_PR_C ;
        RECT 338.855 48.865 339.025 49.035 ;
      LAYER met1 ;
        RECT 338.780 49.020 339.100 49.080 ;
        RECT 338.585 48.880 339.100 49.020 ;
        RECT 338.780 48.820 339.100 48.880 ;
      LAYER via ;
        RECT 338.810 48.820 339.070 49.080 ;
      LAYER met2 ;
        RECT 260.140 49.275 260.420 49.645 ;
        RECT 338.800 49.275 339.080 49.645 ;
        RECT 260.210 34.520 260.350 49.275 ;
        RECT 338.870 49.110 339.010 49.275 ;
        RECT 338.810 48.790 339.070 49.110 ;
        RECT 260.140 32.120 260.490 34.520 ;
      LAYER via2 ;
        RECT 260.140 49.320 260.420 49.600 ;
        RECT 338.800 49.320 339.080 49.600 ;
      LAYER met3 ;
        RECT 260.115 49.610 260.445 49.625 ;
        RECT 338.775 49.610 339.105 49.625 ;
        RECT 260.115 49.310 339.105 49.610 ;
        RECT 260.115 49.295 260.445 49.310 ;
        RECT 338.775 49.295 339.105 49.310 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.810 32.120 58.090 34.520 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.730 32.120 82.010 34.520 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 284.130 32.120 284.410 34.520 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 295.610 46.795 297.270 46.995 ;
      LAYER L1M1_PR_C ;
        RECT 296.995 46.825 297.165 46.995 ;
      LAYER met1 ;
        RECT 296.935 46.795 297.225 47.025 ;
        RECT 297.010 46.640 297.150 46.795 ;
        RECT 301.520 46.640 301.840 46.700 ;
        RECT 297.010 46.500 301.840 46.640 ;
        RECT 301.520 46.440 301.840 46.500 ;
      LAYER via ;
        RECT 301.550 46.440 301.810 46.700 ;
      LAYER met2 ;
        RECT 301.550 46.410 301.810 46.730 ;
        RECT 301.610 34.520 301.750 46.410 ;
        RECT 301.540 32.120 301.890 34.520 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.550 32.120 319.830 34.520 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 380.425 46.635 380.945 48.185 ;
      LAYER L1M1_PR_C ;
        RECT 380.715 47.505 380.885 47.675 ;
      LAYER met1 ;
        RECT 339.240 47.660 339.560 47.720 ;
        RECT 380.655 47.660 380.945 47.705 ;
        RECT 339.240 47.520 380.945 47.660 ;
        RECT 339.240 47.460 339.560 47.520 ;
        RECT 380.655 47.475 380.945 47.520 ;
      LAYER via ;
        RECT 339.270 47.460 339.530 47.720 ;
      LAYER met2 ;
        RECT 339.270 47.430 339.530 47.750 ;
        RECT 339.330 46.810 339.470 47.430 ;
        RECT 337.490 46.670 339.470 46.810 ;
        RECT 337.490 34.520 337.630 46.670 ;
        RECT 337.420 32.120 337.770 34.520 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 355.340 50.720 355.660 50.780 ;
        RECT 366.840 50.720 367.160 50.780 ;
        RECT 355.340 50.580 367.160 50.720 ;
        RECT 355.340 50.520 355.660 50.580 ;
        RECT 366.840 50.520 367.160 50.580 ;
      LAYER via ;
        RECT 355.370 50.520 355.630 50.780 ;
        RECT 366.870 50.520 367.130 50.780 ;
      LAYER met2 ;
        RECT 366.930 50.810 367.070 54.000 ;
        RECT 355.370 50.490 355.630 50.810 ;
        RECT 366.870 50.490 367.130 50.810 ;
        RECT 355.430 34.520 355.570 50.490 ;
        RECT 355.360 32.120 355.710 34.520 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.370 32.120 373.650 34.520 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.850 32.120 391.130 34.520 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.790 32.120 409.070 34.520 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.660 32.120 427.010 34.520 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.670 32.120 444.950 34.520 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.650 32.120 105.930 34.520 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 464.605 46.635 465.125 48.185 ;
      LAYER L1M1_PR_C ;
        RECT 464.895 46.825 465.065 46.995 ;
      LAYER met1 ;
        RECT 462.060 46.980 462.380 47.040 ;
        RECT 464.835 46.980 465.125 47.025 ;
        RECT 462.060 46.840 465.125 46.980 ;
        RECT 462.060 46.780 462.380 46.840 ;
        RECT 464.835 46.795 465.125 46.840 ;
      LAYER via ;
        RECT 462.090 46.780 462.350 47.040 ;
      LAYER met2 ;
        RECT 462.090 46.750 462.350 47.070 ;
        RECT 462.150 34.520 462.290 46.750 ;
        RECT 462.080 32.120 462.430 34.520 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.090 32.120 480.370 34.520 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.030 32.120 498.310 34.520 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.900 32.120 516.250 34.520 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.910 32.120 534.190 34.520 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.320 32.120 551.670 34.520 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.330 32.120 569.610 34.520 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.270 32.120 587.550 34.520 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 604.905 48.695 605.425 50.245 ;
      LAYER L1M1_PR_C ;
        RECT 605.195 48.865 605.365 49.035 ;
      LAYER met1 ;
        RECT 605.120 49.020 605.440 49.080 ;
        RECT 604.925 48.880 605.440 49.020 ;
        RECT 605.120 48.820 605.440 48.880 ;
      LAYER via ;
        RECT 605.150 48.820 605.410 49.080 ;
      LAYER met2 ;
        RECT 605.150 48.790 605.410 49.110 ;
        RECT 605.210 34.520 605.350 48.790 ;
        RECT 605.140 32.120 605.490 34.520 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 623.150 32.120 623.430 34.520 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 175.955 47.355 176.290 48.115 ;
        RECT 176.810 47.355 177.140 48.115 ;
        RECT 175.955 47.185 177.625 47.355 ;
        RECT 177.380 46.620 177.625 47.185 ;
        RECT 175.955 46.450 177.625 46.620 ;
        RECT 175.955 46.025 176.290 46.450 ;
        RECT 176.810 46.025 177.145 46.450 ;
      LAYER L1M1_PR_C ;
        RECT 176.015 47.505 176.185 47.675 ;
      LAYER met1 ;
        RECT 174.100 47.660 174.420 47.720 ;
        RECT 175.955 47.660 176.245 47.705 ;
        RECT 174.100 47.520 176.245 47.660 ;
        RECT 174.100 47.460 174.420 47.520 ;
        RECT 175.955 47.475 176.245 47.520 ;
        RECT 130.860 46.980 131.180 47.040 ;
        RECT 140.520 46.980 140.840 47.040 ;
        RECT 130.860 46.840 140.840 46.980 ;
        RECT 130.860 46.780 131.180 46.840 ;
        RECT 140.520 46.780 140.840 46.840 ;
      LAYER via ;
        RECT 174.130 47.460 174.390 47.720 ;
        RECT 130.890 46.780 131.150 47.040 ;
        RECT 140.550 46.780 140.810 47.040 ;
      LAYER met2 ;
        RECT 173.270 48.170 173.410 54.000 ;
        RECT 173.270 48.030 174.330 48.170 ;
        RECT 174.190 47.750 174.330 48.030 ;
        RECT 174.130 47.430 174.390 47.750 ;
        RECT 130.890 46.750 131.150 47.070 ;
        RECT 140.550 46.750 140.810 47.070 ;
        RECT 130.950 37.970 131.090 46.750 ;
        RECT 140.610 46.245 140.750 46.750 ;
        RECT 174.190 46.245 174.330 47.430 ;
        RECT 140.540 45.875 140.820 46.245 ;
        RECT 174.120 45.875 174.400 46.245 ;
        RECT 129.110 37.830 131.090 37.970 ;
        RECT 129.110 34.520 129.250 37.830 ;
        RECT 129.040 32.120 129.390 34.520 ;
      LAYER via2 ;
        RECT 140.540 45.920 140.820 46.200 ;
        RECT 174.120 45.920 174.400 46.200 ;
      LAYER met3 ;
        RECT 140.515 46.210 140.845 46.225 ;
        RECT 174.095 46.210 174.425 46.225 ;
        RECT 140.515 45.910 174.425 46.210 ;
        RECT 140.515 45.895 140.845 45.910 ;
        RECT 174.095 45.895 174.425 45.910 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.630 32.120 640.910 34.520 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.570 32.120 658.850 34.520 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.030 32.120 153.310 34.520 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.880 32.120 177.230 34.520 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.890 32.120 195.170 34.520 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.300 41.795 212.580 42.165 ;
        RECT 212.370 34.520 212.510 41.795 ;
        RECT 212.300 32.120 212.650 34.520 ;
      LAYER via2 ;
        RECT 212.300 41.840 212.580 42.120 ;
      LAYER met3 ;
        RECT 212.275 42.130 212.605 42.145 ;
        RECT 214.780 42.130 215.160 42.140 ;
        RECT 212.275 41.830 215.160 42.130 ;
        RECT 212.275 41.815 212.605 41.830 ;
        RECT 214.780 41.820 215.160 41.830 ;
      LAYER via3 ;
        RECT 214.810 41.820 215.130 42.140 ;
      LAYER met4 ;
        RECT 214.820 42.145 215.120 54.000 ;
        RECT 214.805 41.815 215.135 42.145 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.310 32.120 230.590 34.520 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.250 32.120 248.530 34.520 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.120 32.120 266.470 34.520 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.710 34.520 87.850 54.000 ;
        RECT 87.640 32.120 87.990 34.520 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 290.110 32.120 290.390 34.520 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.590 32.120 307.870 34.520 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.530 32.120 325.810 34.520 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 298.760 53.440 299.080 53.500 ;
        RECT 298.760 53.300 328.430 53.440 ;
        RECT 298.760 53.240 299.080 53.300 ;
        RECT 328.290 53.100 328.430 53.300 ;
        RECT 340.160 53.100 340.480 53.160 ;
        RECT 328.290 52.960 340.480 53.100 ;
        RECT 340.160 52.900 340.480 52.960 ;
        RECT 340.160 49.360 340.480 49.420 ;
        RECT 340.160 49.220 343.610 49.360 ;
        RECT 340.160 49.160 340.480 49.220 ;
        RECT 343.470 49.080 343.610 49.220 ;
        RECT 343.380 48.820 343.700 49.080 ;
      LAYER via ;
        RECT 298.790 53.240 299.050 53.500 ;
        RECT 340.190 52.900 340.450 53.160 ;
        RECT 340.190 49.160 340.450 49.420 ;
        RECT 343.410 48.820 343.670 49.080 ;
      LAYER met2 ;
        RECT 298.850 53.530 298.990 54.000 ;
        RECT 298.790 53.210 299.050 53.530 ;
        RECT 340.190 52.870 340.450 53.190 ;
        RECT 340.250 49.450 340.390 52.870 ;
        RECT 340.190 49.130 340.450 49.450 ;
        RECT 343.410 48.790 343.670 49.110 ;
        RECT 343.470 34.520 343.610 48.790 ;
        RECT 343.400 32.120 343.750 34.520 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.410 32.120 361.690 34.520 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.890 34.520 379.030 54.000 ;
        RECT 378.820 32.120 379.170 34.520 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.830 32.120 397.110 34.520 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.770 32.120 415.050 34.520 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 436.545 46.635 437.065 48.185 ;
      LAYER L1M1_PR_C ;
        RECT 436.835 46.825 437.005 46.995 ;
      LAYER met1 ;
        RECT 432.620 46.980 432.940 47.040 ;
        RECT 436.775 46.980 437.065 47.025 ;
        RECT 432.620 46.840 437.065 46.980 ;
        RECT 432.620 46.780 432.940 46.840 ;
        RECT 436.775 46.795 437.065 46.840 ;
      LAYER via ;
        RECT 432.650 46.780 432.910 47.040 ;
      LAYER met2 ;
        RECT 432.650 46.750 432.910 47.070 ;
        RECT 432.710 34.520 432.850 46.750 ;
        RECT 432.640 32.120 432.990 34.520 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.650 32.120 450.930 34.520 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.630 32.120 111.910 34.520 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.060 32.120 468.410 34.520 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.070 32.120 486.350 34.520 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 504.010 32.120 504.290 34.520 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.880 32.120 522.230 34.520 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 539.890 32.120 540.170 34.520 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.370 32.120 557.650 34.520 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.310 32.120 575.590 34.520 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.180 32.120 593.530 34.520 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 611.190 32.120 611.470 34.520 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 628.600 32.120 628.950 34.520 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 135.000 39.160 135.320 39.220 ;
        RECT 154.320 39.160 154.640 39.220 ;
        RECT 135.000 39.020 154.640 39.160 ;
        RECT 135.000 38.960 135.320 39.020 ;
        RECT 154.320 38.960 154.640 39.020 ;
      LAYER via ;
        RECT 135.030 38.960 135.290 39.220 ;
        RECT 154.350 38.960 154.610 39.220 ;
      LAYER met2 ;
        RECT 153.490 50.210 153.630 54.000 ;
        RECT 153.490 50.070 154.550 50.210 ;
        RECT 154.410 39.250 154.550 50.070 ;
        RECT 135.030 38.930 135.290 39.250 ;
        RECT 154.350 38.930 154.610 39.250 ;
        RECT 135.090 34.520 135.230 38.930 ;
        RECT 135.020 32.120 135.370 34.520 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.610 32.120 646.890 34.520 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.550 32.120 664.830 34.520 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.010 32.120 159.290 34.520 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 174.100 51.740 174.420 51.800 ;
        RECT 182.840 51.740 183.160 51.800 ;
        RECT 174.100 51.600 183.160 51.740 ;
        RECT 174.100 51.540 174.420 51.600 ;
        RECT 182.840 51.540 183.160 51.600 ;
      LAYER via ;
        RECT 174.130 51.540 174.390 51.800 ;
        RECT 182.870 51.540 183.130 51.800 ;
      LAYER met2 ;
        RECT 174.190 51.830 174.330 54.000 ;
        RECT 174.130 51.510 174.390 51.830 ;
        RECT 182.870 51.510 183.130 51.830 ;
        RECT 182.930 34.520 183.070 51.510 ;
        RECT 182.860 32.120 183.210 34.520 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.870 32.120 201.150 34.520 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.280 32.120 218.630 34.520 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.290 32.120 236.570 34.520 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.160 32.120 254.510 34.520 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 272.100 32.120 272.450 34.520 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.620 32.120 93.970 34.520 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.610 32.120 117.890 34.520 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.070 32.120 141.350 34.520 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.990 32.120 165.270 34.520 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.790 32.120 64.070 34.520 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.770 32.120 70.050 34.520 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.000 28.000 30.000 3555.920 ;
        RECT 42.000 3549.720 44.000 3559.920 ;
        RECT 142.000 3549.720 144.000 3559.920 ;
        RECT 242.000 3549.720 244.000 3559.920 ;
        RECT 342.000 3549.720 344.000 3559.920 ;
        RECT 442.000 3549.720 444.000 3559.920 ;
        RECT 542.000 3549.720 544.000 3559.920 ;
        RECT 642.000 3549.720 644.000 3559.920 ;
        RECT 742.000 3549.720 744.000 3559.920 ;
        RECT 842.000 3549.720 844.000 3559.920 ;
        RECT 942.000 3549.720 944.000 3559.920 ;
        RECT 1042.000 3549.720 1044.000 3559.920 ;
        RECT 1142.000 3549.720 1144.000 3559.920 ;
        RECT 1242.000 3549.720 1244.000 3559.920 ;
        RECT 1342.000 3549.720 1344.000 3559.920 ;
        RECT 1442.000 3549.720 1444.000 3559.920 ;
        RECT 1542.000 3549.720 1544.000 3559.920 ;
        RECT 1642.000 3549.720 1644.000 3559.920 ;
        RECT 1742.000 3549.720 1744.000 3559.920 ;
        RECT 1842.000 3549.720 1844.000 3559.920 ;
        RECT 1942.000 3549.720 1944.000 3559.920 ;
        RECT 2042.000 3549.720 2044.000 3559.920 ;
        RECT 2142.000 3549.720 2144.000 3559.920 ;
        RECT 2242.000 3549.720 2244.000 3559.920 ;
        RECT 2342.000 3549.720 2344.000 3559.920 ;
        RECT 2442.000 3549.720 2444.000 3559.920 ;
        RECT 2542.000 3549.720 2544.000 3559.920 ;
        RECT 2642.000 3549.720 2644.000 3559.920 ;
        RECT 2742.000 3549.720 2744.000 3559.920 ;
        RECT 2842.000 3549.720 2844.000 3559.920 ;
        RECT 2942.000 3549.720 2944.000 3559.920 ;
        RECT 42.000 24.000 44.000 34.520 ;
        RECT 142.000 24.000 144.000 34.520 ;
        RECT 242.000 24.000 244.000 34.520 ;
        RECT 342.000 24.000 344.000 34.520 ;
        RECT 442.000 24.000 444.000 34.520 ;
        RECT 542.000 24.000 544.000 34.520 ;
        RECT 642.000 24.000 644.000 34.520 ;
        RECT 742.000 24.000 744.000 34.520 ;
        RECT 842.000 24.000 844.000 34.520 ;
        RECT 942.000 24.000 944.000 34.520 ;
        RECT 1042.000 24.000 1044.000 34.520 ;
        RECT 1142.000 24.000 1144.000 34.520 ;
        RECT 1242.000 24.000 1244.000 34.520 ;
        RECT 1342.000 24.000 1344.000 34.520 ;
        RECT 1442.000 24.000 1444.000 34.520 ;
        RECT 1542.000 24.000 1544.000 34.520 ;
        RECT 1642.000 24.000 1644.000 34.520 ;
        RECT 1742.000 24.000 1744.000 34.520 ;
        RECT 1842.000 24.000 1844.000 34.520 ;
        RECT 1942.000 24.000 1944.000 34.520 ;
        RECT 2042.000 24.000 2044.000 34.520 ;
        RECT 2142.000 24.000 2144.000 34.520 ;
        RECT 2242.000 24.000 2244.000 34.520 ;
        RECT 2342.000 24.000 2344.000 34.520 ;
        RECT 2442.000 24.000 2444.000 34.520 ;
        RECT 2542.000 24.000 2544.000 34.520 ;
        RECT 2642.000 24.000 2644.000 34.520 ;
        RECT 2742.000 24.000 2744.000 34.520 ;
        RECT 2842.000 24.000 2844.000 34.520 ;
        RECT 2942.000 24.000 2944.000 34.520 ;
        RECT 2964.580 28.000 2966.580 3555.920 ;
      LAYER M4M5_PR_C ;
        RECT 28.410 3554.330 29.590 3555.510 ;
        RECT 42.410 3554.330 43.590 3555.510 ;
        RECT 142.410 3554.330 143.590 3555.510 ;
        RECT 242.410 3554.330 243.590 3555.510 ;
        RECT 342.410 3554.330 343.590 3555.510 ;
        RECT 442.410 3554.330 443.590 3555.510 ;
        RECT 542.410 3554.330 543.590 3555.510 ;
        RECT 642.410 3554.330 643.590 3555.510 ;
        RECT 742.410 3554.330 743.590 3555.510 ;
        RECT 842.410 3554.330 843.590 3555.510 ;
        RECT 942.410 3554.330 943.590 3555.510 ;
        RECT 1042.410 3554.330 1043.590 3555.510 ;
        RECT 1142.410 3554.330 1143.590 3555.510 ;
        RECT 1242.410 3554.330 1243.590 3555.510 ;
        RECT 1342.410 3554.330 1343.590 3555.510 ;
        RECT 1442.410 3554.330 1443.590 3555.510 ;
        RECT 1542.410 3554.330 1543.590 3555.510 ;
        RECT 1642.410 3554.330 1643.590 3555.510 ;
        RECT 1742.410 3554.330 1743.590 3555.510 ;
        RECT 1842.410 3554.330 1843.590 3555.510 ;
        RECT 1942.410 3554.330 1943.590 3555.510 ;
        RECT 2042.410 3554.330 2043.590 3555.510 ;
        RECT 2142.410 3554.330 2143.590 3555.510 ;
        RECT 2242.410 3554.330 2243.590 3555.510 ;
        RECT 2342.410 3554.330 2343.590 3555.510 ;
        RECT 2442.410 3554.330 2443.590 3555.510 ;
        RECT 2542.410 3554.330 2543.590 3555.510 ;
        RECT 2642.410 3554.330 2643.590 3555.510 ;
        RECT 2742.410 3554.330 2743.590 3555.510 ;
        RECT 2842.410 3554.330 2843.590 3555.510 ;
        RECT 2942.410 3554.330 2943.590 3555.510 ;
        RECT 2964.990 3554.330 2966.170 3555.510 ;
        RECT 28.410 3442.410 29.590 3443.590 ;
        RECT 28.410 3342.410 29.590 3343.590 ;
        RECT 28.410 3242.410 29.590 3243.590 ;
        RECT 28.410 3142.410 29.590 3143.590 ;
        RECT 28.410 3042.410 29.590 3043.590 ;
        RECT 28.410 2942.410 29.590 2943.590 ;
        RECT 28.410 2842.410 29.590 2843.590 ;
        RECT 28.410 2742.410 29.590 2743.590 ;
        RECT 28.410 2642.410 29.590 2643.590 ;
        RECT 28.410 2542.410 29.590 2543.590 ;
        RECT 28.410 2442.410 29.590 2443.590 ;
        RECT 28.410 2342.410 29.590 2343.590 ;
        RECT 28.410 2242.410 29.590 2243.590 ;
        RECT 28.410 2142.410 29.590 2143.590 ;
        RECT 28.410 2042.410 29.590 2043.590 ;
        RECT 28.410 1942.410 29.590 1943.590 ;
        RECT 28.410 1842.410 29.590 1843.590 ;
        RECT 28.410 1742.410 29.590 1743.590 ;
        RECT 28.410 1642.410 29.590 1643.590 ;
        RECT 28.410 1542.410 29.590 1543.590 ;
        RECT 28.410 1442.410 29.590 1443.590 ;
        RECT 28.410 1342.410 29.590 1343.590 ;
        RECT 28.410 1242.410 29.590 1243.590 ;
        RECT 28.410 1142.410 29.590 1143.590 ;
        RECT 28.410 1042.410 29.590 1043.590 ;
        RECT 28.410 942.410 29.590 943.590 ;
        RECT 28.410 842.410 29.590 843.590 ;
        RECT 28.410 742.410 29.590 743.590 ;
        RECT 28.410 642.410 29.590 643.590 ;
        RECT 28.410 542.410 29.590 543.590 ;
        RECT 28.410 442.410 29.590 443.590 ;
        RECT 28.410 342.410 29.590 343.590 ;
        RECT 28.410 242.410 29.590 243.590 ;
        RECT 28.410 142.410 29.590 143.590 ;
        RECT 28.410 42.410 29.590 43.590 ;
        RECT 2964.990 3442.410 2966.170 3443.590 ;
        RECT 2964.990 3342.410 2966.170 3343.590 ;
        RECT 2964.990 3242.410 2966.170 3243.590 ;
        RECT 2964.990 3142.410 2966.170 3143.590 ;
        RECT 2964.990 3042.410 2966.170 3043.590 ;
        RECT 2964.990 2942.410 2966.170 2943.590 ;
        RECT 2964.990 2842.410 2966.170 2843.590 ;
        RECT 2964.990 2742.410 2966.170 2743.590 ;
        RECT 2964.990 2642.410 2966.170 2643.590 ;
        RECT 2964.990 2542.410 2966.170 2543.590 ;
        RECT 2964.990 2442.410 2966.170 2443.590 ;
        RECT 2964.990 2342.410 2966.170 2343.590 ;
        RECT 2964.990 2242.410 2966.170 2243.590 ;
        RECT 2964.990 2142.410 2966.170 2143.590 ;
        RECT 2964.990 2042.410 2966.170 2043.590 ;
        RECT 2964.990 1942.410 2966.170 1943.590 ;
        RECT 2964.990 1842.410 2966.170 1843.590 ;
        RECT 2964.990 1742.410 2966.170 1743.590 ;
        RECT 2964.990 1642.410 2966.170 1643.590 ;
        RECT 2964.990 1542.410 2966.170 1543.590 ;
        RECT 2964.990 1442.410 2966.170 1443.590 ;
        RECT 2964.990 1342.410 2966.170 1343.590 ;
        RECT 2964.990 1242.410 2966.170 1243.590 ;
        RECT 2964.990 1142.410 2966.170 1143.590 ;
        RECT 2964.990 1042.410 2966.170 1043.590 ;
        RECT 2964.990 942.410 2966.170 943.590 ;
        RECT 2964.990 842.410 2966.170 843.590 ;
        RECT 2964.990 742.410 2966.170 743.590 ;
        RECT 2964.990 642.410 2966.170 643.590 ;
        RECT 2964.990 542.410 2966.170 543.590 ;
        RECT 2964.990 442.410 2966.170 443.590 ;
        RECT 2964.990 342.410 2966.170 343.590 ;
        RECT 2964.990 242.410 2966.170 243.590 ;
        RECT 2964.990 142.410 2966.170 143.590 ;
        RECT 2964.990 42.410 2966.170 43.590 ;
        RECT 28.410 28.410 29.590 29.590 ;
        RECT 42.410 28.410 43.590 29.590 ;
        RECT 142.410 28.410 143.590 29.590 ;
        RECT 242.410 28.410 243.590 29.590 ;
        RECT 342.410 28.410 343.590 29.590 ;
        RECT 442.410 28.410 443.590 29.590 ;
        RECT 542.410 28.410 543.590 29.590 ;
        RECT 642.410 28.410 643.590 29.590 ;
        RECT 742.410 28.410 743.590 29.590 ;
        RECT 842.410 28.410 843.590 29.590 ;
        RECT 942.410 28.410 943.590 29.590 ;
        RECT 1042.410 28.410 1043.590 29.590 ;
        RECT 1142.410 28.410 1143.590 29.590 ;
        RECT 1242.410 28.410 1243.590 29.590 ;
        RECT 1342.410 28.410 1343.590 29.590 ;
        RECT 1442.410 28.410 1443.590 29.590 ;
        RECT 1542.410 28.410 1543.590 29.590 ;
        RECT 1642.410 28.410 1643.590 29.590 ;
        RECT 1742.410 28.410 1743.590 29.590 ;
        RECT 1842.410 28.410 1843.590 29.590 ;
        RECT 1942.410 28.410 1943.590 29.590 ;
        RECT 2042.410 28.410 2043.590 29.590 ;
        RECT 2142.410 28.410 2143.590 29.590 ;
        RECT 2242.410 28.410 2243.590 29.590 ;
        RECT 2342.410 28.410 2343.590 29.590 ;
        RECT 2442.410 28.410 2443.590 29.590 ;
        RECT 2542.410 28.410 2543.590 29.590 ;
        RECT 2642.410 28.410 2643.590 29.590 ;
        RECT 2742.410 28.410 2743.590 29.590 ;
        RECT 2842.410 28.410 2843.590 29.590 ;
        RECT 2942.410 28.410 2943.590 29.590 ;
        RECT 2964.990 28.410 2966.170 29.590 ;
      LAYER met5 ;
        RECT 28.000 3553.920 2966.580 3555.920 ;
        RECT 24.000 3442.000 39.880 3444.000 ;
        RECT 2955.080 3442.000 2970.580 3444.000 ;
        RECT 24.000 3342.000 39.880 3344.000 ;
        RECT 2955.080 3342.000 2970.580 3344.000 ;
        RECT 24.000 3242.000 39.880 3244.000 ;
        RECT 2955.080 3242.000 2970.580 3244.000 ;
        RECT 24.000 3142.000 39.880 3144.000 ;
        RECT 2955.080 3142.000 2970.580 3144.000 ;
        RECT 24.000 3042.000 39.880 3044.000 ;
        RECT 2955.080 3042.000 2970.580 3044.000 ;
        RECT 24.000 2942.000 39.880 2944.000 ;
        RECT 2955.080 2942.000 2970.580 2944.000 ;
        RECT 24.000 2842.000 39.880 2844.000 ;
        RECT 2955.080 2842.000 2970.580 2844.000 ;
        RECT 24.000 2742.000 39.880 2744.000 ;
        RECT 2955.080 2742.000 2970.580 2744.000 ;
        RECT 24.000 2642.000 39.880 2644.000 ;
        RECT 2955.080 2642.000 2970.580 2644.000 ;
        RECT 24.000 2542.000 39.880 2544.000 ;
        RECT 2955.080 2542.000 2970.580 2544.000 ;
        RECT 24.000 2442.000 39.880 2444.000 ;
        RECT 2955.080 2442.000 2970.580 2444.000 ;
        RECT 24.000 2342.000 39.880 2344.000 ;
        RECT 2955.080 2342.000 2970.580 2344.000 ;
        RECT 24.000 2242.000 39.880 2244.000 ;
        RECT 2955.080 2242.000 2970.580 2244.000 ;
        RECT 24.000 2142.000 39.880 2144.000 ;
        RECT 2955.080 2142.000 2970.580 2144.000 ;
        RECT 24.000 2042.000 39.880 2044.000 ;
        RECT 2955.080 2042.000 2970.580 2044.000 ;
        RECT 24.000 1942.000 39.880 1944.000 ;
        RECT 2955.080 1942.000 2970.580 1944.000 ;
        RECT 24.000 1842.000 39.880 1844.000 ;
        RECT 2955.080 1842.000 2970.580 1844.000 ;
        RECT 24.000 1742.000 39.880 1744.000 ;
        RECT 2955.080 1742.000 2970.580 1744.000 ;
        RECT 24.000 1642.000 39.880 1644.000 ;
        RECT 2955.080 1642.000 2970.580 1644.000 ;
        RECT 24.000 1542.000 39.880 1544.000 ;
        RECT 2955.080 1542.000 2970.580 1544.000 ;
        RECT 24.000 1442.000 39.880 1444.000 ;
        RECT 2955.080 1442.000 2970.580 1444.000 ;
        RECT 24.000 1342.000 39.880 1344.000 ;
        RECT 2955.080 1342.000 2970.580 1344.000 ;
        RECT 24.000 1242.000 39.880 1244.000 ;
        RECT 2955.080 1242.000 2970.580 1244.000 ;
        RECT 24.000 1142.000 39.880 1144.000 ;
        RECT 2955.080 1142.000 2970.580 1144.000 ;
        RECT 24.000 1042.000 39.880 1044.000 ;
        RECT 2955.080 1042.000 2970.580 1044.000 ;
        RECT 24.000 942.000 39.880 944.000 ;
        RECT 2955.080 942.000 2970.580 944.000 ;
        RECT 24.000 842.000 39.880 844.000 ;
        RECT 2955.080 842.000 2970.580 844.000 ;
        RECT 24.000 742.000 39.880 744.000 ;
        RECT 2955.080 742.000 2970.580 744.000 ;
        RECT 24.000 642.000 39.880 644.000 ;
        RECT 2955.080 642.000 2970.580 644.000 ;
        RECT 24.000 542.000 39.880 544.000 ;
        RECT 2955.080 542.000 2970.580 544.000 ;
        RECT 24.000 442.000 39.880 444.000 ;
        RECT 2955.080 442.000 2970.580 444.000 ;
        RECT 24.000 342.000 39.880 344.000 ;
        RECT 2955.080 342.000 2970.580 344.000 ;
        RECT 24.000 242.000 39.880 244.000 ;
        RECT 2955.080 242.000 2970.580 244.000 ;
        RECT 24.000 142.000 39.880 144.000 ;
        RECT 2955.080 142.000 2970.580 144.000 ;
        RECT 24.000 42.000 39.880 44.000 ;
        RECT 2955.080 42.000 2970.580 44.000 ;
        RECT 28.000 28.000 2966.580 30.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 24.000 24.000 26.000 3559.920 ;
        RECT 92.000 3549.720 94.000 3559.920 ;
        RECT 192.000 3549.720 194.000 3559.920 ;
        RECT 292.000 3549.720 294.000 3559.920 ;
        RECT 392.000 3549.720 394.000 3559.920 ;
        RECT 492.000 3549.720 494.000 3559.920 ;
        RECT 592.000 3549.720 594.000 3559.920 ;
        RECT 692.000 3549.720 694.000 3559.920 ;
        RECT 792.000 3549.720 794.000 3559.920 ;
        RECT 892.000 3549.720 894.000 3559.920 ;
        RECT 992.000 3549.720 994.000 3559.920 ;
        RECT 1092.000 3549.720 1094.000 3559.920 ;
        RECT 1192.000 3549.720 1194.000 3559.920 ;
        RECT 1292.000 3549.720 1294.000 3559.920 ;
        RECT 1392.000 3549.720 1394.000 3559.920 ;
        RECT 1492.000 3549.720 1494.000 3559.920 ;
        RECT 1592.000 3549.720 1594.000 3559.920 ;
        RECT 1692.000 3549.720 1694.000 3559.920 ;
        RECT 1792.000 3549.720 1794.000 3559.920 ;
        RECT 1892.000 3549.720 1894.000 3559.920 ;
        RECT 1992.000 3549.720 1994.000 3559.920 ;
        RECT 2092.000 3549.720 2094.000 3559.920 ;
        RECT 2192.000 3549.720 2194.000 3559.920 ;
        RECT 2292.000 3549.720 2294.000 3559.920 ;
        RECT 2392.000 3549.720 2394.000 3559.920 ;
        RECT 2492.000 3549.720 2494.000 3559.920 ;
        RECT 2592.000 3549.720 2594.000 3559.920 ;
        RECT 2692.000 3549.720 2694.000 3559.920 ;
        RECT 2792.000 3549.720 2794.000 3559.920 ;
        RECT 2892.000 3549.720 2894.000 3559.920 ;
        RECT 92.000 24.000 94.000 34.520 ;
        RECT 192.000 24.000 194.000 34.520 ;
        RECT 292.000 24.000 294.000 34.520 ;
        RECT 392.000 24.000 394.000 34.520 ;
        RECT 492.000 24.000 494.000 34.520 ;
        RECT 592.000 24.000 594.000 34.520 ;
        RECT 692.000 24.000 694.000 34.520 ;
        RECT 792.000 24.000 794.000 34.520 ;
        RECT 892.000 24.000 894.000 34.520 ;
        RECT 992.000 24.000 994.000 34.520 ;
        RECT 1092.000 24.000 1094.000 34.520 ;
        RECT 1192.000 24.000 1194.000 34.520 ;
        RECT 1292.000 24.000 1294.000 34.520 ;
        RECT 1392.000 24.000 1394.000 34.520 ;
        RECT 1492.000 24.000 1494.000 34.520 ;
        RECT 1592.000 24.000 1594.000 34.520 ;
        RECT 1692.000 24.000 1694.000 34.520 ;
        RECT 1792.000 24.000 1794.000 34.520 ;
        RECT 1892.000 24.000 1894.000 34.520 ;
        RECT 1992.000 24.000 1994.000 34.520 ;
        RECT 2092.000 24.000 2094.000 34.520 ;
        RECT 2192.000 24.000 2194.000 34.520 ;
        RECT 2292.000 24.000 2294.000 34.520 ;
        RECT 2392.000 24.000 2394.000 34.520 ;
        RECT 2492.000 24.000 2494.000 34.520 ;
        RECT 2592.000 24.000 2594.000 34.520 ;
        RECT 2692.000 24.000 2694.000 34.520 ;
        RECT 2792.000 24.000 2794.000 34.520 ;
        RECT 2892.000 24.000 2894.000 34.520 ;
        RECT 2968.580 24.000 2970.580 3559.920 ;
      LAYER M4M5_PR_C ;
        RECT 24.410 3558.330 25.590 3559.510 ;
        RECT 92.410 3558.330 93.590 3559.510 ;
        RECT 192.410 3558.330 193.590 3559.510 ;
        RECT 292.410 3558.330 293.590 3559.510 ;
        RECT 392.410 3558.330 393.590 3559.510 ;
        RECT 492.410 3558.330 493.590 3559.510 ;
        RECT 592.410 3558.330 593.590 3559.510 ;
        RECT 692.410 3558.330 693.590 3559.510 ;
        RECT 792.410 3558.330 793.590 3559.510 ;
        RECT 892.410 3558.330 893.590 3559.510 ;
        RECT 992.410 3558.330 993.590 3559.510 ;
        RECT 1092.410 3558.330 1093.590 3559.510 ;
        RECT 1192.410 3558.330 1193.590 3559.510 ;
        RECT 1292.410 3558.330 1293.590 3559.510 ;
        RECT 1392.410 3558.330 1393.590 3559.510 ;
        RECT 1492.410 3558.330 1493.590 3559.510 ;
        RECT 1592.410 3558.330 1593.590 3559.510 ;
        RECT 1692.410 3558.330 1693.590 3559.510 ;
        RECT 1792.410 3558.330 1793.590 3559.510 ;
        RECT 1892.410 3558.330 1893.590 3559.510 ;
        RECT 1992.410 3558.330 1993.590 3559.510 ;
        RECT 2092.410 3558.330 2093.590 3559.510 ;
        RECT 2192.410 3558.330 2193.590 3559.510 ;
        RECT 2292.410 3558.330 2293.590 3559.510 ;
        RECT 2392.410 3558.330 2393.590 3559.510 ;
        RECT 2492.410 3558.330 2493.590 3559.510 ;
        RECT 2592.410 3558.330 2593.590 3559.510 ;
        RECT 2692.410 3558.330 2693.590 3559.510 ;
        RECT 2792.410 3558.330 2793.590 3559.510 ;
        RECT 2892.410 3558.330 2893.590 3559.510 ;
        RECT 2968.990 3558.330 2970.170 3559.510 ;
        RECT 24.410 3492.410 25.590 3493.590 ;
        RECT 24.410 3392.410 25.590 3393.590 ;
        RECT 24.410 3292.410 25.590 3293.590 ;
        RECT 24.410 3192.410 25.590 3193.590 ;
        RECT 24.410 3092.410 25.590 3093.590 ;
        RECT 24.410 2992.410 25.590 2993.590 ;
        RECT 24.410 2892.410 25.590 2893.590 ;
        RECT 24.410 2792.410 25.590 2793.590 ;
        RECT 24.410 2692.410 25.590 2693.590 ;
        RECT 24.410 2592.410 25.590 2593.590 ;
        RECT 24.410 2492.410 25.590 2493.590 ;
        RECT 24.410 2392.410 25.590 2393.590 ;
        RECT 24.410 2292.410 25.590 2293.590 ;
        RECT 24.410 2192.410 25.590 2193.590 ;
        RECT 24.410 2092.410 25.590 2093.590 ;
        RECT 24.410 1992.410 25.590 1993.590 ;
        RECT 24.410 1892.410 25.590 1893.590 ;
        RECT 24.410 1792.410 25.590 1793.590 ;
        RECT 24.410 1692.410 25.590 1693.590 ;
        RECT 24.410 1592.410 25.590 1593.590 ;
        RECT 24.410 1492.410 25.590 1493.590 ;
        RECT 24.410 1392.410 25.590 1393.590 ;
        RECT 24.410 1292.410 25.590 1293.590 ;
        RECT 24.410 1192.410 25.590 1193.590 ;
        RECT 24.410 1092.410 25.590 1093.590 ;
        RECT 24.410 992.410 25.590 993.590 ;
        RECT 24.410 892.410 25.590 893.590 ;
        RECT 24.410 792.410 25.590 793.590 ;
        RECT 24.410 692.410 25.590 693.590 ;
        RECT 24.410 592.410 25.590 593.590 ;
        RECT 24.410 492.410 25.590 493.590 ;
        RECT 24.410 392.410 25.590 393.590 ;
        RECT 24.410 292.410 25.590 293.590 ;
        RECT 24.410 192.410 25.590 193.590 ;
        RECT 24.410 92.410 25.590 93.590 ;
        RECT 2968.990 3492.410 2970.170 3493.590 ;
        RECT 2968.990 3392.410 2970.170 3393.590 ;
        RECT 2968.990 3292.410 2970.170 3293.590 ;
        RECT 2968.990 3192.410 2970.170 3193.590 ;
        RECT 2968.990 3092.410 2970.170 3093.590 ;
        RECT 2968.990 2992.410 2970.170 2993.590 ;
        RECT 2968.990 2892.410 2970.170 2893.590 ;
        RECT 2968.990 2792.410 2970.170 2793.590 ;
        RECT 2968.990 2692.410 2970.170 2693.590 ;
        RECT 2968.990 2592.410 2970.170 2593.590 ;
        RECT 2968.990 2492.410 2970.170 2493.590 ;
        RECT 2968.990 2392.410 2970.170 2393.590 ;
        RECT 2968.990 2292.410 2970.170 2293.590 ;
        RECT 2968.990 2192.410 2970.170 2193.590 ;
        RECT 2968.990 2092.410 2970.170 2093.590 ;
        RECT 2968.990 1992.410 2970.170 1993.590 ;
        RECT 2968.990 1892.410 2970.170 1893.590 ;
        RECT 2968.990 1792.410 2970.170 1793.590 ;
        RECT 2968.990 1692.410 2970.170 1693.590 ;
        RECT 2968.990 1592.410 2970.170 1593.590 ;
        RECT 2968.990 1492.410 2970.170 1493.590 ;
        RECT 2968.990 1392.410 2970.170 1393.590 ;
        RECT 2968.990 1292.410 2970.170 1293.590 ;
        RECT 2968.990 1192.410 2970.170 1193.590 ;
        RECT 2968.990 1092.410 2970.170 1093.590 ;
        RECT 2968.990 992.410 2970.170 993.590 ;
        RECT 2968.990 892.410 2970.170 893.590 ;
        RECT 2968.990 792.410 2970.170 793.590 ;
        RECT 2968.990 692.410 2970.170 693.590 ;
        RECT 2968.990 592.410 2970.170 593.590 ;
        RECT 2968.990 492.410 2970.170 493.590 ;
        RECT 2968.990 392.410 2970.170 393.590 ;
        RECT 2968.990 292.410 2970.170 293.590 ;
        RECT 2968.990 192.410 2970.170 193.590 ;
        RECT 2968.990 92.410 2970.170 93.590 ;
        RECT 24.410 24.410 25.590 25.590 ;
        RECT 92.410 24.410 93.590 25.590 ;
        RECT 192.410 24.410 193.590 25.590 ;
        RECT 292.410 24.410 293.590 25.590 ;
        RECT 392.410 24.410 393.590 25.590 ;
        RECT 492.410 24.410 493.590 25.590 ;
        RECT 592.410 24.410 593.590 25.590 ;
        RECT 692.410 24.410 693.590 25.590 ;
        RECT 792.410 24.410 793.590 25.590 ;
        RECT 892.410 24.410 893.590 25.590 ;
        RECT 992.410 24.410 993.590 25.590 ;
        RECT 1092.410 24.410 1093.590 25.590 ;
        RECT 1192.410 24.410 1193.590 25.590 ;
        RECT 1292.410 24.410 1293.590 25.590 ;
        RECT 1392.410 24.410 1393.590 25.590 ;
        RECT 1492.410 24.410 1493.590 25.590 ;
        RECT 1592.410 24.410 1593.590 25.590 ;
        RECT 1692.410 24.410 1693.590 25.590 ;
        RECT 1792.410 24.410 1793.590 25.590 ;
        RECT 1892.410 24.410 1893.590 25.590 ;
        RECT 1992.410 24.410 1993.590 25.590 ;
        RECT 2092.410 24.410 2093.590 25.590 ;
        RECT 2192.410 24.410 2193.590 25.590 ;
        RECT 2292.410 24.410 2293.590 25.590 ;
        RECT 2392.410 24.410 2393.590 25.590 ;
        RECT 2492.410 24.410 2493.590 25.590 ;
        RECT 2592.410 24.410 2593.590 25.590 ;
        RECT 2692.410 24.410 2693.590 25.590 ;
        RECT 2792.410 24.410 2793.590 25.590 ;
        RECT 2892.410 24.410 2893.590 25.590 ;
        RECT 2968.990 24.410 2970.170 25.590 ;
      LAYER met5 ;
        RECT 24.000 3557.920 2970.580 3559.920 ;
        RECT 24.000 3492.000 39.880 3494.000 ;
        RECT 2955.080 3492.000 2970.580 3494.000 ;
        RECT 24.000 3392.000 39.880 3394.000 ;
        RECT 2955.080 3392.000 2970.580 3394.000 ;
        RECT 24.000 3292.000 39.880 3294.000 ;
        RECT 2955.080 3292.000 2970.580 3294.000 ;
        RECT 24.000 3192.000 39.880 3194.000 ;
        RECT 2955.080 3192.000 2970.580 3194.000 ;
        RECT 24.000 3092.000 39.880 3094.000 ;
        RECT 2955.080 3092.000 2970.580 3094.000 ;
        RECT 24.000 2992.000 39.880 2994.000 ;
        RECT 2955.080 2992.000 2970.580 2994.000 ;
        RECT 24.000 2892.000 39.880 2894.000 ;
        RECT 2955.080 2892.000 2970.580 2894.000 ;
        RECT 24.000 2792.000 39.880 2794.000 ;
        RECT 2955.080 2792.000 2970.580 2794.000 ;
        RECT 24.000 2692.000 39.880 2694.000 ;
        RECT 2955.080 2692.000 2970.580 2694.000 ;
        RECT 24.000 2592.000 39.880 2594.000 ;
        RECT 2955.080 2592.000 2970.580 2594.000 ;
        RECT 24.000 2492.000 39.880 2494.000 ;
        RECT 2955.080 2492.000 2970.580 2494.000 ;
        RECT 24.000 2392.000 39.880 2394.000 ;
        RECT 2955.080 2392.000 2970.580 2394.000 ;
        RECT 24.000 2292.000 39.880 2294.000 ;
        RECT 2955.080 2292.000 2970.580 2294.000 ;
        RECT 24.000 2192.000 39.880 2194.000 ;
        RECT 2955.080 2192.000 2970.580 2194.000 ;
        RECT 24.000 2092.000 39.880 2094.000 ;
        RECT 2955.080 2092.000 2970.580 2094.000 ;
        RECT 24.000 1992.000 39.880 1994.000 ;
        RECT 2955.080 1992.000 2970.580 1994.000 ;
        RECT 24.000 1892.000 39.880 1894.000 ;
        RECT 2955.080 1892.000 2970.580 1894.000 ;
        RECT 24.000 1792.000 39.880 1794.000 ;
        RECT 2955.080 1792.000 2970.580 1794.000 ;
        RECT 24.000 1692.000 39.880 1694.000 ;
        RECT 2955.080 1692.000 2970.580 1694.000 ;
        RECT 24.000 1592.000 39.880 1594.000 ;
        RECT 2955.080 1592.000 2970.580 1594.000 ;
        RECT 24.000 1492.000 39.880 1494.000 ;
        RECT 2955.080 1492.000 2970.580 1494.000 ;
        RECT 24.000 1392.000 39.880 1394.000 ;
        RECT 2955.080 1392.000 2970.580 1394.000 ;
        RECT 24.000 1292.000 39.880 1294.000 ;
        RECT 2955.080 1292.000 2970.580 1294.000 ;
        RECT 24.000 1192.000 39.880 1194.000 ;
        RECT 2955.080 1192.000 2970.580 1194.000 ;
        RECT 24.000 1092.000 39.880 1094.000 ;
        RECT 2955.080 1092.000 2970.580 1094.000 ;
        RECT 24.000 992.000 39.880 994.000 ;
        RECT 2955.080 992.000 2970.580 994.000 ;
        RECT 24.000 892.000 39.880 894.000 ;
        RECT 2955.080 892.000 2970.580 894.000 ;
        RECT 24.000 792.000 39.880 794.000 ;
        RECT 2955.080 792.000 2970.580 794.000 ;
        RECT 24.000 692.000 39.880 694.000 ;
        RECT 2955.080 692.000 2970.580 694.000 ;
        RECT 24.000 592.000 39.880 594.000 ;
        RECT 2955.080 592.000 2970.580 594.000 ;
        RECT 24.000 492.000 39.880 494.000 ;
        RECT 2955.080 492.000 2970.580 494.000 ;
        RECT 24.000 392.000 39.880 394.000 ;
        RECT 2955.080 392.000 2970.580 394.000 ;
        RECT 24.000 292.000 39.880 294.000 ;
        RECT 2955.080 292.000 2970.580 294.000 ;
        RECT 24.000 192.000 39.880 194.000 ;
        RECT 2955.080 192.000 2970.580 194.000 ;
        RECT 24.000 92.000 39.880 94.000 ;
        RECT 2955.080 92.000 2970.580 94.000 ;
        RECT 24.000 24.000 2970.580 26.000 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 20.000 20.000 22.000 3563.920 ;
        RECT 51.600 3549.720 53.600 3567.920 ;
        RECT 151.600 3549.720 153.600 3567.920 ;
        RECT 251.600 3549.720 253.600 3567.920 ;
        RECT 351.600 3549.720 353.600 3567.920 ;
        RECT 451.600 3549.720 453.600 3567.920 ;
        RECT 551.600 3549.720 553.600 3567.920 ;
        RECT 651.600 3549.720 653.600 3567.920 ;
        RECT 751.600 3549.720 753.600 3567.920 ;
        RECT 851.600 3549.720 853.600 3567.920 ;
        RECT 951.600 3549.720 953.600 3567.920 ;
        RECT 1051.600 3549.720 1053.600 3567.920 ;
        RECT 1151.600 3549.720 1153.600 3567.920 ;
        RECT 1251.600 3549.720 1253.600 3567.920 ;
        RECT 1351.600 3549.720 1353.600 3567.920 ;
        RECT 1451.600 3549.720 1453.600 3567.920 ;
        RECT 1551.600 3549.720 1553.600 3567.920 ;
        RECT 1651.600 3549.720 1653.600 3567.920 ;
        RECT 1751.600 3549.720 1753.600 3567.920 ;
        RECT 1851.600 3549.720 1853.600 3567.920 ;
        RECT 1951.600 3549.720 1953.600 3567.920 ;
        RECT 2051.600 3549.720 2053.600 3567.920 ;
        RECT 2151.600 3549.720 2153.600 3567.920 ;
        RECT 2251.600 3549.720 2253.600 3567.920 ;
        RECT 2351.600 3549.720 2353.600 3567.920 ;
        RECT 2451.600 3549.720 2453.600 3567.920 ;
        RECT 2551.600 3549.720 2553.600 3567.920 ;
        RECT 2651.600 3549.720 2653.600 3567.920 ;
        RECT 2751.600 3549.720 2753.600 3567.920 ;
        RECT 2851.600 3549.720 2853.600 3567.920 ;
        RECT 51.600 16.000 53.600 34.520 ;
        RECT 151.600 16.000 153.600 34.520 ;
        RECT 251.600 16.000 253.600 34.520 ;
        RECT 351.600 16.000 353.600 34.520 ;
        RECT 451.600 16.000 453.600 34.520 ;
        RECT 551.600 16.000 553.600 34.520 ;
        RECT 651.600 16.000 653.600 34.520 ;
        RECT 751.600 16.000 753.600 34.520 ;
        RECT 851.600 16.000 853.600 34.520 ;
        RECT 951.600 16.000 953.600 34.520 ;
        RECT 1051.600 16.000 1053.600 34.520 ;
        RECT 1151.600 16.000 1153.600 34.520 ;
        RECT 1251.600 16.000 1253.600 34.520 ;
        RECT 1351.600 16.000 1353.600 34.520 ;
        RECT 1451.600 16.000 1453.600 34.520 ;
        RECT 1551.600 16.000 1553.600 34.520 ;
        RECT 1651.600 16.000 1653.600 34.520 ;
        RECT 1751.600 16.000 1753.600 34.520 ;
        RECT 1851.600 16.000 1853.600 34.520 ;
        RECT 1951.600 16.000 1953.600 34.520 ;
        RECT 2051.600 16.000 2053.600 34.520 ;
        RECT 2151.600 16.000 2153.600 34.520 ;
        RECT 2251.600 16.000 2253.600 34.520 ;
        RECT 2351.600 16.000 2353.600 34.520 ;
        RECT 2451.600 16.000 2453.600 34.520 ;
        RECT 2551.600 16.000 2553.600 34.520 ;
        RECT 2651.600 16.000 2653.600 34.520 ;
        RECT 2751.600 16.000 2753.600 34.520 ;
        RECT 2851.600 16.000 2853.600 34.520 ;
        RECT 2972.580 20.000 2974.580 3563.920 ;
      LAYER M4M5_PR_C ;
        RECT 20.410 3562.330 21.590 3563.510 ;
        RECT 52.010 3562.330 53.190 3563.510 ;
        RECT 152.010 3562.330 153.190 3563.510 ;
        RECT 252.010 3562.330 253.190 3563.510 ;
        RECT 352.010 3562.330 353.190 3563.510 ;
        RECT 452.010 3562.330 453.190 3563.510 ;
        RECT 552.010 3562.330 553.190 3563.510 ;
        RECT 652.010 3562.330 653.190 3563.510 ;
        RECT 752.010 3562.330 753.190 3563.510 ;
        RECT 852.010 3562.330 853.190 3563.510 ;
        RECT 952.010 3562.330 953.190 3563.510 ;
        RECT 1052.010 3562.330 1053.190 3563.510 ;
        RECT 1152.010 3562.330 1153.190 3563.510 ;
        RECT 1252.010 3562.330 1253.190 3563.510 ;
        RECT 1352.010 3562.330 1353.190 3563.510 ;
        RECT 1452.010 3562.330 1453.190 3563.510 ;
        RECT 1552.010 3562.330 1553.190 3563.510 ;
        RECT 1652.010 3562.330 1653.190 3563.510 ;
        RECT 1752.010 3562.330 1753.190 3563.510 ;
        RECT 1852.010 3562.330 1853.190 3563.510 ;
        RECT 1952.010 3562.330 1953.190 3563.510 ;
        RECT 2052.010 3562.330 2053.190 3563.510 ;
        RECT 2152.010 3562.330 2153.190 3563.510 ;
        RECT 2252.010 3562.330 2253.190 3563.510 ;
        RECT 2352.010 3562.330 2353.190 3563.510 ;
        RECT 2452.010 3562.330 2453.190 3563.510 ;
        RECT 2552.010 3562.330 2553.190 3563.510 ;
        RECT 2652.010 3562.330 2653.190 3563.510 ;
        RECT 2752.010 3562.330 2753.190 3563.510 ;
        RECT 2852.010 3562.330 2853.190 3563.510 ;
        RECT 2972.990 3562.330 2974.170 3563.510 ;
        RECT 20.410 3452.010 21.590 3453.190 ;
        RECT 20.410 3352.010 21.590 3353.190 ;
        RECT 20.410 3252.010 21.590 3253.190 ;
        RECT 20.410 3152.010 21.590 3153.190 ;
        RECT 20.410 3052.010 21.590 3053.190 ;
        RECT 20.410 2952.010 21.590 2953.190 ;
        RECT 20.410 2852.010 21.590 2853.190 ;
        RECT 20.410 2752.010 21.590 2753.190 ;
        RECT 20.410 2652.010 21.590 2653.190 ;
        RECT 20.410 2552.010 21.590 2553.190 ;
        RECT 20.410 2452.010 21.590 2453.190 ;
        RECT 20.410 2352.010 21.590 2353.190 ;
        RECT 20.410 2252.010 21.590 2253.190 ;
        RECT 20.410 2152.010 21.590 2153.190 ;
        RECT 20.410 2052.010 21.590 2053.190 ;
        RECT 20.410 1952.010 21.590 1953.190 ;
        RECT 20.410 1852.010 21.590 1853.190 ;
        RECT 20.410 1752.010 21.590 1753.190 ;
        RECT 20.410 1652.010 21.590 1653.190 ;
        RECT 20.410 1552.010 21.590 1553.190 ;
        RECT 20.410 1452.010 21.590 1453.190 ;
        RECT 20.410 1352.010 21.590 1353.190 ;
        RECT 20.410 1252.010 21.590 1253.190 ;
        RECT 20.410 1152.010 21.590 1153.190 ;
        RECT 20.410 1052.010 21.590 1053.190 ;
        RECT 20.410 952.010 21.590 953.190 ;
        RECT 20.410 852.010 21.590 853.190 ;
        RECT 20.410 752.010 21.590 753.190 ;
        RECT 20.410 652.010 21.590 653.190 ;
        RECT 20.410 552.010 21.590 553.190 ;
        RECT 20.410 452.010 21.590 453.190 ;
        RECT 20.410 352.010 21.590 353.190 ;
        RECT 20.410 252.010 21.590 253.190 ;
        RECT 20.410 152.010 21.590 153.190 ;
        RECT 20.410 52.010 21.590 53.190 ;
        RECT 2972.990 3452.010 2974.170 3453.190 ;
        RECT 2972.990 3352.010 2974.170 3353.190 ;
        RECT 2972.990 3252.010 2974.170 3253.190 ;
        RECT 2972.990 3152.010 2974.170 3153.190 ;
        RECT 2972.990 3052.010 2974.170 3053.190 ;
        RECT 2972.990 2952.010 2974.170 2953.190 ;
        RECT 2972.990 2852.010 2974.170 2853.190 ;
        RECT 2972.990 2752.010 2974.170 2753.190 ;
        RECT 2972.990 2652.010 2974.170 2653.190 ;
        RECT 2972.990 2552.010 2974.170 2553.190 ;
        RECT 2972.990 2452.010 2974.170 2453.190 ;
        RECT 2972.990 2352.010 2974.170 2353.190 ;
        RECT 2972.990 2252.010 2974.170 2253.190 ;
        RECT 2972.990 2152.010 2974.170 2153.190 ;
        RECT 2972.990 2052.010 2974.170 2053.190 ;
        RECT 2972.990 1952.010 2974.170 1953.190 ;
        RECT 2972.990 1852.010 2974.170 1853.190 ;
        RECT 2972.990 1752.010 2974.170 1753.190 ;
        RECT 2972.990 1652.010 2974.170 1653.190 ;
        RECT 2972.990 1552.010 2974.170 1553.190 ;
        RECT 2972.990 1452.010 2974.170 1453.190 ;
        RECT 2972.990 1352.010 2974.170 1353.190 ;
        RECT 2972.990 1252.010 2974.170 1253.190 ;
        RECT 2972.990 1152.010 2974.170 1153.190 ;
        RECT 2972.990 1052.010 2974.170 1053.190 ;
        RECT 2972.990 952.010 2974.170 953.190 ;
        RECT 2972.990 852.010 2974.170 853.190 ;
        RECT 2972.990 752.010 2974.170 753.190 ;
        RECT 2972.990 652.010 2974.170 653.190 ;
        RECT 2972.990 552.010 2974.170 553.190 ;
        RECT 2972.990 452.010 2974.170 453.190 ;
        RECT 2972.990 352.010 2974.170 353.190 ;
        RECT 2972.990 252.010 2974.170 253.190 ;
        RECT 2972.990 152.010 2974.170 153.190 ;
        RECT 2972.990 52.010 2974.170 53.190 ;
        RECT 20.410 20.410 21.590 21.590 ;
        RECT 52.010 20.410 53.190 21.590 ;
        RECT 152.010 20.410 153.190 21.590 ;
        RECT 252.010 20.410 253.190 21.590 ;
        RECT 352.010 20.410 353.190 21.590 ;
        RECT 452.010 20.410 453.190 21.590 ;
        RECT 552.010 20.410 553.190 21.590 ;
        RECT 652.010 20.410 653.190 21.590 ;
        RECT 752.010 20.410 753.190 21.590 ;
        RECT 852.010 20.410 853.190 21.590 ;
        RECT 952.010 20.410 953.190 21.590 ;
        RECT 1052.010 20.410 1053.190 21.590 ;
        RECT 1152.010 20.410 1153.190 21.590 ;
        RECT 1252.010 20.410 1253.190 21.590 ;
        RECT 1352.010 20.410 1353.190 21.590 ;
        RECT 1452.010 20.410 1453.190 21.590 ;
        RECT 1552.010 20.410 1553.190 21.590 ;
        RECT 1652.010 20.410 1653.190 21.590 ;
        RECT 1752.010 20.410 1753.190 21.590 ;
        RECT 1852.010 20.410 1853.190 21.590 ;
        RECT 1952.010 20.410 1953.190 21.590 ;
        RECT 2052.010 20.410 2053.190 21.590 ;
        RECT 2152.010 20.410 2153.190 21.590 ;
        RECT 2252.010 20.410 2253.190 21.590 ;
        RECT 2352.010 20.410 2353.190 21.590 ;
        RECT 2452.010 20.410 2453.190 21.590 ;
        RECT 2552.010 20.410 2553.190 21.590 ;
        RECT 2652.010 20.410 2653.190 21.590 ;
        RECT 2752.010 20.410 2753.190 21.590 ;
        RECT 2852.010 20.410 2853.190 21.590 ;
        RECT 2972.990 20.410 2974.170 21.590 ;
      LAYER met5 ;
        RECT 20.000 3561.920 2974.580 3563.920 ;
        RECT 16.000 3451.600 39.880 3453.600 ;
        RECT 2955.080 3451.600 2978.580 3453.600 ;
        RECT 16.000 3351.600 39.880 3353.600 ;
        RECT 2955.080 3351.600 2978.580 3353.600 ;
        RECT 16.000 3251.600 39.880 3253.600 ;
        RECT 2955.080 3251.600 2978.580 3253.600 ;
        RECT 16.000 3151.600 39.880 3153.600 ;
        RECT 2955.080 3151.600 2978.580 3153.600 ;
        RECT 16.000 3051.600 39.880 3053.600 ;
        RECT 2955.080 3051.600 2978.580 3053.600 ;
        RECT 16.000 2951.600 39.880 2953.600 ;
        RECT 2955.080 2951.600 2978.580 2953.600 ;
        RECT 16.000 2851.600 39.880 2853.600 ;
        RECT 2955.080 2851.600 2978.580 2853.600 ;
        RECT 16.000 2751.600 39.880 2753.600 ;
        RECT 2955.080 2751.600 2978.580 2753.600 ;
        RECT 16.000 2651.600 39.880 2653.600 ;
        RECT 2955.080 2651.600 2978.580 2653.600 ;
        RECT 16.000 2551.600 39.880 2553.600 ;
        RECT 2955.080 2551.600 2978.580 2553.600 ;
        RECT 16.000 2451.600 39.880 2453.600 ;
        RECT 2955.080 2451.600 2978.580 2453.600 ;
        RECT 16.000 2351.600 39.880 2353.600 ;
        RECT 2955.080 2351.600 2978.580 2353.600 ;
        RECT 16.000 2251.600 39.880 2253.600 ;
        RECT 2955.080 2251.600 2978.580 2253.600 ;
        RECT 16.000 2151.600 39.880 2153.600 ;
        RECT 2955.080 2151.600 2978.580 2153.600 ;
        RECT 16.000 2051.600 39.880 2053.600 ;
        RECT 2955.080 2051.600 2978.580 2053.600 ;
        RECT 16.000 1951.600 39.880 1953.600 ;
        RECT 2955.080 1951.600 2978.580 1953.600 ;
        RECT 16.000 1851.600 39.880 1853.600 ;
        RECT 2955.080 1851.600 2978.580 1853.600 ;
        RECT 16.000 1751.600 39.880 1753.600 ;
        RECT 2955.080 1751.600 2978.580 1753.600 ;
        RECT 16.000 1651.600 39.880 1653.600 ;
        RECT 2955.080 1651.600 2978.580 1653.600 ;
        RECT 16.000 1551.600 39.880 1553.600 ;
        RECT 2955.080 1551.600 2978.580 1553.600 ;
        RECT 16.000 1451.600 39.880 1453.600 ;
        RECT 2955.080 1451.600 2978.580 1453.600 ;
        RECT 16.000 1351.600 39.880 1353.600 ;
        RECT 2955.080 1351.600 2978.580 1353.600 ;
        RECT 16.000 1251.600 39.880 1253.600 ;
        RECT 2955.080 1251.600 2978.580 1253.600 ;
        RECT 16.000 1151.600 39.880 1153.600 ;
        RECT 2955.080 1151.600 2978.580 1153.600 ;
        RECT 16.000 1051.600 39.880 1053.600 ;
        RECT 2955.080 1051.600 2978.580 1053.600 ;
        RECT 16.000 951.600 39.880 953.600 ;
        RECT 2955.080 951.600 2978.580 953.600 ;
        RECT 16.000 851.600 39.880 853.600 ;
        RECT 2955.080 851.600 2978.580 853.600 ;
        RECT 16.000 751.600 39.880 753.600 ;
        RECT 2955.080 751.600 2978.580 753.600 ;
        RECT 16.000 651.600 39.880 653.600 ;
        RECT 2955.080 651.600 2978.580 653.600 ;
        RECT 16.000 551.600 39.880 553.600 ;
        RECT 2955.080 551.600 2978.580 553.600 ;
        RECT 16.000 451.600 39.880 453.600 ;
        RECT 2955.080 451.600 2978.580 453.600 ;
        RECT 16.000 351.600 39.880 353.600 ;
        RECT 2955.080 351.600 2978.580 353.600 ;
        RECT 16.000 251.600 39.880 253.600 ;
        RECT 2955.080 251.600 2978.580 253.600 ;
        RECT 16.000 151.600 39.880 153.600 ;
        RECT 2955.080 151.600 2978.580 153.600 ;
        RECT 16.000 51.600 39.880 53.600 ;
        RECT 2955.080 51.600 2978.580 53.600 ;
        RECT 20.000 20.000 2974.580 22.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 16.000 16.000 18.000 3567.920 ;
        RECT 101.600 3549.720 103.600 3567.920 ;
        RECT 201.600 3549.720 203.600 3567.920 ;
        RECT 301.600 3549.720 303.600 3567.920 ;
        RECT 401.600 3549.720 403.600 3567.920 ;
        RECT 501.600 3549.720 503.600 3567.920 ;
        RECT 601.600 3549.720 603.600 3567.920 ;
        RECT 701.600 3549.720 703.600 3567.920 ;
        RECT 801.600 3549.720 803.600 3567.920 ;
        RECT 901.600 3549.720 903.600 3567.920 ;
        RECT 1001.600 3549.720 1003.600 3567.920 ;
        RECT 1101.600 3549.720 1103.600 3567.920 ;
        RECT 1201.600 3549.720 1203.600 3567.920 ;
        RECT 1301.600 3549.720 1303.600 3567.920 ;
        RECT 1401.600 3549.720 1403.600 3567.920 ;
        RECT 1501.600 3549.720 1503.600 3567.920 ;
        RECT 1601.600 3549.720 1603.600 3567.920 ;
        RECT 1701.600 3549.720 1703.600 3567.920 ;
        RECT 1801.600 3549.720 1803.600 3567.920 ;
        RECT 1901.600 3549.720 1903.600 3567.920 ;
        RECT 2001.600 3549.720 2003.600 3567.920 ;
        RECT 2101.600 3549.720 2103.600 3567.920 ;
        RECT 2201.600 3549.720 2203.600 3567.920 ;
        RECT 2301.600 3549.720 2303.600 3567.920 ;
        RECT 2401.600 3549.720 2403.600 3567.920 ;
        RECT 2501.600 3549.720 2503.600 3567.920 ;
        RECT 2601.600 3549.720 2603.600 3567.920 ;
        RECT 2701.600 3549.720 2703.600 3567.920 ;
        RECT 2801.600 3549.720 2803.600 3567.920 ;
        RECT 2901.600 3549.720 2903.600 3567.920 ;
        RECT 101.600 16.000 103.600 34.520 ;
        RECT 201.600 16.000 203.600 34.520 ;
        RECT 301.600 16.000 303.600 34.520 ;
        RECT 401.600 16.000 403.600 34.520 ;
        RECT 501.600 16.000 503.600 34.520 ;
        RECT 601.600 16.000 603.600 34.520 ;
        RECT 701.600 16.000 703.600 34.520 ;
        RECT 801.600 16.000 803.600 34.520 ;
        RECT 901.600 16.000 903.600 34.520 ;
        RECT 1001.600 16.000 1003.600 34.520 ;
        RECT 1101.600 16.000 1103.600 34.520 ;
        RECT 1201.600 16.000 1203.600 34.520 ;
        RECT 1301.600 16.000 1303.600 34.520 ;
        RECT 1401.600 16.000 1403.600 34.520 ;
        RECT 1501.600 16.000 1503.600 34.520 ;
        RECT 1601.600 16.000 1603.600 34.520 ;
        RECT 1701.600 16.000 1703.600 34.520 ;
        RECT 1801.600 16.000 1803.600 34.520 ;
        RECT 1901.600 16.000 1903.600 34.520 ;
        RECT 2001.600 16.000 2003.600 34.520 ;
        RECT 2101.600 16.000 2103.600 34.520 ;
        RECT 2201.600 16.000 2203.600 34.520 ;
        RECT 2301.600 16.000 2303.600 34.520 ;
        RECT 2401.600 16.000 2403.600 34.520 ;
        RECT 2501.600 16.000 2503.600 34.520 ;
        RECT 2601.600 16.000 2603.600 34.520 ;
        RECT 2701.600 16.000 2703.600 34.520 ;
        RECT 2801.600 16.000 2803.600 34.520 ;
        RECT 2901.600 16.000 2903.600 34.520 ;
        RECT 2976.580 16.000 2978.580 3567.920 ;
      LAYER M4M5_PR_C ;
        RECT 16.410 3566.330 17.590 3567.510 ;
        RECT 102.010 3566.330 103.190 3567.510 ;
        RECT 202.010 3566.330 203.190 3567.510 ;
        RECT 302.010 3566.330 303.190 3567.510 ;
        RECT 402.010 3566.330 403.190 3567.510 ;
        RECT 502.010 3566.330 503.190 3567.510 ;
        RECT 602.010 3566.330 603.190 3567.510 ;
        RECT 702.010 3566.330 703.190 3567.510 ;
        RECT 802.010 3566.330 803.190 3567.510 ;
        RECT 902.010 3566.330 903.190 3567.510 ;
        RECT 1002.010 3566.330 1003.190 3567.510 ;
        RECT 1102.010 3566.330 1103.190 3567.510 ;
        RECT 1202.010 3566.330 1203.190 3567.510 ;
        RECT 1302.010 3566.330 1303.190 3567.510 ;
        RECT 1402.010 3566.330 1403.190 3567.510 ;
        RECT 1502.010 3566.330 1503.190 3567.510 ;
        RECT 1602.010 3566.330 1603.190 3567.510 ;
        RECT 1702.010 3566.330 1703.190 3567.510 ;
        RECT 1802.010 3566.330 1803.190 3567.510 ;
        RECT 1902.010 3566.330 1903.190 3567.510 ;
        RECT 2002.010 3566.330 2003.190 3567.510 ;
        RECT 2102.010 3566.330 2103.190 3567.510 ;
        RECT 2202.010 3566.330 2203.190 3567.510 ;
        RECT 2302.010 3566.330 2303.190 3567.510 ;
        RECT 2402.010 3566.330 2403.190 3567.510 ;
        RECT 2502.010 3566.330 2503.190 3567.510 ;
        RECT 2602.010 3566.330 2603.190 3567.510 ;
        RECT 2702.010 3566.330 2703.190 3567.510 ;
        RECT 2802.010 3566.330 2803.190 3567.510 ;
        RECT 2902.010 3566.330 2903.190 3567.510 ;
        RECT 2976.990 3566.330 2978.170 3567.510 ;
        RECT 16.410 3502.010 17.590 3503.190 ;
        RECT 16.410 3402.010 17.590 3403.190 ;
        RECT 16.410 3302.010 17.590 3303.190 ;
        RECT 16.410 3202.010 17.590 3203.190 ;
        RECT 16.410 3102.010 17.590 3103.190 ;
        RECT 16.410 3002.010 17.590 3003.190 ;
        RECT 16.410 2902.010 17.590 2903.190 ;
        RECT 16.410 2802.010 17.590 2803.190 ;
        RECT 16.410 2702.010 17.590 2703.190 ;
        RECT 16.410 2602.010 17.590 2603.190 ;
        RECT 16.410 2502.010 17.590 2503.190 ;
        RECT 16.410 2402.010 17.590 2403.190 ;
        RECT 16.410 2302.010 17.590 2303.190 ;
        RECT 16.410 2202.010 17.590 2203.190 ;
        RECT 16.410 2102.010 17.590 2103.190 ;
        RECT 16.410 2002.010 17.590 2003.190 ;
        RECT 16.410 1902.010 17.590 1903.190 ;
        RECT 16.410 1802.010 17.590 1803.190 ;
        RECT 16.410 1702.010 17.590 1703.190 ;
        RECT 16.410 1602.010 17.590 1603.190 ;
        RECT 16.410 1502.010 17.590 1503.190 ;
        RECT 16.410 1402.010 17.590 1403.190 ;
        RECT 16.410 1302.010 17.590 1303.190 ;
        RECT 16.410 1202.010 17.590 1203.190 ;
        RECT 16.410 1102.010 17.590 1103.190 ;
        RECT 16.410 1002.010 17.590 1003.190 ;
        RECT 16.410 902.010 17.590 903.190 ;
        RECT 16.410 802.010 17.590 803.190 ;
        RECT 16.410 702.010 17.590 703.190 ;
        RECT 16.410 602.010 17.590 603.190 ;
        RECT 16.410 502.010 17.590 503.190 ;
        RECT 16.410 402.010 17.590 403.190 ;
        RECT 16.410 302.010 17.590 303.190 ;
        RECT 16.410 202.010 17.590 203.190 ;
        RECT 16.410 102.010 17.590 103.190 ;
        RECT 2976.990 3502.010 2978.170 3503.190 ;
        RECT 2976.990 3402.010 2978.170 3403.190 ;
        RECT 2976.990 3302.010 2978.170 3303.190 ;
        RECT 2976.990 3202.010 2978.170 3203.190 ;
        RECT 2976.990 3102.010 2978.170 3103.190 ;
        RECT 2976.990 3002.010 2978.170 3003.190 ;
        RECT 2976.990 2902.010 2978.170 2903.190 ;
        RECT 2976.990 2802.010 2978.170 2803.190 ;
        RECT 2976.990 2702.010 2978.170 2703.190 ;
        RECT 2976.990 2602.010 2978.170 2603.190 ;
        RECT 2976.990 2502.010 2978.170 2503.190 ;
        RECT 2976.990 2402.010 2978.170 2403.190 ;
        RECT 2976.990 2302.010 2978.170 2303.190 ;
        RECT 2976.990 2202.010 2978.170 2203.190 ;
        RECT 2976.990 2102.010 2978.170 2103.190 ;
        RECT 2976.990 2002.010 2978.170 2003.190 ;
        RECT 2976.990 1902.010 2978.170 1903.190 ;
        RECT 2976.990 1802.010 2978.170 1803.190 ;
        RECT 2976.990 1702.010 2978.170 1703.190 ;
        RECT 2976.990 1602.010 2978.170 1603.190 ;
        RECT 2976.990 1502.010 2978.170 1503.190 ;
        RECT 2976.990 1402.010 2978.170 1403.190 ;
        RECT 2976.990 1302.010 2978.170 1303.190 ;
        RECT 2976.990 1202.010 2978.170 1203.190 ;
        RECT 2976.990 1102.010 2978.170 1103.190 ;
        RECT 2976.990 1002.010 2978.170 1003.190 ;
        RECT 2976.990 902.010 2978.170 903.190 ;
        RECT 2976.990 802.010 2978.170 803.190 ;
        RECT 2976.990 702.010 2978.170 703.190 ;
        RECT 2976.990 602.010 2978.170 603.190 ;
        RECT 2976.990 502.010 2978.170 503.190 ;
        RECT 2976.990 402.010 2978.170 403.190 ;
        RECT 2976.990 302.010 2978.170 303.190 ;
        RECT 2976.990 202.010 2978.170 203.190 ;
        RECT 2976.990 102.010 2978.170 103.190 ;
        RECT 16.410 16.410 17.590 17.590 ;
        RECT 102.010 16.410 103.190 17.590 ;
        RECT 202.010 16.410 203.190 17.590 ;
        RECT 302.010 16.410 303.190 17.590 ;
        RECT 402.010 16.410 403.190 17.590 ;
        RECT 502.010 16.410 503.190 17.590 ;
        RECT 602.010 16.410 603.190 17.590 ;
        RECT 702.010 16.410 703.190 17.590 ;
        RECT 802.010 16.410 803.190 17.590 ;
        RECT 902.010 16.410 903.190 17.590 ;
        RECT 1002.010 16.410 1003.190 17.590 ;
        RECT 1102.010 16.410 1103.190 17.590 ;
        RECT 1202.010 16.410 1203.190 17.590 ;
        RECT 1302.010 16.410 1303.190 17.590 ;
        RECT 1402.010 16.410 1403.190 17.590 ;
        RECT 1502.010 16.410 1503.190 17.590 ;
        RECT 1602.010 16.410 1603.190 17.590 ;
        RECT 1702.010 16.410 1703.190 17.590 ;
        RECT 1802.010 16.410 1803.190 17.590 ;
        RECT 1902.010 16.410 1903.190 17.590 ;
        RECT 2002.010 16.410 2003.190 17.590 ;
        RECT 2102.010 16.410 2103.190 17.590 ;
        RECT 2202.010 16.410 2203.190 17.590 ;
        RECT 2302.010 16.410 2303.190 17.590 ;
        RECT 2402.010 16.410 2403.190 17.590 ;
        RECT 2502.010 16.410 2503.190 17.590 ;
        RECT 2602.010 16.410 2603.190 17.590 ;
        RECT 2702.010 16.410 2703.190 17.590 ;
        RECT 2802.010 16.410 2803.190 17.590 ;
        RECT 2902.010 16.410 2903.190 17.590 ;
        RECT 2976.990 16.410 2978.170 17.590 ;
      LAYER met5 ;
        RECT 16.000 3565.920 2978.580 3567.920 ;
        RECT 16.000 3501.600 39.880 3503.600 ;
        RECT 2955.080 3501.600 2978.580 3503.600 ;
        RECT 16.000 3401.600 39.880 3403.600 ;
        RECT 2955.080 3401.600 2978.580 3403.600 ;
        RECT 16.000 3301.600 39.880 3303.600 ;
        RECT 2955.080 3301.600 2978.580 3303.600 ;
        RECT 16.000 3201.600 39.880 3203.600 ;
        RECT 2955.080 3201.600 2978.580 3203.600 ;
        RECT 16.000 3101.600 39.880 3103.600 ;
        RECT 2955.080 3101.600 2978.580 3103.600 ;
        RECT 16.000 3001.600 39.880 3003.600 ;
        RECT 2955.080 3001.600 2978.580 3003.600 ;
        RECT 16.000 2901.600 39.880 2903.600 ;
        RECT 2955.080 2901.600 2978.580 2903.600 ;
        RECT 16.000 2801.600 39.880 2803.600 ;
        RECT 2955.080 2801.600 2978.580 2803.600 ;
        RECT 16.000 2701.600 39.880 2703.600 ;
        RECT 2955.080 2701.600 2978.580 2703.600 ;
        RECT 16.000 2601.600 39.880 2603.600 ;
        RECT 2955.080 2601.600 2978.580 2603.600 ;
        RECT 16.000 2501.600 39.880 2503.600 ;
        RECT 2955.080 2501.600 2978.580 2503.600 ;
        RECT 16.000 2401.600 39.880 2403.600 ;
        RECT 2955.080 2401.600 2978.580 2403.600 ;
        RECT 16.000 2301.600 39.880 2303.600 ;
        RECT 2955.080 2301.600 2978.580 2303.600 ;
        RECT 16.000 2201.600 39.880 2203.600 ;
        RECT 2955.080 2201.600 2978.580 2203.600 ;
        RECT 16.000 2101.600 39.880 2103.600 ;
        RECT 2955.080 2101.600 2978.580 2103.600 ;
        RECT 16.000 2001.600 39.880 2003.600 ;
        RECT 2955.080 2001.600 2978.580 2003.600 ;
        RECT 16.000 1901.600 39.880 1903.600 ;
        RECT 2955.080 1901.600 2978.580 1903.600 ;
        RECT 16.000 1801.600 39.880 1803.600 ;
        RECT 2955.080 1801.600 2978.580 1803.600 ;
        RECT 16.000 1701.600 39.880 1703.600 ;
        RECT 2955.080 1701.600 2978.580 1703.600 ;
        RECT 16.000 1601.600 39.880 1603.600 ;
        RECT 2955.080 1601.600 2978.580 1603.600 ;
        RECT 16.000 1501.600 39.880 1503.600 ;
        RECT 2955.080 1501.600 2978.580 1503.600 ;
        RECT 16.000 1401.600 39.880 1403.600 ;
        RECT 2955.080 1401.600 2978.580 1403.600 ;
        RECT 16.000 1301.600 39.880 1303.600 ;
        RECT 2955.080 1301.600 2978.580 1303.600 ;
        RECT 16.000 1201.600 39.880 1203.600 ;
        RECT 2955.080 1201.600 2978.580 1203.600 ;
        RECT 16.000 1101.600 39.880 1103.600 ;
        RECT 2955.080 1101.600 2978.580 1103.600 ;
        RECT 16.000 1001.600 39.880 1003.600 ;
        RECT 2955.080 1001.600 2978.580 1003.600 ;
        RECT 16.000 901.600 39.880 903.600 ;
        RECT 2955.080 901.600 2978.580 903.600 ;
        RECT 16.000 801.600 39.880 803.600 ;
        RECT 2955.080 801.600 2978.580 803.600 ;
        RECT 16.000 701.600 39.880 703.600 ;
        RECT 2955.080 701.600 2978.580 703.600 ;
        RECT 16.000 601.600 39.880 603.600 ;
        RECT 2955.080 601.600 2978.580 603.600 ;
        RECT 16.000 501.600 39.880 503.600 ;
        RECT 2955.080 501.600 2978.580 503.600 ;
        RECT 16.000 401.600 39.880 403.600 ;
        RECT 2955.080 401.600 2978.580 403.600 ;
        RECT 16.000 301.600 39.880 303.600 ;
        RECT 2955.080 301.600 2978.580 303.600 ;
        RECT 16.000 201.600 39.880 203.600 ;
        RECT 2955.080 201.600 2978.580 203.600 ;
        RECT 16.000 101.600 39.880 103.600 ;
        RECT 2955.080 101.600 2978.580 103.600 ;
        RECT 16.000 16.000 2978.580 18.000 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 12.000 12.000 14.000 3571.920 ;
        RECT 61.200 3549.720 63.200 3575.920 ;
        RECT 161.200 3549.720 163.200 3575.920 ;
        RECT 261.200 3549.720 263.200 3575.920 ;
        RECT 361.200 3549.720 363.200 3575.920 ;
        RECT 461.200 3549.720 463.200 3575.920 ;
        RECT 561.200 3549.720 563.200 3575.920 ;
        RECT 661.200 3549.720 663.200 3575.920 ;
        RECT 761.200 3549.720 763.200 3575.920 ;
        RECT 861.200 3549.720 863.200 3575.920 ;
        RECT 961.200 3549.720 963.200 3575.920 ;
        RECT 1061.200 3549.720 1063.200 3575.920 ;
        RECT 1161.200 3549.720 1163.200 3575.920 ;
        RECT 1261.200 3549.720 1263.200 3575.920 ;
        RECT 1361.200 3549.720 1363.200 3575.920 ;
        RECT 1461.200 3549.720 1463.200 3575.920 ;
        RECT 1561.200 3549.720 1563.200 3575.920 ;
        RECT 1661.200 3549.720 1663.200 3575.920 ;
        RECT 1761.200 3549.720 1763.200 3575.920 ;
        RECT 1861.200 3549.720 1863.200 3575.920 ;
        RECT 1961.200 3549.720 1963.200 3575.920 ;
        RECT 2061.200 3549.720 2063.200 3575.920 ;
        RECT 2161.200 3549.720 2163.200 3575.920 ;
        RECT 2261.200 3549.720 2263.200 3575.920 ;
        RECT 2361.200 3549.720 2363.200 3575.920 ;
        RECT 2461.200 3549.720 2463.200 3575.920 ;
        RECT 2561.200 3549.720 2563.200 3575.920 ;
        RECT 2661.200 3549.720 2663.200 3575.920 ;
        RECT 2761.200 3549.720 2763.200 3575.920 ;
        RECT 2861.200 3549.720 2863.200 3575.920 ;
        RECT 61.200 8.000 63.200 34.520 ;
        RECT 161.200 8.000 163.200 34.520 ;
        RECT 261.200 8.000 263.200 34.520 ;
        RECT 361.200 8.000 363.200 34.520 ;
        RECT 461.200 8.000 463.200 34.520 ;
        RECT 561.200 8.000 563.200 34.520 ;
        RECT 661.200 8.000 663.200 34.520 ;
        RECT 761.200 8.000 763.200 34.520 ;
        RECT 861.200 8.000 863.200 34.520 ;
        RECT 961.200 8.000 963.200 34.520 ;
        RECT 1061.200 8.000 1063.200 34.520 ;
        RECT 1161.200 8.000 1163.200 34.520 ;
        RECT 1261.200 8.000 1263.200 34.520 ;
        RECT 1361.200 8.000 1363.200 34.520 ;
        RECT 1461.200 8.000 1463.200 34.520 ;
        RECT 1561.200 8.000 1563.200 34.520 ;
        RECT 1661.200 8.000 1663.200 34.520 ;
        RECT 1761.200 8.000 1763.200 34.520 ;
        RECT 1861.200 8.000 1863.200 34.520 ;
        RECT 1961.200 8.000 1963.200 34.520 ;
        RECT 2061.200 8.000 2063.200 34.520 ;
        RECT 2161.200 8.000 2163.200 34.520 ;
        RECT 2261.200 8.000 2263.200 34.520 ;
        RECT 2361.200 8.000 2363.200 34.520 ;
        RECT 2461.200 8.000 2463.200 34.520 ;
        RECT 2561.200 8.000 2563.200 34.520 ;
        RECT 2661.200 8.000 2663.200 34.520 ;
        RECT 2761.200 8.000 2763.200 34.520 ;
        RECT 2861.200 8.000 2863.200 34.520 ;
        RECT 2980.580 12.000 2982.580 3571.920 ;
      LAYER M4M5_PR_C ;
        RECT 12.410 3570.330 13.590 3571.510 ;
        RECT 61.610 3570.330 62.790 3571.510 ;
        RECT 161.610 3570.330 162.790 3571.510 ;
        RECT 261.610 3570.330 262.790 3571.510 ;
        RECT 361.610 3570.330 362.790 3571.510 ;
        RECT 461.610 3570.330 462.790 3571.510 ;
        RECT 561.610 3570.330 562.790 3571.510 ;
        RECT 661.610 3570.330 662.790 3571.510 ;
        RECT 761.610 3570.330 762.790 3571.510 ;
        RECT 861.610 3570.330 862.790 3571.510 ;
        RECT 961.610 3570.330 962.790 3571.510 ;
        RECT 1061.610 3570.330 1062.790 3571.510 ;
        RECT 1161.610 3570.330 1162.790 3571.510 ;
        RECT 1261.610 3570.330 1262.790 3571.510 ;
        RECT 1361.610 3570.330 1362.790 3571.510 ;
        RECT 1461.610 3570.330 1462.790 3571.510 ;
        RECT 1561.610 3570.330 1562.790 3571.510 ;
        RECT 1661.610 3570.330 1662.790 3571.510 ;
        RECT 1761.610 3570.330 1762.790 3571.510 ;
        RECT 1861.610 3570.330 1862.790 3571.510 ;
        RECT 1961.610 3570.330 1962.790 3571.510 ;
        RECT 2061.610 3570.330 2062.790 3571.510 ;
        RECT 2161.610 3570.330 2162.790 3571.510 ;
        RECT 2261.610 3570.330 2262.790 3571.510 ;
        RECT 2361.610 3570.330 2362.790 3571.510 ;
        RECT 2461.610 3570.330 2462.790 3571.510 ;
        RECT 2561.610 3570.330 2562.790 3571.510 ;
        RECT 2661.610 3570.330 2662.790 3571.510 ;
        RECT 2761.610 3570.330 2762.790 3571.510 ;
        RECT 2861.610 3570.330 2862.790 3571.510 ;
        RECT 2980.990 3570.330 2982.170 3571.510 ;
        RECT 12.410 3461.610 13.590 3462.790 ;
        RECT 12.410 3361.610 13.590 3362.790 ;
        RECT 12.410 3261.610 13.590 3262.790 ;
        RECT 12.410 3161.610 13.590 3162.790 ;
        RECT 12.410 3061.610 13.590 3062.790 ;
        RECT 12.410 2961.610 13.590 2962.790 ;
        RECT 12.410 2861.610 13.590 2862.790 ;
        RECT 12.410 2761.610 13.590 2762.790 ;
        RECT 12.410 2661.610 13.590 2662.790 ;
        RECT 12.410 2561.610 13.590 2562.790 ;
        RECT 12.410 2461.610 13.590 2462.790 ;
        RECT 12.410 2361.610 13.590 2362.790 ;
        RECT 12.410 2261.610 13.590 2262.790 ;
        RECT 12.410 2161.610 13.590 2162.790 ;
        RECT 12.410 2061.610 13.590 2062.790 ;
        RECT 12.410 1961.610 13.590 1962.790 ;
        RECT 12.410 1861.610 13.590 1862.790 ;
        RECT 12.410 1761.610 13.590 1762.790 ;
        RECT 12.410 1661.610 13.590 1662.790 ;
        RECT 12.410 1561.610 13.590 1562.790 ;
        RECT 12.410 1461.610 13.590 1462.790 ;
        RECT 12.410 1361.610 13.590 1362.790 ;
        RECT 12.410 1261.610 13.590 1262.790 ;
        RECT 12.410 1161.610 13.590 1162.790 ;
        RECT 12.410 1061.610 13.590 1062.790 ;
        RECT 12.410 961.610 13.590 962.790 ;
        RECT 12.410 861.610 13.590 862.790 ;
        RECT 12.410 761.610 13.590 762.790 ;
        RECT 12.410 661.610 13.590 662.790 ;
        RECT 12.410 561.610 13.590 562.790 ;
        RECT 12.410 461.610 13.590 462.790 ;
        RECT 12.410 361.610 13.590 362.790 ;
        RECT 12.410 261.610 13.590 262.790 ;
        RECT 12.410 161.610 13.590 162.790 ;
        RECT 12.410 61.610 13.590 62.790 ;
        RECT 2980.990 3461.610 2982.170 3462.790 ;
        RECT 2980.990 3361.610 2982.170 3362.790 ;
        RECT 2980.990 3261.610 2982.170 3262.790 ;
        RECT 2980.990 3161.610 2982.170 3162.790 ;
        RECT 2980.990 3061.610 2982.170 3062.790 ;
        RECT 2980.990 2961.610 2982.170 2962.790 ;
        RECT 2980.990 2861.610 2982.170 2862.790 ;
        RECT 2980.990 2761.610 2982.170 2762.790 ;
        RECT 2980.990 2661.610 2982.170 2662.790 ;
        RECT 2980.990 2561.610 2982.170 2562.790 ;
        RECT 2980.990 2461.610 2982.170 2462.790 ;
        RECT 2980.990 2361.610 2982.170 2362.790 ;
        RECT 2980.990 2261.610 2982.170 2262.790 ;
        RECT 2980.990 2161.610 2982.170 2162.790 ;
        RECT 2980.990 2061.610 2982.170 2062.790 ;
        RECT 2980.990 1961.610 2982.170 1962.790 ;
        RECT 2980.990 1861.610 2982.170 1862.790 ;
        RECT 2980.990 1761.610 2982.170 1762.790 ;
        RECT 2980.990 1661.610 2982.170 1662.790 ;
        RECT 2980.990 1561.610 2982.170 1562.790 ;
        RECT 2980.990 1461.610 2982.170 1462.790 ;
        RECT 2980.990 1361.610 2982.170 1362.790 ;
        RECT 2980.990 1261.610 2982.170 1262.790 ;
        RECT 2980.990 1161.610 2982.170 1162.790 ;
        RECT 2980.990 1061.610 2982.170 1062.790 ;
        RECT 2980.990 961.610 2982.170 962.790 ;
        RECT 2980.990 861.610 2982.170 862.790 ;
        RECT 2980.990 761.610 2982.170 762.790 ;
        RECT 2980.990 661.610 2982.170 662.790 ;
        RECT 2980.990 561.610 2982.170 562.790 ;
        RECT 2980.990 461.610 2982.170 462.790 ;
        RECT 2980.990 361.610 2982.170 362.790 ;
        RECT 2980.990 261.610 2982.170 262.790 ;
        RECT 2980.990 161.610 2982.170 162.790 ;
        RECT 2980.990 61.610 2982.170 62.790 ;
        RECT 12.410 12.410 13.590 13.590 ;
        RECT 61.610 12.410 62.790 13.590 ;
        RECT 161.610 12.410 162.790 13.590 ;
        RECT 261.610 12.410 262.790 13.590 ;
        RECT 361.610 12.410 362.790 13.590 ;
        RECT 461.610 12.410 462.790 13.590 ;
        RECT 561.610 12.410 562.790 13.590 ;
        RECT 661.610 12.410 662.790 13.590 ;
        RECT 761.610 12.410 762.790 13.590 ;
        RECT 861.610 12.410 862.790 13.590 ;
        RECT 961.610 12.410 962.790 13.590 ;
        RECT 1061.610 12.410 1062.790 13.590 ;
        RECT 1161.610 12.410 1162.790 13.590 ;
        RECT 1261.610 12.410 1262.790 13.590 ;
        RECT 1361.610 12.410 1362.790 13.590 ;
        RECT 1461.610 12.410 1462.790 13.590 ;
        RECT 1561.610 12.410 1562.790 13.590 ;
        RECT 1661.610 12.410 1662.790 13.590 ;
        RECT 1761.610 12.410 1762.790 13.590 ;
        RECT 1861.610 12.410 1862.790 13.590 ;
        RECT 1961.610 12.410 1962.790 13.590 ;
        RECT 2061.610 12.410 2062.790 13.590 ;
        RECT 2161.610 12.410 2162.790 13.590 ;
        RECT 2261.610 12.410 2262.790 13.590 ;
        RECT 2361.610 12.410 2362.790 13.590 ;
        RECT 2461.610 12.410 2462.790 13.590 ;
        RECT 2561.610 12.410 2562.790 13.590 ;
        RECT 2661.610 12.410 2662.790 13.590 ;
        RECT 2761.610 12.410 2762.790 13.590 ;
        RECT 2861.610 12.410 2862.790 13.590 ;
        RECT 2980.990 12.410 2982.170 13.590 ;
      LAYER met5 ;
        RECT 12.000 3569.920 2982.580 3571.920 ;
        RECT 8.000 3461.200 39.880 3463.200 ;
        RECT 2955.080 3461.200 2986.580 3463.200 ;
        RECT 8.000 3361.200 39.880 3363.200 ;
        RECT 2955.080 3361.200 2986.580 3363.200 ;
        RECT 8.000 3261.200 39.880 3263.200 ;
        RECT 2955.080 3261.200 2986.580 3263.200 ;
        RECT 8.000 3161.200 39.880 3163.200 ;
        RECT 2955.080 3161.200 2986.580 3163.200 ;
        RECT 8.000 3061.200 39.880 3063.200 ;
        RECT 2955.080 3061.200 2986.580 3063.200 ;
        RECT 8.000 2961.200 39.880 2963.200 ;
        RECT 2955.080 2961.200 2986.580 2963.200 ;
        RECT 8.000 2861.200 39.880 2863.200 ;
        RECT 2955.080 2861.200 2986.580 2863.200 ;
        RECT 8.000 2761.200 39.880 2763.200 ;
        RECT 2955.080 2761.200 2986.580 2763.200 ;
        RECT 8.000 2661.200 39.880 2663.200 ;
        RECT 2955.080 2661.200 2986.580 2663.200 ;
        RECT 8.000 2561.200 39.880 2563.200 ;
        RECT 2955.080 2561.200 2986.580 2563.200 ;
        RECT 8.000 2461.200 39.880 2463.200 ;
        RECT 2955.080 2461.200 2986.580 2463.200 ;
        RECT 8.000 2361.200 39.880 2363.200 ;
        RECT 2955.080 2361.200 2986.580 2363.200 ;
        RECT 8.000 2261.200 39.880 2263.200 ;
        RECT 2955.080 2261.200 2986.580 2263.200 ;
        RECT 8.000 2161.200 39.880 2163.200 ;
        RECT 2955.080 2161.200 2986.580 2163.200 ;
        RECT 8.000 2061.200 39.880 2063.200 ;
        RECT 2955.080 2061.200 2986.580 2063.200 ;
        RECT 8.000 1961.200 39.880 1963.200 ;
        RECT 2955.080 1961.200 2986.580 1963.200 ;
        RECT 8.000 1861.200 39.880 1863.200 ;
        RECT 2955.080 1861.200 2986.580 1863.200 ;
        RECT 8.000 1761.200 39.880 1763.200 ;
        RECT 2955.080 1761.200 2986.580 1763.200 ;
        RECT 8.000 1661.200 39.880 1663.200 ;
        RECT 2955.080 1661.200 2986.580 1663.200 ;
        RECT 8.000 1561.200 39.880 1563.200 ;
        RECT 2955.080 1561.200 2986.580 1563.200 ;
        RECT 8.000 1461.200 39.880 1463.200 ;
        RECT 2955.080 1461.200 2986.580 1463.200 ;
        RECT 8.000 1361.200 39.880 1363.200 ;
        RECT 2955.080 1361.200 2986.580 1363.200 ;
        RECT 8.000 1261.200 39.880 1263.200 ;
        RECT 2955.080 1261.200 2986.580 1263.200 ;
        RECT 8.000 1161.200 39.880 1163.200 ;
        RECT 2955.080 1161.200 2986.580 1163.200 ;
        RECT 8.000 1061.200 39.880 1063.200 ;
        RECT 2955.080 1061.200 2986.580 1063.200 ;
        RECT 8.000 961.200 39.880 963.200 ;
        RECT 2955.080 961.200 2986.580 963.200 ;
        RECT 8.000 861.200 39.880 863.200 ;
        RECT 2955.080 861.200 2986.580 863.200 ;
        RECT 8.000 761.200 39.880 763.200 ;
        RECT 2955.080 761.200 2986.580 763.200 ;
        RECT 8.000 661.200 39.880 663.200 ;
        RECT 2955.080 661.200 2986.580 663.200 ;
        RECT 8.000 561.200 39.880 563.200 ;
        RECT 2955.080 561.200 2986.580 563.200 ;
        RECT 8.000 461.200 39.880 463.200 ;
        RECT 2955.080 461.200 2986.580 463.200 ;
        RECT 8.000 361.200 39.880 363.200 ;
        RECT 2955.080 361.200 2986.580 363.200 ;
        RECT 8.000 261.200 39.880 263.200 ;
        RECT 2955.080 261.200 2986.580 263.200 ;
        RECT 8.000 161.200 39.880 163.200 ;
        RECT 2955.080 161.200 2986.580 163.200 ;
        RECT 8.000 61.200 39.880 63.200 ;
        RECT 2955.080 61.200 2986.580 63.200 ;
        RECT 12.000 12.000 2982.580 14.000 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 8.000 8.000 10.000 3575.920 ;
        RECT 111.200 3549.720 113.200 3575.920 ;
        RECT 211.200 3549.720 213.200 3575.920 ;
        RECT 311.200 3549.720 313.200 3575.920 ;
        RECT 411.200 3549.720 413.200 3575.920 ;
        RECT 511.200 3549.720 513.200 3575.920 ;
        RECT 611.200 3549.720 613.200 3575.920 ;
        RECT 711.200 3549.720 713.200 3575.920 ;
        RECT 811.200 3549.720 813.200 3575.920 ;
        RECT 911.200 3549.720 913.200 3575.920 ;
        RECT 1011.200 3549.720 1013.200 3575.920 ;
        RECT 1111.200 3549.720 1113.200 3575.920 ;
        RECT 1211.200 3549.720 1213.200 3575.920 ;
        RECT 1311.200 3549.720 1313.200 3575.920 ;
        RECT 1411.200 3549.720 1413.200 3575.920 ;
        RECT 1511.200 3549.720 1513.200 3575.920 ;
        RECT 1611.200 3549.720 1613.200 3575.920 ;
        RECT 1711.200 3549.720 1713.200 3575.920 ;
        RECT 1811.200 3549.720 1813.200 3575.920 ;
        RECT 1911.200 3549.720 1913.200 3575.920 ;
        RECT 2011.200 3549.720 2013.200 3575.920 ;
        RECT 2111.200 3549.720 2113.200 3575.920 ;
        RECT 2211.200 3549.720 2213.200 3575.920 ;
        RECT 2311.200 3549.720 2313.200 3575.920 ;
        RECT 2411.200 3549.720 2413.200 3575.920 ;
        RECT 2511.200 3549.720 2513.200 3575.920 ;
        RECT 2611.200 3549.720 2613.200 3575.920 ;
        RECT 2711.200 3549.720 2713.200 3575.920 ;
        RECT 2811.200 3549.720 2813.200 3575.920 ;
        RECT 2911.200 3549.720 2913.200 3575.920 ;
        RECT 111.200 8.000 113.200 34.520 ;
        RECT 211.200 8.000 213.200 34.520 ;
        RECT 311.200 8.000 313.200 34.520 ;
        RECT 411.200 8.000 413.200 34.520 ;
        RECT 511.200 8.000 513.200 34.520 ;
        RECT 611.200 8.000 613.200 34.520 ;
        RECT 711.200 8.000 713.200 34.520 ;
        RECT 811.200 8.000 813.200 34.520 ;
        RECT 911.200 8.000 913.200 34.520 ;
        RECT 1011.200 8.000 1013.200 34.520 ;
        RECT 1111.200 8.000 1113.200 34.520 ;
        RECT 1211.200 8.000 1213.200 34.520 ;
        RECT 1311.200 8.000 1313.200 34.520 ;
        RECT 1411.200 8.000 1413.200 34.520 ;
        RECT 1511.200 8.000 1513.200 34.520 ;
        RECT 1611.200 8.000 1613.200 34.520 ;
        RECT 1711.200 8.000 1713.200 34.520 ;
        RECT 1811.200 8.000 1813.200 34.520 ;
        RECT 1911.200 8.000 1913.200 34.520 ;
        RECT 2011.200 8.000 2013.200 34.520 ;
        RECT 2111.200 8.000 2113.200 34.520 ;
        RECT 2211.200 8.000 2213.200 34.520 ;
        RECT 2311.200 8.000 2313.200 34.520 ;
        RECT 2411.200 8.000 2413.200 34.520 ;
        RECT 2511.200 8.000 2513.200 34.520 ;
        RECT 2611.200 8.000 2613.200 34.520 ;
        RECT 2711.200 8.000 2713.200 34.520 ;
        RECT 2811.200 8.000 2813.200 34.520 ;
        RECT 2911.200 8.000 2913.200 34.520 ;
        RECT 2984.580 8.000 2986.580 3575.920 ;
      LAYER M4M5_PR_C ;
        RECT 8.410 3574.330 9.590 3575.510 ;
        RECT 111.610 3574.330 112.790 3575.510 ;
        RECT 211.610 3574.330 212.790 3575.510 ;
        RECT 311.610 3574.330 312.790 3575.510 ;
        RECT 411.610 3574.330 412.790 3575.510 ;
        RECT 511.610 3574.330 512.790 3575.510 ;
        RECT 611.610 3574.330 612.790 3575.510 ;
        RECT 711.610 3574.330 712.790 3575.510 ;
        RECT 811.610 3574.330 812.790 3575.510 ;
        RECT 911.610 3574.330 912.790 3575.510 ;
        RECT 1011.610 3574.330 1012.790 3575.510 ;
        RECT 1111.610 3574.330 1112.790 3575.510 ;
        RECT 1211.610 3574.330 1212.790 3575.510 ;
        RECT 1311.610 3574.330 1312.790 3575.510 ;
        RECT 1411.610 3574.330 1412.790 3575.510 ;
        RECT 1511.610 3574.330 1512.790 3575.510 ;
        RECT 1611.610 3574.330 1612.790 3575.510 ;
        RECT 1711.610 3574.330 1712.790 3575.510 ;
        RECT 1811.610 3574.330 1812.790 3575.510 ;
        RECT 1911.610 3574.330 1912.790 3575.510 ;
        RECT 2011.610 3574.330 2012.790 3575.510 ;
        RECT 2111.610 3574.330 2112.790 3575.510 ;
        RECT 2211.610 3574.330 2212.790 3575.510 ;
        RECT 2311.610 3574.330 2312.790 3575.510 ;
        RECT 2411.610 3574.330 2412.790 3575.510 ;
        RECT 2511.610 3574.330 2512.790 3575.510 ;
        RECT 2611.610 3574.330 2612.790 3575.510 ;
        RECT 2711.610 3574.330 2712.790 3575.510 ;
        RECT 2811.610 3574.330 2812.790 3575.510 ;
        RECT 2911.610 3574.330 2912.790 3575.510 ;
        RECT 2984.990 3574.330 2986.170 3575.510 ;
        RECT 8.410 3511.610 9.590 3512.790 ;
        RECT 8.410 3411.610 9.590 3412.790 ;
        RECT 8.410 3311.610 9.590 3312.790 ;
        RECT 8.410 3211.610 9.590 3212.790 ;
        RECT 8.410 3111.610 9.590 3112.790 ;
        RECT 8.410 3011.610 9.590 3012.790 ;
        RECT 8.410 2911.610 9.590 2912.790 ;
        RECT 8.410 2811.610 9.590 2812.790 ;
        RECT 8.410 2711.610 9.590 2712.790 ;
        RECT 8.410 2611.610 9.590 2612.790 ;
        RECT 8.410 2511.610 9.590 2512.790 ;
        RECT 8.410 2411.610 9.590 2412.790 ;
        RECT 8.410 2311.610 9.590 2312.790 ;
        RECT 8.410 2211.610 9.590 2212.790 ;
        RECT 8.410 2111.610 9.590 2112.790 ;
        RECT 8.410 2011.610 9.590 2012.790 ;
        RECT 8.410 1911.610 9.590 1912.790 ;
        RECT 8.410 1811.610 9.590 1812.790 ;
        RECT 8.410 1711.610 9.590 1712.790 ;
        RECT 8.410 1611.610 9.590 1612.790 ;
        RECT 8.410 1511.610 9.590 1512.790 ;
        RECT 8.410 1411.610 9.590 1412.790 ;
        RECT 8.410 1311.610 9.590 1312.790 ;
        RECT 8.410 1211.610 9.590 1212.790 ;
        RECT 8.410 1111.610 9.590 1112.790 ;
        RECT 8.410 1011.610 9.590 1012.790 ;
        RECT 8.410 911.610 9.590 912.790 ;
        RECT 8.410 811.610 9.590 812.790 ;
        RECT 8.410 711.610 9.590 712.790 ;
        RECT 8.410 611.610 9.590 612.790 ;
        RECT 8.410 511.610 9.590 512.790 ;
        RECT 8.410 411.610 9.590 412.790 ;
        RECT 8.410 311.610 9.590 312.790 ;
        RECT 8.410 211.610 9.590 212.790 ;
        RECT 8.410 111.610 9.590 112.790 ;
        RECT 2984.990 3511.610 2986.170 3512.790 ;
        RECT 2984.990 3411.610 2986.170 3412.790 ;
        RECT 2984.990 3311.610 2986.170 3312.790 ;
        RECT 2984.990 3211.610 2986.170 3212.790 ;
        RECT 2984.990 3111.610 2986.170 3112.790 ;
        RECT 2984.990 3011.610 2986.170 3012.790 ;
        RECT 2984.990 2911.610 2986.170 2912.790 ;
        RECT 2984.990 2811.610 2986.170 2812.790 ;
        RECT 2984.990 2711.610 2986.170 2712.790 ;
        RECT 2984.990 2611.610 2986.170 2612.790 ;
        RECT 2984.990 2511.610 2986.170 2512.790 ;
        RECT 2984.990 2411.610 2986.170 2412.790 ;
        RECT 2984.990 2311.610 2986.170 2312.790 ;
        RECT 2984.990 2211.610 2986.170 2212.790 ;
        RECT 2984.990 2111.610 2986.170 2112.790 ;
        RECT 2984.990 2011.610 2986.170 2012.790 ;
        RECT 2984.990 1911.610 2986.170 1912.790 ;
        RECT 2984.990 1811.610 2986.170 1812.790 ;
        RECT 2984.990 1711.610 2986.170 1712.790 ;
        RECT 2984.990 1611.610 2986.170 1612.790 ;
        RECT 2984.990 1511.610 2986.170 1512.790 ;
        RECT 2984.990 1411.610 2986.170 1412.790 ;
        RECT 2984.990 1311.610 2986.170 1312.790 ;
        RECT 2984.990 1211.610 2986.170 1212.790 ;
        RECT 2984.990 1111.610 2986.170 1112.790 ;
        RECT 2984.990 1011.610 2986.170 1012.790 ;
        RECT 2984.990 911.610 2986.170 912.790 ;
        RECT 2984.990 811.610 2986.170 812.790 ;
        RECT 2984.990 711.610 2986.170 712.790 ;
        RECT 2984.990 611.610 2986.170 612.790 ;
        RECT 2984.990 511.610 2986.170 512.790 ;
        RECT 2984.990 411.610 2986.170 412.790 ;
        RECT 2984.990 311.610 2986.170 312.790 ;
        RECT 2984.990 211.610 2986.170 212.790 ;
        RECT 2984.990 111.610 2986.170 112.790 ;
        RECT 8.410 8.410 9.590 9.590 ;
        RECT 111.610 8.410 112.790 9.590 ;
        RECT 211.610 8.410 212.790 9.590 ;
        RECT 311.610 8.410 312.790 9.590 ;
        RECT 411.610 8.410 412.790 9.590 ;
        RECT 511.610 8.410 512.790 9.590 ;
        RECT 611.610 8.410 612.790 9.590 ;
        RECT 711.610 8.410 712.790 9.590 ;
        RECT 811.610 8.410 812.790 9.590 ;
        RECT 911.610 8.410 912.790 9.590 ;
        RECT 1011.610 8.410 1012.790 9.590 ;
        RECT 1111.610 8.410 1112.790 9.590 ;
        RECT 1211.610 8.410 1212.790 9.590 ;
        RECT 1311.610 8.410 1312.790 9.590 ;
        RECT 1411.610 8.410 1412.790 9.590 ;
        RECT 1511.610 8.410 1512.790 9.590 ;
        RECT 1611.610 8.410 1612.790 9.590 ;
        RECT 1711.610 8.410 1712.790 9.590 ;
        RECT 1811.610 8.410 1812.790 9.590 ;
        RECT 1911.610 8.410 1912.790 9.590 ;
        RECT 2011.610 8.410 2012.790 9.590 ;
        RECT 2111.610 8.410 2112.790 9.590 ;
        RECT 2211.610 8.410 2212.790 9.590 ;
        RECT 2311.610 8.410 2312.790 9.590 ;
        RECT 2411.610 8.410 2412.790 9.590 ;
        RECT 2511.610 8.410 2512.790 9.590 ;
        RECT 2611.610 8.410 2612.790 9.590 ;
        RECT 2711.610 8.410 2712.790 9.590 ;
        RECT 2811.610 8.410 2812.790 9.590 ;
        RECT 2911.610 8.410 2912.790 9.590 ;
        RECT 2984.990 8.410 2986.170 9.590 ;
      LAYER met5 ;
        RECT 8.000 3573.920 2986.580 3575.920 ;
        RECT 8.000 3511.200 39.880 3513.200 ;
        RECT 2955.080 3511.200 2986.580 3513.200 ;
        RECT 8.000 3411.200 39.880 3413.200 ;
        RECT 2955.080 3411.200 2986.580 3413.200 ;
        RECT 8.000 3311.200 39.880 3313.200 ;
        RECT 2955.080 3311.200 2986.580 3313.200 ;
        RECT 8.000 3211.200 39.880 3213.200 ;
        RECT 2955.080 3211.200 2986.580 3213.200 ;
        RECT 8.000 3111.200 39.880 3113.200 ;
        RECT 2955.080 3111.200 2986.580 3113.200 ;
        RECT 8.000 3011.200 39.880 3013.200 ;
        RECT 2955.080 3011.200 2986.580 3013.200 ;
        RECT 8.000 2911.200 39.880 2913.200 ;
        RECT 2955.080 2911.200 2986.580 2913.200 ;
        RECT 8.000 2811.200 39.880 2813.200 ;
        RECT 2955.080 2811.200 2986.580 2813.200 ;
        RECT 8.000 2711.200 39.880 2713.200 ;
        RECT 2955.080 2711.200 2986.580 2713.200 ;
        RECT 8.000 2611.200 39.880 2613.200 ;
        RECT 2955.080 2611.200 2986.580 2613.200 ;
        RECT 8.000 2511.200 39.880 2513.200 ;
        RECT 2955.080 2511.200 2986.580 2513.200 ;
        RECT 8.000 2411.200 39.880 2413.200 ;
        RECT 2955.080 2411.200 2986.580 2413.200 ;
        RECT 8.000 2311.200 39.880 2313.200 ;
        RECT 2955.080 2311.200 2986.580 2313.200 ;
        RECT 8.000 2211.200 39.880 2213.200 ;
        RECT 2955.080 2211.200 2986.580 2213.200 ;
        RECT 8.000 2111.200 39.880 2113.200 ;
        RECT 2955.080 2111.200 2986.580 2113.200 ;
        RECT 8.000 2011.200 39.880 2013.200 ;
        RECT 2955.080 2011.200 2986.580 2013.200 ;
        RECT 8.000 1911.200 39.880 1913.200 ;
        RECT 2955.080 1911.200 2986.580 1913.200 ;
        RECT 8.000 1811.200 39.880 1813.200 ;
        RECT 2955.080 1811.200 2986.580 1813.200 ;
        RECT 8.000 1711.200 39.880 1713.200 ;
        RECT 2955.080 1711.200 2986.580 1713.200 ;
        RECT 8.000 1611.200 39.880 1613.200 ;
        RECT 2955.080 1611.200 2986.580 1613.200 ;
        RECT 8.000 1511.200 39.880 1513.200 ;
        RECT 2955.080 1511.200 2986.580 1513.200 ;
        RECT 8.000 1411.200 39.880 1413.200 ;
        RECT 2955.080 1411.200 2986.580 1413.200 ;
        RECT 8.000 1311.200 39.880 1313.200 ;
        RECT 2955.080 1311.200 2986.580 1313.200 ;
        RECT 8.000 1211.200 39.880 1213.200 ;
        RECT 2955.080 1211.200 2986.580 1213.200 ;
        RECT 8.000 1111.200 39.880 1113.200 ;
        RECT 2955.080 1111.200 2986.580 1113.200 ;
        RECT 8.000 1011.200 39.880 1013.200 ;
        RECT 2955.080 1011.200 2986.580 1013.200 ;
        RECT 8.000 911.200 39.880 913.200 ;
        RECT 2955.080 911.200 2986.580 913.200 ;
        RECT 8.000 811.200 39.880 813.200 ;
        RECT 2955.080 811.200 2986.580 813.200 ;
        RECT 8.000 711.200 39.880 713.200 ;
        RECT 2955.080 711.200 2986.580 713.200 ;
        RECT 8.000 611.200 39.880 613.200 ;
        RECT 2955.080 611.200 2986.580 613.200 ;
        RECT 8.000 511.200 39.880 513.200 ;
        RECT 2955.080 511.200 2986.580 513.200 ;
        RECT 8.000 411.200 39.880 413.200 ;
        RECT 2955.080 411.200 2986.580 413.200 ;
        RECT 8.000 311.200 39.880 313.200 ;
        RECT 2955.080 311.200 2986.580 313.200 ;
        RECT 8.000 211.200 39.880 213.200 ;
        RECT 2955.080 211.200 2986.580 213.200 ;
        RECT 8.000 111.200 39.880 113.200 ;
        RECT 2955.080 111.200 2986.580 113.200 ;
        RECT 8.000 8.000 2986.580 10.000 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 4.000 4.000 6.000 3579.920 ;
        RECT 70.800 3549.720 72.800 3583.920 ;
        RECT 170.800 3549.720 172.800 3583.920 ;
        RECT 270.800 3549.720 272.800 3583.920 ;
        RECT 370.800 3549.720 372.800 3583.920 ;
        RECT 470.800 3549.720 472.800 3583.920 ;
        RECT 570.800 3549.720 572.800 3583.920 ;
        RECT 670.800 3549.720 672.800 3583.920 ;
        RECT 770.800 3549.720 772.800 3583.920 ;
        RECT 870.800 3549.720 872.800 3583.920 ;
        RECT 970.800 3549.720 972.800 3583.920 ;
        RECT 1070.800 3549.720 1072.800 3583.920 ;
        RECT 1170.800 3549.720 1172.800 3583.920 ;
        RECT 1270.800 3549.720 1272.800 3583.920 ;
        RECT 1370.800 3549.720 1372.800 3583.920 ;
        RECT 1470.800 3549.720 1472.800 3583.920 ;
        RECT 1570.800 3549.720 1572.800 3583.920 ;
        RECT 1670.800 3549.720 1672.800 3583.920 ;
        RECT 1770.800 3549.720 1772.800 3583.920 ;
        RECT 1870.800 3549.720 1872.800 3583.920 ;
        RECT 1970.800 3549.720 1972.800 3583.920 ;
        RECT 2070.800 3549.720 2072.800 3583.920 ;
        RECT 2170.800 3549.720 2172.800 3583.920 ;
        RECT 2270.800 3549.720 2272.800 3583.920 ;
        RECT 2370.800 3549.720 2372.800 3583.920 ;
        RECT 2470.800 3549.720 2472.800 3583.920 ;
        RECT 2570.800 3549.720 2572.800 3583.920 ;
        RECT 2670.800 3549.720 2672.800 3583.920 ;
        RECT 2770.800 3549.720 2772.800 3583.920 ;
        RECT 2870.800 3549.720 2872.800 3583.920 ;
        RECT 70.800 0.000 72.800 34.520 ;
        RECT 170.800 0.000 172.800 34.520 ;
        RECT 270.800 0.000 272.800 34.520 ;
        RECT 370.800 0.000 372.800 34.520 ;
        RECT 470.800 0.000 472.800 34.520 ;
        RECT 570.800 0.000 572.800 34.520 ;
        RECT 670.800 0.000 672.800 34.520 ;
        RECT 770.800 0.000 772.800 34.520 ;
        RECT 870.800 0.000 872.800 34.520 ;
        RECT 970.800 0.000 972.800 34.520 ;
        RECT 1070.800 0.000 1072.800 34.520 ;
        RECT 1170.800 0.000 1172.800 34.520 ;
        RECT 1270.800 0.000 1272.800 34.520 ;
        RECT 1370.800 0.000 1372.800 34.520 ;
        RECT 1470.800 0.000 1472.800 34.520 ;
        RECT 1570.800 0.000 1572.800 34.520 ;
        RECT 1670.800 0.000 1672.800 34.520 ;
        RECT 1770.800 0.000 1772.800 34.520 ;
        RECT 1870.800 0.000 1872.800 34.520 ;
        RECT 1970.800 0.000 1972.800 34.520 ;
        RECT 2070.800 0.000 2072.800 34.520 ;
        RECT 2170.800 0.000 2172.800 34.520 ;
        RECT 2270.800 0.000 2272.800 34.520 ;
        RECT 2370.800 0.000 2372.800 34.520 ;
        RECT 2470.800 0.000 2472.800 34.520 ;
        RECT 2570.800 0.000 2572.800 34.520 ;
        RECT 2670.800 0.000 2672.800 34.520 ;
        RECT 2770.800 0.000 2772.800 34.520 ;
        RECT 2870.800 0.000 2872.800 34.520 ;
        RECT 2988.580 4.000 2990.580 3579.920 ;
      LAYER M4M5_PR_C ;
        RECT 4.410 3578.330 5.590 3579.510 ;
        RECT 71.210 3578.330 72.390 3579.510 ;
        RECT 171.210 3578.330 172.390 3579.510 ;
        RECT 271.210 3578.330 272.390 3579.510 ;
        RECT 371.210 3578.330 372.390 3579.510 ;
        RECT 471.210 3578.330 472.390 3579.510 ;
        RECT 571.210 3578.330 572.390 3579.510 ;
        RECT 671.210 3578.330 672.390 3579.510 ;
        RECT 771.210 3578.330 772.390 3579.510 ;
        RECT 871.210 3578.330 872.390 3579.510 ;
        RECT 971.210 3578.330 972.390 3579.510 ;
        RECT 1071.210 3578.330 1072.390 3579.510 ;
        RECT 1171.210 3578.330 1172.390 3579.510 ;
        RECT 1271.210 3578.330 1272.390 3579.510 ;
        RECT 1371.210 3578.330 1372.390 3579.510 ;
        RECT 1471.210 3578.330 1472.390 3579.510 ;
        RECT 1571.210 3578.330 1572.390 3579.510 ;
        RECT 1671.210 3578.330 1672.390 3579.510 ;
        RECT 1771.210 3578.330 1772.390 3579.510 ;
        RECT 1871.210 3578.330 1872.390 3579.510 ;
        RECT 1971.210 3578.330 1972.390 3579.510 ;
        RECT 2071.210 3578.330 2072.390 3579.510 ;
        RECT 2171.210 3578.330 2172.390 3579.510 ;
        RECT 2271.210 3578.330 2272.390 3579.510 ;
        RECT 2371.210 3578.330 2372.390 3579.510 ;
        RECT 2471.210 3578.330 2472.390 3579.510 ;
        RECT 2571.210 3578.330 2572.390 3579.510 ;
        RECT 2671.210 3578.330 2672.390 3579.510 ;
        RECT 2771.210 3578.330 2772.390 3579.510 ;
        RECT 2871.210 3578.330 2872.390 3579.510 ;
        RECT 2988.990 3578.330 2990.170 3579.510 ;
        RECT 4.410 3471.210 5.590 3472.390 ;
        RECT 4.410 3371.210 5.590 3372.390 ;
        RECT 4.410 3271.210 5.590 3272.390 ;
        RECT 4.410 3171.210 5.590 3172.390 ;
        RECT 4.410 3071.210 5.590 3072.390 ;
        RECT 4.410 2971.210 5.590 2972.390 ;
        RECT 4.410 2871.210 5.590 2872.390 ;
        RECT 4.410 2771.210 5.590 2772.390 ;
        RECT 4.410 2671.210 5.590 2672.390 ;
        RECT 4.410 2571.210 5.590 2572.390 ;
        RECT 4.410 2471.210 5.590 2472.390 ;
        RECT 4.410 2371.210 5.590 2372.390 ;
        RECT 4.410 2271.210 5.590 2272.390 ;
        RECT 4.410 2171.210 5.590 2172.390 ;
        RECT 4.410 2071.210 5.590 2072.390 ;
        RECT 4.410 1971.210 5.590 1972.390 ;
        RECT 4.410 1871.210 5.590 1872.390 ;
        RECT 4.410 1771.210 5.590 1772.390 ;
        RECT 4.410 1671.210 5.590 1672.390 ;
        RECT 4.410 1571.210 5.590 1572.390 ;
        RECT 4.410 1471.210 5.590 1472.390 ;
        RECT 4.410 1371.210 5.590 1372.390 ;
        RECT 4.410 1271.210 5.590 1272.390 ;
        RECT 4.410 1171.210 5.590 1172.390 ;
        RECT 4.410 1071.210 5.590 1072.390 ;
        RECT 4.410 971.210 5.590 972.390 ;
        RECT 4.410 871.210 5.590 872.390 ;
        RECT 4.410 771.210 5.590 772.390 ;
        RECT 4.410 671.210 5.590 672.390 ;
        RECT 4.410 571.210 5.590 572.390 ;
        RECT 4.410 471.210 5.590 472.390 ;
        RECT 4.410 371.210 5.590 372.390 ;
        RECT 4.410 271.210 5.590 272.390 ;
        RECT 4.410 171.210 5.590 172.390 ;
        RECT 4.410 71.210 5.590 72.390 ;
        RECT 2988.990 3471.210 2990.170 3472.390 ;
        RECT 2988.990 3371.210 2990.170 3372.390 ;
        RECT 2988.990 3271.210 2990.170 3272.390 ;
        RECT 2988.990 3171.210 2990.170 3172.390 ;
        RECT 2988.990 3071.210 2990.170 3072.390 ;
        RECT 2988.990 2971.210 2990.170 2972.390 ;
        RECT 2988.990 2871.210 2990.170 2872.390 ;
        RECT 2988.990 2771.210 2990.170 2772.390 ;
        RECT 2988.990 2671.210 2990.170 2672.390 ;
        RECT 2988.990 2571.210 2990.170 2572.390 ;
        RECT 2988.990 2471.210 2990.170 2472.390 ;
        RECT 2988.990 2371.210 2990.170 2372.390 ;
        RECT 2988.990 2271.210 2990.170 2272.390 ;
        RECT 2988.990 2171.210 2990.170 2172.390 ;
        RECT 2988.990 2071.210 2990.170 2072.390 ;
        RECT 2988.990 1971.210 2990.170 1972.390 ;
        RECT 2988.990 1871.210 2990.170 1872.390 ;
        RECT 2988.990 1771.210 2990.170 1772.390 ;
        RECT 2988.990 1671.210 2990.170 1672.390 ;
        RECT 2988.990 1571.210 2990.170 1572.390 ;
        RECT 2988.990 1471.210 2990.170 1472.390 ;
        RECT 2988.990 1371.210 2990.170 1372.390 ;
        RECT 2988.990 1271.210 2990.170 1272.390 ;
        RECT 2988.990 1171.210 2990.170 1172.390 ;
        RECT 2988.990 1071.210 2990.170 1072.390 ;
        RECT 2988.990 971.210 2990.170 972.390 ;
        RECT 2988.990 871.210 2990.170 872.390 ;
        RECT 2988.990 771.210 2990.170 772.390 ;
        RECT 2988.990 671.210 2990.170 672.390 ;
        RECT 2988.990 571.210 2990.170 572.390 ;
        RECT 2988.990 471.210 2990.170 472.390 ;
        RECT 2988.990 371.210 2990.170 372.390 ;
        RECT 2988.990 271.210 2990.170 272.390 ;
        RECT 2988.990 171.210 2990.170 172.390 ;
        RECT 2988.990 71.210 2990.170 72.390 ;
        RECT 4.410 4.410 5.590 5.590 ;
        RECT 71.210 4.410 72.390 5.590 ;
        RECT 171.210 4.410 172.390 5.590 ;
        RECT 271.210 4.410 272.390 5.590 ;
        RECT 371.210 4.410 372.390 5.590 ;
        RECT 471.210 4.410 472.390 5.590 ;
        RECT 571.210 4.410 572.390 5.590 ;
        RECT 671.210 4.410 672.390 5.590 ;
        RECT 771.210 4.410 772.390 5.590 ;
        RECT 871.210 4.410 872.390 5.590 ;
        RECT 971.210 4.410 972.390 5.590 ;
        RECT 1071.210 4.410 1072.390 5.590 ;
        RECT 1171.210 4.410 1172.390 5.590 ;
        RECT 1271.210 4.410 1272.390 5.590 ;
        RECT 1371.210 4.410 1372.390 5.590 ;
        RECT 1471.210 4.410 1472.390 5.590 ;
        RECT 1571.210 4.410 1572.390 5.590 ;
        RECT 1671.210 4.410 1672.390 5.590 ;
        RECT 1771.210 4.410 1772.390 5.590 ;
        RECT 1871.210 4.410 1872.390 5.590 ;
        RECT 1971.210 4.410 1972.390 5.590 ;
        RECT 2071.210 4.410 2072.390 5.590 ;
        RECT 2171.210 4.410 2172.390 5.590 ;
        RECT 2271.210 4.410 2272.390 5.590 ;
        RECT 2371.210 4.410 2372.390 5.590 ;
        RECT 2471.210 4.410 2472.390 5.590 ;
        RECT 2571.210 4.410 2572.390 5.590 ;
        RECT 2671.210 4.410 2672.390 5.590 ;
        RECT 2771.210 4.410 2772.390 5.590 ;
        RECT 2871.210 4.410 2872.390 5.590 ;
        RECT 2988.990 4.410 2990.170 5.590 ;
      LAYER met5 ;
        RECT 4.000 3577.920 2990.580 3579.920 ;
        RECT 0.000 3470.800 39.880 3472.800 ;
        RECT 2955.080 3470.800 2994.580 3472.800 ;
        RECT 0.000 3370.800 39.880 3372.800 ;
        RECT 2955.080 3370.800 2994.580 3372.800 ;
        RECT 0.000 3270.800 39.880 3272.800 ;
        RECT 2955.080 3270.800 2994.580 3272.800 ;
        RECT 0.000 3170.800 39.880 3172.800 ;
        RECT 2955.080 3170.800 2994.580 3172.800 ;
        RECT 0.000 3070.800 39.880 3072.800 ;
        RECT 2955.080 3070.800 2994.580 3072.800 ;
        RECT 0.000 2970.800 39.880 2972.800 ;
        RECT 2955.080 2970.800 2994.580 2972.800 ;
        RECT 0.000 2870.800 39.880 2872.800 ;
        RECT 2955.080 2870.800 2994.580 2872.800 ;
        RECT 0.000 2770.800 39.880 2772.800 ;
        RECT 2955.080 2770.800 2994.580 2772.800 ;
        RECT 0.000 2670.800 39.880 2672.800 ;
        RECT 2955.080 2670.800 2994.580 2672.800 ;
        RECT 0.000 2570.800 39.880 2572.800 ;
        RECT 2955.080 2570.800 2994.580 2572.800 ;
        RECT 0.000 2470.800 39.880 2472.800 ;
        RECT 2955.080 2470.800 2994.580 2472.800 ;
        RECT 0.000 2370.800 39.880 2372.800 ;
        RECT 2955.080 2370.800 2994.580 2372.800 ;
        RECT 0.000 2270.800 39.880 2272.800 ;
        RECT 2955.080 2270.800 2994.580 2272.800 ;
        RECT 0.000 2170.800 39.880 2172.800 ;
        RECT 2955.080 2170.800 2994.580 2172.800 ;
        RECT 0.000 2070.800 39.880 2072.800 ;
        RECT 2955.080 2070.800 2994.580 2072.800 ;
        RECT 0.000 1970.800 39.880 1972.800 ;
        RECT 2955.080 1970.800 2994.580 1972.800 ;
        RECT 0.000 1870.800 39.880 1872.800 ;
        RECT 2955.080 1870.800 2994.580 1872.800 ;
        RECT 0.000 1770.800 39.880 1772.800 ;
        RECT 2955.080 1770.800 2994.580 1772.800 ;
        RECT 0.000 1670.800 39.880 1672.800 ;
        RECT 2955.080 1670.800 2994.580 1672.800 ;
        RECT 0.000 1570.800 39.880 1572.800 ;
        RECT 2955.080 1570.800 2994.580 1572.800 ;
        RECT 0.000 1470.800 39.880 1472.800 ;
        RECT 2955.080 1470.800 2994.580 1472.800 ;
        RECT 0.000 1370.800 39.880 1372.800 ;
        RECT 2955.080 1370.800 2994.580 1372.800 ;
        RECT 0.000 1270.800 39.880 1272.800 ;
        RECT 2955.080 1270.800 2994.580 1272.800 ;
        RECT 0.000 1170.800 39.880 1172.800 ;
        RECT 2955.080 1170.800 2994.580 1172.800 ;
        RECT 0.000 1070.800 39.880 1072.800 ;
        RECT 2955.080 1070.800 2994.580 1072.800 ;
        RECT 0.000 970.800 39.880 972.800 ;
        RECT 2955.080 970.800 2994.580 972.800 ;
        RECT 0.000 870.800 39.880 872.800 ;
        RECT 2955.080 870.800 2994.580 872.800 ;
        RECT 0.000 770.800 39.880 772.800 ;
        RECT 2955.080 770.800 2994.580 772.800 ;
        RECT 0.000 670.800 39.880 672.800 ;
        RECT 2955.080 670.800 2994.580 672.800 ;
        RECT 0.000 570.800 39.880 572.800 ;
        RECT 2955.080 570.800 2994.580 572.800 ;
        RECT 0.000 470.800 39.880 472.800 ;
        RECT 2955.080 470.800 2994.580 472.800 ;
        RECT 0.000 370.800 39.880 372.800 ;
        RECT 2955.080 370.800 2994.580 372.800 ;
        RECT 0.000 270.800 39.880 272.800 ;
        RECT 2955.080 270.800 2994.580 272.800 ;
        RECT 0.000 170.800 39.880 172.800 ;
        RECT 2955.080 170.800 2994.580 172.800 ;
        RECT 0.000 70.800 39.880 72.800 ;
        RECT 2955.080 70.800 2994.580 72.800 ;
        RECT 4.000 4.000 2990.580 6.000 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 2.000 3583.920 ;
        RECT 120.800 3549.720 122.800 3583.920 ;
        RECT 220.800 3549.720 222.800 3583.920 ;
        RECT 320.800 3549.720 322.800 3583.920 ;
        RECT 420.800 3549.720 422.800 3583.920 ;
        RECT 520.800 3549.720 522.800 3583.920 ;
        RECT 620.800 3549.720 622.800 3583.920 ;
        RECT 720.800 3549.720 722.800 3583.920 ;
        RECT 820.800 3549.720 822.800 3583.920 ;
        RECT 920.800 3549.720 922.800 3583.920 ;
        RECT 1020.800 3549.720 1022.800 3583.920 ;
        RECT 1120.800 3549.720 1122.800 3583.920 ;
        RECT 1220.800 3549.720 1222.800 3583.920 ;
        RECT 1320.800 3549.720 1322.800 3583.920 ;
        RECT 1420.800 3549.720 1422.800 3583.920 ;
        RECT 1520.800 3549.720 1522.800 3583.920 ;
        RECT 1620.800 3549.720 1622.800 3583.920 ;
        RECT 1720.800 3549.720 1722.800 3583.920 ;
        RECT 1820.800 3549.720 1822.800 3583.920 ;
        RECT 1920.800 3549.720 1922.800 3583.920 ;
        RECT 2020.800 3549.720 2022.800 3583.920 ;
        RECT 2120.800 3549.720 2122.800 3583.920 ;
        RECT 2220.800 3549.720 2222.800 3583.920 ;
        RECT 2320.800 3549.720 2322.800 3583.920 ;
        RECT 2420.800 3549.720 2422.800 3583.920 ;
        RECT 2520.800 3549.720 2522.800 3583.920 ;
        RECT 2620.800 3549.720 2622.800 3583.920 ;
        RECT 2720.800 3549.720 2722.800 3583.920 ;
        RECT 2820.800 3549.720 2822.800 3583.920 ;
        RECT 2920.800 3549.720 2922.800 3583.920 ;
        RECT 120.800 0.000 122.800 34.520 ;
        RECT 220.800 0.000 222.800 34.520 ;
        RECT 320.800 0.000 322.800 34.520 ;
        RECT 420.800 0.000 422.800 34.520 ;
        RECT 520.800 0.000 522.800 34.520 ;
        RECT 620.800 0.000 622.800 34.520 ;
        RECT 720.800 0.000 722.800 34.520 ;
        RECT 820.800 0.000 822.800 34.520 ;
        RECT 920.800 0.000 922.800 34.520 ;
        RECT 1020.800 0.000 1022.800 34.520 ;
        RECT 1120.800 0.000 1122.800 34.520 ;
        RECT 1220.800 0.000 1222.800 34.520 ;
        RECT 1320.800 0.000 1322.800 34.520 ;
        RECT 1420.800 0.000 1422.800 34.520 ;
        RECT 1520.800 0.000 1522.800 34.520 ;
        RECT 1620.800 0.000 1622.800 34.520 ;
        RECT 1720.800 0.000 1722.800 34.520 ;
        RECT 1820.800 0.000 1822.800 34.520 ;
        RECT 1920.800 0.000 1922.800 34.520 ;
        RECT 2020.800 0.000 2022.800 34.520 ;
        RECT 2120.800 0.000 2122.800 34.520 ;
        RECT 2220.800 0.000 2222.800 34.520 ;
        RECT 2320.800 0.000 2322.800 34.520 ;
        RECT 2420.800 0.000 2422.800 34.520 ;
        RECT 2520.800 0.000 2522.800 34.520 ;
        RECT 2620.800 0.000 2622.800 34.520 ;
        RECT 2720.800 0.000 2722.800 34.520 ;
        RECT 2820.800 0.000 2822.800 34.520 ;
        RECT 2920.800 0.000 2922.800 34.520 ;
        RECT 2992.580 0.000 2994.580 3583.920 ;
      LAYER M4M5_PR_C ;
        RECT 0.410 3582.330 1.590 3583.510 ;
        RECT 121.210 3582.330 122.390 3583.510 ;
        RECT 221.210 3582.330 222.390 3583.510 ;
        RECT 321.210 3582.330 322.390 3583.510 ;
        RECT 421.210 3582.330 422.390 3583.510 ;
        RECT 521.210 3582.330 522.390 3583.510 ;
        RECT 621.210 3582.330 622.390 3583.510 ;
        RECT 721.210 3582.330 722.390 3583.510 ;
        RECT 821.210 3582.330 822.390 3583.510 ;
        RECT 921.210 3582.330 922.390 3583.510 ;
        RECT 1021.210 3582.330 1022.390 3583.510 ;
        RECT 1121.210 3582.330 1122.390 3583.510 ;
        RECT 1221.210 3582.330 1222.390 3583.510 ;
        RECT 1321.210 3582.330 1322.390 3583.510 ;
        RECT 1421.210 3582.330 1422.390 3583.510 ;
        RECT 1521.210 3582.330 1522.390 3583.510 ;
        RECT 1621.210 3582.330 1622.390 3583.510 ;
        RECT 1721.210 3582.330 1722.390 3583.510 ;
        RECT 1821.210 3582.330 1822.390 3583.510 ;
        RECT 1921.210 3582.330 1922.390 3583.510 ;
        RECT 2021.210 3582.330 2022.390 3583.510 ;
        RECT 2121.210 3582.330 2122.390 3583.510 ;
        RECT 2221.210 3582.330 2222.390 3583.510 ;
        RECT 2321.210 3582.330 2322.390 3583.510 ;
        RECT 2421.210 3582.330 2422.390 3583.510 ;
        RECT 2521.210 3582.330 2522.390 3583.510 ;
        RECT 2621.210 3582.330 2622.390 3583.510 ;
        RECT 2721.210 3582.330 2722.390 3583.510 ;
        RECT 2821.210 3582.330 2822.390 3583.510 ;
        RECT 2921.210 3582.330 2922.390 3583.510 ;
        RECT 2992.990 3582.330 2994.170 3583.510 ;
        RECT 0.410 3521.210 1.590 3522.390 ;
        RECT 0.410 3421.210 1.590 3422.390 ;
        RECT 0.410 3321.210 1.590 3322.390 ;
        RECT 0.410 3221.210 1.590 3222.390 ;
        RECT 0.410 3121.210 1.590 3122.390 ;
        RECT 0.410 3021.210 1.590 3022.390 ;
        RECT 0.410 2921.210 1.590 2922.390 ;
        RECT 0.410 2821.210 1.590 2822.390 ;
        RECT 0.410 2721.210 1.590 2722.390 ;
        RECT 0.410 2621.210 1.590 2622.390 ;
        RECT 0.410 2521.210 1.590 2522.390 ;
        RECT 0.410 2421.210 1.590 2422.390 ;
        RECT 0.410 2321.210 1.590 2322.390 ;
        RECT 0.410 2221.210 1.590 2222.390 ;
        RECT 0.410 2121.210 1.590 2122.390 ;
        RECT 0.410 2021.210 1.590 2022.390 ;
        RECT 0.410 1921.210 1.590 1922.390 ;
        RECT 0.410 1821.210 1.590 1822.390 ;
        RECT 0.410 1721.210 1.590 1722.390 ;
        RECT 0.410 1621.210 1.590 1622.390 ;
        RECT 0.410 1521.210 1.590 1522.390 ;
        RECT 0.410 1421.210 1.590 1422.390 ;
        RECT 0.410 1321.210 1.590 1322.390 ;
        RECT 0.410 1221.210 1.590 1222.390 ;
        RECT 0.410 1121.210 1.590 1122.390 ;
        RECT 0.410 1021.210 1.590 1022.390 ;
        RECT 0.410 921.210 1.590 922.390 ;
        RECT 0.410 821.210 1.590 822.390 ;
        RECT 0.410 721.210 1.590 722.390 ;
        RECT 0.410 621.210 1.590 622.390 ;
        RECT 0.410 521.210 1.590 522.390 ;
        RECT 0.410 421.210 1.590 422.390 ;
        RECT 0.410 321.210 1.590 322.390 ;
        RECT 0.410 221.210 1.590 222.390 ;
        RECT 0.410 121.210 1.590 122.390 ;
        RECT 2992.990 3521.210 2994.170 3522.390 ;
        RECT 2992.990 3421.210 2994.170 3422.390 ;
        RECT 2992.990 3321.210 2994.170 3322.390 ;
        RECT 2992.990 3221.210 2994.170 3222.390 ;
        RECT 2992.990 3121.210 2994.170 3122.390 ;
        RECT 2992.990 3021.210 2994.170 3022.390 ;
        RECT 2992.990 2921.210 2994.170 2922.390 ;
        RECT 2992.990 2821.210 2994.170 2822.390 ;
        RECT 2992.990 2721.210 2994.170 2722.390 ;
        RECT 2992.990 2621.210 2994.170 2622.390 ;
        RECT 2992.990 2521.210 2994.170 2522.390 ;
        RECT 2992.990 2421.210 2994.170 2422.390 ;
        RECT 2992.990 2321.210 2994.170 2322.390 ;
        RECT 2992.990 2221.210 2994.170 2222.390 ;
        RECT 2992.990 2121.210 2994.170 2122.390 ;
        RECT 2992.990 2021.210 2994.170 2022.390 ;
        RECT 2992.990 1921.210 2994.170 1922.390 ;
        RECT 2992.990 1821.210 2994.170 1822.390 ;
        RECT 2992.990 1721.210 2994.170 1722.390 ;
        RECT 2992.990 1621.210 2994.170 1622.390 ;
        RECT 2992.990 1521.210 2994.170 1522.390 ;
        RECT 2992.990 1421.210 2994.170 1422.390 ;
        RECT 2992.990 1321.210 2994.170 1322.390 ;
        RECT 2992.990 1221.210 2994.170 1222.390 ;
        RECT 2992.990 1121.210 2994.170 1122.390 ;
        RECT 2992.990 1021.210 2994.170 1022.390 ;
        RECT 2992.990 921.210 2994.170 922.390 ;
        RECT 2992.990 821.210 2994.170 822.390 ;
        RECT 2992.990 721.210 2994.170 722.390 ;
        RECT 2992.990 621.210 2994.170 622.390 ;
        RECT 2992.990 521.210 2994.170 522.390 ;
        RECT 2992.990 421.210 2994.170 422.390 ;
        RECT 2992.990 321.210 2994.170 322.390 ;
        RECT 2992.990 221.210 2994.170 222.390 ;
        RECT 2992.990 121.210 2994.170 122.390 ;
        RECT 0.410 0.410 1.590 1.590 ;
        RECT 121.210 0.410 122.390 1.590 ;
        RECT 221.210 0.410 222.390 1.590 ;
        RECT 321.210 0.410 322.390 1.590 ;
        RECT 421.210 0.410 422.390 1.590 ;
        RECT 521.210 0.410 522.390 1.590 ;
        RECT 621.210 0.410 622.390 1.590 ;
        RECT 721.210 0.410 722.390 1.590 ;
        RECT 821.210 0.410 822.390 1.590 ;
        RECT 921.210 0.410 922.390 1.590 ;
        RECT 1021.210 0.410 1022.390 1.590 ;
        RECT 1121.210 0.410 1122.390 1.590 ;
        RECT 1221.210 0.410 1222.390 1.590 ;
        RECT 1321.210 0.410 1322.390 1.590 ;
        RECT 1421.210 0.410 1422.390 1.590 ;
        RECT 1521.210 0.410 1522.390 1.590 ;
        RECT 1621.210 0.410 1622.390 1.590 ;
        RECT 1721.210 0.410 1722.390 1.590 ;
        RECT 1821.210 0.410 1822.390 1.590 ;
        RECT 1921.210 0.410 1922.390 1.590 ;
        RECT 2021.210 0.410 2022.390 1.590 ;
        RECT 2121.210 0.410 2122.390 1.590 ;
        RECT 2221.210 0.410 2222.390 1.590 ;
        RECT 2321.210 0.410 2322.390 1.590 ;
        RECT 2421.210 0.410 2422.390 1.590 ;
        RECT 2521.210 0.410 2522.390 1.590 ;
        RECT 2621.210 0.410 2622.390 1.590 ;
        RECT 2721.210 0.410 2722.390 1.590 ;
        RECT 2821.210 0.410 2822.390 1.590 ;
        RECT 2921.210 0.410 2922.390 1.590 ;
        RECT 2992.990 0.410 2994.170 1.590 ;
      LAYER met5 ;
        RECT 0.000 3581.920 2994.580 3583.920 ;
        RECT 0.000 3520.800 39.880 3522.800 ;
        RECT 2955.080 3520.800 2994.580 3522.800 ;
        RECT 0.000 3420.800 39.880 3422.800 ;
        RECT 2955.080 3420.800 2994.580 3422.800 ;
        RECT 0.000 3320.800 39.880 3322.800 ;
        RECT 2955.080 3320.800 2994.580 3322.800 ;
        RECT 0.000 3220.800 39.880 3222.800 ;
        RECT 2955.080 3220.800 2994.580 3222.800 ;
        RECT 0.000 3120.800 39.880 3122.800 ;
        RECT 2955.080 3120.800 2994.580 3122.800 ;
        RECT 0.000 3020.800 39.880 3022.800 ;
        RECT 2955.080 3020.800 2994.580 3022.800 ;
        RECT 0.000 2920.800 39.880 2922.800 ;
        RECT 2955.080 2920.800 2994.580 2922.800 ;
        RECT 0.000 2820.800 39.880 2822.800 ;
        RECT 2955.080 2820.800 2994.580 2822.800 ;
        RECT 0.000 2720.800 39.880 2722.800 ;
        RECT 2955.080 2720.800 2994.580 2722.800 ;
        RECT 0.000 2620.800 39.880 2622.800 ;
        RECT 2955.080 2620.800 2994.580 2622.800 ;
        RECT 0.000 2520.800 39.880 2522.800 ;
        RECT 2955.080 2520.800 2994.580 2522.800 ;
        RECT 0.000 2420.800 39.880 2422.800 ;
        RECT 2955.080 2420.800 2994.580 2422.800 ;
        RECT 0.000 2320.800 39.880 2322.800 ;
        RECT 2955.080 2320.800 2994.580 2322.800 ;
        RECT 0.000 2220.800 39.880 2222.800 ;
        RECT 2955.080 2220.800 2994.580 2222.800 ;
        RECT 0.000 2120.800 39.880 2122.800 ;
        RECT 2955.080 2120.800 2994.580 2122.800 ;
        RECT 0.000 2020.800 39.880 2022.800 ;
        RECT 2955.080 2020.800 2994.580 2022.800 ;
        RECT 0.000 1920.800 39.880 1922.800 ;
        RECT 2955.080 1920.800 2994.580 1922.800 ;
        RECT 0.000 1820.800 39.880 1822.800 ;
        RECT 2955.080 1820.800 2994.580 1822.800 ;
        RECT 0.000 1720.800 39.880 1722.800 ;
        RECT 2955.080 1720.800 2994.580 1722.800 ;
        RECT 0.000 1620.800 39.880 1622.800 ;
        RECT 2955.080 1620.800 2994.580 1622.800 ;
        RECT 0.000 1520.800 39.880 1522.800 ;
        RECT 2955.080 1520.800 2994.580 1522.800 ;
        RECT 0.000 1420.800 39.880 1422.800 ;
        RECT 2955.080 1420.800 2994.580 1422.800 ;
        RECT 0.000 1320.800 39.880 1322.800 ;
        RECT 2955.080 1320.800 2994.580 1322.800 ;
        RECT 0.000 1220.800 39.880 1222.800 ;
        RECT 2955.080 1220.800 2994.580 1222.800 ;
        RECT 0.000 1120.800 39.880 1122.800 ;
        RECT 2955.080 1120.800 2994.580 1122.800 ;
        RECT 0.000 1020.800 39.880 1022.800 ;
        RECT 2955.080 1020.800 2994.580 1022.800 ;
        RECT 0.000 920.800 39.880 922.800 ;
        RECT 2955.080 920.800 2994.580 922.800 ;
        RECT 0.000 820.800 39.880 822.800 ;
        RECT 2955.080 820.800 2994.580 822.800 ;
        RECT 0.000 720.800 39.880 722.800 ;
        RECT 2955.080 720.800 2994.580 722.800 ;
        RECT 0.000 620.800 39.880 622.800 ;
        RECT 2955.080 620.800 2994.580 622.800 ;
        RECT 0.000 520.800 39.880 522.800 ;
        RECT 2955.080 520.800 2994.580 522.800 ;
        RECT 0.000 420.800 39.880 422.800 ;
        RECT 2955.080 420.800 2994.580 422.800 ;
        RECT 0.000 320.800 39.880 322.800 ;
        RECT 2955.080 320.800 2994.580 322.800 ;
        RECT 0.000 220.800 39.880 222.800 ;
        RECT 2955.080 220.800 2994.580 222.800 ;
        RECT 0.000 120.800 39.880 122.800 ;
        RECT 2955.080 120.800 2994.580 122.800 ;
        RECT 0.000 0.000 2994.580 2.000 ;
    END
  END vssa2
  OBS
      LAYER nwell ;
        RECT 42.280 618.225 631.460 619.830 ;
      LAYER pwell ;
        RECT 42.615 616.835 42.785 617.005 ;
        RECT 43.995 616.835 44.165 617.005 ;
        RECT 49.515 616.835 49.685 617.005 ;
      LAYER nwell ;
        RECT 42.280 612.785 631.460 615.615 ;
      LAYER pwell ;
        RECT 42.615 611.395 42.785 611.565 ;
        RECT 43.995 611.395 44.165 611.565 ;
        RECT 49.515 611.395 49.685 611.565 ;
      LAYER nwell ;
        RECT 42.280 607.345 631.460 610.175 ;
      LAYER pwell ;
        RECT 42.615 605.955 42.785 606.125 ;
        RECT 43.995 605.955 44.165 606.125 ;
        RECT 49.515 605.955 49.685 606.125 ;
      LAYER nwell ;
        RECT 42.280 601.905 631.460 604.735 ;
      LAYER pwell ;
        RECT 42.615 600.515 42.785 600.685 ;
        RECT 43.995 600.515 44.165 600.685 ;
        RECT 49.515 600.515 49.685 600.685 ;
      LAYER nwell ;
        RECT 42.280 596.465 631.460 599.295 ;
      LAYER pwell ;
        RECT 42.615 595.075 42.785 595.245 ;
        RECT 43.995 595.075 44.165 595.245 ;
        RECT 49.515 595.075 49.685 595.245 ;
      LAYER nwell ;
        RECT 42.280 591.025 631.460 593.855 ;
      LAYER pwell ;
        RECT 42.615 589.635 42.785 589.805 ;
        RECT 43.995 589.635 44.165 589.805 ;
        RECT 49.515 589.635 49.685 589.805 ;
      LAYER nwell ;
        RECT 42.280 585.585 631.460 588.415 ;
      LAYER pwell ;
        RECT 42.615 584.195 42.785 584.365 ;
        RECT 43.995 584.195 44.165 584.365 ;
        RECT 49.515 584.195 49.685 584.365 ;
      LAYER nwell ;
        RECT 42.280 580.145 631.460 582.975 ;
      LAYER pwell ;
        RECT 42.615 578.755 42.785 578.925 ;
        RECT 43.995 578.755 44.165 578.925 ;
        RECT 49.515 578.755 49.685 578.925 ;
      LAYER nwell ;
        RECT 42.280 574.705 631.460 577.535 ;
      LAYER pwell ;
        RECT 42.615 573.315 42.785 573.485 ;
        RECT 43.995 573.315 44.165 573.485 ;
        RECT 49.515 573.315 49.685 573.485 ;
      LAYER nwell ;
        RECT 42.280 569.265 631.460 572.095 ;
      LAYER pwell ;
        RECT 42.615 567.875 42.785 568.045 ;
        RECT 43.995 567.875 44.165 568.045 ;
        RECT 49.515 567.875 49.685 568.045 ;
      LAYER nwell ;
        RECT 42.280 563.825 631.460 566.655 ;
      LAYER pwell ;
        RECT 42.615 562.435 42.785 562.605 ;
        RECT 43.995 562.435 44.165 562.605 ;
        RECT 49.515 562.435 49.685 562.605 ;
      LAYER nwell ;
        RECT 42.280 558.385 631.460 561.215 ;
      LAYER pwell ;
        RECT 42.615 556.995 42.785 557.165 ;
        RECT 43.995 556.995 44.165 557.165 ;
        RECT 49.515 556.995 49.685 557.165 ;
      LAYER nwell ;
        RECT 42.280 552.945 631.460 555.775 ;
      LAYER pwell ;
        RECT 42.615 551.555 42.785 551.725 ;
        RECT 43.995 551.555 44.165 551.725 ;
        RECT 49.515 551.555 49.685 551.725 ;
      LAYER nwell ;
        RECT 42.280 547.505 631.460 550.335 ;
      LAYER pwell ;
        RECT 42.615 546.115 42.785 546.285 ;
        RECT 43.995 546.115 44.165 546.285 ;
        RECT 49.515 546.115 49.685 546.285 ;
      LAYER nwell ;
        RECT 42.280 542.065 631.460 544.895 ;
      LAYER pwell ;
        RECT 42.615 540.675 42.785 540.845 ;
        RECT 43.995 540.675 44.165 540.845 ;
        RECT 49.515 540.675 49.685 540.845 ;
      LAYER nwell ;
        RECT 42.280 536.625 631.460 539.455 ;
      LAYER pwell ;
        RECT 42.615 535.235 42.785 535.405 ;
        RECT 43.995 535.235 44.165 535.405 ;
        RECT 49.515 535.235 49.685 535.405 ;
      LAYER nwell ;
        RECT 42.280 531.185 631.460 534.015 ;
      LAYER pwell ;
        RECT 42.615 529.795 42.785 529.965 ;
        RECT 43.995 529.795 44.165 529.965 ;
        RECT 49.515 529.795 49.685 529.965 ;
      LAYER nwell ;
        RECT 42.280 525.745 631.460 528.575 ;
      LAYER pwell ;
        RECT 42.615 524.355 42.785 524.525 ;
        RECT 43.995 524.355 44.165 524.525 ;
        RECT 49.515 524.355 49.685 524.525 ;
      LAYER nwell ;
        RECT 42.280 520.305 631.460 523.135 ;
      LAYER pwell ;
        RECT 42.615 518.915 42.785 519.085 ;
        RECT 43.995 518.915 44.165 519.085 ;
        RECT 49.515 518.915 49.685 519.085 ;
      LAYER nwell ;
        RECT 42.280 514.865 631.460 517.695 ;
      LAYER pwell ;
        RECT 42.615 513.475 42.785 513.645 ;
        RECT 43.995 513.475 44.165 513.645 ;
        RECT 49.515 513.475 49.685 513.645 ;
      LAYER nwell ;
        RECT 42.280 509.425 631.460 512.255 ;
      LAYER pwell ;
        RECT 42.615 508.035 42.785 508.205 ;
        RECT 43.995 508.035 44.165 508.205 ;
        RECT 49.515 508.035 49.685 508.205 ;
      LAYER nwell ;
        RECT 42.280 503.985 631.460 506.815 ;
      LAYER pwell ;
        RECT 42.615 502.595 42.785 502.765 ;
        RECT 43.995 502.595 44.165 502.765 ;
        RECT 49.515 502.595 49.685 502.765 ;
      LAYER nwell ;
        RECT 42.280 498.545 631.460 501.375 ;
      LAYER pwell ;
        RECT 42.615 497.155 42.785 497.325 ;
        RECT 43.995 497.155 44.165 497.325 ;
        RECT 49.515 497.155 49.685 497.325 ;
      LAYER nwell ;
        RECT 42.280 493.105 631.460 495.935 ;
      LAYER pwell ;
        RECT 42.615 491.715 42.785 491.885 ;
        RECT 43.995 491.715 44.165 491.885 ;
        RECT 49.515 491.715 49.685 491.885 ;
      LAYER nwell ;
        RECT 42.280 487.665 631.460 490.495 ;
      LAYER pwell ;
        RECT 42.615 486.275 42.785 486.445 ;
        RECT 43.995 486.275 44.165 486.445 ;
        RECT 49.515 486.275 49.685 486.445 ;
      LAYER nwell ;
        RECT 42.280 482.225 631.460 485.055 ;
      LAYER pwell ;
        RECT 42.615 480.835 42.785 481.005 ;
        RECT 43.995 480.835 44.165 481.005 ;
        RECT 49.515 480.835 49.685 481.005 ;
      LAYER nwell ;
        RECT 42.280 476.785 631.460 479.615 ;
      LAYER pwell ;
        RECT 42.615 475.395 42.785 475.565 ;
        RECT 43.995 475.395 44.165 475.565 ;
        RECT 49.515 475.395 49.685 475.565 ;
      LAYER nwell ;
        RECT 42.280 471.345 631.460 474.175 ;
      LAYER pwell ;
        RECT 42.615 469.955 42.785 470.125 ;
        RECT 43.995 469.955 44.165 470.125 ;
        RECT 49.515 469.955 49.685 470.125 ;
      LAYER nwell ;
        RECT 42.280 465.905 631.460 468.735 ;
      LAYER pwell ;
        RECT 42.615 464.515 42.785 464.685 ;
        RECT 43.995 464.515 44.165 464.685 ;
        RECT 49.515 464.515 49.685 464.685 ;
      LAYER nwell ;
        RECT 42.280 460.465 631.460 463.295 ;
      LAYER pwell ;
        RECT 42.615 459.075 42.785 459.245 ;
        RECT 43.995 459.075 44.165 459.245 ;
        RECT 49.515 459.075 49.685 459.245 ;
      LAYER nwell ;
        RECT 42.280 455.025 631.460 457.855 ;
      LAYER pwell ;
        RECT 42.615 453.635 42.785 453.805 ;
        RECT 43.995 453.635 44.165 453.805 ;
        RECT 49.515 453.635 49.685 453.805 ;
      LAYER nwell ;
        RECT 42.280 449.585 631.460 452.415 ;
      LAYER pwell ;
        RECT 42.615 448.195 42.785 448.365 ;
        RECT 43.995 448.195 44.165 448.365 ;
        RECT 49.515 448.195 49.685 448.365 ;
      LAYER nwell ;
        RECT 42.280 444.145 631.460 446.975 ;
      LAYER pwell ;
        RECT 42.615 442.755 42.785 442.925 ;
        RECT 43.995 442.755 44.165 442.925 ;
        RECT 49.515 442.755 49.685 442.925 ;
      LAYER nwell ;
        RECT 42.280 438.705 631.460 441.535 ;
      LAYER pwell ;
        RECT 42.615 437.315 42.785 437.485 ;
        RECT 43.995 437.315 44.165 437.485 ;
        RECT 49.515 437.315 49.685 437.485 ;
      LAYER nwell ;
        RECT 42.280 433.265 631.460 436.095 ;
      LAYER pwell ;
        RECT 42.615 431.875 42.785 432.045 ;
        RECT 43.995 431.875 44.165 432.045 ;
        RECT 49.515 431.875 49.685 432.045 ;
      LAYER nwell ;
        RECT 42.280 427.825 631.460 430.655 ;
      LAYER pwell ;
        RECT 42.615 426.435 42.785 426.605 ;
        RECT 43.995 426.435 44.165 426.605 ;
        RECT 49.515 426.435 49.685 426.605 ;
      LAYER nwell ;
        RECT 42.280 422.385 631.460 425.215 ;
      LAYER pwell ;
        RECT 42.615 420.995 42.785 421.165 ;
        RECT 43.995 420.995 44.165 421.165 ;
        RECT 49.515 420.995 49.685 421.165 ;
      LAYER nwell ;
        RECT 42.280 416.945 631.460 419.775 ;
      LAYER pwell ;
        RECT 42.615 415.555 42.785 415.725 ;
        RECT 43.995 415.555 44.165 415.725 ;
        RECT 49.515 415.555 49.685 415.725 ;
      LAYER nwell ;
        RECT 42.280 411.505 631.460 414.335 ;
      LAYER pwell ;
        RECT 42.615 410.115 42.785 410.285 ;
        RECT 43.995 410.115 44.165 410.285 ;
        RECT 49.515 410.115 49.685 410.285 ;
      LAYER nwell ;
        RECT 42.280 406.065 631.460 408.895 ;
      LAYER pwell ;
        RECT 42.615 404.675 42.785 404.845 ;
        RECT 43.995 404.675 44.165 404.845 ;
        RECT 49.515 404.675 49.685 404.845 ;
      LAYER nwell ;
        RECT 42.280 400.625 631.460 403.455 ;
      LAYER pwell ;
        RECT 42.615 399.235 42.785 399.405 ;
        RECT 43.995 399.235 44.165 399.405 ;
        RECT 49.515 399.235 49.685 399.405 ;
      LAYER nwell ;
        RECT 42.280 395.185 631.460 398.015 ;
      LAYER pwell ;
        RECT 42.615 393.795 42.785 393.965 ;
        RECT 43.995 393.795 44.165 393.965 ;
        RECT 49.515 393.795 49.685 393.965 ;
      LAYER nwell ;
        RECT 42.280 389.745 631.460 392.575 ;
      LAYER pwell ;
        RECT 42.615 388.355 42.785 388.525 ;
        RECT 43.995 388.355 44.165 388.525 ;
        RECT 49.515 388.355 49.685 388.525 ;
      LAYER nwell ;
        RECT 42.280 384.305 631.460 387.135 ;
      LAYER pwell ;
        RECT 42.615 382.915 42.785 383.085 ;
        RECT 43.995 382.915 44.165 383.085 ;
        RECT 49.515 382.915 49.685 383.085 ;
      LAYER nwell ;
        RECT 42.280 378.865 631.460 381.695 ;
      LAYER pwell ;
        RECT 42.615 377.475 42.785 377.645 ;
        RECT 43.995 377.475 44.165 377.645 ;
        RECT 49.515 377.475 49.685 377.645 ;
      LAYER nwell ;
        RECT 42.280 373.425 631.460 376.255 ;
      LAYER pwell ;
        RECT 42.615 372.035 42.785 372.205 ;
        RECT 43.995 372.035 44.165 372.205 ;
        RECT 49.515 372.035 49.685 372.205 ;
      LAYER nwell ;
        RECT 42.280 367.985 631.460 370.815 ;
      LAYER pwell ;
        RECT 42.615 366.595 42.785 366.765 ;
        RECT 43.995 366.595 44.165 366.765 ;
        RECT 49.515 366.595 49.685 366.765 ;
      LAYER nwell ;
        RECT 42.280 362.545 631.460 365.375 ;
      LAYER pwell ;
        RECT 42.615 361.155 42.785 361.325 ;
        RECT 43.995 361.155 44.165 361.325 ;
        RECT 49.515 361.155 49.685 361.325 ;
      LAYER nwell ;
        RECT 42.280 357.105 631.460 359.935 ;
      LAYER pwell ;
        RECT 42.615 355.715 42.785 355.885 ;
        RECT 43.995 355.715 44.165 355.885 ;
        RECT 49.515 355.715 49.685 355.885 ;
      LAYER nwell ;
        RECT 42.280 351.665 631.460 354.495 ;
      LAYER pwell ;
        RECT 42.615 350.275 42.785 350.445 ;
        RECT 43.995 350.275 44.165 350.445 ;
        RECT 49.515 350.275 49.685 350.445 ;
      LAYER nwell ;
        RECT 42.280 346.225 631.460 349.055 ;
      LAYER pwell ;
        RECT 42.615 344.835 42.785 345.005 ;
        RECT 43.995 344.835 44.165 345.005 ;
        RECT 49.515 344.835 49.685 345.005 ;
      LAYER nwell ;
        RECT 42.280 340.785 631.460 343.615 ;
      LAYER pwell ;
        RECT 42.615 339.395 42.785 339.565 ;
        RECT 43.995 339.395 44.165 339.565 ;
        RECT 49.515 339.395 49.685 339.565 ;
      LAYER nwell ;
        RECT 42.280 335.345 631.460 338.175 ;
      LAYER pwell ;
        RECT 42.615 333.955 42.785 334.125 ;
        RECT 43.995 333.955 44.165 334.125 ;
        RECT 49.515 333.955 49.685 334.125 ;
      LAYER nwell ;
        RECT 42.280 329.905 631.460 332.735 ;
      LAYER pwell ;
        RECT 42.615 328.515 42.785 328.685 ;
        RECT 43.995 328.515 44.165 328.685 ;
        RECT 49.515 328.515 49.685 328.685 ;
      LAYER nwell ;
        RECT 42.280 324.465 631.460 327.295 ;
      LAYER pwell ;
        RECT 42.615 323.075 42.785 323.245 ;
        RECT 43.995 323.075 44.165 323.245 ;
        RECT 49.515 323.075 49.685 323.245 ;
      LAYER nwell ;
        RECT 42.280 319.025 631.460 321.855 ;
      LAYER pwell ;
        RECT 42.615 317.635 42.785 317.805 ;
        RECT 43.995 317.635 44.165 317.805 ;
        RECT 49.515 317.635 49.685 317.805 ;
      LAYER nwell ;
        RECT 42.280 313.585 631.460 316.415 ;
      LAYER pwell ;
        RECT 42.615 312.195 42.785 312.365 ;
        RECT 43.995 312.195 44.165 312.365 ;
        RECT 49.515 312.195 49.685 312.365 ;
      LAYER nwell ;
        RECT 42.280 308.145 631.460 310.975 ;
      LAYER pwell ;
        RECT 42.615 306.755 42.785 306.925 ;
        RECT 43.995 306.755 44.165 306.925 ;
        RECT 49.515 306.755 49.685 306.925 ;
      LAYER nwell ;
        RECT 42.280 302.705 631.460 305.535 ;
      LAYER pwell ;
        RECT 42.615 301.315 42.785 301.485 ;
        RECT 43.995 301.315 44.165 301.485 ;
        RECT 49.515 301.315 49.685 301.485 ;
      LAYER nwell ;
        RECT 42.280 297.265 631.460 300.095 ;
      LAYER pwell ;
        RECT 42.615 295.875 42.785 296.045 ;
        RECT 43.995 295.875 44.165 296.045 ;
        RECT 49.515 295.875 49.685 296.045 ;
      LAYER nwell ;
        RECT 42.280 291.825 631.460 294.655 ;
      LAYER pwell ;
        RECT 42.615 290.435 42.785 290.605 ;
        RECT 43.995 290.435 44.165 290.605 ;
        RECT 49.515 290.435 49.685 290.605 ;
      LAYER nwell ;
        RECT 42.280 286.385 631.460 289.215 ;
      LAYER pwell ;
        RECT 42.615 284.995 42.785 285.165 ;
        RECT 43.995 284.995 44.165 285.165 ;
        RECT 49.515 284.995 49.685 285.165 ;
      LAYER nwell ;
        RECT 42.280 280.945 631.460 283.775 ;
      LAYER pwell ;
        RECT 42.615 279.555 42.785 279.725 ;
        RECT 43.995 279.555 44.165 279.725 ;
        RECT 49.515 279.555 49.685 279.725 ;
      LAYER nwell ;
        RECT 42.280 275.505 631.460 278.335 ;
      LAYER pwell ;
        RECT 42.615 274.115 42.785 274.285 ;
        RECT 43.995 274.115 44.165 274.285 ;
        RECT 49.515 274.115 49.685 274.285 ;
      LAYER nwell ;
        RECT 42.280 270.065 631.460 272.895 ;
      LAYER pwell ;
        RECT 42.615 268.675 42.785 268.845 ;
        RECT 43.995 268.675 44.165 268.845 ;
        RECT 49.515 268.675 49.685 268.845 ;
      LAYER nwell ;
        RECT 42.280 264.625 631.460 267.455 ;
      LAYER pwell ;
        RECT 42.615 263.235 42.785 263.405 ;
        RECT 43.995 263.235 44.165 263.405 ;
        RECT 49.515 263.235 49.685 263.405 ;
      LAYER nwell ;
        RECT 42.280 259.185 631.460 262.015 ;
      LAYER pwell ;
        RECT 42.615 257.795 42.785 257.965 ;
        RECT 43.995 257.795 44.165 257.965 ;
        RECT 49.515 257.795 49.685 257.965 ;
      LAYER nwell ;
        RECT 42.280 253.745 631.460 256.575 ;
      LAYER pwell ;
        RECT 42.615 252.355 42.785 252.525 ;
        RECT 43.995 252.355 44.165 252.525 ;
        RECT 49.515 252.355 49.685 252.525 ;
      LAYER nwell ;
        RECT 42.280 248.305 631.460 251.135 ;
      LAYER pwell ;
        RECT 42.615 246.915 42.785 247.085 ;
        RECT 43.995 246.915 44.165 247.085 ;
        RECT 49.515 246.915 49.685 247.085 ;
      LAYER nwell ;
        RECT 42.280 242.865 631.460 245.695 ;
      LAYER pwell ;
        RECT 42.615 241.475 42.785 241.645 ;
        RECT 43.995 241.475 44.165 241.645 ;
        RECT 49.515 241.475 49.685 241.645 ;
      LAYER nwell ;
        RECT 42.280 237.425 631.460 240.255 ;
      LAYER pwell ;
        RECT 42.615 236.035 42.785 236.205 ;
        RECT 43.995 236.035 44.165 236.205 ;
        RECT 49.515 236.035 49.685 236.205 ;
      LAYER nwell ;
        RECT 42.280 231.985 631.460 234.815 ;
      LAYER pwell ;
        RECT 42.615 230.595 42.785 230.765 ;
        RECT 43.995 230.595 44.165 230.765 ;
        RECT 49.515 230.595 49.685 230.765 ;
      LAYER nwell ;
        RECT 42.280 226.545 631.460 229.375 ;
      LAYER pwell ;
        RECT 42.615 225.155 42.785 225.325 ;
        RECT 43.995 225.155 44.165 225.325 ;
        RECT 49.515 225.155 49.685 225.325 ;
      LAYER nwell ;
        RECT 42.280 221.105 631.460 223.935 ;
      LAYER pwell ;
        RECT 42.615 219.715 42.785 219.885 ;
        RECT 43.995 219.715 44.165 219.885 ;
        RECT 49.515 219.715 49.685 219.885 ;
      LAYER nwell ;
        RECT 42.280 215.665 631.460 218.495 ;
      LAYER pwell ;
        RECT 42.615 214.275 42.785 214.445 ;
        RECT 43.995 214.275 44.165 214.445 ;
        RECT 49.515 214.275 49.685 214.445 ;
      LAYER nwell ;
        RECT 42.280 210.225 631.460 213.055 ;
      LAYER pwell ;
        RECT 42.615 208.835 42.785 209.005 ;
        RECT 43.995 208.835 44.165 209.005 ;
        RECT 49.515 208.835 49.685 209.005 ;
      LAYER nwell ;
        RECT 42.280 204.785 631.460 207.615 ;
      LAYER pwell ;
        RECT 42.615 203.395 42.785 203.565 ;
        RECT 43.995 203.395 44.165 203.565 ;
        RECT 49.515 203.395 49.685 203.565 ;
      LAYER nwell ;
        RECT 42.280 199.345 631.460 202.175 ;
      LAYER pwell ;
        RECT 42.615 197.955 42.785 198.125 ;
        RECT 43.995 197.955 44.165 198.125 ;
        RECT 49.515 197.955 49.685 198.125 ;
      LAYER nwell ;
        RECT 42.280 193.905 631.460 196.735 ;
      LAYER pwell ;
        RECT 42.615 192.515 42.785 192.685 ;
        RECT 43.995 192.515 44.165 192.685 ;
        RECT 49.515 192.515 49.685 192.685 ;
      LAYER nwell ;
        RECT 42.280 188.465 631.460 191.295 ;
      LAYER pwell ;
        RECT 42.615 187.075 42.785 187.245 ;
        RECT 43.995 187.075 44.165 187.245 ;
        RECT 49.515 187.075 49.685 187.245 ;
      LAYER nwell ;
        RECT 42.280 183.025 631.460 185.855 ;
      LAYER pwell ;
        RECT 42.615 181.635 42.785 181.805 ;
        RECT 43.995 181.635 44.165 181.805 ;
        RECT 49.515 181.635 49.685 181.805 ;
      LAYER nwell ;
        RECT 42.280 177.585 631.460 180.415 ;
      LAYER pwell ;
        RECT 42.615 176.195 42.785 176.365 ;
        RECT 43.995 176.195 44.165 176.365 ;
        RECT 49.515 176.195 49.685 176.365 ;
      LAYER nwell ;
        RECT 42.280 172.145 631.460 174.975 ;
      LAYER pwell ;
        RECT 42.615 170.755 42.785 170.925 ;
        RECT 43.995 170.755 44.165 170.925 ;
        RECT 49.515 170.755 49.685 170.925 ;
      LAYER nwell ;
        RECT 42.280 166.705 631.460 169.535 ;
      LAYER pwell ;
        RECT 42.615 165.315 42.785 165.485 ;
        RECT 43.995 165.315 44.165 165.485 ;
        RECT 49.515 165.315 49.685 165.485 ;
      LAYER nwell ;
        RECT 42.280 161.265 631.460 164.095 ;
      LAYER pwell ;
        RECT 42.615 159.875 42.785 160.045 ;
        RECT 43.995 159.875 44.165 160.045 ;
        RECT 49.515 159.875 49.685 160.045 ;
      LAYER nwell ;
        RECT 42.280 155.825 631.460 158.655 ;
      LAYER pwell ;
        RECT 42.615 154.435 42.785 154.605 ;
        RECT 43.995 154.435 44.165 154.605 ;
        RECT 49.515 154.435 49.685 154.605 ;
      LAYER nwell ;
        RECT 42.280 150.385 631.460 153.215 ;
      LAYER pwell ;
        RECT 42.615 148.995 42.785 149.165 ;
        RECT 43.995 148.995 44.165 149.165 ;
        RECT 49.515 148.995 49.685 149.165 ;
      LAYER nwell ;
        RECT 42.280 144.945 631.460 147.775 ;
      LAYER pwell ;
        RECT 42.615 143.555 42.785 143.725 ;
        RECT 43.995 143.555 44.165 143.725 ;
        RECT 49.515 143.555 49.685 143.725 ;
      LAYER nwell ;
        RECT 42.280 139.505 631.460 142.335 ;
      LAYER pwell ;
        RECT 42.615 138.115 42.785 138.285 ;
        RECT 43.995 138.115 44.165 138.285 ;
        RECT 49.515 138.115 49.685 138.285 ;
      LAYER nwell ;
        RECT 42.280 134.065 631.460 136.895 ;
      LAYER pwell ;
        RECT 42.615 132.675 42.785 132.845 ;
        RECT 43.995 132.675 44.165 132.845 ;
        RECT 49.515 132.675 49.685 132.845 ;
      LAYER nwell ;
        RECT 42.280 128.625 631.460 131.455 ;
      LAYER pwell ;
        RECT 42.615 127.235 42.785 127.405 ;
        RECT 43.995 127.235 44.165 127.405 ;
        RECT 49.515 127.235 49.685 127.405 ;
      LAYER nwell ;
        RECT 42.280 123.185 631.460 126.015 ;
      LAYER pwell ;
        RECT 42.615 121.795 42.785 121.965 ;
        RECT 43.995 121.795 44.165 121.965 ;
        RECT 49.515 121.795 49.685 121.965 ;
      LAYER nwell ;
        RECT 42.280 117.745 631.460 120.575 ;
      LAYER pwell ;
        RECT 42.615 116.355 42.785 116.525 ;
        RECT 43.995 116.355 44.165 116.525 ;
        RECT 49.515 116.355 49.685 116.525 ;
      LAYER nwell ;
        RECT 42.280 112.305 631.460 115.135 ;
      LAYER pwell ;
        RECT 42.615 110.915 42.785 111.085 ;
        RECT 43.995 110.915 44.165 111.085 ;
        RECT 49.515 110.915 49.685 111.085 ;
      LAYER nwell ;
        RECT 42.280 106.865 631.460 109.695 ;
      LAYER pwell ;
        RECT 42.615 105.475 42.785 105.645 ;
        RECT 43.995 105.475 44.165 105.645 ;
        RECT 49.515 105.475 49.685 105.645 ;
      LAYER nwell ;
        RECT 42.280 101.425 631.460 104.255 ;
      LAYER pwell ;
        RECT 42.615 100.035 42.785 100.205 ;
        RECT 43.995 100.035 44.165 100.205 ;
        RECT 49.515 100.035 49.685 100.205 ;
      LAYER nwell ;
        RECT 42.280 95.985 631.460 98.815 ;
      LAYER pwell ;
        RECT 42.615 94.595 42.785 94.765 ;
        RECT 43.995 94.595 44.165 94.765 ;
        RECT 49.515 94.595 49.685 94.765 ;
      LAYER nwell ;
        RECT 42.280 90.545 631.460 93.375 ;
      LAYER pwell ;
        RECT 42.615 89.155 42.785 89.325 ;
        RECT 43.995 89.155 44.165 89.325 ;
        RECT 49.515 89.155 49.685 89.325 ;
      LAYER nwell ;
        RECT 42.280 85.105 631.460 87.935 ;
      LAYER pwell ;
        RECT 42.615 83.715 42.785 83.885 ;
        RECT 43.995 83.715 44.165 83.885 ;
        RECT 49.515 83.715 49.685 83.885 ;
      LAYER nwell ;
        RECT 42.280 79.665 631.460 82.495 ;
      LAYER pwell ;
        RECT 42.615 78.275 42.785 78.445 ;
        RECT 43.995 78.275 44.165 78.445 ;
        RECT 49.515 78.275 49.685 78.445 ;
      LAYER nwell ;
        RECT 42.280 74.225 631.460 77.055 ;
      LAYER pwell ;
        RECT 42.615 72.835 42.785 73.005 ;
        RECT 43.995 72.835 44.165 73.005 ;
        RECT 49.515 72.835 49.685 73.005 ;
      LAYER nwell ;
        RECT 42.280 68.785 631.460 71.615 ;
      LAYER pwell ;
        RECT 42.615 67.395 42.785 67.565 ;
        RECT 43.995 67.395 44.165 67.565 ;
        RECT 49.515 67.395 49.685 67.565 ;
      LAYER nwell ;
        RECT 42.280 63.345 631.460 66.175 ;
      LAYER pwell ;
        RECT 42.615 61.955 42.785 62.125 ;
        RECT 43.995 61.955 44.165 62.125 ;
        RECT 49.515 61.955 49.685 62.125 ;
      LAYER nwell ;
        RECT 42.280 57.905 631.460 60.735 ;
      LAYER pwell ;
        RECT 42.615 56.515 42.785 56.685 ;
        RECT 43.995 56.515 44.165 56.685 ;
        RECT 49.515 56.515 49.685 56.685 ;
      LAYER nwell ;
        RECT 42.280 52.465 631.460 55.295 ;
      LAYER pwell ;
        RECT 70.675 51.480 70.845 52.005 ;
        RECT 98.735 51.480 98.905 52.005 ;
        RECT 126.795 51.480 126.965 52.005 ;
        RECT 154.855 51.480 155.025 52.005 ;
        RECT 182.915 51.480 183.085 52.005 ;
        RECT 210.975 51.480 211.145 52.005 ;
        RECT 239.035 51.480 239.205 52.005 ;
        RECT 267.095 51.480 267.265 52.005 ;
        RECT 295.155 51.480 295.325 52.005 ;
        RECT 323.215 51.480 323.385 52.005 ;
        RECT 351.275 51.480 351.445 52.005 ;
        RECT 379.335 51.480 379.505 52.005 ;
        RECT 407.395 51.480 407.565 52.005 ;
        RECT 435.455 51.480 435.625 52.005 ;
        RECT 463.515 51.480 463.685 52.005 ;
        RECT 491.575 51.480 491.745 52.005 ;
        RECT 519.635 51.480 519.805 52.005 ;
        RECT 547.695 51.480 547.865 52.005 ;
        RECT 575.755 51.480 575.925 52.005 ;
        RECT 603.815 51.480 603.985 52.005 ;
        RECT 42.615 51.075 42.785 51.245 ;
        RECT 43.995 51.075 44.165 51.245 ;
        RECT 49.515 51.075 49.685 51.245 ;
        RECT 55.035 51.075 55.205 51.245 ;
        RECT 57.335 51.075 57.505 51.245 ;
        RECT 60.555 51.075 60.725 51.245 ;
        RECT 62.855 51.075 63.025 51.245 ;
        RECT 66.075 51.075 66.245 51.245 ;
        RECT 68.375 51.075 68.545 51.245 ;
        RECT 69.765 51.110 69.925 51.220 ;
        RECT 71.135 51.075 71.305 51.245 ;
        RECT 72.065 51.100 72.225 51.210 ;
        RECT 72.975 51.075 73.145 51.245 ;
        RECT 74.355 51.075 74.525 51.245 ;
        RECT 76.665 51.110 76.825 51.220 ;
        RECT 77.575 51.075 77.745 51.245 ;
        RECT 78.040 51.075 78.210 51.245 ;
        RECT 78.955 51.075 79.125 51.245 ;
        RECT 81.255 51.075 81.425 51.245 ;
        RECT 82.635 51.075 82.805 51.245 ;
        RECT 85.390 51.105 85.510 51.215 ;
        RECT 85.855 51.075 86.025 51.245 ;
        RECT 87.695 51.075 87.865 51.245 ;
        RECT 91.375 51.075 91.545 51.245 ;
        RECT 96.895 51.075 97.065 51.245 ;
        RECT 99.195 51.075 99.365 51.245 ;
        RECT 100.115 51.075 100.285 51.245 ;
        RECT 103.795 51.075 103.965 51.245 ;
        RECT 105.180 51.075 105.350 51.245 ;
        RECT 107.935 51.075 108.105 51.245 ;
        RECT 109.315 51.075 109.485 51.245 ;
        RECT 111.615 51.075 111.785 51.245 ;
        RECT 113.455 51.075 113.625 51.245 ;
        RECT 120.355 51.075 120.525 51.245 ;
        RECT 122.195 51.075 122.365 51.245 ;
        RECT 125.875 51.075 126.045 51.245 ;
        RECT 127.255 51.075 127.425 51.245 ;
        RECT 134.615 51.075 134.785 51.245 ;
        RECT 135.995 51.075 136.165 51.245 ;
        RECT 139.675 51.075 139.845 51.245 ;
        RECT 140.145 51.100 140.305 51.210 ;
        RECT 141.515 51.075 141.685 51.245 ;
        RECT 148.415 51.075 148.585 51.245 ;
        RECT 150.255 51.075 150.425 51.245 ;
        RECT 153.935 51.075 154.105 51.245 ;
        RECT 155.315 51.075 155.485 51.245 ;
        RECT 162.675 51.075 162.845 51.245 ;
        RECT 164.055 51.075 164.225 51.245 ;
        RECT 168.205 51.100 168.365 51.210 ;
        RECT 169.575 51.075 169.745 51.245 ;
        RECT 170.495 51.075 170.665 51.245 ;
        RECT 178.315 51.075 178.485 51.245 ;
        RECT 179.235 51.075 179.405 51.245 ;
        RECT 181.995 51.075 182.165 51.245 ;
        RECT 183.375 51.075 183.545 51.245 ;
        RECT 185.215 51.075 185.385 51.245 ;
        RECT 190.735 51.075 190.905 51.245 ;
        RECT 193.955 51.075 194.125 51.245 ;
        RECT 195.335 51.075 195.505 51.245 ;
        RECT 195.795 51.075 195.965 51.245 ;
        RECT 197.635 51.215 197.805 51.245 ;
        RECT 197.630 51.105 197.805 51.215 ;
        RECT 197.635 51.075 197.805 51.105 ;
        RECT 198.095 51.075 198.265 51.245 ;
        RECT 206.375 51.075 206.545 51.245 ;
        RECT 206.835 51.075 207.005 51.245 ;
        RECT 210.060 51.075 210.230 51.245 ;
        RECT 210.510 51.105 210.630 51.215 ;
        RECT 211.445 51.110 211.605 51.220 ;
        RECT 212.360 51.075 212.530 51.245 ;
        RECT 217.415 51.075 217.585 51.245 ;
        RECT 219.715 51.075 219.885 51.245 ;
        RECT 222.935 51.075 223.105 51.245 ;
        RECT 223.400 51.075 223.570 51.245 ;
        RECT 224.770 51.105 224.890 51.215 ;
        RECT 225.695 51.075 225.865 51.245 ;
        RECT 227.535 51.075 227.705 51.245 ;
        RECT 229.370 51.105 229.490 51.215 ;
        RECT 229.835 51.075 230.005 51.245 ;
        RECT 231.215 51.075 231.385 51.245 ;
        RECT 233.975 51.075 234.145 51.245 ;
        RECT 235.355 51.075 235.525 51.245 ;
        RECT 237.660 51.075 237.830 51.245 ;
        RECT 239.495 51.075 239.665 51.245 ;
        RECT 241.335 51.075 241.505 51.245 ;
        RECT 245.015 51.075 245.190 51.245 ;
        RECT 250.535 51.075 250.705 51.245 ;
        RECT 252.375 51.075 252.545 51.245 ;
        RECT 253.760 51.075 253.930 51.245 ;
        RECT 256.060 51.075 256.230 51.245 ;
        RECT 261.115 51.075 261.285 51.245 ;
        RECT 263.415 51.075 263.585 51.245 ;
        RECT 264.795 51.075 264.965 51.245 ;
        RECT 266.635 51.075 266.805 51.245 ;
        RECT 267.555 51.075 267.725 51.245 ;
        RECT 270.320 51.075 270.490 51.245 ;
        RECT 271.240 51.075 271.410 51.245 ;
        RECT 277.675 51.075 277.845 51.245 ;
        RECT 278.595 51.075 278.765 51.245 ;
        RECT 281.820 51.075 281.990 51.245 ;
        RECT 282.280 51.075 282.450 51.245 ;
        RECT 285.955 51.075 286.125 51.245 ;
        RECT 289.635 51.075 289.810 51.245 ;
        RECT 295.620 51.075 295.790 51.245 ;
        RECT 296.995 51.075 297.165 51.245 ;
        RECT 299.755 51.075 299.925 51.245 ;
        RECT 300.680 51.075 300.850 51.245 ;
        RECT 304.815 51.075 304.985 51.245 ;
        RECT 305.285 51.110 305.445 51.220 ;
        RECT 306.200 51.075 306.370 51.245 ;
        RECT 308.505 51.100 308.665 51.210 ;
        RECT 309.875 51.075 310.045 51.245 ;
        RECT 313.555 51.075 313.725 51.245 ;
        RECT 314.480 51.075 314.650 51.245 ;
        RECT 317.235 51.075 317.405 51.245 ;
        RECT 318.615 51.075 318.785 51.245 ;
        RECT 319.075 51.075 319.245 51.245 ;
        RECT 322.305 51.100 322.465 51.210 ;
        RECT 322.750 51.105 322.870 51.215 ;
        RECT 323.220 51.075 323.390 51.245 ;
        RECT 323.675 51.075 323.845 51.245 ;
        RECT 325.515 51.075 325.685 51.245 ;
        RECT 329.200 51.075 329.370 51.245 ;
        RECT 330.575 51.075 330.745 51.245 ;
        RECT 336.095 51.075 336.265 51.245 ;
        RECT 336.555 51.075 336.725 51.245 ;
        RECT 337.935 51.075 338.105 51.245 ;
        RECT 339.775 51.075 339.945 51.245 ;
        RECT 340.240 51.075 340.410 51.245 ;
        RECT 343.460 51.075 343.630 51.245 ;
        RECT 347.595 51.075 347.765 51.245 ;
        RECT 350.815 51.075 350.985 51.245 ;
        RECT 351.740 51.075 351.910 51.245 ;
        RECT 354.500 51.075 354.670 51.245 ;
        RECT 358.635 51.075 358.805 51.245 ;
        RECT 359.095 51.075 359.265 51.245 ;
        RECT 362.780 51.075 362.950 51.245 ;
        RECT 364.155 51.075 364.325 51.245 ;
        RECT 366.000 51.075 366.170 51.245 ;
        RECT 366.915 51.075 367.085 51.245 ;
        RECT 370.135 51.075 370.305 51.245 ;
        RECT 370.600 51.075 370.770 51.245 ;
        RECT 373.820 51.075 373.990 51.245 ;
        RECT 374.735 51.075 374.905 51.245 ;
        RECT 377.955 51.075 378.125 51.245 ;
        RECT 378.425 51.110 378.585 51.220 ;
        RECT 379.795 51.075 379.965 51.245 ;
        RECT 381.175 51.075 381.345 51.245 ;
        RECT 381.635 51.075 381.805 51.245 ;
        RECT 383.015 51.075 383.185 51.245 ;
        RECT 384.855 51.075 385.025 51.245 ;
        RECT 386.235 51.075 386.405 51.245 ;
        RECT 386.695 51.075 386.865 51.245 ;
        RECT 388.075 51.075 388.245 51.245 ;
        RECT 389.915 51.075 390.085 51.245 ;
        RECT 391.295 51.075 391.465 51.245 ;
        RECT 394.055 51.075 394.225 51.245 ;
        RECT 395.435 51.075 395.605 51.245 ;
        RECT 396.815 51.075 396.985 51.245 ;
        RECT 399.115 51.075 399.285 51.245 ;
        RECT 400.495 51.075 400.665 51.245 ;
        RECT 402.335 51.075 402.505 51.245 ;
        RECT 404.175 51.075 404.345 51.245 ;
        RECT 405.555 51.075 405.725 51.245 ;
        RECT 406.015 51.075 406.185 51.245 ;
        RECT 407.855 51.075 408.025 51.245 ;
        RECT 411.075 51.075 411.245 51.245 ;
        RECT 412.910 51.105 413.030 51.215 ;
        RECT 413.375 51.075 413.545 51.245 ;
        RECT 414.755 51.075 414.925 51.245 ;
        RECT 418.895 51.075 419.065 51.245 ;
        RECT 420.275 51.075 420.445 51.245 ;
        RECT 422.115 51.075 422.285 51.245 ;
        RECT 424.415 51.075 424.585 51.245 ;
        RECT 427.630 51.105 427.750 51.215 ;
        RECT 428.095 51.075 428.265 51.245 ;
        RECT 429.475 51.075 429.645 51.245 ;
        RECT 429.935 51.075 430.105 51.245 ;
        RECT 434.990 51.105 435.110 51.215 ;
        RECT 435.455 51.075 435.625 51.245 ;
        RECT 435.915 51.075 436.085 51.245 ;
        RECT 436.835 51.075 437.005 51.245 ;
        RECT 441.435 51.075 441.605 51.245 ;
        RECT 442.355 51.075 442.525 51.245 ;
        RECT 446.955 51.075 447.125 51.245 ;
        RECT 447.875 51.075 448.045 51.245 ;
        RECT 450.175 51.075 450.345 51.245 ;
        RECT 451.555 51.075 451.725 51.245 ;
        RECT 452.475 51.075 452.645 51.245 ;
        RECT 457.070 51.105 457.190 51.215 ;
        RECT 457.535 51.075 457.705 51.245 ;
        RECT 457.995 51.075 458.165 51.245 ;
        RECT 458.915 51.075 459.085 51.245 ;
        RECT 463.975 51.075 464.145 51.245 ;
        RECT 464.435 51.075 464.605 51.245 ;
        RECT 468.110 51.105 468.230 51.215 ;
        RECT 468.575 51.075 468.745 51.245 ;
        RECT 469.495 51.075 469.665 51.245 ;
        RECT 469.955 51.075 470.125 51.245 ;
        RECT 475.015 51.075 475.185 51.245 ;
        RECT 475.475 51.075 475.645 51.245 ;
        RECT 477.310 51.105 477.430 51.215 ;
        RECT 478.235 51.075 478.405 51.245 ;
        RECT 479.615 51.075 479.785 51.245 ;
        RECT 480.535 51.075 480.705 51.245 ;
        RECT 480.995 51.075 481.165 51.245 ;
        RECT 486.055 51.075 486.225 51.245 ;
        RECT 486.510 51.105 486.630 51.215 ;
        RECT 486.975 51.075 487.145 51.245 ;
        RECT 488.355 51.075 488.525 51.245 ;
        RECT 492.035 51.075 492.205 51.245 ;
        RECT 493.875 51.075 494.045 51.245 ;
        RECT 497.555 51.075 497.725 51.245 ;
        RECT 499.395 51.075 499.565 51.245 ;
        RECT 503.075 51.075 503.245 51.245 ;
        RECT 504.925 51.100 505.085 51.210 ;
        RECT 506.295 51.075 506.465 51.245 ;
        RECT 508.595 51.075 508.765 51.245 ;
        RECT 511.825 51.100 511.985 51.210 ;
        RECT 512.735 51.075 512.905 51.245 ;
        RECT 514.115 51.075 514.285 51.245 ;
        RECT 519.630 51.105 519.750 51.215 ;
        RECT 520.095 51.075 520.265 51.245 ;
        RECT 521.475 51.075 521.645 51.245 ;
        RECT 525.615 51.075 525.785 51.245 ;
        RECT 526.995 51.075 527.165 51.245 ;
        RECT 531.135 51.075 531.305 51.245 ;
        RECT 532.515 51.075 532.685 51.245 ;
        RECT 534.350 51.105 534.470 51.215 ;
        RECT 534.815 51.075 534.985 51.245 ;
        RECT 536.195 51.075 536.365 51.245 ;
        RECT 536.655 51.075 536.825 51.245 ;
        RECT 541.710 51.105 541.830 51.215 ;
        RECT 542.175 51.075 542.345 51.245 ;
        RECT 543.555 51.075 543.725 51.245 ;
        RECT 548.155 51.075 548.325 51.245 ;
        RECT 549.075 51.075 549.245 51.245 ;
        RECT 552.750 51.105 552.870 51.215 ;
        RECT 553.215 51.075 553.385 51.245 ;
        RECT 553.675 51.075 553.845 51.245 ;
        RECT 554.595 51.075 554.765 51.245 ;
        RECT 559.195 51.075 559.365 51.245 ;
        RECT 560.115 51.075 560.285 51.245 ;
        RECT 562.415 51.075 562.585 51.245 ;
        RECT 563.795 51.075 563.965 51.245 ;
        RECT 564.715 51.075 564.885 51.245 ;
        RECT 565.175 51.075 565.345 51.245 ;
        RECT 570.235 51.075 570.405 51.245 ;
        RECT 570.690 51.105 570.810 51.215 ;
        RECT 571.155 51.075 571.325 51.245 ;
        RECT 572.535 51.075 572.705 51.245 ;
        RECT 576.215 51.075 576.385 51.245 ;
        RECT 578.055 51.075 578.225 51.245 ;
        RECT 581.735 51.075 581.905 51.245 ;
        RECT 583.575 51.075 583.745 51.245 ;
        RECT 587.255 51.075 587.425 51.245 ;
        RECT 589.105 51.100 589.265 51.210 ;
        RECT 590.475 51.075 590.645 51.245 ;
        RECT 592.775 51.075 592.945 51.245 ;
        RECT 596.005 51.100 596.165 51.210 ;
        RECT 596.915 51.075 597.085 51.245 ;
        RECT 598.295 51.075 598.465 51.245 ;
        RECT 603.810 51.105 603.930 51.215 ;
        RECT 604.275 51.075 604.445 51.245 ;
        RECT 605.655 51.075 605.825 51.245 ;
        RECT 609.795 51.075 609.965 51.245 ;
        RECT 611.175 51.075 611.345 51.245 ;
        RECT 615.315 51.075 615.485 51.245 ;
        RECT 616.695 51.075 616.865 51.245 ;
        RECT 618.530 51.105 618.650 51.215 ;
        RECT 618.995 51.075 619.165 51.245 ;
        RECT 620.375 51.075 620.545 51.245 ;
        RECT 620.835 51.075 621.005 51.245 ;
        RECT 623.590 51.105 623.710 51.215 ;
        RECT 624.055 51.075 624.225 51.245 ;
        RECT 625.435 51.075 625.605 51.245 ;
        RECT 629.125 51.100 629.285 51.220 ;
        RECT 630.955 51.075 631.125 51.245 ;
        RECT 56.875 50.315 57.045 50.840 ;
        RECT 84.935 50.315 85.105 50.840 ;
        RECT 112.995 50.315 113.165 50.840 ;
        RECT 141.055 50.315 141.225 50.840 ;
        RECT 169.115 50.315 169.285 50.840 ;
        RECT 197.175 50.315 197.345 50.840 ;
        RECT 225.235 50.315 225.405 50.840 ;
        RECT 253.295 50.315 253.465 50.840 ;
        RECT 281.355 50.315 281.525 50.840 ;
        RECT 309.415 50.315 309.585 50.840 ;
        RECT 337.475 50.315 337.645 50.840 ;
        RECT 365.535 50.315 365.705 50.840 ;
        RECT 393.595 50.315 393.765 50.840 ;
        RECT 421.655 50.315 421.825 50.840 ;
        RECT 449.715 50.315 449.885 50.840 ;
        RECT 477.775 50.315 477.945 50.840 ;
        RECT 505.835 50.315 506.005 50.840 ;
        RECT 533.895 50.315 534.065 50.840 ;
        RECT 561.955 50.315 562.125 50.840 ;
        RECT 590.015 50.315 590.185 50.840 ;
        RECT 618.075 50.315 618.245 50.840 ;
      LAYER nwell ;
        RECT 42.280 47.025 631.460 49.855 ;
      LAYER pwell ;
        RECT 70.675 46.040 70.845 46.565 ;
        RECT 98.735 46.040 98.905 46.565 ;
        RECT 126.795 46.040 126.965 46.565 ;
        RECT 154.855 46.040 155.025 46.565 ;
        RECT 182.915 46.040 183.085 46.565 ;
        RECT 210.975 46.040 211.145 46.565 ;
        RECT 239.035 46.040 239.205 46.565 ;
        RECT 267.095 46.040 267.265 46.565 ;
        RECT 295.155 46.040 295.325 46.565 ;
        RECT 323.215 46.040 323.385 46.565 ;
        RECT 351.275 46.040 351.445 46.565 ;
        RECT 379.335 46.040 379.505 46.565 ;
        RECT 407.395 46.040 407.565 46.565 ;
        RECT 435.455 46.040 435.625 46.565 ;
        RECT 463.515 46.040 463.685 46.565 ;
        RECT 491.575 46.040 491.745 46.565 ;
        RECT 519.635 46.040 519.805 46.565 ;
        RECT 547.695 46.040 547.865 46.565 ;
        RECT 575.755 46.040 575.925 46.565 ;
        RECT 603.815 46.040 603.985 46.565 ;
        RECT 42.615 45.635 42.785 45.805 ;
        RECT 43.995 45.635 44.165 45.805 ;
        RECT 49.515 45.635 49.685 45.805 ;
        RECT 55.035 45.635 55.205 45.805 ;
        RECT 57.335 45.635 57.505 45.805 ;
        RECT 60.555 45.635 60.725 45.805 ;
        RECT 62.855 45.635 63.025 45.805 ;
        RECT 66.075 45.635 66.245 45.805 ;
        RECT 68.375 45.635 68.545 45.805 ;
        RECT 69.765 45.670 69.925 45.780 ;
        RECT 71.135 45.635 71.305 45.805 ;
        RECT 71.595 45.635 71.765 45.805 ;
        RECT 72.515 45.635 72.685 45.805 ;
        RECT 73.895 45.635 74.065 45.805 ;
        RECT 77.115 45.635 77.285 45.805 ;
        RECT 77.575 45.635 77.745 45.805 ;
        RECT 78.500 45.635 78.670 45.805 ;
        RECT 80.795 45.635 80.965 45.805 ;
        RECT 81.715 45.635 81.885 45.805 ;
        RECT 84.485 45.670 84.645 45.780 ;
        RECT 85.395 45.635 85.565 45.805 ;
        RECT 85.865 45.660 86.025 45.770 ;
        RECT 86.775 45.635 86.945 45.805 ;
        RECT 87.235 45.635 87.405 45.805 ;
        RECT 88.155 45.635 88.325 45.805 ;
        RECT 90.920 45.635 91.090 45.805 ;
        RECT 91.840 45.635 92.010 45.805 ;
        RECT 95.055 45.635 95.225 45.805 ;
        RECT 95.975 45.635 96.145 45.805 ;
        RECT 99.195 45.635 99.365 45.805 ;
        RECT 100.110 45.665 100.230 45.775 ;
        RECT 100.575 45.635 100.745 45.805 ;
        RECT 102.415 45.635 102.585 45.805 ;
        RECT 102.870 45.665 102.990 45.775 ;
        RECT 103.340 45.635 103.510 45.805 ;
        RECT 106.090 45.635 106.260 45.805 ;
        RECT 107.475 45.635 107.645 45.805 ;
        RECT 110.235 45.635 110.405 45.805 ;
        RECT 111.160 45.635 111.330 45.805 ;
        RECT 114.385 45.660 114.545 45.770 ;
        RECT 115.290 45.635 115.465 45.805 ;
        RECT 118.970 45.635 119.140 45.805 ;
        RECT 119.435 45.635 119.605 45.805 ;
        RECT 123.115 45.635 123.285 45.805 ;
        RECT 124.495 45.635 124.665 45.805 ;
        RECT 127.250 45.665 127.370 45.775 ;
        RECT 127.715 45.635 127.885 45.805 ;
        RECT 128.630 45.635 128.800 45.805 ;
        RECT 132.775 45.635 132.945 45.805 ;
        RECT 136.455 45.775 136.625 45.805 ;
        RECT 136.450 45.665 136.625 45.775 ;
        RECT 136.455 45.635 136.625 45.665 ;
        RECT 136.915 45.635 137.085 45.805 ;
        RECT 138.755 45.635 138.925 45.805 ;
        RECT 141.975 45.635 142.145 45.805 ;
        RECT 142.890 45.665 143.010 45.775 ;
        RECT 143.355 45.635 143.525 45.805 ;
        RECT 143.820 45.635 143.990 45.805 ;
        RECT 145.195 45.635 145.365 45.805 ;
        RECT 148.880 45.635 149.050 45.805 ;
        RECT 151.175 45.635 151.345 45.805 ;
        RECT 153.015 45.635 153.185 45.805 ;
        RECT 155.315 45.635 155.485 45.805 ;
        RECT 157.155 45.635 157.325 45.805 ;
        RECT 164.055 45.635 164.225 45.805 ;
        RECT 165.895 45.635 166.065 45.805 ;
        RECT 167.735 45.635 167.905 45.805 ;
        RECT 169.115 45.635 169.285 45.805 ;
        RECT 169.575 45.635 169.745 45.805 ;
        RECT 171.415 45.635 171.585 45.805 ;
        RECT 173.250 45.665 173.370 45.775 ;
        RECT 173.720 45.635 173.890 45.805 ;
        RECT 177.855 45.635 178.025 45.805 ;
        RECT 181.075 45.635 181.245 45.805 ;
        RECT 181.535 45.635 181.705 45.805 ;
        RECT 183.375 45.635 183.545 45.805 ;
        RECT 184.755 45.775 184.925 45.805 ;
        RECT 184.750 45.665 184.925 45.775 ;
        RECT 185.670 45.665 185.790 45.775 ;
        RECT 184.755 45.635 184.925 45.665 ;
        RECT 186.135 45.635 186.305 45.805 ;
        RECT 193.495 45.635 193.665 45.805 ;
        RECT 194.875 45.635 195.045 45.805 ;
        RECT 197.175 45.635 197.345 45.805 ;
        RECT 198.565 45.660 198.725 45.770 ;
        RECT 199.935 45.635 200.105 45.805 ;
        RECT 203.610 45.665 203.730 45.775 ;
        RECT 204.075 45.635 204.245 45.805 ;
        RECT 205.915 45.635 206.085 45.805 ;
        RECT 209.595 45.635 209.765 45.805 ;
        RECT 211.430 45.635 211.600 45.805 ;
        RECT 213.270 45.665 213.390 45.775 ;
        RECT 214.195 45.635 214.365 45.805 ;
        RECT 215.575 45.635 215.745 45.805 ;
        RECT 218.335 45.635 218.505 45.805 ;
        RECT 219.255 45.635 219.425 45.805 ;
        RECT 222.015 45.635 222.185 45.805 ;
        RECT 223.395 45.635 223.565 45.805 ;
        RECT 223.855 45.635 224.025 45.805 ;
        RECT 227.530 45.665 227.650 45.775 ;
        RECT 228.460 45.635 228.630 45.805 ;
        RECT 228.915 45.635 229.085 45.805 ;
        RECT 230.750 45.635 230.920 45.805 ;
        RECT 232.595 45.635 232.765 45.805 ;
        RECT 234.895 45.635 235.065 45.805 ;
        RECT 236.275 45.635 236.445 45.805 ;
        RECT 238.115 45.635 238.285 45.805 ;
        RECT 238.570 45.665 238.690 45.775 ;
        RECT 239.500 45.635 239.670 45.805 ;
        RECT 241.790 45.665 241.910 45.775 ;
        RECT 242.720 45.635 242.890 45.805 ;
        RECT 245.935 45.635 246.105 45.805 ;
        RECT 246.855 45.635 247.025 45.805 ;
        RECT 249.620 45.635 249.790 45.805 ;
        RECT 250.530 45.635 250.700 45.805 ;
        RECT 252.835 45.635 253.005 45.805 ;
        RECT 254.675 45.635 254.845 45.805 ;
        RECT 256.980 45.635 257.150 45.805 ;
        RECT 258.360 45.635 258.530 45.805 ;
        RECT 260.195 45.635 260.365 45.805 ;
        RECT 261.575 45.635 261.745 45.805 ;
        RECT 263.875 45.635 264.045 45.805 ;
        RECT 265.715 45.635 265.885 45.805 ;
        RECT 267.555 45.635 267.725 45.805 ;
        RECT 269.395 45.635 269.565 45.805 ;
        RECT 271.235 45.635 271.405 45.805 ;
        RECT 273.075 45.635 273.250 45.805 ;
        RECT 276.760 45.635 276.930 45.805 ;
        RECT 277.215 45.635 277.385 45.805 ;
        RECT 280.895 45.635 281.065 45.805 ;
        RECT 282.735 45.635 282.905 45.805 ;
        RECT 284.115 45.635 284.285 45.805 ;
        RECT 284.570 45.665 284.690 45.775 ;
        RECT 285.035 45.635 285.205 45.805 ;
        RECT 285.500 45.635 285.670 45.805 ;
        RECT 289.635 45.635 289.805 45.805 ;
        RECT 291.475 45.635 291.645 45.805 ;
        RECT 293.315 45.635 293.485 45.805 ;
        RECT 295.155 45.635 295.325 45.805 ;
        RECT 295.620 45.635 295.790 45.805 ;
        RECT 298.830 45.665 298.950 45.775 ;
        RECT 299.755 45.635 299.930 45.805 ;
        RECT 303.440 45.635 303.610 45.805 ;
        RECT 303.895 45.635 304.065 45.805 ;
        RECT 307.575 45.635 307.745 45.805 ;
        RECT 309.415 45.635 309.585 45.805 ;
        RECT 311.260 45.635 311.430 45.805 ;
        RECT 313.090 45.665 313.210 45.775 ;
        RECT 314.020 45.635 314.190 45.805 ;
        RECT 315.395 45.635 315.565 45.805 ;
        RECT 318.155 45.635 318.325 45.805 ;
        RECT 320.915 45.635 321.085 45.805 ;
        RECT 321.835 45.635 322.005 45.805 ;
        RECT 322.750 45.665 322.870 45.775 ;
        RECT 323.675 45.635 323.850 45.805 ;
        RECT 327.350 45.665 327.470 45.775 ;
        RECT 327.815 45.635 327.985 45.805 ;
        RECT 328.280 45.635 328.450 45.805 ;
        RECT 331.500 45.635 331.670 45.805 ;
        RECT 332.415 45.635 332.585 45.805 ;
        RECT 335.635 45.635 335.805 45.805 ;
        RECT 336.095 45.635 336.265 45.805 ;
        RECT 337.935 45.635 338.105 45.805 ;
        RECT 339.320 45.635 339.490 45.805 ;
        RECT 341.610 45.665 341.730 45.775 ;
        RECT 342.535 45.635 342.705 45.805 ;
        RECT 343.455 45.635 343.625 45.805 ;
        RECT 344.370 45.665 344.490 45.775 ;
        RECT 344.835 45.635 345.005 45.805 ;
        RECT 345.755 45.635 345.925 45.805 ;
        RECT 348.975 45.635 349.145 45.805 ;
        RECT 350.810 45.665 350.930 45.775 ;
        RECT 351.740 45.635 351.910 45.805 ;
        RECT 352.195 45.635 352.365 45.805 ;
        RECT 355.875 45.775 356.045 45.805 ;
        RECT 355.870 45.665 356.045 45.775 ;
        RECT 355.875 45.635 356.045 45.665 ;
        RECT 356.800 45.635 356.970 45.805 ;
        RECT 359.560 45.635 359.730 45.805 ;
        RECT 360.935 45.635 361.105 45.805 ;
        RECT 363.695 45.635 363.865 45.805 ;
        RECT 364.615 45.635 364.785 45.805 ;
        RECT 365.995 45.635 366.165 45.805 ;
        RECT 367.380 45.635 367.550 45.805 ;
        RECT 369.685 45.660 369.845 45.770 ;
        RECT 371.060 45.635 371.230 45.805 ;
        RECT 371.515 45.635 371.685 45.805 ;
        RECT 375.195 45.635 375.365 45.805 ;
        RECT 377.035 45.635 377.205 45.805 ;
        RECT 378.875 45.775 379.045 45.805 ;
        RECT 378.870 45.665 379.045 45.775 ;
        RECT 378.875 45.635 379.045 45.665 ;
        RECT 379.795 45.635 379.965 45.805 ;
        RECT 380.255 45.635 380.425 45.805 ;
        RECT 381.175 45.635 381.345 45.805 ;
        RECT 383.945 45.660 384.105 45.770 ;
        RECT 384.855 45.635 385.025 45.805 ;
        RECT 385.315 45.635 385.485 45.805 ;
        RECT 386.235 45.635 386.405 45.805 ;
        RECT 386.695 45.635 386.865 45.805 ;
        RECT 389.915 45.635 390.085 45.805 ;
        RECT 390.375 45.635 390.545 45.805 ;
        RECT 391.295 45.635 391.465 45.805 ;
        RECT 391.755 45.635 391.925 45.805 ;
        RECT 394.975 45.635 395.145 45.805 ;
        RECT 396.355 45.635 396.525 45.805 ;
        RECT 397.275 45.635 397.445 45.805 ;
        RECT 399.575 45.635 399.745 45.805 ;
        RECT 400.035 45.635 400.205 45.805 ;
        RECT 401.415 45.635 401.585 45.805 ;
        RECT 405.095 45.635 405.265 45.805 ;
        RECT 406.930 45.665 407.050 45.775 ;
        RECT 407.855 45.635 408.025 45.805 ;
        RECT 409.235 45.635 409.405 45.805 ;
        RECT 410.615 45.635 410.785 45.805 ;
        RECT 412.915 45.635 413.085 45.805 ;
        RECT 413.835 45.635 414.005 45.805 ;
        RECT 414.295 45.635 414.465 45.805 ;
        RECT 417.975 45.635 418.145 45.805 ;
        RECT 419.355 45.635 419.525 45.805 ;
        RECT 423.035 45.635 423.205 45.805 ;
        RECT 424.415 45.635 424.585 45.805 ;
        RECT 424.875 45.635 425.045 45.805 ;
        RECT 428.095 45.635 428.265 45.805 ;
        RECT 429.475 45.635 429.645 45.805 ;
        RECT 433.615 45.635 433.785 45.805 ;
        RECT 434.990 45.665 435.110 45.775 ;
        RECT 435.915 45.635 436.085 45.805 ;
        RECT 437.295 45.635 437.465 45.805 ;
        RECT 439.135 45.635 439.305 45.805 ;
        RECT 440.975 45.635 441.145 45.805 ;
        RECT 442.355 45.635 442.525 45.805 ;
        RECT 446.035 45.635 446.205 45.805 ;
        RECT 447.415 45.635 447.585 45.805 ;
        RECT 447.875 45.635 448.045 45.805 ;
        RECT 451.095 45.635 451.265 45.805 ;
        RECT 452.475 45.635 452.645 45.805 ;
        RECT 453.395 45.635 453.565 45.805 ;
        RECT 456.155 45.635 456.325 45.805 ;
        RECT 456.615 45.635 456.785 45.805 ;
        RECT 457.535 45.635 457.705 45.805 ;
        RECT 462.135 45.635 462.305 45.805 ;
        RECT 463.050 45.665 463.170 45.775 ;
        RECT 463.975 45.635 464.145 45.805 ;
        RECT 465.355 45.635 465.525 45.805 ;
        RECT 467.655 45.635 467.825 45.805 ;
        RECT 469.035 45.635 469.205 45.805 ;
        RECT 470.415 45.635 470.585 45.805 ;
        RECT 470.875 45.635 471.045 45.805 ;
        RECT 474.095 45.635 474.265 45.805 ;
        RECT 475.475 45.635 475.645 45.805 ;
        RECT 476.395 45.635 476.565 45.805 ;
        RECT 479.155 45.635 479.325 45.805 ;
        RECT 480.535 45.635 480.705 45.805 ;
        RECT 481.915 45.635 482.085 45.805 ;
        RECT 484.215 45.635 484.385 45.805 ;
        RECT 485.135 45.635 485.305 45.805 ;
        RECT 485.595 45.635 485.765 45.805 ;
        RECT 490.655 45.635 490.825 45.805 ;
        RECT 491.110 45.665 491.230 45.775 ;
        RECT 492.035 45.635 492.205 45.805 ;
        RECT 493.415 45.635 493.585 45.805 ;
        RECT 496.175 45.635 496.345 45.805 ;
        RECT 497.095 45.635 497.265 45.805 ;
        RECT 498.475 45.635 498.645 45.805 ;
        RECT 499.395 45.635 499.565 45.805 ;
        RECT 501.230 45.665 501.350 45.775 ;
        RECT 501.695 45.635 501.865 45.805 ;
        RECT 502.155 45.635 502.325 45.805 ;
        RECT 503.075 45.635 503.245 45.805 ;
        RECT 503.535 45.635 503.705 45.805 ;
        RECT 507.215 45.635 507.385 45.805 ;
        RECT 508.595 45.635 508.765 45.805 ;
        RECT 512.275 45.635 512.445 45.805 ;
        RECT 513.655 45.635 513.825 45.805 ;
        RECT 519.175 45.775 519.345 45.805 ;
        RECT 519.170 45.665 519.345 45.775 ;
        RECT 519.175 45.635 519.345 45.665 ;
        RECT 520.095 45.635 520.265 45.805 ;
        RECT 521.475 45.635 521.645 45.805 ;
        RECT 524.695 45.635 524.865 45.805 ;
        RECT 525.155 45.635 525.325 45.805 ;
        RECT 526.535 45.635 526.705 45.805 ;
        RECT 527.915 45.635 528.085 45.805 ;
        RECT 530.215 45.635 530.385 45.805 ;
        RECT 531.595 45.635 531.765 45.805 ;
        RECT 533.435 45.635 533.605 45.805 ;
        RECT 535.275 45.635 535.445 45.805 ;
        RECT 536.655 45.635 536.825 45.805 ;
        RECT 538.955 45.635 539.125 45.805 ;
        RECT 540.335 45.635 540.505 45.805 ;
        RECT 541.715 45.635 541.885 45.805 ;
        RECT 542.175 45.635 542.345 45.805 ;
        RECT 547.230 45.665 547.350 45.775 ;
        RECT 547.695 45.635 547.865 45.805 ;
        RECT 548.155 45.635 548.325 45.805 ;
        RECT 549.535 45.635 549.705 45.805 ;
        RECT 553.215 45.635 553.385 45.805 ;
        RECT 554.595 45.635 554.765 45.805 ;
        RECT 556.435 45.635 556.605 45.805 ;
        RECT 558.275 45.635 558.445 45.805 ;
        RECT 559.655 45.635 559.825 45.805 ;
        RECT 561.955 45.635 562.125 45.805 ;
        RECT 563.335 45.635 563.505 45.805 ;
        RECT 564.715 45.635 564.885 45.805 ;
        RECT 567.475 45.635 567.645 45.805 ;
        RECT 568.395 45.635 568.565 45.805 ;
        RECT 569.775 45.635 569.945 45.805 ;
        RECT 570.695 45.635 570.865 45.805 ;
        RECT 575.290 45.665 575.410 45.775 ;
        RECT 576.215 45.635 576.385 45.805 ;
        RECT 577.595 45.635 577.765 45.805 ;
        RECT 581.275 45.635 581.445 45.805 ;
        RECT 581.735 45.635 581.905 45.805 ;
        RECT 582.655 45.635 582.825 45.805 ;
        RECT 584.965 45.660 585.125 45.770 ;
        RECT 585.875 45.635 586.045 45.805 ;
        RECT 586.335 45.635 586.505 45.805 ;
        RECT 587.255 45.635 587.425 45.805 ;
        RECT 587.715 45.635 587.885 45.805 ;
        RECT 591.395 45.635 591.565 45.805 ;
        RECT 592.775 45.635 592.945 45.805 ;
        RECT 596.455 45.635 596.625 45.805 ;
        RECT 597.835 45.635 598.005 45.805 ;
        RECT 598.290 45.665 598.410 45.775 ;
        RECT 599.215 45.635 599.385 45.805 ;
        RECT 603.350 45.665 603.470 45.775 ;
        RECT 604.275 45.635 604.445 45.805 ;
        RECT 604.735 45.635 604.905 45.805 ;
        RECT 605.655 45.635 605.825 45.805 ;
        RECT 609.335 45.635 609.505 45.805 ;
        RECT 610.255 45.635 610.425 45.805 ;
        RECT 610.715 45.635 610.885 45.805 ;
        RECT 613.475 45.635 613.645 45.805 ;
        RECT 614.395 45.635 614.565 45.805 ;
        RECT 615.775 45.635 615.945 45.805 ;
        RECT 618.995 45.635 619.165 45.805 ;
        RECT 619.455 45.635 619.625 45.805 ;
        RECT 620.835 45.635 621.005 45.805 ;
        RECT 621.750 45.665 621.870 45.775 ;
        RECT 622.215 45.635 622.385 45.805 ;
        RECT 623.595 45.635 623.765 45.805 ;
        RECT 624.515 45.635 624.685 45.805 ;
        RECT 625.895 45.635 626.065 45.805 ;
        RECT 627.735 45.635 627.905 45.805 ;
        RECT 629.570 45.665 629.690 45.775 ;
        RECT 630.955 45.635 631.125 45.805 ;
        RECT 56.875 44.875 57.045 45.400 ;
        RECT 71.135 44.875 71.305 45.400 ;
        RECT 85.395 44.875 85.565 45.400 ;
        RECT 99.655 44.875 99.825 45.400 ;
        RECT 113.915 44.875 114.085 45.400 ;
        RECT 128.175 44.875 128.345 45.400 ;
        RECT 142.435 44.875 142.605 45.400 ;
        RECT 156.695 44.875 156.865 45.400 ;
        RECT 170.955 44.875 171.125 45.400 ;
        RECT 185.215 44.875 185.385 45.400 ;
        RECT 199.475 44.875 199.645 45.400 ;
        RECT 213.735 44.875 213.905 45.400 ;
        RECT 227.995 44.875 228.165 45.400 ;
        RECT 242.255 44.875 242.425 45.400 ;
        RECT 256.515 44.875 256.685 45.400 ;
        RECT 270.775 44.875 270.945 45.400 ;
        RECT 285.035 44.875 285.205 45.400 ;
        RECT 299.295 44.875 299.465 45.400 ;
        RECT 313.555 44.875 313.725 45.400 ;
        RECT 327.815 44.875 327.985 45.400 ;
        RECT 342.075 44.875 342.245 45.400 ;
        RECT 356.335 44.875 356.505 45.400 ;
        RECT 370.595 44.875 370.765 45.400 ;
        RECT 384.855 44.875 385.025 45.400 ;
        RECT 399.115 44.875 399.285 45.400 ;
        RECT 413.375 44.875 413.545 45.400 ;
        RECT 427.635 44.875 427.805 45.400 ;
        RECT 441.895 44.875 442.065 45.400 ;
        RECT 456.155 44.875 456.325 45.400 ;
        RECT 470.415 44.875 470.585 45.400 ;
        RECT 484.675 44.875 484.845 45.400 ;
        RECT 498.935 44.875 499.105 45.400 ;
        RECT 513.195 44.875 513.365 45.400 ;
        RECT 527.455 44.875 527.625 45.400 ;
        RECT 541.715 44.875 541.885 45.400 ;
        RECT 555.975 44.875 556.145 45.400 ;
        RECT 570.235 44.875 570.405 45.400 ;
        RECT 584.495 44.875 584.665 45.400 ;
        RECT 598.755 44.875 598.925 45.400 ;
        RECT 613.015 44.875 613.185 45.400 ;
        RECT 627.275 44.875 627.445 45.400 ;
      LAYER nwell ;
        RECT 42.280 42.810 631.460 44.415 ;
      LAYER li1 ;
        RECT 42.470 619.555 631.270 619.725 ;
        RECT 42.555 618.465 43.765 619.555 ;
        RECT 43.935 618.465 49.280 619.555 ;
        RECT 49.455 618.465 631.270 619.555 ;
        RECT 42.555 617.755 43.075 618.295 ;
        RECT 43.245 617.925 43.765 618.465 ;
        RECT 43.935 617.775 46.515 618.295 ;
        RECT 46.685 617.945 49.280 618.465 ;
        RECT 49.455 617.775 52.035 618.295 ;
        RECT 52.205 617.945 631.270 618.465 ;
        RECT 54.000 617.775 631.270 617.945 ;
        RECT 42.555 617.005 43.765 617.755 ;
        RECT 43.935 617.005 49.280 617.775 ;
        RECT 49.455 617.005 631.270 617.775 ;
        RECT 42.470 616.835 631.270 617.005 ;
        RECT 42.555 616.085 43.765 616.835 ;
        RECT 42.555 615.545 43.075 616.085 ;
        RECT 43.935 616.065 49.280 616.835 ;
        RECT 49.455 616.065 631.270 616.835 ;
        RECT 43.245 615.375 43.765 615.915 ;
        RECT 43.935 615.545 46.515 616.065 ;
        RECT 46.685 615.375 49.280 615.895 ;
        RECT 49.455 615.545 52.035 616.065 ;
        RECT 54.000 615.895 631.270 616.065 ;
        RECT 52.205 615.375 631.270 615.895 ;
        RECT 42.555 614.285 43.765 615.375 ;
        RECT 43.935 614.285 49.280 615.375 ;
        RECT 49.455 614.285 631.270 615.375 ;
        RECT 42.470 614.115 631.270 614.285 ;
        RECT 42.555 613.025 43.765 614.115 ;
        RECT 43.935 613.025 49.280 614.115 ;
        RECT 49.455 613.025 631.270 614.115 ;
        RECT 42.555 612.315 43.075 612.855 ;
        RECT 43.245 612.485 43.765 613.025 ;
        RECT 43.935 612.335 46.515 612.855 ;
        RECT 46.685 612.505 49.280 613.025 ;
        RECT 49.455 612.335 52.035 612.855 ;
        RECT 52.205 612.505 631.270 613.025 ;
        RECT 54.000 612.335 631.270 612.505 ;
        RECT 42.555 611.565 43.765 612.315 ;
        RECT 43.935 611.565 49.280 612.335 ;
        RECT 49.455 611.565 631.270 612.335 ;
        RECT 42.470 611.395 631.270 611.565 ;
        RECT 42.555 610.645 43.765 611.395 ;
        RECT 42.555 610.105 43.075 610.645 ;
        RECT 43.935 610.625 49.280 611.395 ;
        RECT 49.455 610.625 631.270 611.395 ;
        RECT 43.245 609.935 43.765 610.475 ;
        RECT 43.935 610.105 46.515 610.625 ;
        RECT 46.685 609.935 49.280 610.455 ;
        RECT 49.455 610.105 52.035 610.625 ;
        RECT 54.000 610.455 631.270 610.625 ;
        RECT 52.205 609.935 631.270 610.455 ;
        RECT 42.555 608.845 43.765 609.935 ;
        RECT 43.935 608.845 49.280 609.935 ;
        RECT 49.455 608.845 631.270 609.935 ;
        RECT 42.470 608.675 631.270 608.845 ;
        RECT 42.555 607.585 43.765 608.675 ;
        RECT 43.935 607.585 49.280 608.675 ;
        RECT 49.455 607.585 631.270 608.675 ;
        RECT 42.555 606.875 43.075 607.415 ;
        RECT 43.245 607.045 43.765 607.585 ;
        RECT 43.935 606.895 46.515 607.415 ;
        RECT 46.685 607.065 49.280 607.585 ;
        RECT 49.455 606.895 52.035 607.415 ;
        RECT 52.205 607.065 631.270 607.585 ;
        RECT 54.000 606.895 631.270 607.065 ;
        RECT 42.555 606.125 43.765 606.875 ;
        RECT 43.935 606.125 49.280 606.895 ;
        RECT 49.455 606.125 631.270 606.895 ;
        RECT 42.470 605.955 631.270 606.125 ;
        RECT 42.555 605.205 43.765 605.955 ;
        RECT 42.555 604.665 43.075 605.205 ;
        RECT 43.935 605.185 49.280 605.955 ;
        RECT 49.455 605.185 631.270 605.955 ;
        RECT 43.245 604.495 43.765 605.035 ;
        RECT 43.935 604.665 46.515 605.185 ;
        RECT 46.685 604.495 49.280 605.015 ;
        RECT 49.455 604.665 52.035 605.185 ;
        RECT 54.000 605.015 631.270 605.185 ;
        RECT 52.205 604.495 631.270 605.015 ;
        RECT 42.555 603.405 43.765 604.495 ;
        RECT 43.935 603.405 49.280 604.495 ;
        RECT 49.455 603.405 631.270 604.495 ;
        RECT 42.470 603.235 631.270 603.405 ;
        RECT 42.555 602.145 43.765 603.235 ;
        RECT 43.935 602.145 49.280 603.235 ;
        RECT 49.455 602.145 631.270 603.235 ;
        RECT 42.555 601.435 43.075 601.975 ;
        RECT 43.245 601.605 43.765 602.145 ;
        RECT 43.935 601.455 46.515 601.975 ;
        RECT 46.685 601.625 49.280 602.145 ;
        RECT 49.455 601.455 52.035 601.975 ;
        RECT 52.205 601.625 631.270 602.145 ;
        RECT 54.000 601.455 631.270 601.625 ;
        RECT 42.555 600.685 43.765 601.435 ;
        RECT 43.935 600.685 49.280 601.455 ;
        RECT 49.455 600.685 631.270 601.455 ;
        RECT 42.470 600.515 631.270 600.685 ;
        RECT 42.555 599.765 43.765 600.515 ;
        RECT 42.555 599.225 43.075 599.765 ;
        RECT 43.935 599.745 49.280 600.515 ;
        RECT 49.455 599.745 631.270 600.515 ;
        RECT 43.245 599.055 43.765 599.595 ;
        RECT 43.935 599.225 46.515 599.745 ;
        RECT 46.685 599.055 49.280 599.575 ;
        RECT 49.455 599.225 52.035 599.745 ;
        RECT 54.000 599.575 631.270 599.745 ;
        RECT 52.205 599.055 631.270 599.575 ;
        RECT 42.555 597.965 43.765 599.055 ;
        RECT 43.935 597.965 49.280 599.055 ;
        RECT 49.455 597.965 631.270 599.055 ;
        RECT 42.470 597.795 631.270 597.965 ;
        RECT 42.555 596.705 43.765 597.795 ;
        RECT 43.935 596.705 49.280 597.795 ;
        RECT 49.455 596.705 631.270 597.795 ;
        RECT 42.555 595.995 43.075 596.535 ;
        RECT 43.245 596.165 43.765 596.705 ;
        RECT 43.935 596.015 46.515 596.535 ;
        RECT 46.685 596.185 49.280 596.705 ;
        RECT 49.455 596.015 52.035 596.535 ;
        RECT 52.205 596.185 631.270 596.705 ;
        RECT 54.000 596.015 631.270 596.185 ;
        RECT 42.555 595.245 43.765 595.995 ;
        RECT 43.935 595.245 49.280 596.015 ;
        RECT 49.455 595.245 631.270 596.015 ;
        RECT 42.470 595.075 631.270 595.245 ;
        RECT 42.555 594.325 43.765 595.075 ;
        RECT 42.555 593.785 43.075 594.325 ;
        RECT 43.935 594.305 49.280 595.075 ;
        RECT 49.455 594.305 631.270 595.075 ;
        RECT 43.245 593.615 43.765 594.155 ;
        RECT 43.935 593.785 46.515 594.305 ;
        RECT 46.685 593.615 49.280 594.135 ;
        RECT 49.455 593.785 52.035 594.305 ;
        RECT 54.000 594.135 631.270 594.305 ;
        RECT 52.205 593.615 631.270 594.135 ;
        RECT 42.555 592.525 43.765 593.615 ;
        RECT 43.935 592.525 49.280 593.615 ;
        RECT 49.455 592.525 631.270 593.615 ;
        RECT 42.470 592.355 631.270 592.525 ;
        RECT 42.555 591.265 43.765 592.355 ;
        RECT 43.935 591.265 49.280 592.355 ;
        RECT 49.455 591.265 631.270 592.355 ;
        RECT 42.555 590.555 43.075 591.095 ;
        RECT 43.245 590.725 43.765 591.265 ;
        RECT 43.935 590.575 46.515 591.095 ;
        RECT 46.685 590.745 49.280 591.265 ;
        RECT 49.455 590.575 52.035 591.095 ;
        RECT 52.205 590.745 631.270 591.265 ;
        RECT 54.000 590.575 631.270 590.745 ;
        RECT 42.555 589.805 43.765 590.555 ;
        RECT 43.935 589.805 49.280 590.575 ;
        RECT 49.455 589.805 631.270 590.575 ;
        RECT 42.470 589.635 631.270 589.805 ;
        RECT 42.555 588.885 43.765 589.635 ;
        RECT 42.555 588.345 43.075 588.885 ;
        RECT 43.935 588.865 49.280 589.635 ;
        RECT 49.455 588.865 631.270 589.635 ;
        RECT 43.245 588.175 43.765 588.715 ;
        RECT 43.935 588.345 46.515 588.865 ;
        RECT 46.685 588.175 49.280 588.695 ;
        RECT 49.455 588.345 52.035 588.865 ;
        RECT 54.000 588.695 631.270 588.865 ;
        RECT 52.205 588.175 631.270 588.695 ;
        RECT 42.555 587.085 43.765 588.175 ;
        RECT 43.935 587.085 49.280 588.175 ;
        RECT 49.455 587.085 631.270 588.175 ;
        RECT 42.470 586.915 631.270 587.085 ;
        RECT 42.555 585.825 43.765 586.915 ;
        RECT 43.935 585.825 49.280 586.915 ;
        RECT 49.455 585.825 631.270 586.915 ;
        RECT 42.555 585.115 43.075 585.655 ;
        RECT 43.245 585.285 43.765 585.825 ;
        RECT 43.935 585.135 46.515 585.655 ;
        RECT 46.685 585.305 49.280 585.825 ;
        RECT 49.455 585.135 52.035 585.655 ;
        RECT 52.205 585.305 631.270 585.825 ;
        RECT 54.000 585.135 631.270 585.305 ;
        RECT 42.555 584.365 43.765 585.115 ;
        RECT 43.935 584.365 49.280 585.135 ;
        RECT 49.455 584.365 631.270 585.135 ;
        RECT 42.470 584.195 631.270 584.365 ;
        RECT 42.555 583.445 43.765 584.195 ;
        RECT 42.555 582.905 43.075 583.445 ;
        RECT 43.935 583.425 49.280 584.195 ;
        RECT 49.455 583.425 631.270 584.195 ;
        RECT 43.245 582.735 43.765 583.275 ;
        RECT 43.935 582.905 46.515 583.425 ;
        RECT 46.685 582.735 49.280 583.255 ;
        RECT 49.455 582.905 52.035 583.425 ;
        RECT 54.000 583.255 631.270 583.425 ;
        RECT 52.205 582.735 631.270 583.255 ;
        RECT 42.555 581.645 43.765 582.735 ;
        RECT 43.935 581.645 49.280 582.735 ;
        RECT 49.455 581.645 631.270 582.735 ;
        RECT 42.470 581.475 631.270 581.645 ;
        RECT 42.555 580.385 43.765 581.475 ;
        RECT 43.935 580.385 49.280 581.475 ;
        RECT 49.455 580.385 631.270 581.475 ;
        RECT 42.555 579.675 43.075 580.215 ;
        RECT 43.245 579.845 43.765 580.385 ;
        RECT 43.935 579.695 46.515 580.215 ;
        RECT 46.685 579.865 49.280 580.385 ;
        RECT 49.455 579.695 52.035 580.215 ;
        RECT 52.205 579.865 631.270 580.385 ;
        RECT 54.000 579.695 631.270 579.865 ;
        RECT 42.555 578.925 43.765 579.675 ;
        RECT 43.935 578.925 49.280 579.695 ;
        RECT 49.455 578.925 631.270 579.695 ;
        RECT 42.470 578.755 631.270 578.925 ;
        RECT 42.555 578.005 43.765 578.755 ;
        RECT 42.555 577.465 43.075 578.005 ;
        RECT 43.935 577.985 49.280 578.755 ;
        RECT 49.455 577.985 631.270 578.755 ;
        RECT 43.245 577.295 43.765 577.835 ;
        RECT 43.935 577.465 46.515 577.985 ;
        RECT 46.685 577.295 49.280 577.815 ;
        RECT 49.455 577.465 52.035 577.985 ;
        RECT 54.000 577.815 631.270 577.985 ;
        RECT 52.205 577.295 631.270 577.815 ;
        RECT 42.555 576.205 43.765 577.295 ;
        RECT 43.935 576.205 49.280 577.295 ;
        RECT 49.455 576.205 631.270 577.295 ;
        RECT 42.470 576.035 631.270 576.205 ;
        RECT 42.555 574.945 43.765 576.035 ;
        RECT 43.935 574.945 49.280 576.035 ;
        RECT 49.455 574.945 631.270 576.035 ;
        RECT 42.555 574.235 43.075 574.775 ;
        RECT 43.245 574.405 43.765 574.945 ;
        RECT 43.935 574.255 46.515 574.775 ;
        RECT 46.685 574.425 49.280 574.945 ;
        RECT 49.455 574.255 52.035 574.775 ;
        RECT 52.205 574.425 631.270 574.945 ;
        RECT 54.000 574.255 631.270 574.425 ;
        RECT 42.555 573.485 43.765 574.235 ;
        RECT 43.935 573.485 49.280 574.255 ;
        RECT 49.455 573.485 631.270 574.255 ;
        RECT 42.470 573.315 631.270 573.485 ;
        RECT 42.555 572.565 43.765 573.315 ;
        RECT 42.555 572.025 43.075 572.565 ;
        RECT 43.935 572.545 49.280 573.315 ;
        RECT 49.455 572.545 631.270 573.315 ;
        RECT 43.245 571.855 43.765 572.395 ;
        RECT 43.935 572.025 46.515 572.545 ;
        RECT 46.685 571.855 49.280 572.375 ;
        RECT 49.455 572.025 52.035 572.545 ;
        RECT 54.000 572.375 631.270 572.545 ;
        RECT 52.205 571.855 631.270 572.375 ;
        RECT 42.555 570.765 43.765 571.855 ;
        RECT 43.935 570.765 49.280 571.855 ;
        RECT 49.455 570.765 631.270 571.855 ;
        RECT 42.470 570.595 631.270 570.765 ;
        RECT 42.555 569.505 43.765 570.595 ;
        RECT 43.935 569.505 49.280 570.595 ;
        RECT 49.455 569.505 631.270 570.595 ;
        RECT 42.555 568.795 43.075 569.335 ;
        RECT 43.245 568.965 43.765 569.505 ;
        RECT 43.935 568.815 46.515 569.335 ;
        RECT 46.685 568.985 49.280 569.505 ;
        RECT 49.455 568.815 52.035 569.335 ;
        RECT 52.205 568.985 631.270 569.505 ;
        RECT 54.000 568.815 631.270 568.985 ;
        RECT 42.555 568.045 43.765 568.795 ;
        RECT 43.935 568.045 49.280 568.815 ;
        RECT 49.455 568.045 631.270 568.815 ;
        RECT 42.470 567.875 631.270 568.045 ;
        RECT 42.555 567.125 43.765 567.875 ;
        RECT 42.555 566.585 43.075 567.125 ;
        RECT 43.935 567.105 49.280 567.875 ;
        RECT 49.455 567.105 631.270 567.875 ;
        RECT 43.245 566.415 43.765 566.955 ;
        RECT 43.935 566.585 46.515 567.105 ;
        RECT 46.685 566.415 49.280 566.935 ;
        RECT 49.455 566.585 52.035 567.105 ;
        RECT 54.000 566.935 631.270 567.105 ;
        RECT 52.205 566.415 631.270 566.935 ;
        RECT 42.555 565.325 43.765 566.415 ;
        RECT 43.935 565.325 49.280 566.415 ;
        RECT 49.455 565.325 631.270 566.415 ;
        RECT 42.470 565.155 631.270 565.325 ;
        RECT 42.555 564.065 43.765 565.155 ;
        RECT 43.935 564.065 49.280 565.155 ;
        RECT 49.455 564.065 631.270 565.155 ;
        RECT 42.555 563.355 43.075 563.895 ;
        RECT 43.245 563.525 43.765 564.065 ;
        RECT 43.935 563.375 46.515 563.895 ;
        RECT 46.685 563.545 49.280 564.065 ;
        RECT 49.455 563.375 52.035 563.895 ;
        RECT 52.205 563.545 631.270 564.065 ;
        RECT 54.000 563.375 631.270 563.545 ;
        RECT 42.555 562.605 43.765 563.355 ;
        RECT 43.935 562.605 49.280 563.375 ;
        RECT 49.455 562.605 631.270 563.375 ;
        RECT 42.470 562.435 631.270 562.605 ;
        RECT 42.555 561.685 43.765 562.435 ;
        RECT 42.555 561.145 43.075 561.685 ;
        RECT 43.935 561.665 49.280 562.435 ;
        RECT 49.455 561.665 631.270 562.435 ;
        RECT 43.245 560.975 43.765 561.515 ;
        RECT 43.935 561.145 46.515 561.665 ;
        RECT 46.685 560.975 49.280 561.495 ;
        RECT 49.455 561.145 52.035 561.665 ;
        RECT 54.000 561.495 631.270 561.665 ;
        RECT 52.205 560.975 631.270 561.495 ;
        RECT 42.555 559.885 43.765 560.975 ;
        RECT 43.935 559.885 49.280 560.975 ;
        RECT 49.455 559.885 631.270 560.975 ;
        RECT 42.470 559.715 631.270 559.885 ;
        RECT 42.555 558.625 43.765 559.715 ;
        RECT 43.935 558.625 49.280 559.715 ;
        RECT 49.455 558.625 631.270 559.715 ;
        RECT 42.555 557.915 43.075 558.455 ;
        RECT 43.245 558.085 43.765 558.625 ;
        RECT 43.935 557.935 46.515 558.455 ;
        RECT 46.685 558.105 49.280 558.625 ;
        RECT 49.455 557.935 52.035 558.455 ;
        RECT 52.205 558.105 631.270 558.625 ;
        RECT 54.000 557.935 631.270 558.105 ;
        RECT 42.555 557.165 43.765 557.915 ;
        RECT 43.935 557.165 49.280 557.935 ;
        RECT 49.455 557.165 631.270 557.935 ;
        RECT 42.470 556.995 631.270 557.165 ;
        RECT 42.555 556.245 43.765 556.995 ;
        RECT 42.555 555.705 43.075 556.245 ;
        RECT 43.935 556.225 49.280 556.995 ;
        RECT 49.455 556.225 631.270 556.995 ;
        RECT 43.245 555.535 43.765 556.075 ;
        RECT 43.935 555.705 46.515 556.225 ;
        RECT 46.685 555.535 49.280 556.055 ;
        RECT 49.455 555.705 52.035 556.225 ;
        RECT 54.000 556.055 631.270 556.225 ;
        RECT 52.205 555.535 631.270 556.055 ;
        RECT 42.555 554.445 43.765 555.535 ;
        RECT 43.935 554.445 49.280 555.535 ;
        RECT 49.455 554.445 631.270 555.535 ;
        RECT 42.470 554.275 631.270 554.445 ;
        RECT 42.555 553.185 43.765 554.275 ;
        RECT 43.935 553.185 49.280 554.275 ;
        RECT 49.455 553.185 631.270 554.275 ;
        RECT 42.555 552.475 43.075 553.015 ;
        RECT 43.245 552.645 43.765 553.185 ;
        RECT 43.935 552.495 46.515 553.015 ;
        RECT 46.685 552.665 49.280 553.185 ;
        RECT 49.455 552.495 52.035 553.015 ;
        RECT 52.205 552.665 631.270 553.185 ;
        RECT 54.000 552.495 631.270 552.665 ;
        RECT 42.555 551.725 43.765 552.475 ;
        RECT 43.935 551.725 49.280 552.495 ;
        RECT 49.455 551.725 631.270 552.495 ;
        RECT 42.470 551.555 631.270 551.725 ;
        RECT 42.555 550.805 43.765 551.555 ;
        RECT 42.555 550.265 43.075 550.805 ;
        RECT 43.935 550.785 49.280 551.555 ;
        RECT 49.455 550.785 631.270 551.555 ;
        RECT 43.245 550.095 43.765 550.635 ;
        RECT 43.935 550.265 46.515 550.785 ;
        RECT 46.685 550.095 49.280 550.615 ;
        RECT 49.455 550.265 52.035 550.785 ;
        RECT 54.000 550.615 631.270 550.785 ;
        RECT 52.205 550.095 631.270 550.615 ;
        RECT 42.555 549.005 43.765 550.095 ;
        RECT 43.935 549.005 49.280 550.095 ;
        RECT 49.455 549.005 631.270 550.095 ;
        RECT 42.470 548.835 631.270 549.005 ;
        RECT 42.555 547.745 43.765 548.835 ;
        RECT 43.935 547.745 49.280 548.835 ;
        RECT 49.455 547.745 631.270 548.835 ;
        RECT 42.555 547.035 43.075 547.575 ;
        RECT 43.245 547.205 43.765 547.745 ;
        RECT 43.935 547.055 46.515 547.575 ;
        RECT 46.685 547.225 49.280 547.745 ;
        RECT 49.455 547.055 52.035 547.575 ;
        RECT 52.205 547.225 631.270 547.745 ;
        RECT 54.000 547.055 631.270 547.225 ;
        RECT 42.555 546.285 43.765 547.035 ;
        RECT 43.935 546.285 49.280 547.055 ;
        RECT 49.455 546.285 631.270 547.055 ;
        RECT 42.470 546.115 631.270 546.285 ;
        RECT 42.555 545.365 43.765 546.115 ;
        RECT 42.555 544.825 43.075 545.365 ;
        RECT 43.935 545.345 49.280 546.115 ;
        RECT 49.455 545.345 631.270 546.115 ;
        RECT 43.245 544.655 43.765 545.195 ;
        RECT 43.935 544.825 46.515 545.345 ;
        RECT 46.685 544.655 49.280 545.175 ;
        RECT 49.455 544.825 52.035 545.345 ;
        RECT 54.000 545.175 631.270 545.345 ;
        RECT 52.205 544.655 631.270 545.175 ;
        RECT 42.555 543.565 43.765 544.655 ;
        RECT 43.935 543.565 49.280 544.655 ;
        RECT 49.455 543.565 631.270 544.655 ;
        RECT 42.470 543.395 631.270 543.565 ;
        RECT 42.555 542.305 43.765 543.395 ;
        RECT 43.935 542.305 49.280 543.395 ;
        RECT 49.455 542.305 631.270 543.395 ;
        RECT 42.555 541.595 43.075 542.135 ;
        RECT 43.245 541.765 43.765 542.305 ;
        RECT 43.935 541.615 46.515 542.135 ;
        RECT 46.685 541.785 49.280 542.305 ;
        RECT 49.455 541.615 52.035 542.135 ;
        RECT 52.205 541.785 631.270 542.305 ;
        RECT 54.000 541.615 631.270 541.785 ;
        RECT 42.555 540.845 43.765 541.595 ;
        RECT 43.935 540.845 49.280 541.615 ;
        RECT 49.455 540.845 631.270 541.615 ;
        RECT 42.470 540.675 631.270 540.845 ;
        RECT 42.555 539.925 43.765 540.675 ;
        RECT 42.555 539.385 43.075 539.925 ;
        RECT 43.935 539.905 49.280 540.675 ;
        RECT 49.455 539.905 631.270 540.675 ;
        RECT 43.245 539.215 43.765 539.755 ;
        RECT 43.935 539.385 46.515 539.905 ;
        RECT 46.685 539.215 49.280 539.735 ;
        RECT 49.455 539.385 52.035 539.905 ;
        RECT 54.000 539.735 631.270 539.905 ;
        RECT 52.205 539.215 631.270 539.735 ;
        RECT 42.555 538.125 43.765 539.215 ;
        RECT 43.935 538.125 49.280 539.215 ;
        RECT 49.455 538.125 631.270 539.215 ;
        RECT 42.470 537.955 631.270 538.125 ;
        RECT 42.555 536.865 43.765 537.955 ;
        RECT 43.935 536.865 49.280 537.955 ;
        RECT 49.455 536.865 631.270 537.955 ;
        RECT 42.555 536.155 43.075 536.695 ;
        RECT 43.245 536.325 43.765 536.865 ;
        RECT 43.935 536.175 46.515 536.695 ;
        RECT 46.685 536.345 49.280 536.865 ;
        RECT 49.455 536.175 52.035 536.695 ;
        RECT 52.205 536.345 631.270 536.865 ;
        RECT 54.000 536.175 631.270 536.345 ;
        RECT 42.555 535.405 43.765 536.155 ;
        RECT 43.935 535.405 49.280 536.175 ;
        RECT 49.455 535.405 631.270 536.175 ;
        RECT 42.470 535.235 631.270 535.405 ;
        RECT 42.555 534.485 43.765 535.235 ;
        RECT 42.555 533.945 43.075 534.485 ;
        RECT 43.935 534.465 49.280 535.235 ;
        RECT 49.455 534.465 631.270 535.235 ;
        RECT 43.245 533.775 43.765 534.315 ;
        RECT 43.935 533.945 46.515 534.465 ;
        RECT 46.685 533.775 49.280 534.295 ;
        RECT 49.455 533.945 52.035 534.465 ;
        RECT 54.000 534.295 631.270 534.465 ;
        RECT 52.205 533.775 631.270 534.295 ;
        RECT 42.555 532.685 43.765 533.775 ;
        RECT 43.935 532.685 49.280 533.775 ;
        RECT 49.455 532.685 631.270 533.775 ;
        RECT 42.470 532.515 631.270 532.685 ;
        RECT 42.555 531.425 43.765 532.515 ;
        RECT 43.935 531.425 49.280 532.515 ;
        RECT 49.455 531.425 631.270 532.515 ;
        RECT 42.555 530.715 43.075 531.255 ;
        RECT 43.245 530.885 43.765 531.425 ;
        RECT 43.935 530.735 46.515 531.255 ;
        RECT 46.685 530.905 49.280 531.425 ;
        RECT 49.455 530.735 52.035 531.255 ;
        RECT 52.205 530.905 631.270 531.425 ;
        RECT 54.000 530.735 631.270 530.905 ;
        RECT 42.555 529.965 43.765 530.715 ;
        RECT 43.935 529.965 49.280 530.735 ;
        RECT 49.455 529.965 631.270 530.735 ;
        RECT 42.470 529.795 631.270 529.965 ;
        RECT 42.555 529.045 43.765 529.795 ;
        RECT 42.555 528.505 43.075 529.045 ;
        RECT 43.935 529.025 49.280 529.795 ;
        RECT 49.455 529.025 631.270 529.795 ;
        RECT 43.245 528.335 43.765 528.875 ;
        RECT 43.935 528.505 46.515 529.025 ;
        RECT 46.685 528.335 49.280 528.855 ;
        RECT 49.455 528.505 52.035 529.025 ;
        RECT 54.000 528.855 631.270 529.025 ;
        RECT 52.205 528.335 631.270 528.855 ;
        RECT 42.555 527.245 43.765 528.335 ;
        RECT 43.935 527.245 49.280 528.335 ;
        RECT 49.455 527.245 631.270 528.335 ;
        RECT 42.470 527.075 631.270 527.245 ;
        RECT 42.555 525.985 43.765 527.075 ;
        RECT 43.935 525.985 49.280 527.075 ;
        RECT 49.455 525.985 631.270 527.075 ;
        RECT 42.555 525.275 43.075 525.815 ;
        RECT 43.245 525.445 43.765 525.985 ;
        RECT 43.935 525.295 46.515 525.815 ;
        RECT 46.685 525.465 49.280 525.985 ;
        RECT 49.455 525.295 52.035 525.815 ;
        RECT 52.205 525.465 631.270 525.985 ;
        RECT 54.000 525.295 631.270 525.465 ;
        RECT 42.555 524.525 43.765 525.275 ;
        RECT 43.935 524.525 49.280 525.295 ;
        RECT 49.455 524.525 631.270 525.295 ;
        RECT 42.470 524.355 631.270 524.525 ;
        RECT 42.555 523.605 43.765 524.355 ;
        RECT 42.555 523.065 43.075 523.605 ;
        RECT 43.935 523.585 49.280 524.355 ;
        RECT 49.455 523.585 631.270 524.355 ;
        RECT 43.245 522.895 43.765 523.435 ;
        RECT 43.935 523.065 46.515 523.585 ;
        RECT 46.685 522.895 49.280 523.415 ;
        RECT 49.455 523.065 52.035 523.585 ;
        RECT 54.000 523.415 631.270 523.585 ;
        RECT 52.205 522.895 631.270 523.415 ;
        RECT 42.555 521.805 43.765 522.895 ;
        RECT 43.935 521.805 49.280 522.895 ;
        RECT 49.455 521.805 631.270 522.895 ;
        RECT 42.470 521.635 631.270 521.805 ;
        RECT 42.555 520.545 43.765 521.635 ;
        RECT 43.935 520.545 49.280 521.635 ;
        RECT 49.455 520.545 631.270 521.635 ;
        RECT 42.555 519.835 43.075 520.375 ;
        RECT 43.245 520.005 43.765 520.545 ;
        RECT 43.935 519.855 46.515 520.375 ;
        RECT 46.685 520.025 49.280 520.545 ;
        RECT 49.455 519.855 52.035 520.375 ;
        RECT 52.205 520.025 631.270 520.545 ;
        RECT 54.000 519.855 631.270 520.025 ;
        RECT 42.555 519.085 43.765 519.835 ;
        RECT 43.935 519.085 49.280 519.855 ;
        RECT 49.455 519.085 631.270 519.855 ;
        RECT 42.470 518.915 631.270 519.085 ;
        RECT 42.555 518.165 43.765 518.915 ;
        RECT 42.555 517.625 43.075 518.165 ;
        RECT 43.935 518.145 49.280 518.915 ;
        RECT 49.455 518.145 631.270 518.915 ;
        RECT 43.245 517.455 43.765 517.995 ;
        RECT 43.935 517.625 46.515 518.145 ;
        RECT 46.685 517.455 49.280 517.975 ;
        RECT 49.455 517.625 52.035 518.145 ;
        RECT 54.000 517.975 631.270 518.145 ;
        RECT 52.205 517.455 631.270 517.975 ;
        RECT 42.555 516.365 43.765 517.455 ;
        RECT 43.935 516.365 49.280 517.455 ;
        RECT 49.455 516.365 631.270 517.455 ;
        RECT 42.470 516.195 631.270 516.365 ;
        RECT 42.555 515.105 43.765 516.195 ;
        RECT 43.935 515.105 49.280 516.195 ;
        RECT 49.455 515.105 631.270 516.195 ;
        RECT 42.555 514.395 43.075 514.935 ;
        RECT 43.245 514.565 43.765 515.105 ;
        RECT 43.935 514.415 46.515 514.935 ;
        RECT 46.685 514.585 49.280 515.105 ;
        RECT 49.455 514.415 52.035 514.935 ;
        RECT 52.205 514.585 631.270 515.105 ;
        RECT 54.000 514.415 631.270 514.585 ;
        RECT 42.555 513.645 43.765 514.395 ;
        RECT 43.935 513.645 49.280 514.415 ;
        RECT 49.455 513.645 631.270 514.415 ;
        RECT 42.470 513.475 631.270 513.645 ;
        RECT 42.555 512.725 43.765 513.475 ;
        RECT 42.555 512.185 43.075 512.725 ;
        RECT 43.935 512.705 49.280 513.475 ;
        RECT 49.455 512.705 631.270 513.475 ;
        RECT 43.245 512.015 43.765 512.555 ;
        RECT 43.935 512.185 46.515 512.705 ;
        RECT 46.685 512.015 49.280 512.535 ;
        RECT 49.455 512.185 52.035 512.705 ;
        RECT 54.000 512.535 631.270 512.705 ;
        RECT 52.205 512.015 631.270 512.535 ;
        RECT 42.555 510.925 43.765 512.015 ;
        RECT 43.935 510.925 49.280 512.015 ;
        RECT 49.455 510.925 631.270 512.015 ;
        RECT 42.470 510.755 631.270 510.925 ;
        RECT 42.555 509.665 43.765 510.755 ;
        RECT 43.935 509.665 49.280 510.755 ;
        RECT 49.455 509.665 631.270 510.755 ;
        RECT 42.555 508.955 43.075 509.495 ;
        RECT 43.245 509.125 43.765 509.665 ;
        RECT 43.935 508.975 46.515 509.495 ;
        RECT 46.685 509.145 49.280 509.665 ;
        RECT 49.455 508.975 52.035 509.495 ;
        RECT 52.205 509.145 631.270 509.665 ;
        RECT 54.000 508.975 631.270 509.145 ;
        RECT 42.555 508.205 43.765 508.955 ;
        RECT 43.935 508.205 49.280 508.975 ;
        RECT 49.455 508.205 631.270 508.975 ;
        RECT 42.470 508.035 631.270 508.205 ;
        RECT 42.555 507.285 43.765 508.035 ;
        RECT 42.555 506.745 43.075 507.285 ;
        RECT 43.935 507.265 49.280 508.035 ;
        RECT 49.455 507.265 631.270 508.035 ;
        RECT 43.245 506.575 43.765 507.115 ;
        RECT 43.935 506.745 46.515 507.265 ;
        RECT 46.685 506.575 49.280 507.095 ;
        RECT 49.455 506.745 52.035 507.265 ;
        RECT 54.000 507.095 631.270 507.265 ;
        RECT 52.205 506.575 631.270 507.095 ;
        RECT 42.555 505.485 43.765 506.575 ;
        RECT 43.935 505.485 49.280 506.575 ;
        RECT 49.455 505.485 631.270 506.575 ;
        RECT 42.470 505.315 631.270 505.485 ;
        RECT 42.555 504.225 43.765 505.315 ;
        RECT 43.935 504.225 49.280 505.315 ;
        RECT 49.455 504.225 631.270 505.315 ;
        RECT 42.555 503.515 43.075 504.055 ;
        RECT 43.245 503.685 43.765 504.225 ;
        RECT 43.935 503.535 46.515 504.055 ;
        RECT 46.685 503.705 49.280 504.225 ;
        RECT 49.455 503.535 52.035 504.055 ;
        RECT 52.205 503.705 631.270 504.225 ;
        RECT 54.000 503.535 631.270 503.705 ;
        RECT 42.555 502.765 43.765 503.515 ;
        RECT 43.935 502.765 49.280 503.535 ;
        RECT 49.455 502.765 631.270 503.535 ;
        RECT 42.470 502.595 631.270 502.765 ;
        RECT 42.555 501.845 43.765 502.595 ;
        RECT 42.555 501.305 43.075 501.845 ;
        RECT 43.935 501.825 49.280 502.595 ;
        RECT 49.455 501.825 631.270 502.595 ;
        RECT 43.245 501.135 43.765 501.675 ;
        RECT 43.935 501.305 46.515 501.825 ;
        RECT 46.685 501.135 49.280 501.655 ;
        RECT 49.455 501.305 52.035 501.825 ;
        RECT 54.000 501.655 631.270 501.825 ;
        RECT 52.205 501.135 631.270 501.655 ;
        RECT 42.555 500.045 43.765 501.135 ;
        RECT 43.935 500.045 49.280 501.135 ;
        RECT 49.455 500.045 631.270 501.135 ;
        RECT 42.470 499.875 631.270 500.045 ;
        RECT 42.555 498.785 43.765 499.875 ;
        RECT 43.935 498.785 49.280 499.875 ;
        RECT 49.455 498.785 631.270 499.875 ;
        RECT 42.555 498.075 43.075 498.615 ;
        RECT 43.245 498.245 43.765 498.785 ;
        RECT 43.935 498.095 46.515 498.615 ;
        RECT 46.685 498.265 49.280 498.785 ;
        RECT 49.455 498.095 52.035 498.615 ;
        RECT 52.205 498.265 631.270 498.785 ;
        RECT 54.000 498.095 631.270 498.265 ;
        RECT 42.555 497.325 43.765 498.075 ;
        RECT 43.935 497.325 49.280 498.095 ;
        RECT 49.455 497.325 631.270 498.095 ;
        RECT 42.470 497.155 631.270 497.325 ;
        RECT 42.555 496.405 43.765 497.155 ;
        RECT 42.555 495.865 43.075 496.405 ;
        RECT 43.935 496.385 49.280 497.155 ;
        RECT 49.455 496.385 631.270 497.155 ;
        RECT 43.245 495.695 43.765 496.235 ;
        RECT 43.935 495.865 46.515 496.385 ;
        RECT 46.685 495.695 49.280 496.215 ;
        RECT 49.455 495.865 52.035 496.385 ;
        RECT 54.000 496.215 631.270 496.385 ;
        RECT 52.205 495.695 631.270 496.215 ;
        RECT 42.555 494.605 43.765 495.695 ;
        RECT 43.935 494.605 49.280 495.695 ;
        RECT 49.455 494.605 631.270 495.695 ;
        RECT 42.470 494.435 631.270 494.605 ;
        RECT 42.555 493.345 43.765 494.435 ;
        RECT 43.935 493.345 49.280 494.435 ;
        RECT 49.455 493.345 631.270 494.435 ;
        RECT 42.555 492.635 43.075 493.175 ;
        RECT 43.245 492.805 43.765 493.345 ;
        RECT 43.935 492.655 46.515 493.175 ;
        RECT 46.685 492.825 49.280 493.345 ;
        RECT 49.455 492.655 52.035 493.175 ;
        RECT 52.205 492.825 631.270 493.345 ;
        RECT 54.000 492.655 631.270 492.825 ;
        RECT 42.555 491.885 43.765 492.635 ;
        RECT 43.935 491.885 49.280 492.655 ;
        RECT 49.455 491.885 631.270 492.655 ;
        RECT 42.470 491.715 631.270 491.885 ;
        RECT 42.555 490.965 43.765 491.715 ;
        RECT 42.555 490.425 43.075 490.965 ;
        RECT 43.935 490.945 49.280 491.715 ;
        RECT 49.455 490.945 631.270 491.715 ;
        RECT 43.245 490.255 43.765 490.795 ;
        RECT 43.935 490.425 46.515 490.945 ;
        RECT 46.685 490.255 49.280 490.775 ;
        RECT 49.455 490.425 52.035 490.945 ;
        RECT 54.000 490.775 631.270 490.945 ;
        RECT 52.205 490.255 631.270 490.775 ;
        RECT 42.555 489.165 43.765 490.255 ;
        RECT 43.935 489.165 49.280 490.255 ;
        RECT 49.455 489.165 631.270 490.255 ;
        RECT 42.470 488.995 631.270 489.165 ;
        RECT 42.555 487.905 43.765 488.995 ;
        RECT 43.935 487.905 49.280 488.995 ;
        RECT 49.455 487.905 631.270 488.995 ;
        RECT 42.555 487.195 43.075 487.735 ;
        RECT 43.245 487.365 43.765 487.905 ;
        RECT 43.935 487.215 46.515 487.735 ;
        RECT 46.685 487.385 49.280 487.905 ;
        RECT 49.455 487.215 52.035 487.735 ;
        RECT 52.205 487.385 631.270 487.905 ;
        RECT 54.000 487.215 631.270 487.385 ;
        RECT 42.555 486.445 43.765 487.195 ;
        RECT 43.935 486.445 49.280 487.215 ;
        RECT 49.455 486.445 631.270 487.215 ;
        RECT 42.470 486.275 631.270 486.445 ;
        RECT 42.555 485.525 43.765 486.275 ;
        RECT 42.555 484.985 43.075 485.525 ;
        RECT 43.935 485.505 49.280 486.275 ;
        RECT 49.455 485.505 631.270 486.275 ;
        RECT 43.245 484.815 43.765 485.355 ;
        RECT 43.935 484.985 46.515 485.505 ;
        RECT 46.685 484.815 49.280 485.335 ;
        RECT 49.455 484.985 52.035 485.505 ;
        RECT 54.000 485.335 631.270 485.505 ;
        RECT 52.205 484.815 631.270 485.335 ;
        RECT 42.555 483.725 43.765 484.815 ;
        RECT 43.935 483.725 49.280 484.815 ;
        RECT 49.455 483.725 631.270 484.815 ;
        RECT 42.470 483.555 631.270 483.725 ;
        RECT 42.555 482.465 43.765 483.555 ;
        RECT 43.935 482.465 49.280 483.555 ;
        RECT 49.455 482.465 631.270 483.555 ;
        RECT 42.555 481.755 43.075 482.295 ;
        RECT 43.245 481.925 43.765 482.465 ;
        RECT 43.935 481.775 46.515 482.295 ;
        RECT 46.685 481.945 49.280 482.465 ;
        RECT 49.455 481.775 52.035 482.295 ;
        RECT 52.205 481.945 631.270 482.465 ;
        RECT 54.000 481.775 631.270 481.945 ;
        RECT 42.555 481.005 43.765 481.755 ;
        RECT 43.935 481.005 49.280 481.775 ;
        RECT 49.455 481.005 631.270 481.775 ;
        RECT 42.470 480.835 631.270 481.005 ;
        RECT 42.555 480.085 43.765 480.835 ;
        RECT 42.555 479.545 43.075 480.085 ;
        RECT 43.935 480.065 49.280 480.835 ;
        RECT 49.455 480.065 631.270 480.835 ;
        RECT 43.245 479.375 43.765 479.915 ;
        RECT 43.935 479.545 46.515 480.065 ;
        RECT 46.685 479.375 49.280 479.895 ;
        RECT 49.455 479.545 52.035 480.065 ;
        RECT 54.000 479.895 631.270 480.065 ;
        RECT 52.205 479.375 631.270 479.895 ;
        RECT 42.555 478.285 43.765 479.375 ;
        RECT 43.935 478.285 49.280 479.375 ;
        RECT 49.455 478.285 631.270 479.375 ;
        RECT 42.470 478.115 631.270 478.285 ;
        RECT 42.555 477.025 43.765 478.115 ;
        RECT 43.935 477.025 49.280 478.115 ;
        RECT 49.455 477.025 631.270 478.115 ;
        RECT 42.555 476.315 43.075 476.855 ;
        RECT 43.245 476.485 43.765 477.025 ;
        RECT 43.935 476.335 46.515 476.855 ;
        RECT 46.685 476.505 49.280 477.025 ;
        RECT 49.455 476.335 52.035 476.855 ;
        RECT 52.205 476.505 631.270 477.025 ;
        RECT 54.000 476.335 631.270 476.505 ;
        RECT 42.555 475.565 43.765 476.315 ;
        RECT 43.935 475.565 49.280 476.335 ;
        RECT 49.455 475.565 631.270 476.335 ;
        RECT 42.470 475.395 631.270 475.565 ;
        RECT 42.555 474.645 43.765 475.395 ;
        RECT 42.555 474.105 43.075 474.645 ;
        RECT 43.935 474.625 49.280 475.395 ;
        RECT 49.455 474.625 631.270 475.395 ;
        RECT 43.245 473.935 43.765 474.475 ;
        RECT 43.935 474.105 46.515 474.625 ;
        RECT 46.685 473.935 49.280 474.455 ;
        RECT 49.455 474.105 52.035 474.625 ;
        RECT 54.000 474.455 631.270 474.625 ;
        RECT 52.205 473.935 631.270 474.455 ;
        RECT 42.555 472.845 43.765 473.935 ;
        RECT 43.935 472.845 49.280 473.935 ;
        RECT 49.455 472.845 631.270 473.935 ;
        RECT 42.470 472.675 631.270 472.845 ;
        RECT 42.555 471.585 43.765 472.675 ;
        RECT 43.935 471.585 49.280 472.675 ;
        RECT 49.455 471.585 631.270 472.675 ;
        RECT 42.555 470.875 43.075 471.415 ;
        RECT 43.245 471.045 43.765 471.585 ;
        RECT 43.935 470.895 46.515 471.415 ;
        RECT 46.685 471.065 49.280 471.585 ;
        RECT 49.455 470.895 52.035 471.415 ;
        RECT 52.205 471.065 631.270 471.585 ;
        RECT 54.000 470.895 631.270 471.065 ;
        RECT 42.555 470.125 43.765 470.875 ;
        RECT 43.935 470.125 49.280 470.895 ;
        RECT 49.455 470.125 631.270 470.895 ;
        RECT 42.470 469.955 631.270 470.125 ;
        RECT 42.555 469.205 43.765 469.955 ;
        RECT 42.555 468.665 43.075 469.205 ;
        RECT 43.935 469.185 49.280 469.955 ;
        RECT 49.455 469.185 631.270 469.955 ;
        RECT 43.245 468.495 43.765 469.035 ;
        RECT 43.935 468.665 46.515 469.185 ;
        RECT 46.685 468.495 49.280 469.015 ;
        RECT 49.455 468.665 52.035 469.185 ;
        RECT 54.000 469.015 631.270 469.185 ;
        RECT 52.205 468.495 631.270 469.015 ;
        RECT 42.555 467.405 43.765 468.495 ;
        RECT 43.935 467.405 49.280 468.495 ;
        RECT 49.455 467.405 631.270 468.495 ;
        RECT 42.470 467.235 631.270 467.405 ;
        RECT 42.555 466.145 43.765 467.235 ;
        RECT 43.935 466.145 49.280 467.235 ;
        RECT 49.455 466.145 631.270 467.235 ;
        RECT 42.555 465.435 43.075 465.975 ;
        RECT 43.245 465.605 43.765 466.145 ;
        RECT 43.935 465.455 46.515 465.975 ;
        RECT 46.685 465.625 49.280 466.145 ;
        RECT 49.455 465.455 52.035 465.975 ;
        RECT 52.205 465.625 631.270 466.145 ;
        RECT 54.000 465.455 631.270 465.625 ;
        RECT 42.555 464.685 43.765 465.435 ;
        RECT 43.935 464.685 49.280 465.455 ;
        RECT 49.455 464.685 631.270 465.455 ;
        RECT 42.470 464.515 631.270 464.685 ;
        RECT 42.555 463.765 43.765 464.515 ;
        RECT 42.555 463.225 43.075 463.765 ;
        RECT 43.935 463.745 49.280 464.515 ;
        RECT 49.455 463.745 631.270 464.515 ;
        RECT 43.245 463.055 43.765 463.595 ;
        RECT 43.935 463.225 46.515 463.745 ;
        RECT 46.685 463.055 49.280 463.575 ;
        RECT 49.455 463.225 52.035 463.745 ;
        RECT 54.000 463.575 631.270 463.745 ;
        RECT 52.205 463.055 631.270 463.575 ;
        RECT 42.555 461.965 43.765 463.055 ;
        RECT 43.935 461.965 49.280 463.055 ;
        RECT 49.455 461.965 631.270 463.055 ;
        RECT 42.470 461.795 631.270 461.965 ;
        RECT 42.555 460.705 43.765 461.795 ;
        RECT 43.935 460.705 49.280 461.795 ;
        RECT 49.455 460.705 631.270 461.795 ;
        RECT 42.555 459.995 43.075 460.535 ;
        RECT 43.245 460.165 43.765 460.705 ;
        RECT 43.935 460.015 46.515 460.535 ;
        RECT 46.685 460.185 49.280 460.705 ;
        RECT 49.455 460.015 52.035 460.535 ;
        RECT 52.205 460.185 631.270 460.705 ;
        RECT 54.000 460.015 631.270 460.185 ;
        RECT 42.555 459.245 43.765 459.995 ;
        RECT 43.935 459.245 49.280 460.015 ;
        RECT 49.455 459.245 631.270 460.015 ;
        RECT 42.470 459.075 631.270 459.245 ;
        RECT 42.555 458.325 43.765 459.075 ;
        RECT 42.555 457.785 43.075 458.325 ;
        RECT 43.935 458.305 49.280 459.075 ;
        RECT 49.455 458.305 631.270 459.075 ;
        RECT 43.245 457.615 43.765 458.155 ;
        RECT 43.935 457.785 46.515 458.305 ;
        RECT 46.685 457.615 49.280 458.135 ;
        RECT 49.455 457.785 52.035 458.305 ;
        RECT 54.000 458.135 631.270 458.305 ;
        RECT 52.205 457.615 631.270 458.135 ;
        RECT 42.555 456.525 43.765 457.615 ;
        RECT 43.935 456.525 49.280 457.615 ;
        RECT 49.455 456.525 631.270 457.615 ;
        RECT 42.470 456.355 631.270 456.525 ;
        RECT 42.555 455.265 43.765 456.355 ;
        RECT 43.935 455.265 49.280 456.355 ;
        RECT 49.455 455.265 631.270 456.355 ;
        RECT 42.555 454.555 43.075 455.095 ;
        RECT 43.245 454.725 43.765 455.265 ;
        RECT 43.935 454.575 46.515 455.095 ;
        RECT 46.685 454.745 49.280 455.265 ;
        RECT 49.455 454.575 52.035 455.095 ;
        RECT 52.205 454.745 631.270 455.265 ;
        RECT 54.000 454.575 631.270 454.745 ;
        RECT 42.555 453.805 43.765 454.555 ;
        RECT 43.935 453.805 49.280 454.575 ;
        RECT 49.455 453.805 631.270 454.575 ;
        RECT 42.470 453.635 631.270 453.805 ;
        RECT 42.555 452.885 43.765 453.635 ;
        RECT 42.555 452.345 43.075 452.885 ;
        RECT 43.935 452.865 49.280 453.635 ;
        RECT 49.455 452.865 631.270 453.635 ;
        RECT 43.245 452.175 43.765 452.715 ;
        RECT 43.935 452.345 46.515 452.865 ;
        RECT 46.685 452.175 49.280 452.695 ;
        RECT 49.455 452.345 52.035 452.865 ;
        RECT 54.000 452.695 631.270 452.865 ;
        RECT 52.205 452.175 631.270 452.695 ;
        RECT 42.555 451.085 43.765 452.175 ;
        RECT 43.935 451.085 49.280 452.175 ;
        RECT 49.455 451.085 631.270 452.175 ;
        RECT 42.470 450.915 631.270 451.085 ;
        RECT 42.555 449.825 43.765 450.915 ;
        RECT 43.935 449.825 49.280 450.915 ;
        RECT 49.455 449.825 631.270 450.915 ;
        RECT 42.555 449.115 43.075 449.655 ;
        RECT 43.245 449.285 43.765 449.825 ;
        RECT 43.935 449.135 46.515 449.655 ;
        RECT 46.685 449.305 49.280 449.825 ;
        RECT 49.455 449.135 52.035 449.655 ;
        RECT 52.205 449.305 631.270 449.825 ;
        RECT 54.000 449.135 631.270 449.305 ;
        RECT 42.555 448.365 43.765 449.115 ;
        RECT 43.935 448.365 49.280 449.135 ;
        RECT 49.455 448.365 631.270 449.135 ;
        RECT 42.470 448.195 631.270 448.365 ;
        RECT 42.555 447.445 43.765 448.195 ;
        RECT 42.555 446.905 43.075 447.445 ;
        RECT 43.935 447.425 49.280 448.195 ;
        RECT 49.455 447.425 631.270 448.195 ;
        RECT 43.245 446.735 43.765 447.275 ;
        RECT 43.935 446.905 46.515 447.425 ;
        RECT 46.685 446.735 49.280 447.255 ;
        RECT 49.455 446.905 52.035 447.425 ;
        RECT 54.000 447.255 631.270 447.425 ;
        RECT 52.205 446.735 631.270 447.255 ;
        RECT 42.555 445.645 43.765 446.735 ;
        RECT 43.935 445.645 49.280 446.735 ;
        RECT 49.455 445.645 631.270 446.735 ;
        RECT 42.470 445.475 631.270 445.645 ;
        RECT 42.555 444.385 43.765 445.475 ;
        RECT 43.935 444.385 49.280 445.475 ;
        RECT 49.455 444.385 631.270 445.475 ;
        RECT 42.555 443.675 43.075 444.215 ;
        RECT 43.245 443.845 43.765 444.385 ;
        RECT 43.935 443.695 46.515 444.215 ;
        RECT 46.685 443.865 49.280 444.385 ;
        RECT 49.455 443.695 52.035 444.215 ;
        RECT 52.205 443.865 631.270 444.385 ;
        RECT 54.000 443.695 631.270 443.865 ;
        RECT 42.555 442.925 43.765 443.675 ;
        RECT 43.935 442.925 49.280 443.695 ;
        RECT 49.455 442.925 631.270 443.695 ;
        RECT 42.470 442.755 631.270 442.925 ;
        RECT 42.555 442.005 43.765 442.755 ;
        RECT 42.555 441.465 43.075 442.005 ;
        RECT 43.935 441.985 49.280 442.755 ;
        RECT 49.455 441.985 631.270 442.755 ;
        RECT 43.245 441.295 43.765 441.835 ;
        RECT 43.935 441.465 46.515 441.985 ;
        RECT 46.685 441.295 49.280 441.815 ;
        RECT 49.455 441.465 52.035 441.985 ;
        RECT 54.000 441.815 631.270 441.985 ;
        RECT 52.205 441.295 631.270 441.815 ;
        RECT 42.555 440.205 43.765 441.295 ;
        RECT 43.935 440.205 49.280 441.295 ;
        RECT 49.455 440.205 631.270 441.295 ;
        RECT 42.470 440.035 631.270 440.205 ;
        RECT 42.555 438.945 43.765 440.035 ;
        RECT 43.935 438.945 49.280 440.035 ;
        RECT 49.455 438.945 631.270 440.035 ;
        RECT 42.555 438.235 43.075 438.775 ;
        RECT 43.245 438.405 43.765 438.945 ;
        RECT 43.935 438.255 46.515 438.775 ;
        RECT 46.685 438.425 49.280 438.945 ;
        RECT 49.455 438.255 52.035 438.775 ;
        RECT 52.205 438.425 631.270 438.945 ;
        RECT 54.000 438.255 631.270 438.425 ;
        RECT 42.555 437.485 43.765 438.235 ;
        RECT 43.935 437.485 49.280 438.255 ;
        RECT 49.455 437.485 631.270 438.255 ;
        RECT 42.470 437.315 631.270 437.485 ;
        RECT 42.555 436.565 43.765 437.315 ;
        RECT 42.555 436.025 43.075 436.565 ;
        RECT 43.935 436.545 49.280 437.315 ;
        RECT 49.455 436.545 631.270 437.315 ;
        RECT 43.245 435.855 43.765 436.395 ;
        RECT 43.935 436.025 46.515 436.545 ;
        RECT 46.685 435.855 49.280 436.375 ;
        RECT 49.455 436.025 52.035 436.545 ;
        RECT 54.000 436.375 631.270 436.545 ;
        RECT 52.205 435.855 631.270 436.375 ;
        RECT 42.555 434.765 43.765 435.855 ;
        RECT 43.935 434.765 49.280 435.855 ;
        RECT 49.455 434.765 631.270 435.855 ;
        RECT 42.470 434.595 631.270 434.765 ;
        RECT 42.555 433.505 43.765 434.595 ;
        RECT 43.935 433.505 49.280 434.595 ;
        RECT 49.455 433.505 631.270 434.595 ;
        RECT 42.555 432.795 43.075 433.335 ;
        RECT 43.245 432.965 43.765 433.505 ;
        RECT 43.935 432.815 46.515 433.335 ;
        RECT 46.685 432.985 49.280 433.505 ;
        RECT 49.455 432.815 52.035 433.335 ;
        RECT 52.205 432.985 631.270 433.505 ;
        RECT 54.000 432.815 631.270 432.985 ;
        RECT 42.555 432.045 43.765 432.795 ;
        RECT 43.935 432.045 49.280 432.815 ;
        RECT 49.455 432.045 631.270 432.815 ;
        RECT 42.470 431.875 631.270 432.045 ;
        RECT 42.555 431.125 43.765 431.875 ;
        RECT 42.555 430.585 43.075 431.125 ;
        RECT 43.935 431.105 49.280 431.875 ;
        RECT 49.455 431.105 631.270 431.875 ;
        RECT 43.245 430.415 43.765 430.955 ;
        RECT 43.935 430.585 46.515 431.105 ;
        RECT 46.685 430.415 49.280 430.935 ;
        RECT 49.455 430.585 52.035 431.105 ;
        RECT 54.000 430.935 631.270 431.105 ;
        RECT 52.205 430.415 631.270 430.935 ;
        RECT 42.555 429.325 43.765 430.415 ;
        RECT 43.935 429.325 49.280 430.415 ;
        RECT 49.455 429.325 631.270 430.415 ;
        RECT 42.470 429.155 631.270 429.325 ;
        RECT 42.555 428.065 43.765 429.155 ;
        RECT 43.935 428.065 49.280 429.155 ;
        RECT 49.455 428.065 631.270 429.155 ;
        RECT 42.555 427.355 43.075 427.895 ;
        RECT 43.245 427.525 43.765 428.065 ;
        RECT 43.935 427.375 46.515 427.895 ;
        RECT 46.685 427.545 49.280 428.065 ;
        RECT 49.455 427.375 52.035 427.895 ;
        RECT 52.205 427.545 631.270 428.065 ;
        RECT 54.000 427.375 631.270 427.545 ;
        RECT 42.555 426.605 43.765 427.355 ;
        RECT 43.935 426.605 49.280 427.375 ;
        RECT 49.455 426.605 631.270 427.375 ;
        RECT 42.470 426.435 631.270 426.605 ;
        RECT 42.555 425.685 43.765 426.435 ;
        RECT 42.555 425.145 43.075 425.685 ;
        RECT 43.935 425.665 49.280 426.435 ;
        RECT 49.455 425.665 631.270 426.435 ;
        RECT 43.245 424.975 43.765 425.515 ;
        RECT 43.935 425.145 46.515 425.665 ;
        RECT 46.685 424.975 49.280 425.495 ;
        RECT 49.455 425.145 52.035 425.665 ;
        RECT 54.000 425.495 631.270 425.665 ;
        RECT 52.205 424.975 631.270 425.495 ;
        RECT 42.555 423.885 43.765 424.975 ;
        RECT 43.935 423.885 49.280 424.975 ;
        RECT 49.455 423.885 631.270 424.975 ;
        RECT 42.470 423.715 631.270 423.885 ;
        RECT 42.555 422.625 43.765 423.715 ;
        RECT 43.935 422.625 49.280 423.715 ;
        RECT 49.455 422.625 631.270 423.715 ;
        RECT 42.555 421.915 43.075 422.455 ;
        RECT 43.245 422.085 43.765 422.625 ;
        RECT 43.935 421.935 46.515 422.455 ;
        RECT 46.685 422.105 49.280 422.625 ;
        RECT 49.455 421.935 52.035 422.455 ;
        RECT 52.205 422.105 631.270 422.625 ;
        RECT 54.000 421.935 631.270 422.105 ;
        RECT 42.555 421.165 43.765 421.915 ;
        RECT 43.935 421.165 49.280 421.935 ;
        RECT 49.455 421.165 631.270 421.935 ;
        RECT 42.470 420.995 631.270 421.165 ;
        RECT 42.555 420.245 43.765 420.995 ;
        RECT 42.555 419.705 43.075 420.245 ;
        RECT 43.935 420.225 49.280 420.995 ;
        RECT 49.455 420.225 631.270 420.995 ;
        RECT 43.245 419.535 43.765 420.075 ;
        RECT 43.935 419.705 46.515 420.225 ;
        RECT 46.685 419.535 49.280 420.055 ;
        RECT 49.455 419.705 52.035 420.225 ;
        RECT 54.000 420.055 631.270 420.225 ;
        RECT 52.205 419.535 631.270 420.055 ;
        RECT 42.555 418.445 43.765 419.535 ;
        RECT 43.935 418.445 49.280 419.535 ;
        RECT 49.455 418.445 631.270 419.535 ;
        RECT 42.470 418.275 631.270 418.445 ;
        RECT 42.555 417.185 43.765 418.275 ;
        RECT 43.935 417.185 49.280 418.275 ;
        RECT 49.455 417.185 631.270 418.275 ;
        RECT 42.555 416.475 43.075 417.015 ;
        RECT 43.245 416.645 43.765 417.185 ;
        RECT 43.935 416.495 46.515 417.015 ;
        RECT 46.685 416.665 49.280 417.185 ;
        RECT 49.455 416.495 52.035 417.015 ;
        RECT 52.205 416.665 631.270 417.185 ;
        RECT 54.000 416.495 631.270 416.665 ;
        RECT 42.555 415.725 43.765 416.475 ;
        RECT 43.935 415.725 49.280 416.495 ;
        RECT 49.455 415.725 631.270 416.495 ;
        RECT 42.470 415.555 631.270 415.725 ;
        RECT 42.555 414.805 43.765 415.555 ;
        RECT 42.555 414.265 43.075 414.805 ;
        RECT 43.935 414.785 49.280 415.555 ;
        RECT 49.455 414.785 631.270 415.555 ;
        RECT 43.245 414.095 43.765 414.635 ;
        RECT 43.935 414.265 46.515 414.785 ;
        RECT 46.685 414.095 49.280 414.615 ;
        RECT 49.455 414.265 52.035 414.785 ;
        RECT 54.000 414.615 631.270 414.785 ;
        RECT 52.205 414.095 631.270 414.615 ;
        RECT 42.555 413.005 43.765 414.095 ;
        RECT 43.935 413.005 49.280 414.095 ;
        RECT 49.455 413.005 631.270 414.095 ;
        RECT 42.470 412.835 631.270 413.005 ;
        RECT 42.555 411.745 43.765 412.835 ;
        RECT 43.935 411.745 49.280 412.835 ;
        RECT 49.455 411.745 631.270 412.835 ;
        RECT 42.555 411.035 43.075 411.575 ;
        RECT 43.245 411.205 43.765 411.745 ;
        RECT 43.935 411.055 46.515 411.575 ;
        RECT 46.685 411.225 49.280 411.745 ;
        RECT 49.455 411.055 52.035 411.575 ;
        RECT 52.205 411.225 631.270 411.745 ;
        RECT 54.000 411.055 631.270 411.225 ;
        RECT 42.555 410.285 43.765 411.035 ;
        RECT 43.935 410.285 49.280 411.055 ;
        RECT 49.455 410.285 631.270 411.055 ;
        RECT 42.470 410.115 631.270 410.285 ;
        RECT 42.555 409.365 43.765 410.115 ;
        RECT 42.555 408.825 43.075 409.365 ;
        RECT 43.935 409.345 49.280 410.115 ;
        RECT 49.455 409.345 631.270 410.115 ;
        RECT 43.245 408.655 43.765 409.195 ;
        RECT 43.935 408.825 46.515 409.345 ;
        RECT 46.685 408.655 49.280 409.175 ;
        RECT 49.455 408.825 52.035 409.345 ;
        RECT 54.000 409.175 631.270 409.345 ;
        RECT 52.205 408.655 631.270 409.175 ;
        RECT 42.555 407.565 43.765 408.655 ;
        RECT 43.935 407.565 49.280 408.655 ;
        RECT 49.455 407.565 631.270 408.655 ;
        RECT 42.470 407.395 631.270 407.565 ;
        RECT 42.555 406.305 43.765 407.395 ;
        RECT 43.935 406.305 49.280 407.395 ;
        RECT 49.455 406.305 631.270 407.395 ;
        RECT 42.555 405.595 43.075 406.135 ;
        RECT 43.245 405.765 43.765 406.305 ;
        RECT 43.935 405.615 46.515 406.135 ;
        RECT 46.685 405.785 49.280 406.305 ;
        RECT 49.455 405.615 52.035 406.135 ;
        RECT 52.205 405.785 631.270 406.305 ;
        RECT 54.000 405.615 631.270 405.785 ;
        RECT 42.555 404.845 43.765 405.595 ;
        RECT 43.935 404.845 49.280 405.615 ;
        RECT 49.455 404.845 631.270 405.615 ;
        RECT 42.470 404.675 631.270 404.845 ;
        RECT 42.555 403.925 43.765 404.675 ;
        RECT 42.555 403.385 43.075 403.925 ;
        RECT 43.935 403.905 49.280 404.675 ;
        RECT 49.455 403.905 631.270 404.675 ;
        RECT 43.245 403.215 43.765 403.755 ;
        RECT 43.935 403.385 46.515 403.905 ;
        RECT 46.685 403.215 49.280 403.735 ;
        RECT 49.455 403.385 52.035 403.905 ;
        RECT 54.000 403.735 631.270 403.905 ;
        RECT 52.205 403.215 631.270 403.735 ;
        RECT 42.555 402.125 43.765 403.215 ;
        RECT 43.935 402.125 49.280 403.215 ;
        RECT 49.455 402.125 631.270 403.215 ;
        RECT 42.470 401.955 631.270 402.125 ;
        RECT 42.555 400.865 43.765 401.955 ;
        RECT 43.935 400.865 49.280 401.955 ;
        RECT 49.455 400.865 631.270 401.955 ;
        RECT 42.555 400.155 43.075 400.695 ;
        RECT 43.245 400.325 43.765 400.865 ;
        RECT 43.935 400.175 46.515 400.695 ;
        RECT 46.685 400.345 49.280 400.865 ;
        RECT 49.455 400.175 52.035 400.695 ;
        RECT 52.205 400.345 631.270 400.865 ;
        RECT 54.000 400.175 631.270 400.345 ;
        RECT 42.555 399.405 43.765 400.155 ;
        RECT 43.935 399.405 49.280 400.175 ;
        RECT 49.455 399.405 631.270 400.175 ;
        RECT 42.470 399.235 631.270 399.405 ;
        RECT 42.555 398.485 43.765 399.235 ;
        RECT 42.555 397.945 43.075 398.485 ;
        RECT 43.935 398.465 49.280 399.235 ;
        RECT 49.455 398.465 631.270 399.235 ;
        RECT 43.245 397.775 43.765 398.315 ;
        RECT 43.935 397.945 46.515 398.465 ;
        RECT 46.685 397.775 49.280 398.295 ;
        RECT 49.455 397.945 52.035 398.465 ;
        RECT 54.000 398.295 631.270 398.465 ;
        RECT 52.205 397.775 631.270 398.295 ;
        RECT 42.555 396.685 43.765 397.775 ;
        RECT 43.935 396.685 49.280 397.775 ;
        RECT 49.455 396.685 631.270 397.775 ;
        RECT 42.470 396.515 631.270 396.685 ;
        RECT 42.555 395.425 43.765 396.515 ;
        RECT 43.935 395.425 49.280 396.515 ;
        RECT 49.455 395.425 631.270 396.515 ;
        RECT 42.555 394.715 43.075 395.255 ;
        RECT 43.245 394.885 43.765 395.425 ;
        RECT 43.935 394.735 46.515 395.255 ;
        RECT 46.685 394.905 49.280 395.425 ;
        RECT 49.455 394.735 52.035 395.255 ;
        RECT 52.205 394.905 631.270 395.425 ;
        RECT 54.000 394.735 631.270 394.905 ;
        RECT 42.555 393.965 43.765 394.715 ;
        RECT 43.935 393.965 49.280 394.735 ;
        RECT 49.455 393.965 631.270 394.735 ;
        RECT 42.470 393.795 631.270 393.965 ;
        RECT 42.555 393.045 43.765 393.795 ;
        RECT 42.555 392.505 43.075 393.045 ;
        RECT 43.935 393.025 49.280 393.795 ;
        RECT 49.455 393.025 631.270 393.795 ;
        RECT 43.245 392.335 43.765 392.875 ;
        RECT 43.935 392.505 46.515 393.025 ;
        RECT 46.685 392.335 49.280 392.855 ;
        RECT 49.455 392.505 52.035 393.025 ;
        RECT 54.000 392.855 631.270 393.025 ;
        RECT 52.205 392.335 631.270 392.855 ;
        RECT 42.555 391.245 43.765 392.335 ;
        RECT 43.935 391.245 49.280 392.335 ;
        RECT 49.455 391.245 631.270 392.335 ;
        RECT 42.470 391.075 631.270 391.245 ;
        RECT 42.555 389.985 43.765 391.075 ;
        RECT 43.935 389.985 49.280 391.075 ;
        RECT 49.455 389.985 631.270 391.075 ;
        RECT 42.555 389.275 43.075 389.815 ;
        RECT 43.245 389.445 43.765 389.985 ;
        RECT 43.935 389.295 46.515 389.815 ;
        RECT 46.685 389.465 49.280 389.985 ;
        RECT 49.455 389.295 52.035 389.815 ;
        RECT 52.205 389.465 631.270 389.985 ;
        RECT 54.000 389.295 631.270 389.465 ;
        RECT 42.555 388.525 43.765 389.275 ;
        RECT 43.935 388.525 49.280 389.295 ;
        RECT 49.455 388.525 631.270 389.295 ;
        RECT 42.470 388.355 631.270 388.525 ;
        RECT 42.555 387.605 43.765 388.355 ;
        RECT 42.555 387.065 43.075 387.605 ;
        RECT 43.935 387.585 49.280 388.355 ;
        RECT 49.455 387.585 631.270 388.355 ;
        RECT 43.245 386.895 43.765 387.435 ;
        RECT 43.935 387.065 46.515 387.585 ;
        RECT 46.685 386.895 49.280 387.415 ;
        RECT 49.455 387.065 52.035 387.585 ;
        RECT 54.000 387.415 631.270 387.585 ;
        RECT 52.205 386.895 631.270 387.415 ;
        RECT 42.555 385.805 43.765 386.895 ;
        RECT 43.935 385.805 49.280 386.895 ;
        RECT 49.455 385.805 631.270 386.895 ;
        RECT 42.470 385.635 631.270 385.805 ;
        RECT 42.555 384.545 43.765 385.635 ;
        RECT 43.935 384.545 49.280 385.635 ;
        RECT 49.455 384.545 631.270 385.635 ;
        RECT 42.555 383.835 43.075 384.375 ;
        RECT 43.245 384.005 43.765 384.545 ;
        RECT 43.935 383.855 46.515 384.375 ;
        RECT 46.685 384.025 49.280 384.545 ;
        RECT 49.455 383.855 52.035 384.375 ;
        RECT 52.205 384.025 631.270 384.545 ;
        RECT 54.000 383.855 631.270 384.025 ;
        RECT 42.555 383.085 43.765 383.835 ;
        RECT 43.935 383.085 49.280 383.855 ;
        RECT 49.455 383.085 631.270 383.855 ;
        RECT 42.470 382.915 631.270 383.085 ;
        RECT 42.555 382.165 43.765 382.915 ;
        RECT 42.555 381.625 43.075 382.165 ;
        RECT 43.935 382.145 49.280 382.915 ;
        RECT 49.455 382.145 631.270 382.915 ;
        RECT 43.245 381.455 43.765 381.995 ;
        RECT 43.935 381.625 46.515 382.145 ;
        RECT 46.685 381.455 49.280 381.975 ;
        RECT 49.455 381.625 52.035 382.145 ;
        RECT 54.000 381.975 631.270 382.145 ;
        RECT 52.205 381.455 631.270 381.975 ;
        RECT 42.555 380.365 43.765 381.455 ;
        RECT 43.935 380.365 49.280 381.455 ;
        RECT 49.455 380.365 631.270 381.455 ;
        RECT 42.470 380.195 631.270 380.365 ;
        RECT 42.555 379.105 43.765 380.195 ;
        RECT 43.935 379.105 49.280 380.195 ;
        RECT 49.455 379.105 631.270 380.195 ;
        RECT 42.555 378.395 43.075 378.935 ;
        RECT 43.245 378.565 43.765 379.105 ;
        RECT 43.935 378.415 46.515 378.935 ;
        RECT 46.685 378.585 49.280 379.105 ;
        RECT 49.455 378.415 52.035 378.935 ;
        RECT 52.205 378.585 631.270 379.105 ;
        RECT 54.000 378.415 631.270 378.585 ;
        RECT 42.555 377.645 43.765 378.395 ;
        RECT 43.935 377.645 49.280 378.415 ;
        RECT 49.455 377.645 631.270 378.415 ;
        RECT 42.470 377.475 631.270 377.645 ;
        RECT 42.555 376.725 43.765 377.475 ;
        RECT 42.555 376.185 43.075 376.725 ;
        RECT 43.935 376.705 49.280 377.475 ;
        RECT 49.455 376.705 631.270 377.475 ;
        RECT 43.245 376.015 43.765 376.555 ;
        RECT 43.935 376.185 46.515 376.705 ;
        RECT 46.685 376.015 49.280 376.535 ;
        RECT 49.455 376.185 52.035 376.705 ;
        RECT 54.000 376.535 631.270 376.705 ;
        RECT 52.205 376.015 631.270 376.535 ;
        RECT 42.555 374.925 43.765 376.015 ;
        RECT 43.935 374.925 49.280 376.015 ;
        RECT 49.455 374.925 631.270 376.015 ;
        RECT 42.470 374.755 631.270 374.925 ;
        RECT 42.555 373.665 43.765 374.755 ;
        RECT 43.935 373.665 49.280 374.755 ;
        RECT 49.455 373.665 631.270 374.755 ;
        RECT 42.555 372.955 43.075 373.495 ;
        RECT 43.245 373.125 43.765 373.665 ;
        RECT 43.935 372.975 46.515 373.495 ;
        RECT 46.685 373.145 49.280 373.665 ;
        RECT 49.455 372.975 52.035 373.495 ;
        RECT 52.205 373.145 631.270 373.665 ;
        RECT 54.000 372.975 631.270 373.145 ;
        RECT 42.555 372.205 43.765 372.955 ;
        RECT 43.935 372.205 49.280 372.975 ;
        RECT 49.455 372.205 631.270 372.975 ;
        RECT 42.470 372.035 631.270 372.205 ;
        RECT 42.555 371.285 43.765 372.035 ;
        RECT 42.555 370.745 43.075 371.285 ;
        RECT 43.935 371.265 49.280 372.035 ;
        RECT 49.455 371.265 631.270 372.035 ;
        RECT 43.245 370.575 43.765 371.115 ;
        RECT 43.935 370.745 46.515 371.265 ;
        RECT 46.685 370.575 49.280 371.095 ;
        RECT 49.455 370.745 52.035 371.265 ;
        RECT 54.000 371.095 631.270 371.265 ;
        RECT 52.205 370.575 631.270 371.095 ;
        RECT 42.555 369.485 43.765 370.575 ;
        RECT 43.935 369.485 49.280 370.575 ;
        RECT 49.455 369.485 631.270 370.575 ;
        RECT 42.470 369.315 631.270 369.485 ;
        RECT 42.555 368.225 43.765 369.315 ;
        RECT 43.935 368.225 49.280 369.315 ;
        RECT 49.455 368.225 631.270 369.315 ;
        RECT 42.555 367.515 43.075 368.055 ;
        RECT 43.245 367.685 43.765 368.225 ;
        RECT 43.935 367.535 46.515 368.055 ;
        RECT 46.685 367.705 49.280 368.225 ;
        RECT 49.455 367.535 52.035 368.055 ;
        RECT 52.205 367.705 631.270 368.225 ;
        RECT 54.000 367.535 631.270 367.705 ;
        RECT 42.555 366.765 43.765 367.515 ;
        RECT 43.935 366.765 49.280 367.535 ;
        RECT 49.455 366.765 631.270 367.535 ;
        RECT 42.470 366.595 631.270 366.765 ;
        RECT 42.555 365.845 43.765 366.595 ;
        RECT 42.555 365.305 43.075 365.845 ;
        RECT 43.935 365.825 49.280 366.595 ;
        RECT 49.455 365.825 631.270 366.595 ;
        RECT 43.245 365.135 43.765 365.675 ;
        RECT 43.935 365.305 46.515 365.825 ;
        RECT 46.685 365.135 49.280 365.655 ;
        RECT 49.455 365.305 52.035 365.825 ;
        RECT 54.000 365.655 631.270 365.825 ;
        RECT 52.205 365.135 631.270 365.655 ;
        RECT 42.555 364.045 43.765 365.135 ;
        RECT 43.935 364.045 49.280 365.135 ;
        RECT 49.455 364.045 631.270 365.135 ;
        RECT 42.470 363.875 631.270 364.045 ;
        RECT 42.555 362.785 43.765 363.875 ;
        RECT 43.935 362.785 49.280 363.875 ;
        RECT 49.455 362.785 631.270 363.875 ;
        RECT 42.555 362.075 43.075 362.615 ;
        RECT 43.245 362.245 43.765 362.785 ;
        RECT 43.935 362.095 46.515 362.615 ;
        RECT 46.685 362.265 49.280 362.785 ;
        RECT 49.455 362.095 52.035 362.615 ;
        RECT 52.205 362.265 631.270 362.785 ;
        RECT 54.000 362.095 631.270 362.265 ;
        RECT 42.555 361.325 43.765 362.075 ;
        RECT 43.935 361.325 49.280 362.095 ;
        RECT 49.455 361.325 631.270 362.095 ;
        RECT 42.470 361.155 631.270 361.325 ;
        RECT 42.555 360.405 43.765 361.155 ;
        RECT 42.555 359.865 43.075 360.405 ;
        RECT 43.935 360.385 49.280 361.155 ;
        RECT 49.455 360.385 631.270 361.155 ;
        RECT 43.245 359.695 43.765 360.235 ;
        RECT 43.935 359.865 46.515 360.385 ;
        RECT 46.685 359.695 49.280 360.215 ;
        RECT 49.455 359.865 52.035 360.385 ;
        RECT 54.000 360.215 631.270 360.385 ;
        RECT 52.205 359.695 631.270 360.215 ;
        RECT 42.555 358.605 43.765 359.695 ;
        RECT 43.935 358.605 49.280 359.695 ;
        RECT 49.455 358.605 631.270 359.695 ;
        RECT 42.470 358.435 631.270 358.605 ;
        RECT 42.555 357.345 43.765 358.435 ;
        RECT 43.935 357.345 49.280 358.435 ;
        RECT 49.455 357.345 631.270 358.435 ;
        RECT 42.555 356.635 43.075 357.175 ;
        RECT 43.245 356.805 43.765 357.345 ;
        RECT 43.935 356.655 46.515 357.175 ;
        RECT 46.685 356.825 49.280 357.345 ;
        RECT 49.455 356.655 52.035 357.175 ;
        RECT 52.205 356.825 631.270 357.345 ;
        RECT 54.000 356.655 631.270 356.825 ;
        RECT 42.555 355.885 43.765 356.635 ;
        RECT 43.935 355.885 49.280 356.655 ;
        RECT 49.455 355.885 631.270 356.655 ;
        RECT 42.470 355.715 631.270 355.885 ;
        RECT 42.555 354.965 43.765 355.715 ;
        RECT 42.555 354.425 43.075 354.965 ;
        RECT 43.935 354.945 49.280 355.715 ;
        RECT 49.455 354.945 631.270 355.715 ;
        RECT 43.245 354.255 43.765 354.795 ;
        RECT 43.935 354.425 46.515 354.945 ;
        RECT 46.685 354.255 49.280 354.775 ;
        RECT 49.455 354.425 52.035 354.945 ;
        RECT 54.000 354.775 631.270 354.945 ;
        RECT 52.205 354.255 631.270 354.775 ;
        RECT 42.555 353.165 43.765 354.255 ;
        RECT 43.935 353.165 49.280 354.255 ;
        RECT 49.455 353.165 631.270 354.255 ;
        RECT 42.470 352.995 631.270 353.165 ;
        RECT 42.555 351.905 43.765 352.995 ;
        RECT 43.935 351.905 49.280 352.995 ;
        RECT 49.455 351.905 631.270 352.995 ;
        RECT 42.555 351.195 43.075 351.735 ;
        RECT 43.245 351.365 43.765 351.905 ;
        RECT 43.935 351.215 46.515 351.735 ;
        RECT 46.685 351.385 49.280 351.905 ;
        RECT 49.455 351.215 52.035 351.735 ;
        RECT 52.205 351.385 631.270 351.905 ;
        RECT 54.000 351.215 631.270 351.385 ;
        RECT 42.555 350.445 43.765 351.195 ;
        RECT 43.935 350.445 49.280 351.215 ;
        RECT 49.455 350.445 631.270 351.215 ;
        RECT 42.470 350.275 631.270 350.445 ;
        RECT 42.555 349.525 43.765 350.275 ;
        RECT 42.555 348.985 43.075 349.525 ;
        RECT 43.935 349.505 49.280 350.275 ;
        RECT 49.455 349.505 631.270 350.275 ;
        RECT 43.245 348.815 43.765 349.355 ;
        RECT 43.935 348.985 46.515 349.505 ;
        RECT 46.685 348.815 49.280 349.335 ;
        RECT 49.455 348.985 52.035 349.505 ;
        RECT 54.000 349.335 631.270 349.505 ;
        RECT 52.205 348.815 631.270 349.335 ;
        RECT 42.555 347.725 43.765 348.815 ;
        RECT 43.935 347.725 49.280 348.815 ;
        RECT 49.455 347.725 631.270 348.815 ;
        RECT 42.470 347.555 631.270 347.725 ;
        RECT 42.555 346.465 43.765 347.555 ;
        RECT 43.935 346.465 49.280 347.555 ;
        RECT 49.455 346.465 631.270 347.555 ;
        RECT 42.555 345.755 43.075 346.295 ;
        RECT 43.245 345.925 43.765 346.465 ;
        RECT 43.935 345.775 46.515 346.295 ;
        RECT 46.685 345.945 49.280 346.465 ;
        RECT 49.455 345.775 52.035 346.295 ;
        RECT 52.205 345.945 631.270 346.465 ;
        RECT 54.000 345.775 631.270 345.945 ;
        RECT 42.555 345.005 43.765 345.755 ;
        RECT 43.935 345.005 49.280 345.775 ;
        RECT 49.455 345.005 631.270 345.775 ;
        RECT 42.470 344.835 631.270 345.005 ;
        RECT 42.555 344.085 43.765 344.835 ;
        RECT 42.555 343.545 43.075 344.085 ;
        RECT 43.935 344.065 49.280 344.835 ;
        RECT 49.455 344.065 631.270 344.835 ;
        RECT 43.245 343.375 43.765 343.915 ;
        RECT 43.935 343.545 46.515 344.065 ;
        RECT 46.685 343.375 49.280 343.895 ;
        RECT 49.455 343.545 52.035 344.065 ;
        RECT 54.000 343.895 631.270 344.065 ;
        RECT 52.205 343.375 631.270 343.895 ;
        RECT 42.555 342.285 43.765 343.375 ;
        RECT 43.935 342.285 49.280 343.375 ;
        RECT 49.455 342.285 631.270 343.375 ;
        RECT 42.470 342.115 631.270 342.285 ;
        RECT 42.555 341.025 43.765 342.115 ;
        RECT 43.935 341.025 49.280 342.115 ;
        RECT 49.455 341.025 631.270 342.115 ;
        RECT 42.555 340.315 43.075 340.855 ;
        RECT 43.245 340.485 43.765 341.025 ;
        RECT 43.935 340.335 46.515 340.855 ;
        RECT 46.685 340.505 49.280 341.025 ;
        RECT 49.455 340.335 52.035 340.855 ;
        RECT 52.205 340.505 631.270 341.025 ;
        RECT 54.000 340.335 631.270 340.505 ;
        RECT 42.555 339.565 43.765 340.315 ;
        RECT 43.935 339.565 49.280 340.335 ;
        RECT 49.455 339.565 631.270 340.335 ;
        RECT 42.470 339.395 631.270 339.565 ;
        RECT 42.555 338.645 43.765 339.395 ;
        RECT 42.555 338.105 43.075 338.645 ;
        RECT 43.935 338.625 49.280 339.395 ;
        RECT 49.455 338.625 631.270 339.395 ;
        RECT 43.245 337.935 43.765 338.475 ;
        RECT 43.935 338.105 46.515 338.625 ;
        RECT 46.685 337.935 49.280 338.455 ;
        RECT 49.455 338.105 52.035 338.625 ;
        RECT 54.000 338.455 631.270 338.625 ;
        RECT 52.205 337.935 631.270 338.455 ;
        RECT 42.555 336.845 43.765 337.935 ;
        RECT 43.935 336.845 49.280 337.935 ;
        RECT 49.455 336.845 631.270 337.935 ;
        RECT 42.470 336.675 631.270 336.845 ;
        RECT 42.555 335.585 43.765 336.675 ;
        RECT 43.935 335.585 49.280 336.675 ;
        RECT 49.455 335.585 631.270 336.675 ;
        RECT 42.555 334.875 43.075 335.415 ;
        RECT 43.245 335.045 43.765 335.585 ;
        RECT 43.935 334.895 46.515 335.415 ;
        RECT 46.685 335.065 49.280 335.585 ;
        RECT 49.455 334.895 52.035 335.415 ;
        RECT 52.205 335.065 631.270 335.585 ;
        RECT 54.000 334.895 631.270 335.065 ;
        RECT 42.555 334.125 43.765 334.875 ;
        RECT 43.935 334.125 49.280 334.895 ;
        RECT 49.455 334.125 631.270 334.895 ;
        RECT 42.470 333.955 631.270 334.125 ;
        RECT 42.555 333.205 43.765 333.955 ;
        RECT 42.555 332.665 43.075 333.205 ;
        RECT 43.935 333.185 49.280 333.955 ;
        RECT 49.455 333.185 631.270 333.955 ;
        RECT 43.245 332.495 43.765 333.035 ;
        RECT 43.935 332.665 46.515 333.185 ;
        RECT 46.685 332.495 49.280 333.015 ;
        RECT 49.455 332.665 52.035 333.185 ;
        RECT 54.000 333.015 631.270 333.185 ;
        RECT 52.205 332.495 631.270 333.015 ;
        RECT 42.555 331.405 43.765 332.495 ;
        RECT 43.935 331.405 49.280 332.495 ;
        RECT 49.455 331.405 631.270 332.495 ;
        RECT 42.470 331.235 631.270 331.405 ;
        RECT 42.555 330.145 43.765 331.235 ;
        RECT 43.935 330.145 49.280 331.235 ;
        RECT 49.455 330.145 631.270 331.235 ;
        RECT 42.555 329.435 43.075 329.975 ;
        RECT 43.245 329.605 43.765 330.145 ;
        RECT 43.935 329.455 46.515 329.975 ;
        RECT 46.685 329.625 49.280 330.145 ;
        RECT 49.455 329.455 52.035 329.975 ;
        RECT 52.205 329.625 631.270 330.145 ;
        RECT 54.000 329.455 631.270 329.625 ;
        RECT 42.555 328.685 43.765 329.435 ;
        RECT 43.935 328.685 49.280 329.455 ;
        RECT 49.455 328.685 631.270 329.455 ;
        RECT 42.470 328.515 631.270 328.685 ;
        RECT 42.555 327.765 43.765 328.515 ;
        RECT 42.555 327.225 43.075 327.765 ;
        RECT 43.935 327.745 49.280 328.515 ;
        RECT 49.455 327.745 631.270 328.515 ;
        RECT 43.245 327.055 43.765 327.595 ;
        RECT 43.935 327.225 46.515 327.745 ;
        RECT 46.685 327.055 49.280 327.575 ;
        RECT 49.455 327.225 52.035 327.745 ;
        RECT 54.000 327.575 631.270 327.745 ;
        RECT 52.205 327.055 631.270 327.575 ;
        RECT 42.555 325.965 43.765 327.055 ;
        RECT 43.935 325.965 49.280 327.055 ;
        RECT 49.455 325.965 631.270 327.055 ;
        RECT 42.470 325.795 631.270 325.965 ;
        RECT 42.555 324.705 43.765 325.795 ;
        RECT 43.935 324.705 49.280 325.795 ;
        RECT 49.455 324.705 631.270 325.795 ;
        RECT 42.555 323.995 43.075 324.535 ;
        RECT 43.245 324.165 43.765 324.705 ;
        RECT 43.935 324.015 46.515 324.535 ;
        RECT 46.685 324.185 49.280 324.705 ;
        RECT 49.455 324.015 52.035 324.535 ;
        RECT 52.205 324.185 631.270 324.705 ;
        RECT 54.000 324.015 631.270 324.185 ;
        RECT 42.555 323.245 43.765 323.995 ;
        RECT 43.935 323.245 49.280 324.015 ;
        RECT 49.455 323.245 631.270 324.015 ;
        RECT 42.470 323.075 631.270 323.245 ;
        RECT 42.555 322.325 43.765 323.075 ;
        RECT 42.555 321.785 43.075 322.325 ;
        RECT 43.935 322.305 49.280 323.075 ;
        RECT 49.455 322.305 631.270 323.075 ;
        RECT 43.245 321.615 43.765 322.155 ;
        RECT 43.935 321.785 46.515 322.305 ;
        RECT 46.685 321.615 49.280 322.135 ;
        RECT 49.455 321.785 52.035 322.305 ;
        RECT 54.000 322.135 631.270 322.305 ;
        RECT 52.205 321.615 631.270 322.135 ;
        RECT 42.555 320.525 43.765 321.615 ;
        RECT 43.935 320.525 49.280 321.615 ;
        RECT 49.455 320.525 631.270 321.615 ;
        RECT 42.470 320.355 631.270 320.525 ;
        RECT 42.555 319.265 43.765 320.355 ;
        RECT 43.935 319.265 49.280 320.355 ;
        RECT 49.455 319.265 631.270 320.355 ;
        RECT 42.555 318.555 43.075 319.095 ;
        RECT 43.245 318.725 43.765 319.265 ;
        RECT 43.935 318.575 46.515 319.095 ;
        RECT 46.685 318.745 49.280 319.265 ;
        RECT 49.455 318.575 52.035 319.095 ;
        RECT 52.205 318.745 631.270 319.265 ;
        RECT 54.000 318.575 631.270 318.745 ;
        RECT 42.555 317.805 43.765 318.555 ;
        RECT 43.935 317.805 49.280 318.575 ;
        RECT 49.455 317.805 631.270 318.575 ;
        RECT 42.470 317.635 631.270 317.805 ;
        RECT 42.555 316.885 43.765 317.635 ;
        RECT 42.555 316.345 43.075 316.885 ;
        RECT 43.935 316.865 49.280 317.635 ;
        RECT 49.455 316.865 631.270 317.635 ;
        RECT 43.245 316.175 43.765 316.715 ;
        RECT 43.935 316.345 46.515 316.865 ;
        RECT 46.685 316.175 49.280 316.695 ;
        RECT 49.455 316.345 52.035 316.865 ;
        RECT 54.000 316.695 631.270 316.865 ;
        RECT 52.205 316.175 631.270 316.695 ;
        RECT 42.555 315.085 43.765 316.175 ;
        RECT 43.935 315.085 49.280 316.175 ;
        RECT 49.455 315.085 631.270 316.175 ;
        RECT 42.470 314.915 631.270 315.085 ;
        RECT 42.555 313.825 43.765 314.915 ;
        RECT 43.935 313.825 49.280 314.915 ;
        RECT 49.455 313.825 631.270 314.915 ;
        RECT 42.555 313.115 43.075 313.655 ;
        RECT 43.245 313.285 43.765 313.825 ;
        RECT 43.935 313.135 46.515 313.655 ;
        RECT 46.685 313.305 49.280 313.825 ;
        RECT 49.455 313.135 52.035 313.655 ;
        RECT 52.205 313.305 631.270 313.825 ;
        RECT 54.000 313.135 631.270 313.305 ;
        RECT 42.555 312.365 43.765 313.115 ;
        RECT 43.935 312.365 49.280 313.135 ;
        RECT 49.455 312.365 631.270 313.135 ;
        RECT 42.470 312.195 631.270 312.365 ;
        RECT 42.555 311.445 43.765 312.195 ;
        RECT 42.555 310.905 43.075 311.445 ;
        RECT 43.935 311.425 49.280 312.195 ;
        RECT 49.455 311.425 631.270 312.195 ;
        RECT 43.245 310.735 43.765 311.275 ;
        RECT 43.935 310.905 46.515 311.425 ;
        RECT 46.685 310.735 49.280 311.255 ;
        RECT 49.455 310.905 52.035 311.425 ;
        RECT 54.000 311.255 631.270 311.425 ;
        RECT 52.205 310.735 631.270 311.255 ;
        RECT 42.555 309.645 43.765 310.735 ;
        RECT 43.935 309.645 49.280 310.735 ;
        RECT 49.455 309.645 631.270 310.735 ;
        RECT 42.470 309.475 631.270 309.645 ;
        RECT 42.555 308.385 43.765 309.475 ;
        RECT 43.935 308.385 49.280 309.475 ;
        RECT 49.455 308.385 631.270 309.475 ;
        RECT 42.555 307.675 43.075 308.215 ;
        RECT 43.245 307.845 43.765 308.385 ;
        RECT 43.935 307.695 46.515 308.215 ;
        RECT 46.685 307.865 49.280 308.385 ;
        RECT 49.455 307.695 52.035 308.215 ;
        RECT 52.205 307.865 631.270 308.385 ;
        RECT 54.000 307.695 631.270 307.865 ;
        RECT 42.555 306.925 43.765 307.675 ;
        RECT 43.935 306.925 49.280 307.695 ;
        RECT 49.455 306.925 631.270 307.695 ;
        RECT 42.470 306.755 631.270 306.925 ;
        RECT 42.555 306.005 43.765 306.755 ;
        RECT 42.555 305.465 43.075 306.005 ;
        RECT 43.935 305.985 49.280 306.755 ;
        RECT 49.455 305.985 631.270 306.755 ;
        RECT 43.245 305.295 43.765 305.835 ;
        RECT 43.935 305.465 46.515 305.985 ;
        RECT 46.685 305.295 49.280 305.815 ;
        RECT 49.455 305.465 52.035 305.985 ;
        RECT 54.000 305.815 631.270 305.985 ;
        RECT 52.205 305.295 631.270 305.815 ;
        RECT 42.555 304.205 43.765 305.295 ;
        RECT 43.935 304.205 49.280 305.295 ;
        RECT 49.455 304.205 631.270 305.295 ;
        RECT 42.470 304.035 631.270 304.205 ;
        RECT 42.555 302.945 43.765 304.035 ;
        RECT 43.935 302.945 49.280 304.035 ;
        RECT 49.455 302.945 631.270 304.035 ;
        RECT 42.555 302.235 43.075 302.775 ;
        RECT 43.245 302.405 43.765 302.945 ;
        RECT 43.935 302.255 46.515 302.775 ;
        RECT 46.685 302.425 49.280 302.945 ;
        RECT 49.455 302.255 52.035 302.775 ;
        RECT 52.205 302.425 631.270 302.945 ;
        RECT 54.000 302.255 631.270 302.425 ;
        RECT 42.555 301.485 43.765 302.235 ;
        RECT 43.935 301.485 49.280 302.255 ;
        RECT 49.455 301.485 631.270 302.255 ;
        RECT 42.470 301.315 631.270 301.485 ;
        RECT 42.555 300.565 43.765 301.315 ;
        RECT 42.555 300.025 43.075 300.565 ;
        RECT 43.935 300.545 49.280 301.315 ;
        RECT 49.455 300.545 631.270 301.315 ;
        RECT 43.245 299.855 43.765 300.395 ;
        RECT 43.935 300.025 46.515 300.545 ;
        RECT 46.685 299.855 49.280 300.375 ;
        RECT 49.455 300.025 52.035 300.545 ;
        RECT 54.000 300.375 631.270 300.545 ;
        RECT 52.205 299.855 631.270 300.375 ;
        RECT 42.555 298.765 43.765 299.855 ;
        RECT 43.935 298.765 49.280 299.855 ;
        RECT 49.455 298.765 631.270 299.855 ;
        RECT 42.470 298.595 631.270 298.765 ;
        RECT 42.555 297.505 43.765 298.595 ;
        RECT 43.935 297.505 49.280 298.595 ;
        RECT 49.455 297.505 631.270 298.595 ;
        RECT 42.555 296.795 43.075 297.335 ;
        RECT 43.245 296.965 43.765 297.505 ;
        RECT 43.935 296.815 46.515 297.335 ;
        RECT 46.685 296.985 49.280 297.505 ;
        RECT 49.455 296.815 52.035 297.335 ;
        RECT 52.205 296.985 631.270 297.505 ;
        RECT 54.000 296.815 631.270 296.985 ;
        RECT 42.555 296.045 43.765 296.795 ;
        RECT 43.935 296.045 49.280 296.815 ;
        RECT 49.455 296.045 631.270 296.815 ;
        RECT 42.470 295.875 631.270 296.045 ;
        RECT 42.555 295.125 43.765 295.875 ;
        RECT 42.555 294.585 43.075 295.125 ;
        RECT 43.935 295.105 49.280 295.875 ;
        RECT 49.455 295.105 631.270 295.875 ;
        RECT 43.245 294.415 43.765 294.955 ;
        RECT 43.935 294.585 46.515 295.105 ;
        RECT 46.685 294.415 49.280 294.935 ;
        RECT 49.455 294.585 52.035 295.105 ;
        RECT 54.000 294.935 631.270 295.105 ;
        RECT 52.205 294.415 631.270 294.935 ;
        RECT 42.555 293.325 43.765 294.415 ;
        RECT 43.935 293.325 49.280 294.415 ;
        RECT 49.455 293.325 631.270 294.415 ;
        RECT 42.470 293.155 631.270 293.325 ;
        RECT 42.555 292.065 43.765 293.155 ;
        RECT 43.935 292.065 49.280 293.155 ;
        RECT 49.455 292.065 631.270 293.155 ;
        RECT 42.555 291.355 43.075 291.895 ;
        RECT 43.245 291.525 43.765 292.065 ;
        RECT 43.935 291.375 46.515 291.895 ;
        RECT 46.685 291.545 49.280 292.065 ;
        RECT 49.455 291.375 52.035 291.895 ;
        RECT 52.205 291.545 631.270 292.065 ;
        RECT 54.000 291.375 631.270 291.545 ;
        RECT 42.555 290.605 43.765 291.355 ;
        RECT 43.935 290.605 49.280 291.375 ;
        RECT 49.455 290.605 631.270 291.375 ;
        RECT 42.470 290.435 631.270 290.605 ;
        RECT 42.555 289.685 43.765 290.435 ;
        RECT 42.555 289.145 43.075 289.685 ;
        RECT 43.935 289.665 49.280 290.435 ;
        RECT 49.455 289.665 631.270 290.435 ;
        RECT 43.245 288.975 43.765 289.515 ;
        RECT 43.935 289.145 46.515 289.665 ;
        RECT 46.685 288.975 49.280 289.495 ;
        RECT 49.455 289.145 52.035 289.665 ;
        RECT 54.000 289.495 631.270 289.665 ;
        RECT 52.205 288.975 631.270 289.495 ;
        RECT 42.555 287.885 43.765 288.975 ;
        RECT 43.935 287.885 49.280 288.975 ;
        RECT 49.455 287.885 631.270 288.975 ;
        RECT 42.470 287.715 631.270 287.885 ;
        RECT 42.555 286.625 43.765 287.715 ;
        RECT 43.935 286.625 49.280 287.715 ;
        RECT 49.455 286.625 631.270 287.715 ;
        RECT 42.555 285.915 43.075 286.455 ;
        RECT 43.245 286.085 43.765 286.625 ;
        RECT 43.935 285.935 46.515 286.455 ;
        RECT 46.685 286.105 49.280 286.625 ;
        RECT 49.455 285.935 52.035 286.455 ;
        RECT 52.205 286.105 631.270 286.625 ;
        RECT 54.000 285.935 631.270 286.105 ;
        RECT 42.555 285.165 43.765 285.915 ;
        RECT 43.935 285.165 49.280 285.935 ;
        RECT 49.455 285.165 631.270 285.935 ;
        RECT 42.470 284.995 631.270 285.165 ;
        RECT 42.555 284.245 43.765 284.995 ;
        RECT 42.555 283.705 43.075 284.245 ;
        RECT 43.935 284.225 49.280 284.995 ;
        RECT 49.455 284.225 631.270 284.995 ;
        RECT 43.245 283.535 43.765 284.075 ;
        RECT 43.935 283.705 46.515 284.225 ;
        RECT 46.685 283.535 49.280 284.055 ;
        RECT 49.455 283.705 52.035 284.225 ;
        RECT 54.000 284.055 631.270 284.225 ;
        RECT 52.205 283.535 631.270 284.055 ;
        RECT 42.555 282.445 43.765 283.535 ;
        RECT 43.935 282.445 49.280 283.535 ;
        RECT 49.455 282.445 631.270 283.535 ;
        RECT 42.470 282.275 631.270 282.445 ;
        RECT 42.555 281.185 43.765 282.275 ;
        RECT 43.935 281.185 49.280 282.275 ;
        RECT 49.455 281.185 631.270 282.275 ;
        RECT 42.555 280.475 43.075 281.015 ;
        RECT 43.245 280.645 43.765 281.185 ;
        RECT 43.935 280.495 46.515 281.015 ;
        RECT 46.685 280.665 49.280 281.185 ;
        RECT 49.455 280.495 52.035 281.015 ;
        RECT 52.205 280.665 631.270 281.185 ;
        RECT 54.000 280.495 631.270 280.665 ;
        RECT 42.555 279.725 43.765 280.475 ;
        RECT 43.935 279.725 49.280 280.495 ;
        RECT 49.455 279.725 631.270 280.495 ;
        RECT 42.470 279.555 631.270 279.725 ;
        RECT 42.555 278.805 43.765 279.555 ;
        RECT 42.555 278.265 43.075 278.805 ;
        RECT 43.935 278.785 49.280 279.555 ;
        RECT 49.455 278.785 631.270 279.555 ;
        RECT 43.245 278.095 43.765 278.635 ;
        RECT 43.935 278.265 46.515 278.785 ;
        RECT 46.685 278.095 49.280 278.615 ;
        RECT 49.455 278.265 52.035 278.785 ;
        RECT 54.000 278.615 631.270 278.785 ;
        RECT 52.205 278.095 631.270 278.615 ;
        RECT 42.555 277.005 43.765 278.095 ;
        RECT 43.935 277.005 49.280 278.095 ;
        RECT 49.455 277.005 631.270 278.095 ;
        RECT 42.470 276.835 631.270 277.005 ;
        RECT 42.555 275.745 43.765 276.835 ;
        RECT 43.935 275.745 49.280 276.835 ;
        RECT 49.455 275.745 631.270 276.835 ;
        RECT 42.555 275.035 43.075 275.575 ;
        RECT 43.245 275.205 43.765 275.745 ;
        RECT 43.935 275.055 46.515 275.575 ;
        RECT 46.685 275.225 49.280 275.745 ;
        RECT 49.455 275.055 52.035 275.575 ;
        RECT 52.205 275.225 631.270 275.745 ;
        RECT 54.000 275.055 631.270 275.225 ;
        RECT 42.555 274.285 43.765 275.035 ;
        RECT 43.935 274.285 49.280 275.055 ;
        RECT 49.455 274.285 631.270 275.055 ;
        RECT 42.470 274.115 631.270 274.285 ;
        RECT 42.555 273.365 43.765 274.115 ;
        RECT 42.555 272.825 43.075 273.365 ;
        RECT 43.935 273.345 49.280 274.115 ;
        RECT 49.455 273.345 631.270 274.115 ;
        RECT 43.245 272.655 43.765 273.195 ;
        RECT 43.935 272.825 46.515 273.345 ;
        RECT 46.685 272.655 49.280 273.175 ;
        RECT 49.455 272.825 52.035 273.345 ;
        RECT 54.000 273.175 631.270 273.345 ;
        RECT 52.205 272.655 631.270 273.175 ;
        RECT 42.555 271.565 43.765 272.655 ;
        RECT 43.935 271.565 49.280 272.655 ;
        RECT 49.455 271.565 631.270 272.655 ;
        RECT 42.470 271.395 631.270 271.565 ;
        RECT 42.555 270.305 43.765 271.395 ;
        RECT 43.935 270.305 49.280 271.395 ;
        RECT 49.455 270.305 631.270 271.395 ;
        RECT 42.555 269.595 43.075 270.135 ;
        RECT 43.245 269.765 43.765 270.305 ;
        RECT 43.935 269.615 46.515 270.135 ;
        RECT 46.685 269.785 49.280 270.305 ;
        RECT 49.455 269.615 52.035 270.135 ;
        RECT 52.205 269.785 631.270 270.305 ;
        RECT 54.000 269.615 631.270 269.785 ;
        RECT 42.555 268.845 43.765 269.595 ;
        RECT 43.935 268.845 49.280 269.615 ;
        RECT 49.455 268.845 631.270 269.615 ;
        RECT 42.470 268.675 631.270 268.845 ;
        RECT 42.555 267.925 43.765 268.675 ;
        RECT 42.555 267.385 43.075 267.925 ;
        RECT 43.935 267.905 49.280 268.675 ;
        RECT 49.455 267.905 631.270 268.675 ;
        RECT 43.245 267.215 43.765 267.755 ;
        RECT 43.935 267.385 46.515 267.905 ;
        RECT 46.685 267.215 49.280 267.735 ;
        RECT 49.455 267.385 52.035 267.905 ;
        RECT 54.000 267.735 631.270 267.905 ;
        RECT 52.205 267.215 631.270 267.735 ;
        RECT 42.555 266.125 43.765 267.215 ;
        RECT 43.935 266.125 49.280 267.215 ;
        RECT 49.455 266.125 631.270 267.215 ;
        RECT 42.470 265.955 631.270 266.125 ;
        RECT 42.555 264.865 43.765 265.955 ;
        RECT 43.935 264.865 49.280 265.955 ;
        RECT 49.455 264.865 631.270 265.955 ;
        RECT 42.555 264.155 43.075 264.695 ;
        RECT 43.245 264.325 43.765 264.865 ;
        RECT 43.935 264.175 46.515 264.695 ;
        RECT 46.685 264.345 49.280 264.865 ;
        RECT 49.455 264.175 52.035 264.695 ;
        RECT 52.205 264.345 631.270 264.865 ;
        RECT 54.000 264.175 631.270 264.345 ;
        RECT 42.555 263.405 43.765 264.155 ;
        RECT 43.935 263.405 49.280 264.175 ;
        RECT 49.455 263.405 631.270 264.175 ;
        RECT 42.470 263.235 631.270 263.405 ;
        RECT 42.555 262.485 43.765 263.235 ;
        RECT 42.555 261.945 43.075 262.485 ;
        RECT 43.935 262.465 49.280 263.235 ;
        RECT 49.455 262.465 631.270 263.235 ;
        RECT 43.245 261.775 43.765 262.315 ;
        RECT 43.935 261.945 46.515 262.465 ;
        RECT 46.685 261.775 49.280 262.295 ;
        RECT 49.455 261.945 52.035 262.465 ;
        RECT 54.000 262.295 631.270 262.465 ;
        RECT 52.205 261.775 631.270 262.295 ;
        RECT 42.555 260.685 43.765 261.775 ;
        RECT 43.935 260.685 49.280 261.775 ;
        RECT 49.455 260.685 631.270 261.775 ;
        RECT 42.470 260.515 631.270 260.685 ;
        RECT 42.555 259.425 43.765 260.515 ;
        RECT 43.935 259.425 49.280 260.515 ;
        RECT 49.455 259.425 631.270 260.515 ;
        RECT 42.555 258.715 43.075 259.255 ;
        RECT 43.245 258.885 43.765 259.425 ;
        RECT 43.935 258.735 46.515 259.255 ;
        RECT 46.685 258.905 49.280 259.425 ;
        RECT 49.455 258.735 52.035 259.255 ;
        RECT 52.205 258.905 631.270 259.425 ;
        RECT 54.000 258.735 631.270 258.905 ;
        RECT 42.555 257.965 43.765 258.715 ;
        RECT 43.935 257.965 49.280 258.735 ;
        RECT 49.455 257.965 631.270 258.735 ;
        RECT 42.470 257.795 631.270 257.965 ;
        RECT 42.555 257.045 43.765 257.795 ;
        RECT 42.555 256.505 43.075 257.045 ;
        RECT 43.935 257.025 49.280 257.795 ;
        RECT 49.455 257.025 631.270 257.795 ;
        RECT 43.245 256.335 43.765 256.875 ;
        RECT 43.935 256.505 46.515 257.025 ;
        RECT 46.685 256.335 49.280 256.855 ;
        RECT 49.455 256.505 52.035 257.025 ;
        RECT 54.000 256.855 631.270 257.025 ;
        RECT 52.205 256.335 631.270 256.855 ;
        RECT 42.555 255.245 43.765 256.335 ;
        RECT 43.935 255.245 49.280 256.335 ;
        RECT 49.455 255.245 631.270 256.335 ;
        RECT 42.470 255.075 631.270 255.245 ;
        RECT 42.555 253.985 43.765 255.075 ;
        RECT 43.935 253.985 49.280 255.075 ;
        RECT 49.455 253.985 631.270 255.075 ;
        RECT 42.555 253.275 43.075 253.815 ;
        RECT 43.245 253.445 43.765 253.985 ;
        RECT 43.935 253.295 46.515 253.815 ;
        RECT 46.685 253.465 49.280 253.985 ;
        RECT 49.455 253.295 52.035 253.815 ;
        RECT 52.205 253.465 631.270 253.985 ;
        RECT 54.000 253.295 631.270 253.465 ;
        RECT 42.555 252.525 43.765 253.275 ;
        RECT 43.935 252.525 49.280 253.295 ;
        RECT 49.455 252.525 631.270 253.295 ;
        RECT 42.470 252.355 631.270 252.525 ;
        RECT 42.555 251.605 43.765 252.355 ;
        RECT 42.555 251.065 43.075 251.605 ;
        RECT 43.935 251.585 49.280 252.355 ;
        RECT 49.455 251.585 631.270 252.355 ;
        RECT 43.245 250.895 43.765 251.435 ;
        RECT 43.935 251.065 46.515 251.585 ;
        RECT 46.685 250.895 49.280 251.415 ;
        RECT 49.455 251.065 52.035 251.585 ;
        RECT 54.000 251.415 631.270 251.585 ;
        RECT 52.205 250.895 631.270 251.415 ;
        RECT 42.555 249.805 43.765 250.895 ;
        RECT 43.935 249.805 49.280 250.895 ;
        RECT 49.455 249.805 631.270 250.895 ;
        RECT 42.470 249.635 631.270 249.805 ;
        RECT 42.555 248.545 43.765 249.635 ;
        RECT 43.935 248.545 49.280 249.635 ;
        RECT 49.455 248.545 631.270 249.635 ;
        RECT 42.555 247.835 43.075 248.375 ;
        RECT 43.245 248.005 43.765 248.545 ;
        RECT 43.935 247.855 46.515 248.375 ;
        RECT 46.685 248.025 49.280 248.545 ;
        RECT 49.455 247.855 52.035 248.375 ;
        RECT 52.205 248.025 631.270 248.545 ;
        RECT 54.000 247.855 631.270 248.025 ;
        RECT 42.555 247.085 43.765 247.835 ;
        RECT 43.935 247.085 49.280 247.855 ;
        RECT 49.455 247.085 631.270 247.855 ;
        RECT 42.470 246.915 631.270 247.085 ;
        RECT 42.555 246.165 43.765 246.915 ;
        RECT 42.555 245.625 43.075 246.165 ;
        RECT 43.935 246.145 49.280 246.915 ;
        RECT 49.455 246.145 631.270 246.915 ;
        RECT 43.245 245.455 43.765 245.995 ;
        RECT 43.935 245.625 46.515 246.145 ;
        RECT 46.685 245.455 49.280 245.975 ;
        RECT 49.455 245.625 52.035 246.145 ;
        RECT 54.000 245.975 631.270 246.145 ;
        RECT 52.205 245.455 631.270 245.975 ;
        RECT 42.555 244.365 43.765 245.455 ;
        RECT 43.935 244.365 49.280 245.455 ;
        RECT 49.455 244.365 631.270 245.455 ;
        RECT 42.470 244.195 631.270 244.365 ;
        RECT 42.555 243.105 43.765 244.195 ;
        RECT 43.935 243.105 49.280 244.195 ;
        RECT 49.455 243.105 631.270 244.195 ;
        RECT 42.555 242.395 43.075 242.935 ;
        RECT 43.245 242.565 43.765 243.105 ;
        RECT 43.935 242.415 46.515 242.935 ;
        RECT 46.685 242.585 49.280 243.105 ;
        RECT 49.455 242.415 52.035 242.935 ;
        RECT 52.205 242.585 631.270 243.105 ;
        RECT 54.000 242.415 631.270 242.585 ;
        RECT 42.555 241.645 43.765 242.395 ;
        RECT 43.935 241.645 49.280 242.415 ;
        RECT 49.455 241.645 631.270 242.415 ;
        RECT 42.470 241.475 631.270 241.645 ;
        RECT 42.555 240.725 43.765 241.475 ;
        RECT 42.555 240.185 43.075 240.725 ;
        RECT 43.935 240.705 49.280 241.475 ;
        RECT 49.455 240.705 631.270 241.475 ;
        RECT 43.245 240.015 43.765 240.555 ;
        RECT 43.935 240.185 46.515 240.705 ;
        RECT 46.685 240.015 49.280 240.535 ;
        RECT 49.455 240.185 52.035 240.705 ;
        RECT 54.000 240.535 631.270 240.705 ;
        RECT 52.205 240.015 631.270 240.535 ;
        RECT 42.555 238.925 43.765 240.015 ;
        RECT 43.935 238.925 49.280 240.015 ;
        RECT 49.455 238.925 631.270 240.015 ;
        RECT 42.470 238.755 631.270 238.925 ;
        RECT 42.555 237.665 43.765 238.755 ;
        RECT 43.935 237.665 49.280 238.755 ;
        RECT 49.455 237.665 631.270 238.755 ;
        RECT 42.555 236.955 43.075 237.495 ;
        RECT 43.245 237.125 43.765 237.665 ;
        RECT 43.935 236.975 46.515 237.495 ;
        RECT 46.685 237.145 49.280 237.665 ;
        RECT 49.455 236.975 52.035 237.495 ;
        RECT 52.205 237.145 631.270 237.665 ;
        RECT 54.000 236.975 631.270 237.145 ;
        RECT 42.555 236.205 43.765 236.955 ;
        RECT 43.935 236.205 49.280 236.975 ;
        RECT 49.455 236.205 631.270 236.975 ;
        RECT 42.470 236.035 631.270 236.205 ;
        RECT 42.555 235.285 43.765 236.035 ;
        RECT 42.555 234.745 43.075 235.285 ;
        RECT 43.935 235.265 49.280 236.035 ;
        RECT 49.455 235.265 631.270 236.035 ;
        RECT 43.245 234.575 43.765 235.115 ;
        RECT 43.935 234.745 46.515 235.265 ;
        RECT 46.685 234.575 49.280 235.095 ;
        RECT 49.455 234.745 52.035 235.265 ;
        RECT 54.000 235.095 631.270 235.265 ;
        RECT 52.205 234.575 631.270 235.095 ;
        RECT 42.555 233.485 43.765 234.575 ;
        RECT 43.935 233.485 49.280 234.575 ;
        RECT 49.455 233.485 631.270 234.575 ;
        RECT 42.470 233.315 631.270 233.485 ;
        RECT 42.555 232.225 43.765 233.315 ;
        RECT 43.935 232.225 49.280 233.315 ;
        RECT 49.455 232.225 631.270 233.315 ;
        RECT 42.555 231.515 43.075 232.055 ;
        RECT 43.245 231.685 43.765 232.225 ;
        RECT 43.935 231.535 46.515 232.055 ;
        RECT 46.685 231.705 49.280 232.225 ;
        RECT 49.455 231.535 52.035 232.055 ;
        RECT 52.205 231.705 631.270 232.225 ;
        RECT 54.000 231.535 631.270 231.705 ;
        RECT 42.555 230.765 43.765 231.515 ;
        RECT 43.935 230.765 49.280 231.535 ;
        RECT 49.455 230.765 631.270 231.535 ;
        RECT 42.470 230.595 631.270 230.765 ;
        RECT 42.555 229.845 43.765 230.595 ;
        RECT 42.555 229.305 43.075 229.845 ;
        RECT 43.935 229.825 49.280 230.595 ;
        RECT 49.455 229.825 631.270 230.595 ;
        RECT 43.245 229.135 43.765 229.675 ;
        RECT 43.935 229.305 46.515 229.825 ;
        RECT 46.685 229.135 49.280 229.655 ;
        RECT 49.455 229.305 52.035 229.825 ;
        RECT 54.000 229.655 631.270 229.825 ;
        RECT 52.205 229.135 631.270 229.655 ;
        RECT 42.555 228.045 43.765 229.135 ;
        RECT 43.935 228.045 49.280 229.135 ;
        RECT 49.455 228.045 631.270 229.135 ;
        RECT 42.470 227.875 631.270 228.045 ;
        RECT 42.555 226.785 43.765 227.875 ;
        RECT 43.935 226.785 49.280 227.875 ;
        RECT 49.455 226.785 631.270 227.875 ;
        RECT 42.555 226.075 43.075 226.615 ;
        RECT 43.245 226.245 43.765 226.785 ;
        RECT 43.935 226.095 46.515 226.615 ;
        RECT 46.685 226.265 49.280 226.785 ;
        RECT 49.455 226.095 52.035 226.615 ;
        RECT 52.205 226.265 631.270 226.785 ;
        RECT 54.000 226.095 631.270 226.265 ;
        RECT 42.555 225.325 43.765 226.075 ;
        RECT 43.935 225.325 49.280 226.095 ;
        RECT 49.455 225.325 631.270 226.095 ;
        RECT 42.470 225.155 631.270 225.325 ;
        RECT 42.555 224.405 43.765 225.155 ;
        RECT 42.555 223.865 43.075 224.405 ;
        RECT 43.935 224.385 49.280 225.155 ;
        RECT 49.455 224.385 631.270 225.155 ;
        RECT 43.245 223.695 43.765 224.235 ;
        RECT 43.935 223.865 46.515 224.385 ;
        RECT 46.685 223.695 49.280 224.215 ;
        RECT 49.455 223.865 52.035 224.385 ;
        RECT 54.000 224.215 631.270 224.385 ;
        RECT 52.205 223.695 631.270 224.215 ;
        RECT 42.555 222.605 43.765 223.695 ;
        RECT 43.935 222.605 49.280 223.695 ;
        RECT 49.455 222.605 631.270 223.695 ;
        RECT 42.470 222.435 631.270 222.605 ;
        RECT 42.555 221.345 43.765 222.435 ;
        RECT 43.935 221.345 49.280 222.435 ;
        RECT 49.455 221.345 631.270 222.435 ;
        RECT 42.555 220.635 43.075 221.175 ;
        RECT 43.245 220.805 43.765 221.345 ;
        RECT 43.935 220.655 46.515 221.175 ;
        RECT 46.685 220.825 49.280 221.345 ;
        RECT 49.455 220.655 52.035 221.175 ;
        RECT 52.205 220.825 631.270 221.345 ;
        RECT 54.000 220.655 631.270 220.825 ;
        RECT 42.555 219.885 43.765 220.635 ;
        RECT 43.935 219.885 49.280 220.655 ;
        RECT 49.455 219.885 631.270 220.655 ;
        RECT 42.470 219.715 631.270 219.885 ;
        RECT 42.555 218.965 43.765 219.715 ;
        RECT 42.555 218.425 43.075 218.965 ;
        RECT 43.935 218.945 49.280 219.715 ;
        RECT 49.455 218.945 631.270 219.715 ;
        RECT 43.245 218.255 43.765 218.795 ;
        RECT 43.935 218.425 46.515 218.945 ;
        RECT 46.685 218.255 49.280 218.775 ;
        RECT 49.455 218.425 52.035 218.945 ;
        RECT 54.000 218.775 631.270 218.945 ;
        RECT 52.205 218.255 631.270 218.775 ;
        RECT 42.555 217.165 43.765 218.255 ;
        RECT 43.935 217.165 49.280 218.255 ;
        RECT 49.455 217.165 631.270 218.255 ;
        RECT 42.470 216.995 631.270 217.165 ;
        RECT 42.555 215.905 43.765 216.995 ;
        RECT 43.935 215.905 49.280 216.995 ;
        RECT 49.455 215.905 631.270 216.995 ;
        RECT 42.555 215.195 43.075 215.735 ;
        RECT 43.245 215.365 43.765 215.905 ;
        RECT 43.935 215.215 46.515 215.735 ;
        RECT 46.685 215.385 49.280 215.905 ;
        RECT 49.455 215.215 52.035 215.735 ;
        RECT 52.205 215.385 631.270 215.905 ;
        RECT 54.000 215.215 631.270 215.385 ;
        RECT 42.555 214.445 43.765 215.195 ;
        RECT 43.935 214.445 49.280 215.215 ;
        RECT 49.455 214.445 631.270 215.215 ;
        RECT 42.470 214.275 631.270 214.445 ;
        RECT 42.555 213.525 43.765 214.275 ;
        RECT 42.555 212.985 43.075 213.525 ;
        RECT 43.935 213.505 49.280 214.275 ;
        RECT 49.455 213.505 631.270 214.275 ;
        RECT 43.245 212.815 43.765 213.355 ;
        RECT 43.935 212.985 46.515 213.505 ;
        RECT 46.685 212.815 49.280 213.335 ;
        RECT 49.455 212.985 52.035 213.505 ;
        RECT 54.000 213.335 631.270 213.505 ;
        RECT 52.205 212.815 631.270 213.335 ;
        RECT 42.555 211.725 43.765 212.815 ;
        RECT 43.935 211.725 49.280 212.815 ;
        RECT 49.455 211.725 631.270 212.815 ;
        RECT 42.470 211.555 631.270 211.725 ;
        RECT 42.555 210.465 43.765 211.555 ;
        RECT 43.935 210.465 49.280 211.555 ;
        RECT 49.455 210.465 631.270 211.555 ;
        RECT 42.555 209.755 43.075 210.295 ;
        RECT 43.245 209.925 43.765 210.465 ;
        RECT 43.935 209.775 46.515 210.295 ;
        RECT 46.685 209.945 49.280 210.465 ;
        RECT 49.455 209.775 52.035 210.295 ;
        RECT 52.205 209.945 631.270 210.465 ;
        RECT 54.000 209.775 631.270 209.945 ;
        RECT 42.555 209.005 43.765 209.755 ;
        RECT 43.935 209.005 49.280 209.775 ;
        RECT 49.455 209.005 631.270 209.775 ;
        RECT 42.470 208.835 631.270 209.005 ;
        RECT 42.555 208.085 43.765 208.835 ;
        RECT 42.555 207.545 43.075 208.085 ;
        RECT 43.935 208.065 49.280 208.835 ;
        RECT 49.455 208.065 631.270 208.835 ;
        RECT 43.245 207.375 43.765 207.915 ;
        RECT 43.935 207.545 46.515 208.065 ;
        RECT 46.685 207.375 49.280 207.895 ;
        RECT 49.455 207.545 52.035 208.065 ;
        RECT 54.000 207.895 631.270 208.065 ;
        RECT 52.205 207.375 631.270 207.895 ;
        RECT 42.555 206.285 43.765 207.375 ;
        RECT 43.935 206.285 49.280 207.375 ;
        RECT 49.455 206.285 631.270 207.375 ;
        RECT 42.470 206.115 631.270 206.285 ;
        RECT 42.555 205.025 43.765 206.115 ;
        RECT 43.935 205.025 49.280 206.115 ;
        RECT 49.455 205.025 631.270 206.115 ;
        RECT 42.555 204.315 43.075 204.855 ;
        RECT 43.245 204.485 43.765 205.025 ;
        RECT 43.935 204.335 46.515 204.855 ;
        RECT 46.685 204.505 49.280 205.025 ;
        RECT 49.455 204.335 52.035 204.855 ;
        RECT 52.205 204.505 631.270 205.025 ;
        RECT 54.000 204.335 631.270 204.505 ;
        RECT 42.555 203.565 43.765 204.315 ;
        RECT 43.935 203.565 49.280 204.335 ;
        RECT 49.455 203.565 631.270 204.335 ;
        RECT 42.470 203.395 631.270 203.565 ;
        RECT 42.555 202.645 43.765 203.395 ;
        RECT 42.555 202.105 43.075 202.645 ;
        RECT 43.935 202.625 49.280 203.395 ;
        RECT 49.455 202.625 631.270 203.395 ;
        RECT 43.245 201.935 43.765 202.475 ;
        RECT 43.935 202.105 46.515 202.625 ;
        RECT 46.685 201.935 49.280 202.455 ;
        RECT 49.455 202.105 52.035 202.625 ;
        RECT 54.000 202.455 631.270 202.625 ;
        RECT 52.205 201.935 631.270 202.455 ;
        RECT 42.555 200.845 43.765 201.935 ;
        RECT 43.935 200.845 49.280 201.935 ;
        RECT 49.455 200.845 631.270 201.935 ;
        RECT 42.470 200.675 631.270 200.845 ;
        RECT 42.555 199.585 43.765 200.675 ;
        RECT 43.935 199.585 49.280 200.675 ;
        RECT 49.455 199.585 631.270 200.675 ;
        RECT 42.555 198.875 43.075 199.415 ;
        RECT 43.245 199.045 43.765 199.585 ;
        RECT 43.935 198.895 46.515 199.415 ;
        RECT 46.685 199.065 49.280 199.585 ;
        RECT 49.455 198.895 52.035 199.415 ;
        RECT 52.205 199.065 631.270 199.585 ;
        RECT 54.000 198.895 631.270 199.065 ;
        RECT 42.555 198.125 43.765 198.875 ;
        RECT 43.935 198.125 49.280 198.895 ;
        RECT 49.455 198.125 631.270 198.895 ;
        RECT 42.470 197.955 631.270 198.125 ;
        RECT 42.555 197.205 43.765 197.955 ;
        RECT 42.555 196.665 43.075 197.205 ;
        RECT 43.935 197.185 49.280 197.955 ;
        RECT 49.455 197.185 631.270 197.955 ;
        RECT 43.245 196.495 43.765 197.035 ;
        RECT 43.935 196.665 46.515 197.185 ;
        RECT 46.685 196.495 49.280 197.015 ;
        RECT 49.455 196.665 52.035 197.185 ;
        RECT 54.000 197.015 631.270 197.185 ;
        RECT 52.205 196.495 631.270 197.015 ;
        RECT 42.555 195.405 43.765 196.495 ;
        RECT 43.935 195.405 49.280 196.495 ;
        RECT 49.455 195.405 631.270 196.495 ;
        RECT 42.470 195.235 631.270 195.405 ;
        RECT 42.555 194.145 43.765 195.235 ;
        RECT 43.935 194.145 49.280 195.235 ;
        RECT 49.455 194.145 631.270 195.235 ;
        RECT 42.555 193.435 43.075 193.975 ;
        RECT 43.245 193.605 43.765 194.145 ;
        RECT 43.935 193.455 46.515 193.975 ;
        RECT 46.685 193.625 49.280 194.145 ;
        RECT 49.455 193.455 52.035 193.975 ;
        RECT 52.205 193.625 631.270 194.145 ;
        RECT 54.000 193.455 631.270 193.625 ;
        RECT 42.555 192.685 43.765 193.435 ;
        RECT 43.935 192.685 49.280 193.455 ;
        RECT 49.455 192.685 631.270 193.455 ;
        RECT 42.470 192.515 631.270 192.685 ;
        RECT 42.555 191.765 43.765 192.515 ;
        RECT 42.555 191.225 43.075 191.765 ;
        RECT 43.935 191.745 49.280 192.515 ;
        RECT 49.455 191.745 631.270 192.515 ;
        RECT 43.245 191.055 43.765 191.595 ;
        RECT 43.935 191.225 46.515 191.745 ;
        RECT 46.685 191.055 49.280 191.575 ;
        RECT 49.455 191.225 52.035 191.745 ;
        RECT 54.000 191.575 631.270 191.745 ;
        RECT 52.205 191.055 631.270 191.575 ;
        RECT 42.555 189.965 43.765 191.055 ;
        RECT 43.935 189.965 49.280 191.055 ;
        RECT 49.455 189.965 631.270 191.055 ;
        RECT 42.470 189.795 631.270 189.965 ;
        RECT 42.555 188.705 43.765 189.795 ;
        RECT 43.935 188.705 49.280 189.795 ;
        RECT 49.455 188.705 631.270 189.795 ;
        RECT 42.555 187.995 43.075 188.535 ;
        RECT 43.245 188.165 43.765 188.705 ;
        RECT 43.935 188.015 46.515 188.535 ;
        RECT 46.685 188.185 49.280 188.705 ;
        RECT 49.455 188.015 52.035 188.535 ;
        RECT 52.205 188.185 631.270 188.705 ;
        RECT 54.000 188.015 631.270 188.185 ;
        RECT 42.555 187.245 43.765 187.995 ;
        RECT 43.935 187.245 49.280 188.015 ;
        RECT 49.455 187.245 631.270 188.015 ;
        RECT 42.470 187.075 631.270 187.245 ;
        RECT 42.555 186.325 43.765 187.075 ;
        RECT 42.555 185.785 43.075 186.325 ;
        RECT 43.935 186.305 49.280 187.075 ;
        RECT 49.455 186.305 631.270 187.075 ;
        RECT 43.245 185.615 43.765 186.155 ;
        RECT 43.935 185.785 46.515 186.305 ;
        RECT 46.685 185.615 49.280 186.135 ;
        RECT 49.455 185.785 52.035 186.305 ;
        RECT 54.000 186.135 631.270 186.305 ;
        RECT 52.205 185.615 631.270 186.135 ;
        RECT 42.555 184.525 43.765 185.615 ;
        RECT 43.935 184.525 49.280 185.615 ;
        RECT 49.455 184.525 631.270 185.615 ;
        RECT 42.470 184.355 631.270 184.525 ;
        RECT 42.555 183.265 43.765 184.355 ;
        RECT 43.935 183.265 49.280 184.355 ;
        RECT 49.455 183.265 631.270 184.355 ;
        RECT 42.555 182.555 43.075 183.095 ;
        RECT 43.245 182.725 43.765 183.265 ;
        RECT 43.935 182.575 46.515 183.095 ;
        RECT 46.685 182.745 49.280 183.265 ;
        RECT 49.455 182.575 52.035 183.095 ;
        RECT 52.205 182.745 631.270 183.265 ;
        RECT 54.000 182.575 631.270 182.745 ;
        RECT 42.555 181.805 43.765 182.555 ;
        RECT 43.935 181.805 49.280 182.575 ;
        RECT 49.455 181.805 631.270 182.575 ;
        RECT 42.470 181.635 631.270 181.805 ;
        RECT 42.555 180.885 43.765 181.635 ;
        RECT 42.555 180.345 43.075 180.885 ;
        RECT 43.935 180.865 49.280 181.635 ;
        RECT 49.455 180.865 631.270 181.635 ;
        RECT 43.245 180.175 43.765 180.715 ;
        RECT 43.935 180.345 46.515 180.865 ;
        RECT 46.685 180.175 49.280 180.695 ;
        RECT 49.455 180.345 52.035 180.865 ;
        RECT 54.000 180.695 631.270 180.865 ;
        RECT 52.205 180.175 631.270 180.695 ;
        RECT 42.555 179.085 43.765 180.175 ;
        RECT 43.935 179.085 49.280 180.175 ;
        RECT 49.455 179.085 631.270 180.175 ;
        RECT 42.470 178.915 631.270 179.085 ;
        RECT 42.555 177.825 43.765 178.915 ;
        RECT 43.935 177.825 49.280 178.915 ;
        RECT 49.455 177.825 631.270 178.915 ;
        RECT 42.555 177.115 43.075 177.655 ;
        RECT 43.245 177.285 43.765 177.825 ;
        RECT 43.935 177.135 46.515 177.655 ;
        RECT 46.685 177.305 49.280 177.825 ;
        RECT 49.455 177.135 52.035 177.655 ;
        RECT 52.205 177.305 631.270 177.825 ;
        RECT 54.000 177.135 631.270 177.305 ;
        RECT 42.555 176.365 43.765 177.115 ;
        RECT 43.935 176.365 49.280 177.135 ;
        RECT 49.455 176.365 631.270 177.135 ;
        RECT 42.470 176.195 631.270 176.365 ;
        RECT 42.555 175.445 43.765 176.195 ;
        RECT 42.555 174.905 43.075 175.445 ;
        RECT 43.935 175.425 49.280 176.195 ;
        RECT 49.455 175.425 631.270 176.195 ;
        RECT 43.245 174.735 43.765 175.275 ;
        RECT 43.935 174.905 46.515 175.425 ;
        RECT 46.685 174.735 49.280 175.255 ;
        RECT 49.455 174.905 52.035 175.425 ;
        RECT 54.000 175.255 631.270 175.425 ;
        RECT 52.205 174.735 631.270 175.255 ;
        RECT 42.555 173.645 43.765 174.735 ;
        RECT 43.935 173.645 49.280 174.735 ;
        RECT 49.455 173.645 631.270 174.735 ;
        RECT 42.470 173.475 631.270 173.645 ;
        RECT 42.555 172.385 43.765 173.475 ;
        RECT 43.935 172.385 49.280 173.475 ;
        RECT 49.455 172.385 631.270 173.475 ;
        RECT 42.555 171.675 43.075 172.215 ;
        RECT 43.245 171.845 43.765 172.385 ;
        RECT 43.935 171.695 46.515 172.215 ;
        RECT 46.685 171.865 49.280 172.385 ;
        RECT 49.455 171.695 52.035 172.215 ;
        RECT 52.205 171.865 631.270 172.385 ;
        RECT 54.000 171.695 631.270 171.865 ;
        RECT 42.555 170.925 43.765 171.675 ;
        RECT 43.935 170.925 49.280 171.695 ;
        RECT 49.455 170.925 631.270 171.695 ;
        RECT 42.470 170.755 631.270 170.925 ;
        RECT 42.555 170.005 43.765 170.755 ;
        RECT 42.555 169.465 43.075 170.005 ;
        RECT 43.935 169.985 49.280 170.755 ;
        RECT 49.455 169.985 631.270 170.755 ;
        RECT 43.245 169.295 43.765 169.835 ;
        RECT 43.935 169.465 46.515 169.985 ;
        RECT 46.685 169.295 49.280 169.815 ;
        RECT 49.455 169.465 52.035 169.985 ;
        RECT 54.000 169.815 631.270 169.985 ;
        RECT 52.205 169.295 631.270 169.815 ;
        RECT 42.555 168.205 43.765 169.295 ;
        RECT 43.935 168.205 49.280 169.295 ;
        RECT 49.455 168.205 631.270 169.295 ;
        RECT 42.470 168.035 631.270 168.205 ;
        RECT 42.555 166.945 43.765 168.035 ;
        RECT 43.935 166.945 49.280 168.035 ;
        RECT 49.455 166.945 631.270 168.035 ;
        RECT 42.555 166.235 43.075 166.775 ;
        RECT 43.245 166.405 43.765 166.945 ;
        RECT 43.935 166.255 46.515 166.775 ;
        RECT 46.685 166.425 49.280 166.945 ;
        RECT 49.455 166.255 52.035 166.775 ;
        RECT 52.205 166.425 631.270 166.945 ;
        RECT 54.000 166.255 631.270 166.425 ;
        RECT 42.555 165.485 43.765 166.235 ;
        RECT 43.935 165.485 49.280 166.255 ;
        RECT 49.455 165.485 631.270 166.255 ;
        RECT 42.470 165.315 631.270 165.485 ;
        RECT 42.555 164.565 43.765 165.315 ;
        RECT 42.555 164.025 43.075 164.565 ;
        RECT 43.935 164.545 49.280 165.315 ;
        RECT 49.455 164.545 631.270 165.315 ;
        RECT 43.245 163.855 43.765 164.395 ;
        RECT 43.935 164.025 46.515 164.545 ;
        RECT 46.685 163.855 49.280 164.375 ;
        RECT 49.455 164.025 52.035 164.545 ;
        RECT 54.000 164.375 631.270 164.545 ;
        RECT 52.205 163.855 631.270 164.375 ;
        RECT 42.555 162.765 43.765 163.855 ;
        RECT 43.935 162.765 49.280 163.855 ;
        RECT 49.455 162.765 631.270 163.855 ;
        RECT 42.470 162.595 631.270 162.765 ;
        RECT 42.555 161.505 43.765 162.595 ;
        RECT 43.935 161.505 49.280 162.595 ;
        RECT 49.455 161.505 631.270 162.595 ;
        RECT 42.555 160.795 43.075 161.335 ;
        RECT 43.245 160.965 43.765 161.505 ;
        RECT 43.935 160.815 46.515 161.335 ;
        RECT 46.685 160.985 49.280 161.505 ;
        RECT 49.455 160.815 52.035 161.335 ;
        RECT 52.205 160.985 631.270 161.505 ;
        RECT 54.000 160.815 631.270 160.985 ;
        RECT 42.555 160.045 43.765 160.795 ;
        RECT 43.935 160.045 49.280 160.815 ;
        RECT 49.455 160.045 631.270 160.815 ;
        RECT 42.470 159.875 631.270 160.045 ;
        RECT 42.555 159.125 43.765 159.875 ;
        RECT 42.555 158.585 43.075 159.125 ;
        RECT 43.935 159.105 49.280 159.875 ;
        RECT 49.455 159.105 631.270 159.875 ;
        RECT 43.245 158.415 43.765 158.955 ;
        RECT 43.935 158.585 46.515 159.105 ;
        RECT 46.685 158.415 49.280 158.935 ;
        RECT 49.455 158.585 52.035 159.105 ;
        RECT 54.000 158.935 631.270 159.105 ;
        RECT 52.205 158.415 631.270 158.935 ;
        RECT 42.555 157.325 43.765 158.415 ;
        RECT 43.935 157.325 49.280 158.415 ;
        RECT 49.455 157.325 631.270 158.415 ;
        RECT 42.470 157.155 631.270 157.325 ;
        RECT 42.555 156.065 43.765 157.155 ;
        RECT 43.935 156.065 49.280 157.155 ;
        RECT 49.455 156.065 631.270 157.155 ;
        RECT 42.555 155.355 43.075 155.895 ;
        RECT 43.245 155.525 43.765 156.065 ;
        RECT 43.935 155.375 46.515 155.895 ;
        RECT 46.685 155.545 49.280 156.065 ;
        RECT 49.455 155.375 52.035 155.895 ;
        RECT 52.205 155.545 631.270 156.065 ;
        RECT 54.000 155.375 631.270 155.545 ;
        RECT 42.555 154.605 43.765 155.355 ;
        RECT 43.935 154.605 49.280 155.375 ;
        RECT 49.455 154.605 631.270 155.375 ;
        RECT 42.470 154.435 631.270 154.605 ;
        RECT 42.555 153.685 43.765 154.435 ;
        RECT 42.555 153.145 43.075 153.685 ;
        RECT 43.935 153.665 49.280 154.435 ;
        RECT 49.455 153.665 631.270 154.435 ;
        RECT 43.245 152.975 43.765 153.515 ;
        RECT 43.935 153.145 46.515 153.665 ;
        RECT 46.685 152.975 49.280 153.495 ;
        RECT 49.455 153.145 52.035 153.665 ;
        RECT 54.000 153.495 631.270 153.665 ;
        RECT 52.205 152.975 631.270 153.495 ;
        RECT 42.555 151.885 43.765 152.975 ;
        RECT 43.935 151.885 49.280 152.975 ;
        RECT 49.455 151.885 631.270 152.975 ;
        RECT 42.470 151.715 631.270 151.885 ;
        RECT 42.555 150.625 43.765 151.715 ;
        RECT 43.935 150.625 49.280 151.715 ;
        RECT 49.455 150.625 631.270 151.715 ;
        RECT 42.555 149.915 43.075 150.455 ;
        RECT 43.245 150.085 43.765 150.625 ;
        RECT 43.935 149.935 46.515 150.455 ;
        RECT 46.685 150.105 49.280 150.625 ;
        RECT 49.455 149.935 52.035 150.455 ;
        RECT 52.205 150.105 631.270 150.625 ;
        RECT 54.000 149.935 631.270 150.105 ;
        RECT 42.555 149.165 43.765 149.915 ;
        RECT 43.935 149.165 49.280 149.935 ;
        RECT 49.455 149.165 631.270 149.935 ;
        RECT 42.470 148.995 631.270 149.165 ;
        RECT 42.555 148.245 43.765 148.995 ;
        RECT 42.555 147.705 43.075 148.245 ;
        RECT 43.935 148.225 49.280 148.995 ;
        RECT 49.455 148.225 631.270 148.995 ;
        RECT 43.245 147.535 43.765 148.075 ;
        RECT 43.935 147.705 46.515 148.225 ;
        RECT 46.685 147.535 49.280 148.055 ;
        RECT 49.455 147.705 52.035 148.225 ;
        RECT 54.000 148.055 631.270 148.225 ;
        RECT 52.205 147.535 631.270 148.055 ;
        RECT 42.555 146.445 43.765 147.535 ;
        RECT 43.935 146.445 49.280 147.535 ;
        RECT 49.455 146.445 631.270 147.535 ;
        RECT 42.470 146.275 631.270 146.445 ;
        RECT 42.555 145.185 43.765 146.275 ;
        RECT 43.935 145.185 49.280 146.275 ;
        RECT 49.455 145.185 631.270 146.275 ;
        RECT 42.555 144.475 43.075 145.015 ;
        RECT 43.245 144.645 43.765 145.185 ;
        RECT 43.935 144.495 46.515 145.015 ;
        RECT 46.685 144.665 49.280 145.185 ;
        RECT 49.455 144.495 52.035 145.015 ;
        RECT 52.205 144.665 631.270 145.185 ;
        RECT 54.000 144.495 631.270 144.665 ;
        RECT 42.555 143.725 43.765 144.475 ;
        RECT 43.935 143.725 49.280 144.495 ;
        RECT 49.455 143.725 631.270 144.495 ;
        RECT 42.470 143.555 631.270 143.725 ;
        RECT 42.555 142.805 43.765 143.555 ;
        RECT 42.555 142.265 43.075 142.805 ;
        RECT 43.935 142.785 49.280 143.555 ;
        RECT 49.455 142.785 631.270 143.555 ;
        RECT 43.245 142.095 43.765 142.635 ;
        RECT 43.935 142.265 46.515 142.785 ;
        RECT 46.685 142.095 49.280 142.615 ;
        RECT 49.455 142.265 52.035 142.785 ;
        RECT 54.000 142.615 631.270 142.785 ;
        RECT 52.205 142.095 631.270 142.615 ;
        RECT 42.555 141.005 43.765 142.095 ;
        RECT 43.935 141.005 49.280 142.095 ;
        RECT 49.455 141.005 631.270 142.095 ;
        RECT 42.470 140.835 631.270 141.005 ;
        RECT 42.555 139.745 43.765 140.835 ;
        RECT 43.935 139.745 49.280 140.835 ;
        RECT 49.455 139.745 631.270 140.835 ;
        RECT 42.555 139.035 43.075 139.575 ;
        RECT 43.245 139.205 43.765 139.745 ;
        RECT 43.935 139.055 46.515 139.575 ;
        RECT 46.685 139.225 49.280 139.745 ;
        RECT 49.455 139.055 52.035 139.575 ;
        RECT 52.205 139.225 631.270 139.745 ;
        RECT 54.000 139.055 631.270 139.225 ;
        RECT 42.555 138.285 43.765 139.035 ;
        RECT 43.935 138.285 49.280 139.055 ;
        RECT 49.455 138.285 631.270 139.055 ;
        RECT 42.470 138.115 631.270 138.285 ;
        RECT 42.555 137.365 43.765 138.115 ;
        RECT 42.555 136.825 43.075 137.365 ;
        RECT 43.935 137.345 49.280 138.115 ;
        RECT 49.455 137.345 631.270 138.115 ;
        RECT 43.245 136.655 43.765 137.195 ;
        RECT 43.935 136.825 46.515 137.345 ;
        RECT 46.685 136.655 49.280 137.175 ;
        RECT 49.455 136.825 52.035 137.345 ;
        RECT 54.000 137.175 631.270 137.345 ;
        RECT 52.205 136.655 631.270 137.175 ;
        RECT 42.555 135.565 43.765 136.655 ;
        RECT 43.935 135.565 49.280 136.655 ;
        RECT 49.455 135.565 631.270 136.655 ;
        RECT 42.470 135.395 631.270 135.565 ;
        RECT 42.555 134.305 43.765 135.395 ;
        RECT 43.935 134.305 49.280 135.395 ;
        RECT 49.455 134.305 631.270 135.395 ;
        RECT 42.555 133.595 43.075 134.135 ;
        RECT 43.245 133.765 43.765 134.305 ;
        RECT 43.935 133.615 46.515 134.135 ;
        RECT 46.685 133.785 49.280 134.305 ;
        RECT 49.455 133.615 52.035 134.135 ;
        RECT 52.205 133.785 631.270 134.305 ;
        RECT 54.000 133.615 631.270 133.785 ;
        RECT 42.555 132.845 43.765 133.595 ;
        RECT 43.935 132.845 49.280 133.615 ;
        RECT 49.455 132.845 631.270 133.615 ;
        RECT 42.470 132.675 631.270 132.845 ;
        RECT 42.555 131.925 43.765 132.675 ;
        RECT 42.555 131.385 43.075 131.925 ;
        RECT 43.935 131.905 49.280 132.675 ;
        RECT 49.455 131.905 631.270 132.675 ;
        RECT 43.245 131.215 43.765 131.755 ;
        RECT 43.935 131.385 46.515 131.905 ;
        RECT 46.685 131.215 49.280 131.735 ;
        RECT 49.455 131.385 52.035 131.905 ;
        RECT 54.000 131.735 631.270 131.905 ;
        RECT 52.205 131.215 631.270 131.735 ;
        RECT 42.555 130.125 43.765 131.215 ;
        RECT 43.935 130.125 49.280 131.215 ;
        RECT 49.455 130.125 631.270 131.215 ;
        RECT 42.470 129.955 631.270 130.125 ;
        RECT 42.555 128.865 43.765 129.955 ;
        RECT 43.935 128.865 49.280 129.955 ;
        RECT 49.455 128.865 631.270 129.955 ;
        RECT 42.555 128.155 43.075 128.695 ;
        RECT 43.245 128.325 43.765 128.865 ;
        RECT 43.935 128.175 46.515 128.695 ;
        RECT 46.685 128.345 49.280 128.865 ;
        RECT 49.455 128.175 52.035 128.695 ;
        RECT 52.205 128.345 631.270 128.865 ;
        RECT 54.000 128.175 631.270 128.345 ;
        RECT 42.555 127.405 43.765 128.155 ;
        RECT 43.935 127.405 49.280 128.175 ;
        RECT 49.455 127.405 631.270 128.175 ;
        RECT 42.470 127.235 631.270 127.405 ;
        RECT 42.555 126.485 43.765 127.235 ;
        RECT 42.555 125.945 43.075 126.485 ;
        RECT 43.935 126.465 49.280 127.235 ;
        RECT 49.455 126.465 631.270 127.235 ;
        RECT 43.245 125.775 43.765 126.315 ;
        RECT 43.935 125.945 46.515 126.465 ;
        RECT 46.685 125.775 49.280 126.295 ;
        RECT 49.455 125.945 52.035 126.465 ;
        RECT 54.000 126.295 631.270 126.465 ;
        RECT 52.205 125.775 631.270 126.295 ;
        RECT 42.555 124.685 43.765 125.775 ;
        RECT 43.935 124.685 49.280 125.775 ;
        RECT 49.455 124.685 631.270 125.775 ;
        RECT 42.470 124.515 631.270 124.685 ;
        RECT 42.555 123.425 43.765 124.515 ;
        RECT 43.935 123.425 49.280 124.515 ;
        RECT 49.455 123.425 631.270 124.515 ;
        RECT 42.555 122.715 43.075 123.255 ;
        RECT 43.245 122.885 43.765 123.425 ;
        RECT 43.935 122.735 46.515 123.255 ;
        RECT 46.685 122.905 49.280 123.425 ;
        RECT 49.455 122.735 52.035 123.255 ;
        RECT 52.205 122.905 631.270 123.425 ;
        RECT 54.000 122.735 631.270 122.905 ;
        RECT 42.555 121.965 43.765 122.715 ;
        RECT 43.935 121.965 49.280 122.735 ;
        RECT 49.455 121.965 631.270 122.735 ;
        RECT 42.470 121.795 631.270 121.965 ;
        RECT 42.555 121.045 43.765 121.795 ;
        RECT 42.555 120.505 43.075 121.045 ;
        RECT 43.935 121.025 49.280 121.795 ;
        RECT 49.455 121.025 631.270 121.795 ;
        RECT 43.245 120.335 43.765 120.875 ;
        RECT 43.935 120.505 46.515 121.025 ;
        RECT 46.685 120.335 49.280 120.855 ;
        RECT 49.455 120.505 52.035 121.025 ;
        RECT 54.000 120.855 631.270 121.025 ;
        RECT 52.205 120.335 631.270 120.855 ;
        RECT 42.555 119.245 43.765 120.335 ;
        RECT 43.935 119.245 49.280 120.335 ;
        RECT 49.455 119.245 631.270 120.335 ;
        RECT 42.470 119.075 631.270 119.245 ;
        RECT 42.555 117.985 43.765 119.075 ;
        RECT 43.935 117.985 49.280 119.075 ;
        RECT 49.455 117.985 631.270 119.075 ;
        RECT 42.555 117.275 43.075 117.815 ;
        RECT 43.245 117.445 43.765 117.985 ;
        RECT 43.935 117.295 46.515 117.815 ;
        RECT 46.685 117.465 49.280 117.985 ;
        RECT 49.455 117.295 52.035 117.815 ;
        RECT 52.205 117.465 631.270 117.985 ;
        RECT 54.000 117.295 631.270 117.465 ;
        RECT 42.555 116.525 43.765 117.275 ;
        RECT 43.935 116.525 49.280 117.295 ;
        RECT 49.455 116.525 631.270 117.295 ;
        RECT 42.470 116.355 631.270 116.525 ;
        RECT 42.555 115.605 43.765 116.355 ;
        RECT 42.555 115.065 43.075 115.605 ;
        RECT 43.935 115.585 49.280 116.355 ;
        RECT 49.455 115.585 631.270 116.355 ;
        RECT 43.245 114.895 43.765 115.435 ;
        RECT 43.935 115.065 46.515 115.585 ;
        RECT 46.685 114.895 49.280 115.415 ;
        RECT 49.455 115.065 52.035 115.585 ;
        RECT 54.000 115.415 631.270 115.585 ;
        RECT 52.205 114.895 631.270 115.415 ;
        RECT 42.555 113.805 43.765 114.895 ;
        RECT 43.935 113.805 49.280 114.895 ;
        RECT 49.455 113.805 631.270 114.895 ;
        RECT 42.470 113.635 631.270 113.805 ;
        RECT 42.555 112.545 43.765 113.635 ;
        RECT 43.935 112.545 49.280 113.635 ;
        RECT 49.455 112.545 631.270 113.635 ;
        RECT 42.555 111.835 43.075 112.375 ;
        RECT 43.245 112.005 43.765 112.545 ;
        RECT 43.935 111.855 46.515 112.375 ;
        RECT 46.685 112.025 49.280 112.545 ;
        RECT 49.455 111.855 52.035 112.375 ;
        RECT 52.205 112.025 631.270 112.545 ;
        RECT 54.000 111.855 631.270 112.025 ;
        RECT 42.555 111.085 43.765 111.835 ;
        RECT 43.935 111.085 49.280 111.855 ;
        RECT 49.455 111.085 631.270 111.855 ;
        RECT 42.470 110.915 631.270 111.085 ;
        RECT 42.555 110.165 43.765 110.915 ;
        RECT 42.555 109.625 43.075 110.165 ;
        RECT 43.935 110.145 49.280 110.915 ;
        RECT 49.455 110.145 631.270 110.915 ;
        RECT 43.245 109.455 43.765 109.995 ;
        RECT 43.935 109.625 46.515 110.145 ;
        RECT 46.685 109.455 49.280 109.975 ;
        RECT 49.455 109.625 52.035 110.145 ;
        RECT 54.000 109.975 631.270 110.145 ;
        RECT 52.205 109.455 631.270 109.975 ;
        RECT 42.555 108.365 43.765 109.455 ;
        RECT 43.935 108.365 49.280 109.455 ;
        RECT 49.455 108.365 631.270 109.455 ;
        RECT 42.470 108.195 631.270 108.365 ;
        RECT 42.555 107.105 43.765 108.195 ;
        RECT 43.935 107.105 49.280 108.195 ;
        RECT 49.455 107.105 631.270 108.195 ;
        RECT 42.555 106.395 43.075 106.935 ;
        RECT 43.245 106.565 43.765 107.105 ;
        RECT 43.935 106.415 46.515 106.935 ;
        RECT 46.685 106.585 49.280 107.105 ;
        RECT 49.455 106.415 52.035 106.935 ;
        RECT 52.205 106.585 631.270 107.105 ;
        RECT 54.000 106.415 631.270 106.585 ;
        RECT 42.555 105.645 43.765 106.395 ;
        RECT 43.935 105.645 49.280 106.415 ;
        RECT 49.455 105.645 631.270 106.415 ;
        RECT 42.470 105.475 631.270 105.645 ;
        RECT 42.555 104.725 43.765 105.475 ;
        RECT 42.555 104.185 43.075 104.725 ;
        RECT 43.935 104.705 49.280 105.475 ;
        RECT 49.455 104.705 631.270 105.475 ;
        RECT 43.245 104.015 43.765 104.555 ;
        RECT 43.935 104.185 46.515 104.705 ;
        RECT 46.685 104.015 49.280 104.535 ;
        RECT 49.455 104.185 52.035 104.705 ;
        RECT 54.000 104.535 631.270 104.705 ;
        RECT 52.205 104.015 631.270 104.535 ;
        RECT 42.555 102.925 43.765 104.015 ;
        RECT 43.935 102.925 49.280 104.015 ;
        RECT 49.455 102.925 631.270 104.015 ;
        RECT 42.470 102.755 631.270 102.925 ;
        RECT 42.555 101.665 43.765 102.755 ;
        RECT 43.935 101.665 49.280 102.755 ;
        RECT 49.455 101.665 631.270 102.755 ;
        RECT 42.555 100.955 43.075 101.495 ;
        RECT 43.245 101.125 43.765 101.665 ;
        RECT 43.935 100.975 46.515 101.495 ;
        RECT 46.685 101.145 49.280 101.665 ;
        RECT 49.455 100.975 52.035 101.495 ;
        RECT 52.205 101.145 631.270 101.665 ;
        RECT 54.000 100.975 631.270 101.145 ;
        RECT 42.555 100.205 43.765 100.955 ;
        RECT 43.935 100.205 49.280 100.975 ;
        RECT 49.455 100.205 631.270 100.975 ;
        RECT 42.470 100.035 631.270 100.205 ;
        RECT 42.555 99.285 43.765 100.035 ;
        RECT 42.555 98.745 43.075 99.285 ;
        RECT 43.935 99.265 49.280 100.035 ;
        RECT 49.455 99.265 631.270 100.035 ;
        RECT 43.245 98.575 43.765 99.115 ;
        RECT 43.935 98.745 46.515 99.265 ;
        RECT 46.685 98.575 49.280 99.095 ;
        RECT 49.455 98.745 52.035 99.265 ;
        RECT 54.000 99.095 631.270 99.265 ;
        RECT 52.205 98.575 631.270 99.095 ;
        RECT 42.555 97.485 43.765 98.575 ;
        RECT 43.935 97.485 49.280 98.575 ;
        RECT 49.455 97.485 631.270 98.575 ;
        RECT 42.470 97.315 631.270 97.485 ;
        RECT 42.555 96.225 43.765 97.315 ;
        RECT 43.935 96.225 49.280 97.315 ;
        RECT 49.455 96.225 631.270 97.315 ;
        RECT 42.555 95.515 43.075 96.055 ;
        RECT 43.245 95.685 43.765 96.225 ;
        RECT 43.935 95.535 46.515 96.055 ;
        RECT 46.685 95.705 49.280 96.225 ;
        RECT 49.455 95.535 52.035 96.055 ;
        RECT 52.205 95.705 631.270 96.225 ;
        RECT 54.000 95.535 631.270 95.705 ;
        RECT 42.555 94.765 43.765 95.515 ;
        RECT 43.935 94.765 49.280 95.535 ;
        RECT 49.455 94.765 631.270 95.535 ;
        RECT 42.470 94.595 631.270 94.765 ;
        RECT 42.555 93.845 43.765 94.595 ;
        RECT 42.555 93.305 43.075 93.845 ;
        RECT 43.935 93.825 49.280 94.595 ;
        RECT 49.455 93.825 631.270 94.595 ;
        RECT 43.245 93.135 43.765 93.675 ;
        RECT 43.935 93.305 46.515 93.825 ;
        RECT 46.685 93.135 49.280 93.655 ;
        RECT 49.455 93.305 52.035 93.825 ;
        RECT 54.000 93.655 631.270 93.825 ;
        RECT 52.205 93.135 631.270 93.655 ;
        RECT 42.555 92.045 43.765 93.135 ;
        RECT 43.935 92.045 49.280 93.135 ;
        RECT 49.455 92.045 631.270 93.135 ;
        RECT 42.470 91.875 631.270 92.045 ;
        RECT 42.555 90.785 43.765 91.875 ;
        RECT 43.935 90.785 49.280 91.875 ;
        RECT 49.455 90.785 631.270 91.875 ;
        RECT 42.555 90.075 43.075 90.615 ;
        RECT 43.245 90.245 43.765 90.785 ;
        RECT 43.935 90.095 46.515 90.615 ;
        RECT 46.685 90.265 49.280 90.785 ;
        RECT 49.455 90.095 52.035 90.615 ;
        RECT 52.205 90.265 631.270 90.785 ;
        RECT 54.000 90.095 631.270 90.265 ;
        RECT 42.555 89.325 43.765 90.075 ;
        RECT 43.935 89.325 49.280 90.095 ;
        RECT 49.455 89.325 631.270 90.095 ;
        RECT 42.470 89.155 631.270 89.325 ;
        RECT 42.555 88.405 43.765 89.155 ;
        RECT 42.555 87.865 43.075 88.405 ;
        RECT 43.935 88.385 49.280 89.155 ;
        RECT 49.455 88.385 631.270 89.155 ;
        RECT 43.245 87.695 43.765 88.235 ;
        RECT 43.935 87.865 46.515 88.385 ;
        RECT 46.685 87.695 49.280 88.215 ;
        RECT 49.455 87.865 52.035 88.385 ;
        RECT 54.000 88.215 631.270 88.385 ;
        RECT 52.205 87.695 631.270 88.215 ;
        RECT 42.555 86.605 43.765 87.695 ;
        RECT 43.935 86.605 49.280 87.695 ;
        RECT 49.455 86.605 631.270 87.695 ;
        RECT 42.470 86.435 631.270 86.605 ;
        RECT 42.555 85.345 43.765 86.435 ;
        RECT 43.935 85.345 49.280 86.435 ;
        RECT 49.455 85.345 631.270 86.435 ;
        RECT 42.555 84.635 43.075 85.175 ;
        RECT 43.245 84.805 43.765 85.345 ;
        RECT 43.935 84.655 46.515 85.175 ;
        RECT 46.685 84.825 49.280 85.345 ;
        RECT 49.455 84.655 52.035 85.175 ;
        RECT 52.205 84.825 631.270 85.345 ;
        RECT 54.000 84.655 631.270 84.825 ;
        RECT 42.555 83.885 43.765 84.635 ;
        RECT 43.935 83.885 49.280 84.655 ;
        RECT 49.455 83.885 631.270 84.655 ;
        RECT 42.470 83.715 631.270 83.885 ;
        RECT 42.555 82.965 43.765 83.715 ;
        RECT 42.555 82.425 43.075 82.965 ;
        RECT 43.935 82.945 49.280 83.715 ;
        RECT 49.455 82.945 631.270 83.715 ;
        RECT 43.245 82.255 43.765 82.795 ;
        RECT 43.935 82.425 46.515 82.945 ;
        RECT 46.685 82.255 49.280 82.775 ;
        RECT 49.455 82.425 52.035 82.945 ;
        RECT 54.000 82.775 631.270 82.945 ;
        RECT 52.205 82.255 631.270 82.775 ;
        RECT 42.555 81.165 43.765 82.255 ;
        RECT 43.935 81.165 49.280 82.255 ;
        RECT 49.455 81.165 631.270 82.255 ;
        RECT 42.470 80.995 631.270 81.165 ;
        RECT 42.555 79.905 43.765 80.995 ;
        RECT 43.935 79.905 49.280 80.995 ;
        RECT 49.455 79.905 631.270 80.995 ;
        RECT 42.555 79.195 43.075 79.735 ;
        RECT 43.245 79.365 43.765 79.905 ;
        RECT 43.935 79.215 46.515 79.735 ;
        RECT 46.685 79.385 49.280 79.905 ;
        RECT 49.455 79.215 52.035 79.735 ;
        RECT 52.205 79.385 631.270 79.905 ;
        RECT 54.000 79.215 631.270 79.385 ;
        RECT 42.555 78.445 43.765 79.195 ;
        RECT 43.935 78.445 49.280 79.215 ;
        RECT 49.455 78.445 631.270 79.215 ;
        RECT 42.470 78.275 631.270 78.445 ;
        RECT 42.555 77.525 43.765 78.275 ;
        RECT 42.555 76.985 43.075 77.525 ;
        RECT 43.935 77.505 49.280 78.275 ;
        RECT 49.455 77.505 631.270 78.275 ;
        RECT 43.245 76.815 43.765 77.355 ;
        RECT 43.935 76.985 46.515 77.505 ;
        RECT 46.685 76.815 49.280 77.335 ;
        RECT 49.455 76.985 52.035 77.505 ;
        RECT 54.000 77.335 631.270 77.505 ;
        RECT 52.205 76.815 631.270 77.335 ;
        RECT 42.555 75.725 43.765 76.815 ;
        RECT 43.935 75.725 49.280 76.815 ;
        RECT 49.455 75.725 631.270 76.815 ;
        RECT 42.470 75.555 631.270 75.725 ;
        RECT 42.555 74.465 43.765 75.555 ;
        RECT 43.935 74.465 49.280 75.555 ;
        RECT 49.455 74.465 631.270 75.555 ;
        RECT 42.555 73.755 43.075 74.295 ;
        RECT 43.245 73.925 43.765 74.465 ;
        RECT 43.935 73.775 46.515 74.295 ;
        RECT 46.685 73.945 49.280 74.465 ;
        RECT 49.455 73.775 52.035 74.295 ;
        RECT 52.205 73.945 631.270 74.465 ;
        RECT 54.000 73.775 631.270 73.945 ;
        RECT 42.555 73.005 43.765 73.755 ;
        RECT 43.935 73.005 49.280 73.775 ;
        RECT 49.455 73.005 631.270 73.775 ;
        RECT 42.470 72.835 631.270 73.005 ;
        RECT 42.555 72.085 43.765 72.835 ;
        RECT 42.555 71.545 43.075 72.085 ;
        RECT 43.935 72.065 49.280 72.835 ;
        RECT 49.455 72.065 631.270 72.835 ;
        RECT 43.245 71.375 43.765 71.915 ;
        RECT 43.935 71.545 46.515 72.065 ;
        RECT 46.685 71.375 49.280 71.895 ;
        RECT 49.455 71.545 52.035 72.065 ;
        RECT 54.000 71.895 631.270 72.065 ;
        RECT 52.205 71.375 631.270 71.895 ;
        RECT 42.555 70.285 43.765 71.375 ;
        RECT 43.935 70.285 49.280 71.375 ;
        RECT 49.455 70.285 631.270 71.375 ;
        RECT 42.470 70.115 631.270 70.285 ;
        RECT 42.555 69.025 43.765 70.115 ;
        RECT 43.935 69.025 49.280 70.115 ;
        RECT 49.455 69.025 631.270 70.115 ;
        RECT 42.555 68.315 43.075 68.855 ;
        RECT 43.245 68.485 43.765 69.025 ;
        RECT 43.935 68.335 46.515 68.855 ;
        RECT 46.685 68.505 49.280 69.025 ;
        RECT 49.455 68.335 52.035 68.855 ;
        RECT 52.205 68.505 631.270 69.025 ;
        RECT 54.000 68.335 631.270 68.505 ;
        RECT 42.555 67.565 43.765 68.315 ;
        RECT 43.935 67.565 49.280 68.335 ;
        RECT 49.455 67.565 631.270 68.335 ;
        RECT 42.470 67.395 631.270 67.565 ;
        RECT 42.555 66.645 43.765 67.395 ;
        RECT 42.555 66.105 43.075 66.645 ;
        RECT 43.935 66.625 49.280 67.395 ;
        RECT 49.455 66.625 631.270 67.395 ;
        RECT 43.245 65.935 43.765 66.475 ;
        RECT 43.935 66.105 46.515 66.625 ;
        RECT 46.685 65.935 49.280 66.455 ;
        RECT 49.455 66.105 52.035 66.625 ;
        RECT 54.000 66.455 631.270 66.625 ;
        RECT 52.205 65.935 631.270 66.455 ;
        RECT 42.555 64.845 43.765 65.935 ;
        RECT 43.935 64.845 49.280 65.935 ;
        RECT 49.455 64.845 631.270 65.935 ;
        RECT 42.470 64.675 631.270 64.845 ;
        RECT 42.555 63.585 43.765 64.675 ;
        RECT 43.935 63.585 49.280 64.675 ;
        RECT 49.455 63.585 631.270 64.675 ;
        RECT 42.555 62.875 43.075 63.415 ;
        RECT 43.245 63.045 43.765 63.585 ;
        RECT 43.935 62.895 46.515 63.415 ;
        RECT 46.685 63.065 49.280 63.585 ;
        RECT 49.455 62.895 52.035 63.415 ;
        RECT 52.205 63.065 631.270 63.585 ;
        RECT 54.000 62.895 631.270 63.065 ;
        RECT 42.555 62.125 43.765 62.875 ;
        RECT 43.935 62.125 49.280 62.895 ;
        RECT 49.455 62.125 631.270 62.895 ;
        RECT 42.470 61.955 631.270 62.125 ;
        RECT 42.555 61.205 43.765 61.955 ;
        RECT 42.555 60.665 43.075 61.205 ;
        RECT 43.935 61.185 49.280 61.955 ;
        RECT 49.455 61.185 631.270 61.955 ;
        RECT 43.245 60.495 43.765 61.035 ;
        RECT 43.935 60.665 46.515 61.185 ;
        RECT 46.685 60.495 49.280 61.015 ;
        RECT 49.455 60.665 52.035 61.185 ;
        RECT 54.000 61.015 631.270 61.185 ;
        RECT 52.205 60.495 631.270 61.015 ;
        RECT 42.555 59.405 43.765 60.495 ;
        RECT 43.935 59.405 49.280 60.495 ;
        RECT 49.455 59.405 631.270 60.495 ;
        RECT 42.470 59.235 631.270 59.405 ;
        RECT 42.555 58.145 43.765 59.235 ;
        RECT 43.935 58.145 49.280 59.235 ;
        RECT 49.455 58.145 631.270 59.235 ;
        RECT 42.555 57.435 43.075 57.975 ;
        RECT 43.245 57.605 43.765 58.145 ;
        RECT 43.935 57.455 46.515 57.975 ;
        RECT 46.685 57.625 49.280 58.145 ;
        RECT 49.455 57.455 52.035 57.975 ;
        RECT 52.205 57.625 631.270 58.145 ;
        RECT 54.000 57.455 631.270 57.625 ;
        RECT 42.555 56.685 43.765 57.435 ;
        RECT 43.935 56.685 49.280 57.455 ;
        RECT 49.455 56.685 631.270 57.455 ;
        RECT 42.470 56.515 631.270 56.685 ;
        RECT 42.555 55.765 43.765 56.515 ;
        RECT 42.555 55.225 43.075 55.765 ;
        RECT 43.935 55.745 49.280 56.515 ;
        RECT 49.455 55.745 631.270 56.515 ;
        RECT 43.245 55.055 43.765 55.595 ;
        RECT 43.935 55.225 46.515 55.745 ;
        RECT 46.685 55.055 49.280 55.575 ;
        RECT 49.455 55.225 52.035 55.745 ;
        RECT 54.000 55.575 631.270 55.745 ;
        RECT 52.205 55.055 631.270 55.575 ;
        RECT 42.555 53.965 43.765 55.055 ;
        RECT 43.935 53.965 49.280 55.055 ;
        RECT 49.455 54.000 631.270 55.055 ;
        RECT 49.455 53.965 54.800 54.000 ;
        RECT 54.975 53.965 56.645 54.000 ;
        RECT 56.815 53.965 57.105 54.000 ;
        RECT 57.275 53.965 62.620 54.000 ;
        RECT 62.795 53.965 68.140 54.000 ;
        RECT 68.315 53.965 73.660 54.000 ;
        RECT 73.835 53.965 79.180 54.000 ;
        RECT 79.855 53.965 80.085 54.000 ;
        RECT 80.755 53.965 80.965 54.000 ;
        RECT 81.195 53.965 84.705 54.000 ;
        RECT 84.875 53.965 85.165 54.000 ;
        RECT 86.225 53.965 86.555 54.000 ;
        RECT 87.150 53.965 87.415 54.000 ;
        RECT 89.320 53.965 89.490 54.000 ;
        RECT 91.200 53.965 91.415 54.000 ;
        RECT 92.335 53.965 92.515 54.000 ;
        RECT 93.210 53.965 93.380 54.000 ;
        RECT 94.050 53.965 94.220 54.000 ;
        RECT 94.535 53.965 99.880 54.000 ;
        RECT 100.945 53.965 101.275 54.000 ;
        RECT 101.870 53.965 102.135 54.000 ;
        RECT 104.040 53.965 104.210 54.000 ;
        RECT 105.920 53.965 106.135 54.000 ;
        RECT 107.055 53.965 107.235 54.000 ;
        RECT 107.930 53.965 108.100 54.000 ;
        RECT 108.770 53.965 108.940 54.000 ;
        RECT 109.255 53.965 112.765 54.000 ;
        RECT 112.935 53.965 113.225 54.000 ;
        RECT 113.825 53.965 114.155 54.000 ;
        RECT 114.750 53.965 115.015 54.000 ;
        RECT 116.920 53.965 117.090 54.000 ;
        RECT 118.800 53.965 119.015 54.000 ;
        RECT 119.935 53.965 120.115 54.000 ;
        RECT 120.810 53.965 120.980 54.000 ;
        RECT 121.650 53.965 121.820 54.000 ;
        RECT 122.135 53.965 127.480 54.000 ;
        RECT 127.655 53.965 129.325 54.000 ;
        RECT 130.425 53.965 130.675 54.000 ;
        RECT 131.265 53.965 131.515 54.000 ;
        RECT 133.045 53.965 133.295 54.000 ;
        RECT 134.725 53.965 134.975 54.000 ;
        RECT 135.565 53.965 135.815 54.000 ;
        RECT 136.405 53.965 136.655 54.000 ;
        RECT 137.315 53.965 140.825 54.000 ;
        RECT 140.995 53.965 141.285 54.000 ;
        RECT 141.885 53.965 142.215 54.000 ;
        RECT 142.810 53.965 143.075 54.000 ;
        RECT 144.980 53.965 145.150 54.000 ;
        RECT 146.860 53.965 147.075 54.000 ;
        RECT 147.995 53.965 148.175 54.000 ;
        RECT 148.870 53.965 149.040 54.000 ;
        RECT 149.710 53.965 149.880 54.000 ;
        RECT 150.195 53.965 153.705 54.000 ;
        RECT 154.305 53.965 154.635 54.000 ;
        RECT 155.230 53.965 155.495 54.000 ;
        RECT 157.400 53.965 157.570 54.000 ;
        RECT 159.280 53.965 159.495 54.000 ;
        RECT 160.415 53.965 160.595 54.000 ;
        RECT 161.290 53.965 161.460 54.000 ;
        RECT 162.130 53.965 162.300 54.000 ;
        RECT 162.615 53.965 167.960 54.000 ;
        RECT 169.055 53.965 169.345 54.000 ;
        RECT 170.425 53.965 170.755 54.000 ;
        RECT 171.265 53.965 171.515 54.000 ;
        RECT 174.115 53.965 177.625 54.000 ;
        RECT 178.225 53.965 178.555 54.000 ;
        RECT 179.150 53.965 179.415 54.000 ;
        RECT 181.320 53.965 181.490 54.000 ;
        RECT 183.200 53.965 183.415 54.000 ;
        RECT 184.335 53.965 184.515 54.000 ;
        RECT 185.210 53.965 185.380 54.000 ;
        RECT 186.050 53.965 186.220 54.000 ;
        RECT 186.535 53.965 190.045 54.000 ;
        RECT 191.190 53.965 191.360 54.000 ;
        RECT 192.070 53.965 192.240 54.000 ;
        RECT 192.910 53.965 193.080 54.000 ;
        RECT 193.435 53.965 196.945 54.000 ;
        RECT 197.115 53.965 197.405 54.000 ;
        RECT 197.575 53.965 199.245 54.000 ;
        RECT 200.305 53.965 200.635 54.000 ;
        RECT 201.230 53.965 201.495 54.000 ;
        RECT 203.400 53.965 203.570 54.000 ;
        RECT 205.280 53.965 205.495 54.000 ;
        RECT 206.415 53.965 206.595 54.000 ;
        RECT 207.290 53.965 207.460 54.000 ;
        RECT 208.130 53.965 208.300 54.000 ;
        RECT 208.615 53.965 212.125 54.000 ;
        RECT 212.765 53.965 213.015 54.000 ;
        RECT 213.605 53.965 213.855 54.000 ;
        RECT 215.385 53.965 215.635 54.000 ;
        RECT 217.065 53.965 217.315 54.000 ;
        RECT 217.905 53.965 218.155 54.000 ;
        RECT 218.745 53.965 218.995 54.000 ;
        RECT 219.655 53.965 225.000 54.000 ;
        RECT 225.175 53.965 225.465 54.000 ;
        RECT 225.670 53.965 225.955 54.000 ;
        RECT 226.530 53.965 226.860 54.000 ;
        RECT 229.180 53.965 229.460 54.000 ;
        RECT 230.010 53.965 230.340 54.000 ;
        RECT 230.870 53.965 231.200 54.000 ;
        RECT 231.615 53.965 235.125 54.000 ;
        RECT 235.335 53.965 235.565 54.000 ;
        RECT 236.235 53.965 236.445 54.000 ;
        RECT 236.675 53.965 240.185 54.000 ;
        RECT 240.825 53.965 241.075 54.000 ;
        RECT 241.665 53.965 241.915 54.000 ;
        RECT 243.445 53.965 243.695 54.000 ;
        RECT 245.125 53.965 245.375 54.000 ;
        RECT 245.965 53.965 246.215 54.000 ;
        RECT 246.805 53.965 247.055 54.000 ;
        RECT 247.715 53.965 253.060 54.000 ;
        RECT 253.235 53.965 253.525 54.000 ;
        RECT 254.165 53.965 254.415 54.000 ;
        RECT 255.005 53.965 255.255 54.000 ;
        RECT 256.785 53.965 257.035 54.000 ;
        RECT 258.465 53.965 258.715 54.000 ;
        RECT 259.305 53.965 259.555 54.000 ;
        RECT 260.145 53.965 260.395 54.000 ;
        RECT 261.055 53.965 264.565 54.000 ;
        RECT 265.210 53.965 265.540 54.000 ;
        RECT 266.140 53.965 266.400 54.000 ;
        RECT 266.575 53.965 270.085 54.000 ;
        RECT 270.725 53.965 270.975 54.000 ;
        RECT 271.565 53.965 271.815 54.000 ;
        RECT 273.345 53.965 273.595 54.000 ;
        RECT 275.025 53.965 275.275 54.000 ;
        RECT 275.865 53.965 276.115 54.000 ;
        RECT 276.705 53.965 276.955 54.000 ;
        RECT 277.615 53.965 281.125 54.000 ;
        RECT 281.295 53.965 281.585 54.000 ;
        RECT 281.755 53.965 284.345 54.000 ;
        RECT 284.985 53.965 285.235 54.000 ;
        RECT 285.825 53.965 286.075 54.000 ;
        RECT 287.605 53.965 287.855 54.000 ;
        RECT 289.285 53.965 289.535 54.000 ;
        RECT 290.125 53.965 290.375 54.000 ;
        RECT 290.965 53.965 291.215 54.000 ;
        RECT 291.875 53.965 297.220 54.000 ;
        RECT 298.785 53.965 299.035 54.000 ;
        RECT 299.625 53.965 299.875 54.000 ;
        RECT 301.405 53.965 301.655 54.000 ;
        RECT 303.085 53.965 303.335 54.000 ;
        RECT 303.925 53.965 304.175 54.000 ;
        RECT 304.765 53.965 305.015 54.000 ;
        RECT 305.675 53.965 309.185 54.000 ;
        RECT 309.355 53.965 309.645 54.000 ;
        RECT 310.285 53.965 310.535 54.000 ;
        RECT 311.125 53.965 311.375 54.000 ;
        RECT 312.905 53.965 313.155 54.000 ;
        RECT 314.585 53.965 314.835 54.000 ;
        RECT 315.425 53.965 315.675 54.000 ;
        RECT 316.265 53.965 316.515 54.000 ;
        RECT 317.175 53.965 322.520 54.000 ;
        RECT 322.695 53.965 324.365 54.000 ;
        RECT 325.465 53.965 325.715 54.000 ;
        RECT 326.305 53.965 326.555 54.000 ;
        RECT 328.085 53.965 328.335 54.000 ;
        RECT 329.765 53.965 330.015 54.000 ;
        RECT 330.605 53.965 330.855 54.000 ;
        RECT 331.445 53.965 331.695 54.000 ;
        RECT 332.355 53.965 335.865 54.000 ;
        RECT 336.035 53.965 337.245 54.000 ;
        RECT 337.415 53.965 337.705 54.000 ;
        RECT 337.915 53.965 338.145 54.000 ;
        RECT 338.815 53.965 339.025 54.000 ;
        RECT 339.255 53.965 342.765 54.000 ;
        RECT 343.865 53.965 344.115 54.000 ;
        RECT 344.705 53.965 344.955 54.000 ;
        RECT 346.485 53.965 346.735 54.000 ;
        RECT 348.165 53.965 348.415 54.000 ;
        RECT 349.005 53.965 349.255 54.000 ;
        RECT 349.845 53.965 350.095 54.000 ;
        RECT 350.755 53.965 354.265 54.000 ;
        RECT 354.905 53.965 355.155 54.000 ;
        RECT 355.745 53.965 355.995 54.000 ;
        RECT 357.525 53.965 357.775 54.000 ;
        RECT 359.205 53.965 359.455 54.000 ;
        RECT 360.045 53.965 360.295 54.000 ;
        RECT 360.885 53.965 361.135 54.000 ;
        RECT 361.795 53.965 365.305 54.000 ;
        RECT 365.475 53.965 365.765 54.000 ;
        RECT 366.385 53.965 366.715 54.000 ;
        RECT 367.225 53.965 367.475 54.000 ;
        RECT 370.075 53.965 373.585 54.000 ;
        RECT 373.755 53.965 374.965 54.000 ;
        RECT 375.605 53.965 375.855 54.000 ;
        RECT 376.445 53.965 376.695 54.000 ;
        RECT 378.225 53.965 378.475 54.000 ;
        RECT 379.905 53.965 380.155 54.000 ;
        RECT 380.745 53.965 380.995 54.000 ;
        RECT 381.585 53.965 381.835 54.000 ;
        RECT 382.495 53.965 387.840 54.000 ;
        RECT 388.015 53.965 393.360 54.000 ;
        RECT 393.535 53.965 393.825 54.000 ;
        RECT 393.995 53.965 399.340 54.000 ;
        RECT 399.515 53.965 404.860 54.000 ;
        RECT 405.035 53.965 410.380 54.000 ;
        RECT 410.555 53.965 415.900 54.000 ;
        RECT 416.075 53.965 421.420 54.000 ;
        RECT 421.595 53.965 421.885 54.000 ;
        RECT 422.055 53.965 427.400 54.000 ;
        RECT 427.575 53.965 432.920 54.000 ;
        RECT 433.095 53.965 438.440 54.000 ;
        RECT 438.615 53.965 443.960 54.000 ;
        RECT 444.135 53.965 449.480 54.000 ;
        RECT 449.655 53.965 449.945 54.000 ;
        RECT 450.115 53.965 455.460 54.000 ;
        RECT 455.635 53.965 460.980 54.000 ;
        RECT 461.155 53.965 466.500 54.000 ;
        RECT 466.675 53.965 472.020 54.000 ;
        RECT 472.195 53.965 477.540 54.000 ;
        RECT 477.715 53.965 478.005 54.000 ;
        RECT 478.175 53.965 483.520 54.000 ;
        RECT 483.695 53.965 489.040 54.000 ;
        RECT 489.215 53.965 494.560 54.000 ;
        RECT 494.735 53.965 500.080 54.000 ;
        RECT 500.255 53.965 505.600 54.000 ;
        RECT 505.775 53.965 506.065 54.000 ;
        RECT 506.235 53.965 511.580 54.000 ;
        RECT 511.755 53.965 517.100 54.000 ;
        RECT 517.275 53.965 522.620 54.000 ;
        RECT 522.795 53.965 528.140 54.000 ;
        RECT 528.315 53.965 533.660 54.000 ;
        RECT 533.835 53.965 534.125 54.000 ;
        RECT 534.295 53.965 539.640 54.000 ;
        RECT 539.815 53.965 545.160 54.000 ;
        RECT 545.335 53.965 550.680 54.000 ;
        RECT 550.855 53.965 556.200 54.000 ;
        RECT 556.375 53.965 561.720 54.000 ;
        RECT 561.895 53.965 562.185 54.000 ;
        RECT 562.355 53.965 567.700 54.000 ;
        RECT 567.875 53.965 573.220 54.000 ;
        RECT 573.395 53.965 578.740 54.000 ;
        RECT 578.915 53.965 584.260 54.000 ;
        RECT 584.435 53.965 589.780 54.000 ;
        RECT 589.955 53.965 590.245 54.000 ;
        RECT 590.415 53.965 595.760 54.000 ;
        RECT 595.935 53.965 601.280 54.000 ;
        RECT 601.455 53.965 606.800 54.000 ;
        RECT 606.975 53.965 612.320 54.000 ;
        RECT 612.495 53.965 617.840 54.000 ;
        RECT 618.015 53.965 618.305 54.000 ;
        RECT 618.475 53.965 623.820 54.000 ;
        RECT 623.995 53.965 629.340 54.000 ;
        RECT 629.975 53.965 631.185 54.000 ;
        RECT 42.470 53.795 631.270 53.965 ;
        RECT 42.555 52.705 43.765 53.795 ;
        RECT 43.935 52.705 49.280 53.795 ;
        RECT 49.455 52.705 54.800 53.795 ;
        RECT 54.975 52.705 60.320 53.795 ;
        RECT 60.495 52.705 65.840 53.795 ;
        RECT 66.015 52.705 69.525 53.795 ;
        RECT 42.555 51.995 43.075 52.535 ;
        RECT 43.245 52.165 43.765 52.705 ;
        RECT 43.935 52.015 46.515 52.535 ;
        RECT 46.685 52.185 49.280 52.705 ;
        RECT 49.455 52.015 52.035 52.535 ;
        RECT 52.205 52.185 54.800 52.705 ;
        RECT 54.975 52.015 57.555 52.535 ;
        RECT 57.725 52.185 60.320 52.705 ;
        RECT 60.495 52.015 63.075 52.535 ;
        RECT 63.245 52.185 65.840 52.705 ;
        RECT 66.015 52.015 67.665 52.535 ;
        RECT 67.835 52.185 69.525 52.705 ;
        RECT 70.615 52.630 70.905 53.795 ;
        RECT 71.075 52.705 76.420 53.795 ;
        RECT 71.075 52.015 73.655 52.535 ;
        RECT 73.825 52.185 76.420 52.705 ;
        RECT 77.555 52.655 77.785 53.795 ;
        RECT 77.955 52.645 78.285 53.625 ;
        RECT 78.455 52.655 78.665 53.795 ;
        RECT 78.895 52.705 82.405 53.795 ;
        RECT 82.665 53.125 82.835 53.625 ;
        RECT 83.005 53.295 83.335 53.795 ;
        RECT 82.665 52.955 83.330 53.125 ;
        RECT 77.535 52.235 77.865 52.485 ;
        RECT 42.555 51.245 43.765 51.995 ;
        RECT 43.935 51.245 49.280 52.015 ;
        RECT 49.455 51.245 54.800 52.015 ;
        RECT 54.975 51.245 60.320 52.015 ;
        RECT 60.495 51.245 65.840 52.015 ;
        RECT 66.015 51.245 69.525 52.015 ;
        RECT 70.615 51.245 70.905 51.970 ;
        RECT 71.075 51.245 76.420 52.015 ;
        RECT 77.555 51.245 77.785 52.065 ;
        RECT 78.035 52.045 78.285 52.645 ;
        RECT 77.955 51.415 78.285 52.045 ;
        RECT 78.455 51.245 78.665 52.065 ;
        RECT 78.895 52.015 80.545 52.535 ;
        RECT 80.715 52.185 82.405 52.705 ;
        RECT 82.580 52.135 82.930 52.785 ;
        RECT 78.895 51.245 82.405 52.015 ;
        RECT 83.100 51.965 83.330 52.955 ;
        RECT 82.665 51.795 83.330 51.965 ;
        RECT 82.665 51.505 82.835 51.795 ;
        RECT 83.005 51.245 83.335 51.625 ;
        RECT 83.505 51.505 83.730 53.625 ;
        RECT 83.930 53.335 84.195 53.795 ;
        RECT 84.380 53.225 84.615 53.600 ;
        RECT 84.860 53.350 85.930 53.520 ;
        RECT 83.930 52.225 84.210 52.825 ;
        RECT 83.945 51.245 84.195 51.705 ;
        RECT 84.380 51.695 84.550 53.225 ;
        RECT 84.720 52.195 84.960 53.065 ;
        RECT 85.150 52.815 85.590 53.170 ;
        RECT 85.760 52.735 85.930 53.350 ;
        RECT 86.100 52.995 86.270 53.795 ;
        RECT 86.440 53.295 86.690 53.625 ;
        RECT 86.915 53.325 87.800 53.495 ;
        RECT 85.760 52.645 86.270 52.735 ;
        RECT 85.470 52.475 86.270 52.645 ;
        RECT 84.720 51.865 85.300 52.195 ;
        RECT 85.470 51.695 85.640 52.475 ;
        RECT 86.100 52.405 86.270 52.475 ;
        RECT 85.810 52.225 85.980 52.255 ;
        RECT 86.440 52.225 86.610 53.295 ;
        RECT 86.780 52.405 86.970 53.125 ;
        RECT 87.140 52.735 87.460 53.065 ;
        RECT 85.810 51.925 86.610 52.225 ;
        RECT 87.140 52.195 87.330 52.735 ;
        RECT 84.380 51.525 84.710 51.695 ;
        RECT 84.890 51.525 85.640 51.695 ;
        RECT 85.890 51.245 86.260 51.745 ;
        RECT 86.440 51.695 86.610 51.925 ;
        RECT 86.780 51.865 87.330 52.195 ;
        RECT 87.630 52.405 87.800 53.325 ;
        RECT 87.980 53.295 88.195 53.795 ;
        RECT 88.660 52.990 88.830 53.615 ;
        RECT 89.115 53.015 89.295 53.795 ;
        RECT 87.970 52.830 88.830 52.990 ;
        RECT 87.970 52.660 89.080 52.830 ;
        RECT 88.910 52.405 89.080 52.660 ;
        RECT 89.475 52.795 89.810 53.555 ;
        RECT 89.990 52.965 90.160 53.795 ;
        RECT 90.330 52.795 90.660 53.555 ;
        RECT 90.830 52.965 91.000 53.795 ;
        RECT 89.475 52.625 91.145 52.795 ;
        RECT 91.315 52.705 96.660 53.795 ;
        RECT 96.835 52.705 98.505 53.795 ;
        RECT 87.630 52.235 88.720 52.405 ;
        RECT 88.910 52.235 90.730 52.405 ;
        RECT 87.630 51.695 87.800 52.235 ;
        RECT 88.910 52.065 89.080 52.235 ;
        RECT 88.580 51.895 89.080 52.065 ;
        RECT 90.900 52.060 91.145 52.625 ;
        RECT 86.440 51.525 86.900 51.695 ;
        RECT 87.130 51.525 87.800 51.695 ;
        RECT 88.115 51.245 88.285 51.775 ;
        RECT 88.580 51.455 88.940 51.895 ;
        RECT 89.475 51.890 91.145 52.060 ;
        RECT 91.315 52.015 93.895 52.535 ;
        RECT 94.065 52.185 96.660 52.705 ;
        RECT 96.835 52.015 97.585 52.535 ;
        RECT 97.755 52.185 98.505 52.705 ;
        RECT 98.675 52.630 98.965 53.795 ;
        RECT 99.225 53.125 99.395 53.625 ;
        RECT 99.565 53.295 99.895 53.795 ;
        RECT 99.225 52.955 99.890 53.125 ;
        RECT 99.140 52.135 99.490 52.785 ;
        RECT 89.115 51.245 89.285 51.725 ;
        RECT 89.475 51.465 89.810 51.890 ;
        RECT 89.985 51.245 90.155 51.720 ;
        RECT 90.330 51.465 90.665 51.890 ;
        RECT 90.835 51.245 91.005 51.720 ;
        RECT 91.315 51.245 96.660 52.015 ;
        RECT 96.835 51.245 98.505 52.015 ;
        RECT 98.675 51.245 98.965 51.970 ;
        RECT 99.660 51.965 99.890 52.955 ;
        RECT 99.225 51.795 99.890 51.965 ;
        RECT 99.225 51.505 99.395 51.795 ;
        RECT 99.565 51.245 99.895 51.625 ;
        RECT 100.065 51.505 100.290 53.625 ;
        RECT 100.490 53.335 100.755 53.795 ;
        RECT 100.940 53.225 101.175 53.600 ;
        RECT 101.420 53.350 102.490 53.520 ;
        RECT 100.490 52.225 100.770 52.825 ;
        RECT 100.505 51.245 100.755 51.705 ;
        RECT 100.940 51.695 101.110 53.225 ;
        RECT 101.280 52.195 101.520 53.065 ;
        RECT 101.710 52.815 102.150 53.170 ;
        RECT 102.320 52.735 102.490 53.350 ;
        RECT 102.660 52.995 102.830 53.795 ;
        RECT 103.000 53.295 103.250 53.625 ;
        RECT 103.475 53.325 104.360 53.495 ;
        RECT 102.320 52.645 102.830 52.735 ;
        RECT 102.030 52.475 102.830 52.645 ;
        RECT 101.280 51.865 101.860 52.195 ;
        RECT 102.030 51.695 102.200 52.475 ;
        RECT 102.660 52.405 102.830 52.475 ;
        RECT 102.370 52.225 102.540 52.255 ;
        RECT 103.000 52.225 103.170 53.295 ;
        RECT 103.340 52.405 103.530 53.125 ;
        RECT 103.700 52.735 104.020 53.065 ;
        RECT 102.370 51.925 103.170 52.225 ;
        RECT 103.700 52.195 103.890 52.735 ;
        RECT 100.940 51.525 101.270 51.695 ;
        RECT 101.450 51.525 102.200 51.695 ;
        RECT 102.450 51.245 102.820 51.745 ;
        RECT 103.000 51.695 103.170 51.925 ;
        RECT 103.340 51.865 103.890 52.195 ;
        RECT 104.190 52.405 104.360 53.325 ;
        RECT 104.540 53.295 104.755 53.795 ;
        RECT 105.220 52.990 105.390 53.615 ;
        RECT 105.675 53.015 105.855 53.795 ;
        RECT 104.530 52.830 105.390 52.990 ;
        RECT 104.530 52.660 105.640 52.830 ;
        RECT 105.470 52.405 105.640 52.660 ;
        RECT 106.035 52.795 106.370 53.555 ;
        RECT 106.550 52.965 106.720 53.795 ;
        RECT 106.890 52.795 107.220 53.555 ;
        RECT 107.390 52.965 107.560 53.795 ;
        RECT 106.035 52.625 107.705 52.795 ;
        RECT 107.875 52.705 111.385 53.795 ;
        RECT 111.645 53.125 111.815 53.625 ;
        RECT 111.985 53.295 112.315 53.795 ;
        RECT 111.645 52.955 112.310 53.125 ;
        RECT 104.190 52.235 105.280 52.405 ;
        RECT 105.470 52.235 107.290 52.405 ;
        RECT 104.190 51.695 104.360 52.235 ;
        RECT 105.470 52.065 105.640 52.235 ;
        RECT 105.140 51.895 105.640 52.065 ;
        RECT 107.460 52.060 107.705 52.625 ;
        RECT 103.000 51.525 103.460 51.695 ;
        RECT 103.690 51.525 104.360 51.695 ;
        RECT 104.675 51.245 104.845 51.775 ;
        RECT 105.140 51.455 105.500 51.895 ;
        RECT 106.035 51.890 107.705 52.060 ;
        RECT 107.875 52.015 109.525 52.535 ;
        RECT 109.695 52.185 111.385 52.705 ;
        RECT 111.560 52.135 111.910 52.785 ;
        RECT 105.675 51.245 105.845 51.725 ;
        RECT 106.035 51.465 106.370 51.890 ;
        RECT 106.545 51.245 106.715 51.720 ;
        RECT 106.890 51.465 107.225 51.890 ;
        RECT 107.395 51.245 107.565 51.720 ;
        RECT 107.875 51.245 111.385 52.015 ;
        RECT 112.080 51.965 112.310 52.955 ;
        RECT 111.645 51.795 112.310 51.965 ;
        RECT 111.645 51.505 111.815 51.795 ;
        RECT 111.985 51.245 112.315 51.625 ;
        RECT 112.485 51.505 112.710 53.625 ;
        RECT 112.910 53.335 113.175 53.795 ;
        RECT 113.360 53.225 113.595 53.600 ;
        RECT 113.840 53.350 114.910 53.520 ;
        RECT 112.910 52.225 113.190 52.825 ;
        RECT 112.925 51.245 113.175 51.705 ;
        RECT 113.360 51.695 113.530 53.225 ;
        RECT 113.700 52.195 113.940 53.065 ;
        RECT 114.130 52.815 114.570 53.170 ;
        RECT 114.740 52.735 114.910 53.350 ;
        RECT 115.080 52.995 115.250 53.795 ;
        RECT 115.420 53.295 115.670 53.625 ;
        RECT 115.895 53.325 116.780 53.495 ;
        RECT 114.740 52.645 115.250 52.735 ;
        RECT 114.450 52.475 115.250 52.645 ;
        RECT 113.700 51.865 114.280 52.195 ;
        RECT 114.450 51.695 114.620 52.475 ;
        RECT 115.080 52.405 115.250 52.475 ;
        RECT 114.790 52.225 114.960 52.255 ;
        RECT 115.420 52.225 115.590 53.295 ;
        RECT 115.760 52.405 115.950 53.125 ;
        RECT 116.120 52.735 116.440 53.065 ;
        RECT 114.790 51.925 115.590 52.225 ;
        RECT 116.120 52.195 116.310 52.735 ;
        RECT 113.360 51.525 113.690 51.695 ;
        RECT 113.870 51.525 114.620 51.695 ;
        RECT 114.870 51.245 115.240 51.745 ;
        RECT 115.420 51.695 115.590 51.925 ;
        RECT 115.760 51.865 116.310 52.195 ;
        RECT 116.610 52.405 116.780 53.325 ;
        RECT 116.960 53.295 117.175 53.795 ;
        RECT 117.640 52.990 117.810 53.615 ;
        RECT 118.095 53.015 118.275 53.795 ;
        RECT 116.950 52.830 117.810 52.990 ;
        RECT 116.950 52.660 118.060 52.830 ;
        RECT 117.890 52.405 118.060 52.660 ;
        RECT 118.455 52.795 118.790 53.555 ;
        RECT 118.970 52.965 119.140 53.795 ;
        RECT 119.310 52.795 119.640 53.555 ;
        RECT 119.810 52.965 119.980 53.795 ;
        RECT 118.455 52.625 120.125 52.795 ;
        RECT 120.295 52.705 125.640 53.795 ;
        RECT 116.610 52.235 117.700 52.405 ;
        RECT 117.890 52.235 119.710 52.405 ;
        RECT 116.610 51.695 116.780 52.235 ;
        RECT 117.890 52.065 118.060 52.235 ;
        RECT 117.560 51.895 118.060 52.065 ;
        RECT 119.880 52.060 120.125 52.625 ;
        RECT 115.420 51.525 115.880 51.695 ;
        RECT 116.110 51.525 116.780 51.695 ;
        RECT 117.095 51.245 117.265 51.775 ;
        RECT 117.560 51.455 117.920 51.895 ;
        RECT 118.455 51.890 120.125 52.060 ;
        RECT 120.295 52.015 122.875 52.535 ;
        RECT 123.045 52.185 125.640 52.705 ;
        RECT 126.735 52.630 127.025 53.795 ;
        RECT 127.285 53.125 127.455 53.625 ;
        RECT 127.625 53.295 127.955 53.795 ;
        RECT 127.285 52.955 127.950 53.125 ;
        RECT 127.200 52.135 127.550 52.785 ;
        RECT 118.095 51.245 118.265 51.725 ;
        RECT 118.455 51.465 118.790 51.890 ;
        RECT 118.965 51.245 119.135 51.720 ;
        RECT 119.310 51.465 119.645 51.890 ;
        RECT 119.815 51.245 119.985 51.720 ;
        RECT 120.295 51.245 125.640 52.015 ;
        RECT 126.735 51.245 127.025 51.970 ;
        RECT 127.720 51.965 127.950 52.955 ;
        RECT 127.285 51.795 127.950 51.965 ;
        RECT 127.285 51.505 127.455 51.795 ;
        RECT 127.625 51.245 127.955 51.625 ;
        RECT 128.125 51.505 128.350 53.625 ;
        RECT 128.550 53.335 128.815 53.795 ;
        RECT 129.000 53.225 129.235 53.600 ;
        RECT 129.480 53.350 130.550 53.520 ;
        RECT 128.550 52.225 128.830 52.825 ;
        RECT 128.565 51.245 128.815 51.705 ;
        RECT 129.000 51.695 129.170 53.225 ;
        RECT 129.340 52.195 129.580 53.065 ;
        RECT 129.770 52.815 130.210 53.170 ;
        RECT 130.380 52.735 130.550 53.350 ;
        RECT 130.720 52.995 130.890 53.795 ;
        RECT 131.060 53.295 131.310 53.625 ;
        RECT 131.535 53.325 132.420 53.495 ;
        RECT 130.380 52.645 130.890 52.735 ;
        RECT 130.090 52.475 130.890 52.645 ;
        RECT 129.340 51.865 129.920 52.195 ;
        RECT 130.090 51.695 130.260 52.475 ;
        RECT 130.720 52.405 130.890 52.475 ;
        RECT 130.430 52.225 130.600 52.255 ;
        RECT 131.060 52.225 131.230 53.295 ;
        RECT 131.400 52.405 131.590 53.125 ;
        RECT 131.760 52.735 132.080 53.065 ;
        RECT 130.430 51.925 131.230 52.225 ;
        RECT 131.760 52.195 131.950 52.735 ;
        RECT 129.000 51.525 129.330 51.695 ;
        RECT 129.510 51.525 130.260 51.695 ;
        RECT 130.510 51.245 130.880 51.745 ;
        RECT 131.060 51.695 131.230 51.925 ;
        RECT 131.400 51.865 131.950 52.195 ;
        RECT 132.250 52.405 132.420 53.325 ;
        RECT 132.600 53.295 132.815 53.795 ;
        RECT 133.280 52.990 133.450 53.615 ;
        RECT 133.735 53.015 133.915 53.795 ;
        RECT 132.590 52.830 133.450 52.990 ;
        RECT 132.590 52.660 133.700 52.830 ;
        RECT 133.530 52.405 133.700 52.660 ;
        RECT 134.095 52.795 134.430 53.555 ;
        RECT 134.610 52.965 134.780 53.795 ;
        RECT 134.950 52.795 135.280 53.555 ;
        RECT 135.450 52.965 135.620 53.795 ;
        RECT 134.095 52.625 135.765 52.795 ;
        RECT 135.935 52.705 139.445 53.795 ;
        RECT 139.705 53.125 139.875 53.625 ;
        RECT 140.045 53.295 140.375 53.795 ;
        RECT 139.705 52.955 140.370 53.125 ;
        RECT 134.155 52.605 134.325 52.625 ;
        RECT 132.250 52.235 133.340 52.405 ;
        RECT 133.530 52.235 135.350 52.405 ;
        RECT 132.250 51.695 132.420 52.235 ;
        RECT 133.530 52.065 133.700 52.235 ;
        RECT 133.200 51.895 133.700 52.065 ;
        RECT 135.520 52.060 135.765 52.625 ;
        RECT 131.060 51.525 131.520 51.695 ;
        RECT 131.750 51.525 132.420 51.695 ;
        RECT 132.735 51.245 132.905 51.775 ;
        RECT 133.200 51.455 133.560 51.895 ;
        RECT 134.095 51.890 135.765 52.060 ;
        RECT 135.935 52.015 137.585 52.535 ;
        RECT 137.755 52.185 139.445 52.705 ;
        RECT 139.620 52.135 139.970 52.785 ;
        RECT 133.735 51.245 133.905 51.725 ;
        RECT 134.095 51.465 134.430 51.890 ;
        RECT 134.605 51.245 134.775 51.720 ;
        RECT 134.950 51.465 135.285 51.890 ;
        RECT 135.455 51.245 135.625 51.720 ;
        RECT 135.935 51.245 139.445 52.015 ;
        RECT 140.140 51.965 140.370 52.955 ;
        RECT 139.705 51.795 140.370 51.965 ;
        RECT 139.705 51.505 139.875 51.795 ;
        RECT 140.045 51.245 140.375 51.625 ;
        RECT 140.545 51.505 140.770 53.625 ;
        RECT 140.970 53.335 141.235 53.795 ;
        RECT 141.420 53.225 141.655 53.600 ;
        RECT 141.900 53.350 142.970 53.520 ;
        RECT 140.970 52.225 141.250 52.825 ;
        RECT 140.985 51.245 141.235 51.705 ;
        RECT 141.420 51.695 141.590 53.225 ;
        RECT 141.760 52.195 142.000 53.065 ;
        RECT 142.190 52.815 142.630 53.170 ;
        RECT 142.800 52.735 142.970 53.350 ;
        RECT 143.140 52.995 143.310 53.795 ;
        RECT 143.480 53.295 143.730 53.625 ;
        RECT 143.955 53.325 144.840 53.495 ;
        RECT 142.800 52.645 143.310 52.735 ;
        RECT 142.510 52.475 143.310 52.645 ;
        RECT 141.760 51.865 142.340 52.195 ;
        RECT 142.510 51.695 142.680 52.475 ;
        RECT 143.140 52.405 143.310 52.475 ;
        RECT 142.850 52.225 143.020 52.255 ;
        RECT 143.480 52.225 143.650 53.295 ;
        RECT 143.820 52.405 144.010 53.125 ;
        RECT 144.180 52.735 144.500 53.065 ;
        RECT 142.850 51.925 143.650 52.225 ;
        RECT 144.180 52.195 144.370 52.735 ;
        RECT 141.420 51.525 141.750 51.695 ;
        RECT 141.930 51.525 142.680 51.695 ;
        RECT 142.930 51.245 143.300 51.745 ;
        RECT 143.480 51.695 143.650 51.925 ;
        RECT 143.820 51.865 144.370 52.195 ;
        RECT 144.670 52.405 144.840 53.325 ;
        RECT 145.020 53.295 145.235 53.795 ;
        RECT 145.700 52.990 145.870 53.615 ;
        RECT 146.155 53.015 146.335 53.795 ;
        RECT 145.010 52.830 145.870 52.990 ;
        RECT 145.010 52.660 146.120 52.830 ;
        RECT 145.950 52.405 146.120 52.660 ;
        RECT 146.515 52.795 146.850 53.555 ;
        RECT 147.030 52.965 147.200 53.795 ;
        RECT 147.370 52.795 147.700 53.555 ;
        RECT 147.870 52.965 148.040 53.795 ;
        RECT 146.515 52.625 148.185 52.795 ;
        RECT 148.355 52.705 153.700 53.795 ;
        RECT 146.575 52.605 146.745 52.625 ;
        RECT 144.670 52.235 145.760 52.405 ;
        RECT 145.950 52.235 147.770 52.405 ;
        RECT 144.670 51.695 144.840 52.235 ;
        RECT 145.950 52.065 146.120 52.235 ;
        RECT 145.620 51.895 146.120 52.065 ;
        RECT 147.940 52.060 148.185 52.625 ;
        RECT 143.480 51.525 143.940 51.695 ;
        RECT 144.170 51.525 144.840 51.695 ;
        RECT 145.155 51.245 145.325 51.775 ;
        RECT 145.620 51.455 145.980 51.895 ;
        RECT 146.515 51.890 148.185 52.060 ;
        RECT 148.355 52.015 150.935 52.535 ;
        RECT 151.105 52.185 153.700 52.705 ;
        RECT 154.795 52.630 155.085 53.795 ;
        RECT 155.345 53.125 155.515 53.625 ;
        RECT 155.685 53.295 156.015 53.795 ;
        RECT 155.345 52.955 156.010 53.125 ;
        RECT 155.260 52.135 155.610 52.785 ;
        RECT 146.155 51.245 146.325 51.725 ;
        RECT 146.515 51.465 146.850 51.890 ;
        RECT 147.025 51.245 147.195 51.720 ;
        RECT 147.370 51.465 147.705 51.890 ;
        RECT 147.875 51.245 148.045 51.720 ;
        RECT 148.355 51.245 153.700 52.015 ;
        RECT 154.795 51.245 155.085 51.970 ;
        RECT 155.780 51.965 156.010 52.955 ;
        RECT 155.345 51.795 156.010 51.965 ;
        RECT 155.345 51.505 155.515 51.795 ;
        RECT 155.685 51.245 156.015 51.625 ;
        RECT 156.185 51.505 156.410 53.625 ;
        RECT 156.610 53.335 156.875 53.795 ;
        RECT 157.060 53.225 157.295 53.600 ;
        RECT 157.540 53.350 158.610 53.520 ;
        RECT 156.610 52.225 156.890 52.825 ;
        RECT 156.625 51.245 156.875 51.705 ;
        RECT 157.060 51.695 157.230 53.225 ;
        RECT 157.400 52.195 157.640 53.065 ;
        RECT 157.830 52.815 158.270 53.170 ;
        RECT 158.440 52.735 158.610 53.350 ;
        RECT 158.780 52.995 158.950 53.795 ;
        RECT 159.120 53.295 159.370 53.625 ;
        RECT 159.595 53.325 160.480 53.495 ;
        RECT 158.440 52.645 158.950 52.735 ;
        RECT 158.150 52.475 158.950 52.645 ;
        RECT 157.400 51.865 157.980 52.195 ;
        RECT 158.150 51.695 158.320 52.475 ;
        RECT 158.780 52.405 158.950 52.475 ;
        RECT 158.490 52.225 158.660 52.255 ;
        RECT 159.120 52.225 159.290 53.295 ;
        RECT 159.460 52.405 159.650 53.125 ;
        RECT 159.820 52.735 160.140 53.065 ;
        RECT 158.490 51.925 159.290 52.225 ;
        RECT 159.820 52.195 160.010 52.735 ;
        RECT 157.060 51.525 157.390 51.695 ;
        RECT 157.570 51.525 158.320 51.695 ;
        RECT 158.570 51.245 158.940 51.745 ;
        RECT 159.120 51.695 159.290 51.925 ;
        RECT 159.460 51.865 160.010 52.195 ;
        RECT 160.310 52.405 160.480 53.325 ;
        RECT 160.660 53.295 160.875 53.795 ;
        RECT 161.340 52.990 161.510 53.615 ;
        RECT 161.795 53.015 161.975 53.795 ;
        RECT 160.650 52.830 161.510 52.990 ;
        RECT 160.650 52.660 161.760 52.830 ;
        RECT 161.590 52.405 161.760 52.660 ;
        RECT 162.155 52.795 162.490 53.555 ;
        RECT 162.670 52.965 162.840 53.795 ;
        RECT 163.010 52.795 163.340 53.555 ;
        RECT 163.510 52.965 163.680 53.795 ;
        RECT 162.155 52.625 163.825 52.795 ;
        RECT 163.995 52.705 169.340 53.795 ;
        RECT 170.525 53.125 170.695 53.625 ;
        RECT 170.865 53.295 171.195 53.795 ;
        RECT 170.525 52.955 171.190 53.125 ;
        RECT 160.310 52.235 161.400 52.405 ;
        RECT 161.590 52.235 163.410 52.405 ;
        RECT 160.310 51.695 160.480 52.235 ;
        RECT 161.590 52.065 161.760 52.235 ;
        RECT 161.260 51.895 161.760 52.065 ;
        RECT 163.580 52.060 163.825 52.625 ;
        RECT 159.120 51.525 159.580 51.695 ;
        RECT 159.810 51.525 160.480 51.695 ;
        RECT 160.795 51.245 160.965 51.775 ;
        RECT 161.260 51.455 161.620 51.895 ;
        RECT 162.155 51.890 163.825 52.060 ;
        RECT 163.995 52.015 166.575 52.535 ;
        RECT 166.745 52.185 169.340 52.705 ;
        RECT 170.440 52.135 170.790 52.785 ;
        RECT 161.795 51.245 161.965 51.725 ;
        RECT 162.155 51.465 162.490 51.890 ;
        RECT 162.665 51.245 162.835 51.720 ;
        RECT 163.010 51.465 163.345 51.890 ;
        RECT 163.515 51.245 163.685 51.720 ;
        RECT 163.995 51.245 169.340 52.015 ;
        RECT 170.960 51.965 171.190 52.955 ;
        RECT 170.525 51.795 171.190 51.965 ;
        RECT 170.525 51.505 170.695 51.795 ;
        RECT 170.865 51.245 171.195 51.625 ;
        RECT 171.365 51.505 171.590 53.625 ;
        RECT 171.790 53.335 172.055 53.795 ;
        RECT 172.240 53.225 172.475 53.600 ;
        RECT 172.720 53.350 173.790 53.520 ;
        RECT 171.790 52.225 172.070 52.825 ;
        RECT 171.805 51.245 172.055 51.705 ;
        RECT 172.240 51.695 172.410 53.225 ;
        RECT 172.580 52.195 172.820 53.065 ;
        RECT 173.010 52.815 173.450 53.170 ;
        RECT 173.620 52.735 173.790 53.350 ;
        RECT 173.960 52.995 174.130 53.795 ;
        RECT 174.300 53.295 174.550 53.625 ;
        RECT 174.775 53.325 175.660 53.495 ;
        RECT 173.620 52.645 174.130 52.735 ;
        RECT 173.330 52.475 174.130 52.645 ;
        RECT 172.580 51.865 173.160 52.195 ;
        RECT 173.330 51.695 173.500 52.475 ;
        RECT 173.960 52.405 174.130 52.475 ;
        RECT 173.670 52.225 173.840 52.255 ;
        RECT 174.300 52.225 174.470 53.295 ;
        RECT 174.640 52.405 174.830 53.125 ;
        RECT 175.000 52.735 175.320 53.065 ;
        RECT 173.670 51.925 174.470 52.225 ;
        RECT 175.000 52.195 175.190 52.735 ;
        RECT 172.240 51.525 172.570 51.695 ;
        RECT 172.750 51.525 173.500 51.695 ;
        RECT 173.750 51.245 174.120 51.745 ;
        RECT 174.300 51.695 174.470 51.925 ;
        RECT 174.640 51.865 175.190 52.195 ;
        RECT 175.490 52.405 175.660 53.325 ;
        RECT 175.840 53.295 176.055 53.795 ;
        RECT 176.520 52.990 176.690 53.615 ;
        RECT 176.975 53.015 177.155 53.795 ;
        RECT 175.830 52.830 176.690 52.990 ;
        RECT 175.830 52.660 176.940 52.830 ;
        RECT 176.770 52.405 176.940 52.660 ;
        RECT 177.335 52.795 177.670 53.555 ;
        RECT 177.850 52.965 178.020 53.795 ;
        RECT 178.190 52.795 178.520 53.555 ;
        RECT 178.690 52.965 178.860 53.795 ;
        RECT 177.335 52.625 179.005 52.795 ;
        RECT 179.175 52.705 182.685 53.795 ;
        RECT 177.395 52.605 177.565 52.625 ;
        RECT 175.490 52.235 176.580 52.405 ;
        RECT 176.770 52.235 178.590 52.405 ;
        RECT 175.490 51.695 175.660 52.235 ;
        RECT 176.770 52.065 176.940 52.235 ;
        RECT 176.440 51.895 176.940 52.065 ;
        RECT 178.760 52.060 179.005 52.625 ;
        RECT 174.300 51.525 174.760 51.695 ;
        RECT 174.990 51.525 175.660 51.695 ;
        RECT 175.975 51.245 176.145 51.775 ;
        RECT 176.440 51.455 176.800 51.895 ;
        RECT 177.335 51.890 179.005 52.060 ;
        RECT 179.175 52.015 180.825 52.535 ;
        RECT 180.995 52.185 182.685 52.705 ;
        RECT 182.855 52.630 183.145 53.795 ;
        RECT 183.315 52.705 184.985 53.795 ;
        RECT 185.245 53.125 185.415 53.625 ;
        RECT 185.585 53.295 185.915 53.795 ;
        RECT 185.245 52.955 185.910 53.125 ;
        RECT 183.315 52.015 184.065 52.535 ;
        RECT 184.235 52.185 184.985 52.705 ;
        RECT 185.160 52.135 185.510 52.785 ;
        RECT 176.975 51.245 177.145 51.725 ;
        RECT 177.335 51.465 177.670 51.890 ;
        RECT 177.845 51.245 178.015 51.720 ;
        RECT 178.190 51.465 178.525 51.890 ;
        RECT 178.695 51.245 178.865 51.720 ;
        RECT 179.175 51.245 182.685 52.015 ;
        RECT 182.855 51.245 183.145 51.970 ;
        RECT 183.315 51.245 184.985 52.015 ;
        RECT 185.680 51.965 185.910 52.955 ;
        RECT 185.245 51.795 185.910 51.965 ;
        RECT 185.245 51.505 185.415 51.795 ;
        RECT 185.585 51.245 185.915 51.625 ;
        RECT 186.085 51.505 186.310 53.625 ;
        RECT 186.510 53.335 186.775 53.795 ;
        RECT 186.960 53.225 187.195 53.600 ;
        RECT 187.440 53.350 188.510 53.520 ;
        RECT 186.510 52.225 186.790 52.825 ;
        RECT 186.525 51.245 186.775 51.705 ;
        RECT 186.960 51.695 187.130 53.225 ;
        RECT 187.300 52.195 187.540 53.065 ;
        RECT 187.730 52.815 188.170 53.170 ;
        RECT 188.340 52.735 188.510 53.350 ;
        RECT 188.680 52.995 188.850 53.795 ;
        RECT 189.020 53.295 189.270 53.625 ;
        RECT 189.495 53.325 190.380 53.495 ;
        RECT 188.340 52.645 188.850 52.735 ;
        RECT 188.050 52.475 188.850 52.645 ;
        RECT 187.300 51.865 187.880 52.195 ;
        RECT 188.050 51.695 188.220 52.475 ;
        RECT 188.680 52.405 188.850 52.475 ;
        RECT 188.390 52.225 188.560 52.255 ;
        RECT 189.020 52.225 189.190 53.295 ;
        RECT 189.360 52.405 189.550 53.125 ;
        RECT 189.720 52.735 190.040 53.065 ;
        RECT 188.390 51.925 189.190 52.225 ;
        RECT 189.720 52.195 189.910 52.735 ;
        RECT 186.960 51.525 187.290 51.695 ;
        RECT 187.470 51.525 188.220 51.695 ;
        RECT 188.470 51.245 188.840 51.745 ;
        RECT 189.020 51.695 189.190 51.925 ;
        RECT 189.360 51.865 189.910 52.195 ;
        RECT 190.210 52.405 190.380 53.325 ;
        RECT 190.560 53.295 190.775 53.795 ;
        RECT 191.240 52.990 191.410 53.615 ;
        RECT 191.695 53.015 191.875 53.795 ;
        RECT 190.550 52.830 191.410 52.990 ;
        RECT 190.550 52.660 191.660 52.830 ;
        RECT 191.490 52.405 191.660 52.660 ;
        RECT 192.055 52.795 192.390 53.555 ;
        RECT 192.570 52.965 192.740 53.795 ;
        RECT 192.910 52.795 193.240 53.555 ;
        RECT 193.410 52.965 193.580 53.795 ;
        RECT 192.055 52.625 193.725 52.795 ;
        RECT 193.895 52.705 197.405 53.795 ;
        RECT 198.125 53.125 198.295 53.625 ;
        RECT 198.465 53.295 198.795 53.795 ;
        RECT 198.125 52.955 198.790 53.125 ;
        RECT 190.210 52.235 191.300 52.405 ;
        RECT 191.490 52.235 193.310 52.405 ;
        RECT 190.210 51.695 190.380 52.235 ;
        RECT 191.490 52.065 191.660 52.235 ;
        RECT 191.160 51.895 191.660 52.065 ;
        RECT 193.480 52.060 193.725 52.625 ;
        RECT 189.020 51.525 189.480 51.695 ;
        RECT 189.710 51.525 190.380 51.695 ;
        RECT 190.695 51.245 190.865 51.775 ;
        RECT 191.160 51.455 191.520 51.895 ;
        RECT 192.055 51.890 193.725 52.060 ;
        RECT 193.895 52.015 195.545 52.535 ;
        RECT 195.715 52.185 197.405 52.705 ;
        RECT 198.040 52.135 198.390 52.785 ;
        RECT 191.695 51.245 191.865 51.725 ;
        RECT 192.055 51.465 192.390 51.890 ;
        RECT 192.565 51.245 192.735 51.720 ;
        RECT 192.910 51.465 193.245 51.890 ;
        RECT 193.415 51.245 193.585 51.720 ;
        RECT 193.895 51.245 197.405 52.015 ;
        RECT 198.560 51.965 198.790 52.955 ;
        RECT 198.125 51.795 198.790 51.965 ;
        RECT 198.125 51.505 198.295 51.795 ;
        RECT 198.465 51.245 198.795 51.625 ;
        RECT 198.965 51.505 199.190 53.625 ;
        RECT 199.390 53.335 199.655 53.795 ;
        RECT 199.840 53.225 200.075 53.600 ;
        RECT 200.320 53.350 201.390 53.520 ;
        RECT 199.390 52.225 199.670 52.825 ;
        RECT 199.405 51.245 199.655 51.705 ;
        RECT 199.840 51.695 200.010 53.225 ;
        RECT 200.180 52.195 200.420 53.065 ;
        RECT 200.610 52.815 201.050 53.170 ;
        RECT 201.220 52.735 201.390 53.350 ;
        RECT 201.560 52.995 201.730 53.795 ;
        RECT 201.900 53.295 202.150 53.625 ;
        RECT 202.375 53.325 203.260 53.495 ;
        RECT 201.220 52.645 201.730 52.735 ;
        RECT 200.930 52.475 201.730 52.645 ;
        RECT 200.180 51.865 200.760 52.195 ;
        RECT 200.930 51.695 201.100 52.475 ;
        RECT 201.560 52.405 201.730 52.475 ;
        RECT 201.270 52.225 201.440 52.255 ;
        RECT 201.900 52.225 202.070 53.295 ;
        RECT 202.240 52.405 202.430 53.125 ;
        RECT 202.600 52.735 202.920 53.065 ;
        RECT 201.270 51.925 202.070 52.225 ;
        RECT 202.600 52.195 202.790 52.735 ;
        RECT 199.840 51.525 200.170 51.695 ;
        RECT 200.350 51.525 201.100 51.695 ;
        RECT 201.350 51.245 201.720 51.745 ;
        RECT 201.900 51.695 202.070 51.925 ;
        RECT 202.240 51.865 202.790 52.195 ;
        RECT 203.090 52.405 203.260 53.325 ;
        RECT 203.440 53.295 203.655 53.795 ;
        RECT 204.120 52.990 204.290 53.615 ;
        RECT 204.575 53.015 204.755 53.795 ;
        RECT 203.430 52.830 204.290 52.990 ;
        RECT 203.430 52.660 204.540 52.830 ;
        RECT 204.370 52.405 204.540 52.660 ;
        RECT 204.935 52.795 205.270 53.555 ;
        RECT 205.450 52.965 205.620 53.795 ;
        RECT 205.790 52.795 206.120 53.555 ;
        RECT 206.290 52.965 206.460 53.795 ;
        RECT 204.935 52.625 206.605 52.795 ;
        RECT 206.775 52.705 210.285 53.795 ;
        RECT 203.090 52.235 204.180 52.405 ;
        RECT 204.370 52.235 206.190 52.405 ;
        RECT 203.090 51.695 203.260 52.235 ;
        RECT 204.370 52.065 204.540 52.235 ;
        RECT 204.040 51.895 204.540 52.065 ;
        RECT 206.360 52.060 206.605 52.625 ;
        RECT 201.900 51.525 202.360 51.695 ;
        RECT 202.590 51.525 203.260 51.695 ;
        RECT 203.575 51.245 203.745 51.775 ;
        RECT 204.040 51.455 204.400 51.895 ;
        RECT 204.935 51.890 206.605 52.060 ;
        RECT 206.775 52.015 208.425 52.535 ;
        RECT 208.595 52.185 210.285 52.705 ;
        RECT 204.575 51.245 204.745 51.725 ;
        RECT 204.935 51.465 205.270 51.890 ;
        RECT 205.445 51.245 205.615 51.720 ;
        RECT 205.790 51.465 206.125 51.890 ;
        RECT 206.295 51.245 206.465 51.720 ;
        RECT 206.775 51.245 210.285 52.015 ;
        RECT 210.515 51.925 210.685 52.775 ;
        RECT 210.915 52.630 211.205 53.795 ;
        RECT 212.345 53.115 212.595 53.625 ;
        RECT 212.765 53.285 213.015 53.795 ;
        RECT 213.185 53.115 213.435 53.625 ;
        RECT 213.605 53.285 213.855 53.795 ;
        RECT 214.025 53.455 215.115 53.625 ;
        RECT 214.025 53.115 214.275 53.455 ;
        RECT 214.865 53.295 215.115 53.455 ;
        RECT 215.385 53.295 215.635 53.795 ;
        RECT 215.805 53.455 216.895 53.625 ;
        RECT 215.805 53.295 216.055 53.455 ;
        RECT 212.345 52.945 214.275 53.115 ;
        RECT 212.295 52.605 213.895 52.775 ;
        RECT 214.065 52.615 214.275 52.945 ;
        RECT 214.445 53.125 214.695 53.285 ;
        RECT 216.225 53.125 216.475 53.285 ;
        RECT 212.295 52.235 212.785 52.605 ;
        RECT 213.015 52.235 213.555 52.435 ;
        RECT 213.725 52.405 213.895 52.605 ;
        RECT 214.445 52.575 214.830 53.125 ;
        RECT 215.345 52.945 216.475 53.125 ;
        RECT 216.645 52.945 216.895 53.455 ;
        RECT 217.065 52.955 217.315 53.795 ;
        RECT 217.485 53.115 217.735 53.625 ;
        RECT 217.905 53.325 218.155 53.795 ;
        RECT 218.325 53.115 218.575 53.625 ;
        RECT 217.485 52.945 218.575 53.115 ;
        RECT 218.745 52.985 218.995 53.795 ;
        RECT 215.345 52.825 215.515 52.945 ;
        RECT 215.165 52.655 215.515 52.825 ;
        RECT 218.325 52.815 218.575 52.945 ;
        RECT 213.725 52.235 214.105 52.405 ;
        RECT 214.445 52.065 214.655 52.575 ;
        RECT 215.165 52.405 215.355 52.655 ;
        RECT 215.685 52.605 217.175 52.775 ;
        RECT 215.685 52.485 215.855 52.605 ;
        RECT 214.825 52.235 215.355 52.405 ;
        RECT 215.525 52.235 215.855 52.485 ;
        RECT 216.025 52.235 216.645 52.435 ;
        RECT 216.815 52.235 217.175 52.605 ;
        RECT 217.345 52.405 217.670 52.775 ;
        RECT 218.325 52.575 219.130 52.815 ;
        RECT 219.655 52.705 223.165 53.795 ;
        RECT 217.345 52.235 218.650 52.405 ;
        RECT 215.165 52.065 215.355 52.235 ;
        RECT 218.820 52.065 219.130 52.575 ;
        RECT 210.915 51.245 211.205 51.970 ;
        RECT 212.385 51.245 212.555 52.055 ;
        RECT 212.725 51.635 212.975 52.065 ;
        RECT 213.145 51.895 214.735 52.065 ;
        RECT 213.145 51.805 213.480 51.895 ;
        RECT 212.725 51.415 213.895 51.635 ;
        RECT 214.065 51.245 214.235 51.715 ;
        RECT 214.405 51.415 214.735 51.895 ;
        RECT 215.165 51.885 216.935 52.065 ;
        RECT 214.905 51.245 215.595 51.715 ;
        RECT 215.765 51.415 216.095 51.885 ;
        RECT 216.265 51.245 216.435 51.715 ;
        RECT 216.605 51.415 216.935 51.885 ;
        RECT 217.105 51.245 217.275 52.055 ;
        RECT 217.445 51.885 219.130 52.065 ;
        RECT 219.655 52.015 221.305 52.535 ;
        RECT 221.475 52.185 223.165 52.705 ;
        RECT 223.340 52.825 223.615 53.625 ;
        RECT 223.785 52.995 224.115 53.795 ;
        RECT 224.285 52.825 224.455 53.625 ;
        RECT 224.625 52.995 224.875 53.795 ;
        RECT 225.045 53.455 227.140 53.625 ;
        RECT 225.045 52.825 225.375 53.455 ;
        RECT 223.340 52.615 225.375 52.825 ;
        RECT 225.545 52.905 225.715 53.285 ;
        RECT 225.885 53.095 226.215 53.455 ;
        RECT 226.385 52.905 226.555 53.285 ;
        RECT 226.725 53.075 227.140 53.455 ;
        RECT 225.545 52.605 227.305 52.905 ;
        RECT 227.475 52.705 230.985 53.795 ;
        RECT 223.390 52.235 225.050 52.435 ;
        RECT 225.370 52.235 226.735 52.435 ;
        RECT 226.905 52.065 227.305 52.605 ;
        RECT 217.445 51.435 217.775 51.885 ;
        RECT 217.945 51.245 218.115 51.715 ;
        RECT 218.285 51.435 218.615 51.885 ;
        RECT 218.785 51.245 218.955 51.715 ;
        RECT 219.655 51.245 223.165 52.015 ;
        RECT 223.340 51.245 223.615 52.065 ;
        RECT 223.785 51.885 227.305 52.065 ;
        RECT 227.475 52.015 229.125 52.535 ;
        RECT 229.295 52.185 230.985 52.705 ;
        RECT 231.185 52.500 231.435 53.495 ;
        RECT 231.615 52.910 231.795 53.625 ;
        RECT 231.965 53.095 232.415 53.795 ;
        RECT 232.590 52.910 232.770 53.625 ;
        RECT 232.980 53.095 233.310 53.795 ;
        RECT 233.520 52.920 233.710 53.625 ;
        RECT 233.880 53.095 234.210 53.795 ;
        RECT 234.380 52.925 234.570 53.625 ;
        RECT 234.740 53.095 235.070 53.795 ;
        RECT 234.380 52.920 235.125 52.925 ;
        RECT 231.615 52.740 233.350 52.910 ;
        RECT 233.140 52.515 233.350 52.740 ;
        RECT 233.520 52.695 235.125 52.920 ;
        RECT 235.295 52.705 238.805 53.795 ;
        RECT 231.185 52.155 231.945 52.500 ;
        RECT 223.785 51.415 224.115 51.885 ;
        RECT 224.285 51.245 224.455 51.715 ;
        RECT 224.625 51.415 224.955 51.885 ;
        RECT 225.125 51.245 225.295 51.715 ;
        RECT 225.465 51.415 225.795 51.885 ;
        RECT 225.965 51.245 226.135 51.715 ;
        RECT 226.305 51.415 226.635 51.885 ;
        RECT 226.805 51.245 227.090 51.715 ;
        RECT 227.475 51.245 230.985 52.015 ;
        RECT 231.535 51.725 231.870 51.965 ;
        RECT 232.135 51.905 232.425 52.500 ;
        RECT 232.595 52.155 232.970 52.485 ;
        RECT 233.140 52.180 234.675 52.515 ;
        RECT 233.140 51.965 233.350 52.180 ;
        RECT 234.845 52.005 235.125 52.695 ;
        RECT 232.605 51.775 233.350 51.965 ;
        RECT 233.520 51.775 235.125 52.005 ;
        RECT 235.295 52.015 236.945 52.535 ;
        RECT 237.115 52.185 238.805 52.705 ;
        RECT 238.975 52.630 239.265 53.795 ;
        RECT 239.525 52.865 239.695 53.625 ;
        RECT 239.910 53.035 240.240 53.795 ;
        RECT 239.525 52.695 240.240 52.865 ;
        RECT 240.410 52.720 240.665 53.625 ;
        RECT 239.435 52.145 239.790 52.515 ;
        RECT 240.070 52.485 240.240 52.695 ;
        RECT 240.070 52.155 240.325 52.485 ;
        RECT 232.605 51.725 232.795 51.775 ;
        RECT 231.535 51.535 232.795 51.725 ;
        RECT 233.520 51.675 233.710 51.775 ;
        RECT 231.535 51.415 231.870 51.535 ;
        RECT 232.975 51.245 233.305 51.605 ;
        RECT 233.880 51.245 234.210 51.605 ;
        RECT 234.380 51.415 234.570 51.775 ;
        RECT 234.740 51.245 235.070 51.605 ;
        RECT 235.295 51.245 238.805 52.015 ;
        RECT 238.975 51.245 239.265 51.970 ;
        RECT 240.070 51.965 240.240 52.155 ;
        RECT 240.495 51.990 240.665 52.720 ;
        RECT 240.840 52.645 241.100 53.795 ;
        RECT 241.275 52.705 244.785 53.795 ;
        RECT 245.005 53.115 245.255 53.625 ;
        RECT 245.425 53.285 245.675 53.795 ;
        RECT 245.845 53.115 246.095 53.625 ;
        RECT 246.265 53.285 246.515 53.795 ;
        RECT 246.685 53.455 247.775 53.625 ;
        RECT 246.685 53.115 246.935 53.455 ;
        RECT 247.525 53.295 247.775 53.455 ;
        RECT 248.045 53.295 248.295 53.795 ;
        RECT 248.465 53.455 249.555 53.625 ;
        RECT 248.465 53.295 248.715 53.455 ;
        RECT 245.005 52.945 246.935 53.115 ;
        RECT 239.525 51.795 240.240 51.965 ;
        RECT 239.525 51.415 239.695 51.795 ;
        RECT 239.910 51.245 240.240 51.625 ;
        RECT 240.410 51.415 240.665 51.990 ;
        RECT 240.840 51.245 241.100 52.085 ;
        RECT 241.275 52.015 242.925 52.535 ;
        RECT 243.095 52.185 244.785 52.705 ;
        RECT 244.955 52.605 246.555 52.775 ;
        RECT 246.725 52.615 246.935 52.945 ;
        RECT 247.105 53.125 247.355 53.285 ;
        RECT 248.885 53.125 249.135 53.285 ;
        RECT 244.955 52.235 245.445 52.605 ;
        RECT 245.675 52.235 246.215 52.435 ;
        RECT 246.385 52.405 246.555 52.605 ;
        RECT 247.105 52.575 247.490 53.125 ;
        RECT 248.005 52.945 249.135 53.125 ;
        RECT 249.305 52.945 249.555 53.455 ;
        RECT 249.725 52.955 249.975 53.795 ;
        RECT 250.145 53.115 250.395 53.625 ;
        RECT 250.565 53.325 250.815 53.795 ;
        RECT 250.985 53.115 251.235 53.625 ;
        RECT 250.145 52.945 251.235 53.115 ;
        RECT 251.405 52.985 251.655 53.795 ;
        RECT 248.005 52.825 248.175 52.945 ;
        RECT 247.825 52.655 248.175 52.825 ;
        RECT 250.985 52.815 251.235 52.945 ;
        RECT 246.385 52.235 246.765 52.405 ;
        RECT 247.105 52.065 247.315 52.575 ;
        RECT 247.825 52.405 248.015 52.655 ;
        RECT 248.345 52.605 249.835 52.775 ;
        RECT 248.345 52.485 248.515 52.605 ;
        RECT 247.485 52.235 248.015 52.405 ;
        RECT 248.185 52.235 248.515 52.485 ;
        RECT 248.685 52.235 249.305 52.435 ;
        RECT 249.475 52.235 249.835 52.605 ;
        RECT 250.005 52.405 250.330 52.775 ;
        RECT 250.985 52.575 251.790 52.815 ;
        RECT 252.315 52.705 255.825 53.795 ;
        RECT 256.045 53.115 256.295 53.625 ;
        RECT 256.465 53.285 256.715 53.795 ;
        RECT 256.885 53.115 257.135 53.625 ;
        RECT 257.305 53.285 257.555 53.795 ;
        RECT 257.725 53.455 258.815 53.625 ;
        RECT 257.725 53.115 257.975 53.455 ;
        RECT 258.565 53.295 258.815 53.455 ;
        RECT 259.085 53.295 259.335 53.795 ;
        RECT 259.505 53.455 260.595 53.625 ;
        RECT 259.505 53.295 259.755 53.455 ;
        RECT 256.045 52.945 257.975 53.115 ;
        RECT 250.005 52.235 251.310 52.405 ;
        RECT 247.825 52.065 248.015 52.235 ;
        RECT 251.480 52.065 251.790 52.575 ;
        RECT 241.275 51.245 244.785 52.015 ;
        RECT 245.045 51.245 245.215 52.055 ;
        RECT 245.385 51.635 245.635 52.065 ;
        RECT 245.805 51.895 247.395 52.065 ;
        RECT 245.805 51.805 246.140 51.895 ;
        RECT 245.385 51.415 246.555 51.635 ;
        RECT 246.725 51.245 246.895 51.715 ;
        RECT 247.065 51.415 247.395 51.895 ;
        RECT 247.825 51.885 249.595 52.065 ;
        RECT 247.565 51.245 248.255 51.715 ;
        RECT 248.425 51.415 248.755 51.885 ;
        RECT 248.925 51.245 249.095 51.715 ;
        RECT 249.265 51.415 249.595 51.885 ;
        RECT 249.765 51.245 249.935 52.055 ;
        RECT 250.105 51.885 251.790 52.065 ;
        RECT 252.315 52.015 253.965 52.535 ;
        RECT 254.135 52.185 255.825 52.705 ;
        RECT 255.995 52.605 257.595 52.775 ;
        RECT 257.765 52.615 257.975 52.945 ;
        RECT 258.145 53.125 258.395 53.285 ;
        RECT 259.925 53.125 260.175 53.285 ;
        RECT 255.995 52.235 256.485 52.605 ;
        RECT 256.715 52.235 257.255 52.435 ;
        RECT 257.425 52.405 257.595 52.605 ;
        RECT 258.145 52.575 258.530 53.125 ;
        RECT 259.045 52.945 260.175 53.125 ;
        RECT 260.345 52.945 260.595 53.455 ;
        RECT 260.765 52.955 261.015 53.795 ;
        RECT 261.185 53.115 261.435 53.625 ;
        RECT 261.605 53.325 261.855 53.795 ;
        RECT 262.025 53.115 262.275 53.625 ;
        RECT 261.185 52.945 262.275 53.115 ;
        RECT 262.445 52.985 262.695 53.795 ;
        RECT 259.045 52.825 259.215 52.945 ;
        RECT 258.865 52.655 259.215 52.825 ;
        RECT 262.025 52.815 262.275 52.945 ;
        RECT 257.425 52.235 257.805 52.405 ;
        RECT 258.145 52.065 258.355 52.575 ;
        RECT 258.865 52.405 259.055 52.655 ;
        RECT 259.385 52.605 260.875 52.775 ;
        RECT 259.385 52.485 259.555 52.605 ;
        RECT 258.525 52.235 259.055 52.405 ;
        RECT 259.225 52.235 259.555 52.485 ;
        RECT 259.725 52.235 260.345 52.435 ;
        RECT 260.515 52.235 260.875 52.605 ;
        RECT 261.045 52.405 261.370 52.775 ;
        RECT 262.025 52.575 262.830 52.815 ;
        RECT 263.355 52.705 266.865 53.795 ;
        RECT 261.045 52.235 262.350 52.405 ;
        RECT 258.865 52.065 259.055 52.235 ;
        RECT 262.520 52.065 262.830 52.575 ;
        RECT 250.105 51.435 250.435 51.885 ;
        RECT 250.605 51.245 250.775 51.715 ;
        RECT 250.945 51.435 251.275 51.885 ;
        RECT 251.445 51.245 251.615 51.715 ;
        RECT 252.315 51.245 255.825 52.015 ;
        RECT 256.085 51.245 256.255 52.055 ;
        RECT 256.425 51.635 256.675 52.065 ;
        RECT 256.845 51.895 258.435 52.065 ;
        RECT 256.845 51.805 257.180 51.895 ;
        RECT 256.425 51.415 257.595 51.635 ;
        RECT 257.765 51.245 257.935 51.715 ;
        RECT 258.105 51.415 258.435 51.895 ;
        RECT 258.865 51.885 260.635 52.065 ;
        RECT 258.605 51.245 259.295 51.715 ;
        RECT 259.465 51.415 259.795 51.885 ;
        RECT 259.965 51.245 260.135 51.715 ;
        RECT 260.305 51.415 260.635 51.885 ;
        RECT 260.805 51.245 260.975 52.055 ;
        RECT 261.145 51.885 262.830 52.065 ;
        RECT 263.355 52.015 265.005 52.535 ;
        RECT 265.175 52.185 266.865 52.705 ;
        RECT 267.035 52.630 267.325 53.795 ;
        RECT 267.495 52.705 271.005 53.795 ;
        RECT 271.225 53.115 271.475 53.625 ;
        RECT 271.645 53.285 271.895 53.795 ;
        RECT 272.065 53.115 272.315 53.625 ;
        RECT 272.485 53.285 272.735 53.795 ;
        RECT 272.905 53.455 273.995 53.625 ;
        RECT 272.905 53.115 273.155 53.455 ;
        RECT 273.745 53.295 273.995 53.455 ;
        RECT 274.265 53.295 274.515 53.795 ;
        RECT 274.685 53.455 275.775 53.625 ;
        RECT 274.685 53.295 274.935 53.455 ;
        RECT 271.225 52.945 273.155 53.115 ;
        RECT 267.495 52.015 269.145 52.535 ;
        RECT 269.315 52.185 271.005 52.705 ;
        RECT 271.175 52.605 272.775 52.775 ;
        RECT 272.945 52.615 273.155 52.945 ;
        RECT 273.325 53.125 273.575 53.285 ;
        RECT 275.105 53.125 275.355 53.285 ;
        RECT 271.175 52.235 271.665 52.605 ;
        RECT 272.605 52.435 272.775 52.605 ;
        RECT 273.325 52.575 273.710 53.125 ;
        RECT 274.225 52.945 275.355 53.125 ;
        RECT 275.525 52.945 275.775 53.455 ;
        RECT 275.945 52.955 276.195 53.795 ;
        RECT 276.365 53.115 276.615 53.625 ;
        RECT 276.785 53.325 277.035 53.795 ;
        RECT 277.205 53.115 277.455 53.625 ;
        RECT 276.365 52.945 277.455 53.115 ;
        RECT 277.625 52.985 277.875 53.795 ;
        RECT 274.225 52.825 274.395 52.945 ;
        RECT 274.045 52.655 274.395 52.825 ;
        RECT 277.205 52.815 277.455 52.945 ;
        RECT 271.895 52.235 272.435 52.435 ;
        RECT 272.605 52.405 272.785 52.435 ;
        RECT 272.605 52.235 272.985 52.405 ;
        RECT 273.325 52.065 273.535 52.575 ;
        RECT 274.045 52.405 274.235 52.655 ;
        RECT 274.565 52.605 276.055 52.775 ;
        RECT 274.565 52.485 274.735 52.605 ;
        RECT 273.705 52.235 274.235 52.405 ;
        RECT 274.405 52.235 274.735 52.485 ;
        RECT 274.905 52.235 275.525 52.435 ;
        RECT 275.695 52.235 276.055 52.605 ;
        RECT 276.225 52.405 276.550 52.775 ;
        RECT 277.205 52.575 278.010 52.815 ;
        RECT 278.535 52.705 282.045 53.795 ;
        RECT 282.265 53.115 282.515 53.625 ;
        RECT 282.685 53.285 282.935 53.795 ;
        RECT 283.105 53.115 283.355 53.625 ;
        RECT 283.525 53.285 283.775 53.795 ;
        RECT 283.945 53.455 285.035 53.625 ;
        RECT 283.945 53.115 284.195 53.455 ;
        RECT 284.785 53.295 285.035 53.455 ;
        RECT 285.305 53.295 285.555 53.795 ;
        RECT 285.725 53.455 286.815 53.625 ;
        RECT 285.725 53.295 285.975 53.455 ;
        RECT 282.265 52.945 284.195 53.115 ;
        RECT 276.225 52.235 277.530 52.405 ;
        RECT 274.045 52.065 274.235 52.235 ;
        RECT 277.700 52.065 278.010 52.575 ;
        RECT 261.145 51.435 261.475 51.885 ;
        RECT 261.645 51.245 261.815 51.715 ;
        RECT 261.985 51.435 262.315 51.885 ;
        RECT 262.485 51.245 262.655 51.715 ;
        RECT 263.355 51.245 266.865 52.015 ;
        RECT 267.035 51.245 267.325 51.970 ;
        RECT 267.495 51.245 271.005 52.015 ;
        RECT 271.265 51.245 271.435 52.055 ;
        RECT 271.605 51.635 271.855 52.065 ;
        RECT 272.025 51.895 273.615 52.065 ;
        RECT 272.025 51.805 272.360 51.895 ;
        RECT 271.605 51.415 272.775 51.635 ;
        RECT 272.945 51.245 273.115 51.715 ;
        RECT 273.285 51.415 273.615 51.895 ;
        RECT 274.045 51.885 275.815 52.065 ;
        RECT 273.785 51.245 274.475 51.715 ;
        RECT 274.645 51.415 274.975 51.885 ;
        RECT 275.145 51.245 275.315 51.715 ;
        RECT 275.485 51.415 275.815 51.885 ;
        RECT 275.985 51.245 276.155 52.055 ;
        RECT 276.325 51.885 278.010 52.065 ;
        RECT 278.535 52.015 280.185 52.535 ;
        RECT 280.355 52.185 282.045 52.705 ;
        RECT 282.215 52.605 283.815 52.775 ;
        RECT 283.985 52.615 284.195 52.945 ;
        RECT 284.365 53.125 284.615 53.285 ;
        RECT 286.145 53.125 286.395 53.285 ;
        RECT 282.215 52.235 282.705 52.605 ;
        RECT 283.645 52.435 283.815 52.605 ;
        RECT 284.365 52.575 284.750 53.125 ;
        RECT 285.265 52.945 286.395 53.125 ;
        RECT 286.565 52.945 286.815 53.455 ;
        RECT 286.985 52.955 287.235 53.795 ;
        RECT 287.405 53.115 287.655 53.625 ;
        RECT 287.825 53.325 288.075 53.795 ;
        RECT 288.245 53.115 288.495 53.625 ;
        RECT 287.405 52.945 288.495 53.115 ;
        RECT 288.665 52.985 288.915 53.795 ;
        RECT 285.265 52.825 285.435 52.945 ;
        RECT 285.085 52.655 285.435 52.825 ;
        RECT 288.245 52.815 288.495 52.945 ;
        RECT 282.935 52.235 283.475 52.435 ;
        RECT 283.645 52.405 283.825 52.435 ;
        RECT 283.645 52.235 284.025 52.405 ;
        RECT 284.365 52.065 284.575 52.575 ;
        RECT 285.085 52.405 285.275 52.655 ;
        RECT 285.605 52.605 287.095 52.775 ;
        RECT 285.605 52.485 285.775 52.605 ;
        RECT 284.745 52.235 285.275 52.405 ;
        RECT 285.445 52.235 285.775 52.485 ;
        RECT 285.945 52.235 286.565 52.435 ;
        RECT 286.735 52.235 287.095 52.605 ;
        RECT 287.265 52.405 287.590 52.775 ;
        RECT 288.245 52.575 289.050 52.815 ;
        RECT 289.575 52.705 294.920 53.795 ;
        RECT 287.265 52.235 288.570 52.405 ;
        RECT 285.085 52.065 285.275 52.235 ;
        RECT 288.740 52.065 289.050 52.575 ;
        RECT 276.325 51.435 276.655 51.885 ;
        RECT 276.825 51.245 276.995 51.715 ;
        RECT 277.165 51.435 277.495 51.885 ;
        RECT 277.665 51.245 277.835 51.715 ;
        RECT 278.535 51.245 282.045 52.015 ;
        RECT 282.305 51.245 282.475 52.055 ;
        RECT 282.645 51.635 282.895 52.065 ;
        RECT 283.065 51.895 284.655 52.065 ;
        RECT 283.065 51.805 283.400 51.895 ;
        RECT 282.645 51.415 283.815 51.635 ;
        RECT 283.985 51.245 284.155 51.715 ;
        RECT 284.325 51.415 284.655 51.895 ;
        RECT 285.085 51.885 286.855 52.065 ;
        RECT 284.825 51.245 285.515 51.715 ;
        RECT 285.685 51.415 286.015 51.885 ;
        RECT 286.185 51.245 286.355 51.715 ;
        RECT 286.525 51.415 286.855 51.885 ;
        RECT 287.025 51.245 287.195 52.055 ;
        RECT 287.365 51.885 289.050 52.065 ;
        RECT 289.575 52.015 292.155 52.535 ;
        RECT 292.325 52.185 294.920 52.705 ;
        RECT 295.095 52.630 295.385 53.795 ;
        RECT 295.560 52.825 295.835 53.625 ;
        RECT 296.005 52.995 296.335 53.795 ;
        RECT 296.505 52.825 296.675 53.625 ;
        RECT 296.845 52.995 297.095 53.795 ;
        RECT 297.265 53.455 299.360 53.625 ;
        RECT 297.265 52.825 297.595 53.455 ;
        RECT 295.560 52.615 297.595 52.825 ;
        RECT 297.765 52.905 297.935 53.285 ;
        RECT 298.105 53.095 298.435 53.455 ;
        RECT 298.605 52.905 298.775 53.285 ;
        RECT 298.945 53.075 299.360 53.455 ;
        RECT 297.765 52.605 299.525 52.905 ;
        RECT 299.695 52.705 305.040 53.795 ;
        RECT 306.185 53.115 306.435 53.625 ;
        RECT 306.605 53.285 306.855 53.795 ;
        RECT 307.025 53.115 307.275 53.625 ;
        RECT 307.445 53.285 307.695 53.795 ;
        RECT 307.865 53.455 308.955 53.625 ;
        RECT 307.865 53.115 308.115 53.455 ;
        RECT 308.705 53.295 308.955 53.455 ;
        RECT 309.225 53.295 309.475 53.795 ;
        RECT 309.645 53.455 310.735 53.625 ;
        RECT 309.645 53.295 309.895 53.455 ;
        RECT 306.185 52.945 308.115 53.115 ;
        RECT 295.610 52.235 297.270 52.435 ;
        RECT 297.590 52.235 298.955 52.435 ;
        RECT 299.125 52.065 299.525 52.605 ;
        RECT 287.365 51.435 287.695 51.885 ;
        RECT 287.865 51.245 288.035 51.715 ;
        RECT 288.205 51.435 288.535 51.885 ;
        RECT 288.705 51.245 288.875 51.715 ;
        RECT 289.575 51.245 294.920 52.015 ;
        RECT 295.095 51.245 295.385 51.970 ;
        RECT 295.560 51.245 295.835 52.065 ;
        RECT 296.005 51.885 299.525 52.065 ;
        RECT 299.695 52.015 302.275 52.535 ;
        RECT 302.445 52.185 305.040 52.705 ;
        RECT 306.135 52.605 307.735 52.775 ;
        RECT 307.905 52.615 308.115 52.945 ;
        RECT 308.285 53.125 308.535 53.285 ;
        RECT 310.065 53.125 310.315 53.285 ;
        RECT 306.135 52.235 306.625 52.605 ;
        RECT 307.565 52.435 307.735 52.605 ;
        RECT 308.285 52.575 308.670 53.125 ;
        RECT 309.185 52.945 310.315 53.125 ;
        RECT 310.485 52.945 310.735 53.455 ;
        RECT 310.905 52.955 311.155 53.795 ;
        RECT 311.325 53.115 311.575 53.625 ;
        RECT 311.745 53.325 311.995 53.795 ;
        RECT 312.165 53.115 312.415 53.625 ;
        RECT 311.325 52.945 312.415 53.115 ;
        RECT 312.585 52.985 312.835 53.795 ;
        RECT 309.185 52.825 309.355 52.945 ;
        RECT 309.005 52.655 309.355 52.825 ;
        RECT 312.165 52.815 312.415 52.945 ;
        RECT 306.855 52.235 307.395 52.435 ;
        RECT 307.565 52.405 307.745 52.435 ;
        RECT 307.565 52.235 307.945 52.405 ;
        RECT 308.285 52.065 308.495 52.575 ;
        RECT 309.005 52.405 309.195 52.655 ;
        RECT 309.525 52.605 311.015 52.775 ;
        RECT 309.525 52.485 309.695 52.605 ;
        RECT 308.665 52.235 309.195 52.405 ;
        RECT 309.365 52.235 309.695 52.485 ;
        RECT 309.865 52.235 310.485 52.435 ;
        RECT 310.655 52.235 311.015 52.605 ;
        RECT 311.185 52.405 311.510 52.775 ;
        RECT 312.165 52.575 312.970 52.815 ;
        RECT 313.495 52.705 317.005 53.795 ;
        RECT 311.185 52.235 312.490 52.405 ;
        RECT 309.005 52.065 309.195 52.235 ;
        RECT 312.660 52.065 312.970 52.575 ;
        RECT 296.005 51.415 296.335 51.885 ;
        RECT 296.505 51.245 296.675 51.715 ;
        RECT 296.845 51.415 297.175 51.885 ;
        RECT 297.345 51.245 297.515 51.715 ;
        RECT 297.685 51.415 298.015 51.885 ;
        RECT 298.185 51.245 298.355 51.715 ;
        RECT 298.525 51.415 298.855 51.885 ;
        RECT 299.025 51.245 299.310 51.715 ;
        RECT 299.695 51.245 305.040 52.015 ;
        RECT 306.225 51.245 306.395 52.055 ;
        RECT 306.565 51.635 306.815 52.065 ;
        RECT 306.985 51.895 308.575 52.065 ;
        RECT 306.985 51.805 307.320 51.895 ;
        RECT 306.565 51.415 307.735 51.635 ;
        RECT 307.905 51.245 308.075 51.715 ;
        RECT 308.245 51.415 308.575 51.895 ;
        RECT 309.005 51.885 310.775 52.065 ;
        RECT 308.745 51.245 309.435 51.715 ;
        RECT 309.605 51.415 309.935 51.885 ;
        RECT 310.105 51.245 310.275 51.715 ;
        RECT 310.445 51.415 310.775 51.885 ;
        RECT 310.945 51.245 311.115 52.055 ;
        RECT 311.285 51.885 312.970 52.065 ;
        RECT 313.495 52.015 315.145 52.535 ;
        RECT 315.315 52.185 317.005 52.705 ;
        RECT 317.265 52.865 317.435 53.625 ;
        RECT 317.650 53.035 317.980 53.795 ;
        RECT 317.265 52.695 317.980 52.865 ;
        RECT 318.150 52.720 318.405 53.625 ;
        RECT 317.175 52.145 317.530 52.515 ;
        RECT 317.810 52.485 317.980 52.695 ;
        RECT 317.810 52.155 318.065 52.485 ;
        RECT 311.285 51.435 311.615 51.885 ;
        RECT 311.785 51.245 311.955 51.715 ;
        RECT 312.125 51.435 312.455 51.885 ;
        RECT 312.625 51.245 312.795 51.715 ;
        RECT 313.495 51.245 317.005 52.015 ;
        RECT 317.810 51.965 317.980 52.155 ;
        RECT 318.235 51.990 318.405 52.720 ;
        RECT 318.580 52.645 318.840 53.795 ;
        RECT 319.015 52.705 322.525 53.795 ;
        RECT 317.265 51.795 317.980 51.965 ;
        RECT 317.265 51.415 317.435 51.795 ;
        RECT 317.650 51.245 317.980 51.625 ;
        RECT 318.150 51.415 318.405 51.990 ;
        RECT 318.580 51.245 318.840 52.085 ;
        RECT 319.015 52.015 320.665 52.535 ;
        RECT 320.835 52.185 322.525 52.705 ;
        RECT 323.155 52.630 323.445 53.795 ;
        RECT 323.705 52.865 323.875 53.625 ;
        RECT 324.090 53.035 324.420 53.795 ;
        RECT 323.705 52.695 324.420 52.865 ;
        RECT 324.590 52.720 324.845 53.625 ;
        RECT 323.615 52.145 323.970 52.515 ;
        RECT 324.250 52.485 324.420 52.695 ;
        RECT 324.250 52.155 324.505 52.485 ;
        RECT 319.015 51.245 322.525 52.015 ;
        RECT 323.155 51.245 323.445 51.970 ;
        RECT 324.250 51.965 324.420 52.155 ;
        RECT 324.675 51.990 324.845 52.720 ;
        RECT 325.020 52.645 325.280 53.795 ;
        RECT 325.455 52.705 328.965 53.795 ;
        RECT 329.185 53.115 329.435 53.625 ;
        RECT 329.605 53.285 329.855 53.795 ;
        RECT 330.025 53.115 330.275 53.625 ;
        RECT 330.445 53.285 330.695 53.795 ;
        RECT 330.865 53.455 331.955 53.625 ;
        RECT 330.865 53.115 331.115 53.455 ;
        RECT 331.705 53.295 331.955 53.455 ;
        RECT 332.225 53.295 332.475 53.795 ;
        RECT 332.645 53.455 333.735 53.625 ;
        RECT 332.645 53.295 332.895 53.455 ;
        RECT 329.185 52.945 331.115 53.115 ;
        RECT 323.705 51.795 324.420 51.965 ;
        RECT 323.705 51.415 323.875 51.795 ;
        RECT 324.090 51.245 324.420 51.625 ;
        RECT 324.590 51.415 324.845 51.990 ;
        RECT 325.020 51.245 325.280 52.085 ;
        RECT 325.455 52.015 327.105 52.535 ;
        RECT 327.275 52.185 328.965 52.705 ;
        RECT 329.135 52.605 330.735 52.775 ;
        RECT 330.905 52.615 331.115 52.945 ;
        RECT 331.285 53.125 331.535 53.285 ;
        RECT 333.065 53.125 333.315 53.285 ;
        RECT 329.135 52.235 329.625 52.605 ;
        RECT 329.855 52.235 330.395 52.435 ;
        RECT 330.565 52.405 330.735 52.605 ;
        RECT 331.285 52.575 331.670 53.125 ;
        RECT 332.185 52.945 333.315 53.125 ;
        RECT 333.485 52.945 333.735 53.455 ;
        RECT 333.905 52.955 334.155 53.795 ;
        RECT 334.325 53.115 334.575 53.625 ;
        RECT 334.745 53.325 334.995 53.795 ;
        RECT 335.165 53.115 335.415 53.625 ;
        RECT 334.325 52.945 335.415 53.115 ;
        RECT 335.585 52.985 335.835 53.795 ;
        RECT 332.185 52.825 332.355 52.945 ;
        RECT 332.005 52.655 332.355 52.825 ;
        RECT 335.165 52.815 335.415 52.945 ;
        RECT 330.565 52.235 330.945 52.405 ;
        RECT 331.285 52.065 331.495 52.575 ;
        RECT 332.005 52.405 332.195 52.655 ;
        RECT 332.525 52.605 334.015 52.775 ;
        RECT 332.525 52.485 332.695 52.605 ;
        RECT 331.665 52.235 332.195 52.405 ;
        RECT 332.365 52.235 332.695 52.485 ;
        RECT 332.865 52.235 333.485 52.435 ;
        RECT 333.655 52.235 334.015 52.605 ;
        RECT 334.185 52.405 334.510 52.775 ;
        RECT 335.165 52.575 335.970 52.815 ;
        RECT 336.495 52.705 340.005 53.795 ;
        RECT 340.225 53.115 340.475 53.625 ;
        RECT 340.645 53.285 340.895 53.795 ;
        RECT 341.065 53.115 341.315 53.625 ;
        RECT 341.485 53.285 341.735 53.795 ;
        RECT 341.905 53.455 342.995 53.625 ;
        RECT 341.905 53.115 342.155 53.455 ;
        RECT 342.745 53.295 342.995 53.455 ;
        RECT 343.265 53.295 343.515 53.795 ;
        RECT 343.685 53.455 344.775 53.625 ;
        RECT 343.685 53.295 343.935 53.455 ;
        RECT 340.225 52.945 342.155 53.115 ;
        RECT 334.185 52.235 335.490 52.405 ;
        RECT 332.005 52.065 332.195 52.235 ;
        RECT 335.660 52.065 335.970 52.575 ;
        RECT 325.455 51.245 328.965 52.015 ;
        RECT 329.225 51.245 329.395 52.055 ;
        RECT 329.565 51.635 329.815 52.065 ;
        RECT 329.985 51.895 331.575 52.065 ;
        RECT 329.985 51.805 330.320 51.895 ;
        RECT 329.565 51.415 330.735 51.635 ;
        RECT 330.905 51.245 331.075 51.715 ;
        RECT 331.245 51.415 331.575 51.895 ;
        RECT 332.005 51.885 333.775 52.065 ;
        RECT 331.745 51.245 332.435 51.715 ;
        RECT 332.605 51.415 332.935 51.885 ;
        RECT 333.105 51.245 333.275 51.715 ;
        RECT 333.445 51.415 333.775 51.885 ;
        RECT 333.945 51.245 334.115 52.055 ;
        RECT 334.285 51.885 335.970 52.065 ;
        RECT 336.495 52.015 338.145 52.535 ;
        RECT 338.315 52.185 340.005 52.705 ;
        RECT 340.175 52.605 341.775 52.775 ;
        RECT 341.945 52.615 342.155 52.945 ;
        RECT 342.325 53.125 342.575 53.285 ;
        RECT 344.105 53.125 344.355 53.285 ;
        RECT 340.175 52.235 340.665 52.605 ;
        RECT 340.895 52.235 341.435 52.435 ;
        RECT 341.605 52.405 341.775 52.605 ;
        RECT 342.325 52.575 342.710 53.125 ;
        RECT 343.225 52.945 344.355 53.125 ;
        RECT 344.525 52.945 344.775 53.455 ;
        RECT 344.945 52.955 345.195 53.795 ;
        RECT 345.365 53.115 345.615 53.625 ;
        RECT 345.785 53.325 346.035 53.795 ;
        RECT 346.205 53.115 346.455 53.625 ;
        RECT 345.365 52.945 346.455 53.115 ;
        RECT 346.625 52.985 346.875 53.795 ;
        RECT 343.225 52.825 343.395 52.945 ;
        RECT 343.045 52.655 343.395 52.825 ;
        RECT 346.205 52.815 346.455 52.945 ;
        RECT 341.605 52.235 341.985 52.405 ;
        RECT 342.325 52.065 342.535 52.575 ;
        RECT 343.045 52.405 343.235 52.655 ;
        RECT 343.565 52.605 345.055 52.775 ;
        RECT 343.565 52.485 343.735 52.605 ;
        RECT 342.705 52.235 343.235 52.405 ;
        RECT 343.405 52.235 343.735 52.485 ;
        RECT 343.905 52.235 344.525 52.435 ;
        RECT 344.695 52.235 345.055 52.605 ;
        RECT 345.225 52.405 345.550 52.775 ;
        RECT 346.205 52.575 347.010 52.815 ;
        RECT 347.535 52.705 351.045 53.795 ;
        RECT 345.225 52.235 346.530 52.405 ;
        RECT 343.045 52.065 343.235 52.235 ;
        RECT 346.700 52.065 347.010 52.575 ;
        RECT 334.285 51.435 334.615 51.885 ;
        RECT 334.785 51.245 334.955 51.715 ;
        RECT 335.125 51.435 335.455 51.885 ;
        RECT 335.625 51.245 335.795 51.715 ;
        RECT 336.495 51.245 340.005 52.015 ;
        RECT 340.265 51.245 340.435 52.055 ;
        RECT 340.605 51.635 340.855 52.065 ;
        RECT 341.025 51.895 342.615 52.065 ;
        RECT 341.025 51.805 341.360 51.895 ;
        RECT 340.605 51.415 341.775 51.635 ;
        RECT 341.945 51.245 342.115 51.715 ;
        RECT 342.285 51.415 342.615 51.895 ;
        RECT 343.045 51.885 344.815 52.065 ;
        RECT 342.785 51.245 343.475 51.715 ;
        RECT 343.645 51.415 343.975 51.885 ;
        RECT 344.145 51.245 344.315 51.715 ;
        RECT 344.485 51.415 344.815 51.885 ;
        RECT 344.985 51.245 345.155 52.055 ;
        RECT 345.325 51.885 347.010 52.065 ;
        RECT 347.535 52.015 349.185 52.535 ;
        RECT 349.355 52.185 351.045 52.705 ;
        RECT 351.215 52.630 351.505 53.795 ;
        RECT 351.725 53.115 351.975 53.625 ;
        RECT 352.145 53.285 352.395 53.795 ;
        RECT 352.565 53.115 352.815 53.625 ;
        RECT 352.985 53.285 353.235 53.795 ;
        RECT 353.405 53.455 354.495 53.625 ;
        RECT 353.405 53.115 353.655 53.455 ;
        RECT 354.245 53.295 354.495 53.455 ;
        RECT 354.765 53.295 355.015 53.795 ;
        RECT 355.185 53.455 356.275 53.625 ;
        RECT 355.185 53.295 355.435 53.455 ;
        RECT 351.725 52.945 353.655 53.115 ;
        RECT 351.675 52.605 353.275 52.775 ;
        RECT 353.445 52.615 353.655 52.945 ;
        RECT 353.825 53.125 354.075 53.285 ;
        RECT 355.605 53.125 355.855 53.285 ;
        RECT 351.675 52.235 352.165 52.605 ;
        RECT 352.395 52.235 352.935 52.435 ;
        RECT 353.105 52.405 353.275 52.605 ;
        RECT 353.825 52.575 354.210 53.125 ;
        RECT 354.725 52.945 355.855 53.125 ;
        RECT 356.025 52.945 356.275 53.455 ;
        RECT 356.445 52.955 356.695 53.795 ;
        RECT 356.865 53.115 357.115 53.625 ;
        RECT 357.285 53.325 357.535 53.795 ;
        RECT 357.705 53.115 357.955 53.625 ;
        RECT 356.865 52.945 357.955 53.115 ;
        RECT 358.125 52.985 358.375 53.795 ;
        RECT 354.725 52.825 354.895 52.945 ;
        RECT 354.545 52.655 354.895 52.825 ;
        RECT 357.705 52.815 357.955 52.945 ;
        RECT 353.105 52.235 353.485 52.405 ;
        RECT 353.825 52.065 354.035 52.575 ;
        RECT 354.545 52.405 354.735 52.655 ;
        RECT 355.065 52.605 356.555 52.775 ;
        RECT 355.065 52.485 355.235 52.605 ;
        RECT 354.205 52.235 354.735 52.405 ;
        RECT 354.905 52.235 355.235 52.485 ;
        RECT 355.405 52.235 356.025 52.435 ;
        RECT 356.195 52.235 356.555 52.605 ;
        RECT 356.725 52.405 357.050 52.775 ;
        RECT 357.705 52.575 358.510 52.815 ;
        RECT 359.035 52.705 362.545 53.795 ;
        RECT 356.725 52.235 358.030 52.405 ;
        RECT 354.545 52.065 354.735 52.235 ;
        RECT 358.200 52.065 358.510 52.575 ;
        RECT 345.325 51.435 345.655 51.885 ;
        RECT 345.825 51.245 345.995 51.715 ;
        RECT 346.165 51.435 346.495 51.885 ;
        RECT 346.665 51.245 346.835 51.715 ;
        RECT 347.535 51.245 351.045 52.015 ;
        RECT 351.215 51.245 351.505 51.970 ;
        RECT 351.765 51.245 351.935 52.055 ;
        RECT 352.105 51.635 352.355 52.065 ;
        RECT 352.525 51.895 354.115 52.065 ;
        RECT 352.525 51.805 352.860 51.895 ;
        RECT 352.105 51.415 353.275 51.635 ;
        RECT 353.445 51.245 353.615 51.715 ;
        RECT 353.785 51.415 354.115 51.895 ;
        RECT 354.545 51.885 356.315 52.065 ;
        RECT 354.285 51.245 354.975 51.715 ;
        RECT 355.145 51.415 355.475 51.885 ;
        RECT 355.645 51.245 355.815 51.715 ;
        RECT 355.985 51.415 356.315 51.885 ;
        RECT 356.485 51.245 356.655 52.055 ;
        RECT 356.825 51.885 358.510 52.065 ;
        RECT 359.035 52.015 360.685 52.535 ;
        RECT 360.855 52.185 362.545 52.705 ;
        RECT 362.720 52.825 362.995 53.625 ;
        RECT 363.165 52.995 363.495 53.795 ;
        RECT 363.665 52.825 363.835 53.625 ;
        RECT 364.005 52.995 364.255 53.795 ;
        RECT 364.425 53.455 366.520 53.625 ;
        RECT 364.425 52.825 364.755 53.455 ;
        RECT 362.720 52.615 364.755 52.825 ;
        RECT 364.925 52.905 365.095 53.285 ;
        RECT 365.265 53.095 365.595 53.455 ;
        RECT 365.765 52.905 365.935 53.285 ;
        RECT 366.105 53.075 366.520 53.455 ;
        RECT 364.925 52.605 366.685 52.905 ;
        RECT 366.855 52.705 370.365 53.795 ;
        RECT 362.770 52.235 364.430 52.435 ;
        RECT 364.750 52.235 366.115 52.435 ;
        RECT 366.285 52.065 366.685 52.605 ;
        RECT 356.825 51.435 357.155 51.885 ;
        RECT 357.325 51.245 357.495 51.715 ;
        RECT 357.665 51.435 357.995 51.885 ;
        RECT 358.165 51.245 358.335 51.715 ;
        RECT 359.035 51.245 362.545 52.015 ;
        RECT 362.720 51.245 362.995 52.065 ;
        RECT 363.165 51.885 366.685 52.065 ;
        RECT 366.855 52.015 368.505 52.535 ;
        RECT 368.675 52.185 370.365 52.705 ;
        RECT 370.540 52.825 370.815 53.625 ;
        RECT 370.985 52.995 371.315 53.795 ;
        RECT 371.485 52.825 371.655 53.625 ;
        RECT 371.825 52.995 372.075 53.795 ;
        RECT 372.245 53.455 374.340 53.625 ;
        RECT 372.245 52.825 372.575 53.455 ;
        RECT 370.540 52.615 372.575 52.825 ;
        RECT 372.745 52.905 372.915 53.285 ;
        RECT 373.085 53.095 373.415 53.455 ;
        RECT 373.585 52.905 373.755 53.285 ;
        RECT 373.925 53.075 374.340 53.455 ;
        RECT 372.745 52.605 374.505 52.905 ;
        RECT 374.675 52.705 378.185 53.795 ;
        RECT 370.590 52.235 372.250 52.435 ;
        RECT 372.570 52.235 373.935 52.435 ;
        RECT 374.105 52.065 374.505 52.605 ;
        RECT 363.165 51.415 363.495 51.885 ;
        RECT 363.665 51.245 363.835 51.715 ;
        RECT 364.005 51.415 364.335 51.885 ;
        RECT 364.505 51.245 364.675 51.715 ;
        RECT 364.845 51.415 365.175 51.885 ;
        RECT 365.345 51.245 365.515 51.715 ;
        RECT 365.685 51.415 366.015 51.885 ;
        RECT 366.185 51.245 366.470 51.715 ;
        RECT 366.855 51.245 370.365 52.015 ;
        RECT 370.540 51.245 370.815 52.065 ;
        RECT 370.985 51.885 374.505 52.065 ;
        RECT 374.675 52.015 376.325 52.535 ;
        RECT 376.495 52.185 378.185 52.705 ;
        RECT 379.275 52.630 379.565 53.795 ;
        RECT 379.925 53.070 380.255 53.795 ;
        RECT 370.985 51.415 371.315 51.885 ;
        RECT 371.485 51.245 371.655 51.715 ;
        RECT 371.825 51.415 372.155 51.885 ;
        RECT 372.325 51.245 372.495 51.715 ;
        RECT 372.665 51.415 372.995 51.885 ;
        RECT 373.165 51.245 373.335 51.715 ;
        RECT 373.505 51.415 373.835 51.885 ;
        RECT 374.005 51.245 374.290 51.715 ;
        RECT 374.675 51.245 378.185 52.015 ;
        RECT 379.275 51.245 379.565 51.970 ;
        RECT 379.735 51.415 380.255 52.900 ;
        RECT 380.425 52.075 380.945 53.625 ;
        RECT 381.115 52.705 384.625 53.795 ;
        RECT 384.985 53.070 385.315 53.795 ;
        RECT 381.115 52.015 382.765 52.535 ;
        RECT 382.935 52.185 384.625 52.705 ;
        RECT 380.425 51.245 380.765 51.905 ;
        RECT 381.115 51.245 384.625 52.015 ;
        RECT 384.795 51.415 385.315 52.900 ;
        RECT 385.485 52.075 386.005 53.625 ;
        RECT 386.175 52.705 389.685 53.795 ;
        RECT 390.045 53.070 390.375 53.795 ;
        RECT 386.175 52.015 387.825 52.535 ;
        RECT 387.995 52.185 389.685 52.705 ;
        RECT 385.485 51.245 385.825 51.905 ;
        RECT 386.175 51.245 389.685 52.015 ;
        RECT 389.855 51.415 390.375 52.900 ;
        RECT 390.545 52.075 391.065 53.625 ;
        RECT 391.235 52.705 396.580 53.795 ;
        RECT 396.755 52.705 402.100 53.795 ;
        RECT 402.275 52.705 405.785 53.795 ;
        RECT 405.955 52.705 407.165 53.795 ;
        RECT 391.235 52.015 393.815 52.535 ;
        RECT 393.985 52.185 396.580 52.705 ;
        RECT 396.755 52.015 399.335 52.535 ;
        RECT 399.505 52.185 402.100 52.705 ;
        RECT 402.275 52.015 403.925 52.535 ;
        RECT 404.095 52.185 405.785 52.705 ;
        RECT 390.545 51.245 390.885 51.905 ;
        RECT 391.235 51.245 396.580 52.015 ;
        RECT 396.755 51.245 402.100 52.015 ;
        RECT 402.275 51.245 405.785 52.015 ;
        RECT 405.955 51.995 406.475 52.535 ;
        RECT 406.645 52.165 407.165 52.705 ;
        RECT 407.335 52.630 407.625 53.795 ;
        RECT 407.795 52.705 413.140 53.795 ;
        RECT 413.315 52.705 418.660 53.795 ;
        RECT 418.835 52.705 424.180 53.795 ;
        RECT 424.355 52.705 429.700 53.795 ;
        RECT 429.875 52.705 435.220 53.795 ;
        RECT 407.795 52.015 410.375 52.535 ;
        RECT 410.545 52.185 413.140 52.705 ;
        RECT 413.315 52.015 415.895 52.535 ;
        RECT 416.065 52.185 418.660 52.705 ;
        RECT 418.835 52.015 421.415 52.535 ;
        RECT 421.585 52.185 424.180 52.705 ;
        RECT 424.355 52.015 426.935 52.535 ;
        RECT 427.105 52.185 429.700 52.705 ;
        RECT 429.875 52.015 432.455 52.535 ;
        RECT 432.625 52.185 435.220 52.705 ;
        RECT 435.395 52.630 435.685 53.795 ;
        RECT 435.855 52.705 441.200 53.795 ;
        RECT 441.375 52.705 446.720 53.795 ;
        RECT 446.895 52.705 452.240 53.795 ;
        RECT 452.415 52.705 457.760 53.795 ;
        RECT 457.935 52.705 463.280 53.795 ;
        RECT 435.855 52.015 438.435 52.535 ;
        RECT 438.605 52.185 441.200 52.705 ;
        RECT 441.375 52.015 443.955 52.535 ;
        RECT 444.125 52.185 446.720 52.705 ;
        RECT 446.895 52.015 449.475 52.535 ;
        RECT 449.645 52.185 452.240 52.705 ;
        RECT 452.415 52.015 454.995 52.535 ;
        RECT 455.165 52.185 457.760 52.705 ;
        RECT 457.935 52.015 460.515 52.535 ;
        RECT 460.685 52.185 463.280 52.705 ;
        RECT 463.455 52.630 463.745 53.795 ;
        RECT 463.915 52.705 469.260 53.795 ;
        RECT 469.435 52.705 474.780 53.795 ;
        RECT 474.955 52.705 480.300 53.795 ;
        RECT 480.475 52.705 485.820 53.795 ;
        RECT 485.995 52.705 491.340 53.795 ;
        RECT 463.915 52.015 466.495 52.535 ;
        RECT 466.665 52.185 469.260 52.705 ;
        RECT 469.435 52.015 472.015 52.535 ;
        RECT 472.185 52.185 474.780 52.705 ;
        RECT 474.955 52.015 477.535 52.535 ;
        RECT 477.705 52.185 480.300 52.705 ;
        RECT 480.475 52.015 483.055 52.535 ;
        RECT 483.225 52.185 485.820 52.705 ;
        RECT 485.995 52.015 488.575 52.535 ;
        RECT 488.745 52.185 491.340 52.705 ;
        RECT 491.515 52.630 491.805 53.795 ;
        RECT 491.975 52.705 497.320 53.795 ;
        RECT 497.495 52.705 502.840 53.795 ;
        RECT 503.015 52.705 508.360 53.795 ;
        RECT 508.535 52.705 513.880 53.795 ;
        RECT 514.055 52.705 519.400 53.795 ;
        RECT 491.975 52.015 494.555 52.535 ;
        RECT 494.725 52.185 497.320 52.705 ;
        RECT 497.495 52.015 500.075 52.535 ;
        RECT 500.245 52.185 502.840 52.705 ;
        RECT 503.015 52.015 505.595 52.535 ;
        RECT 505.765 52.185 508.360 52.705 ;
        RECT 508.535 52.015 511.115 52.535 ;
        RECT 511.285 52.185 513.880 52.705 ;
        RECT 514.055 52.015 516.635 52.535 ;
        RECT 516.805 52.185 519.400 52.705 ;
        RECT 519.575 52.630 519.865 53.795 ;
        RECT 520.035 52.705 525.380 53.795 ;
        RECT 525.555 52.705 530.900 53.795 ;
        RECT 531.075 52.705 536.420 53.795 ;
        RECT 536.595 52.705 541.940 53.795 ;
        RECT 542.115 52.705 547.460 53.795 ;
        RECT 520.035 52.015 522.615 52.535 ;
        RECT 522.785 52.185 525.380 52.705 ;
        RECT 525.555 52.015 528.135 52.535 ;
        RECT 528.305 52.185 530.900 52.705 ;
        RECT 531.075 52.015 533.655 52.535 ;
        RECT 533.825 52.185 536.420 52.705 ;
        RECT 536.595 52.015 539.175 52.535 ;
        RECT 539.345 52.185 541.940 52.705 ;
        RECT 542.115 52.015 544.695 52.535 ;
        RECT 544.865 52.185 547.460 52.705 ;
        RECT 547.635 52.630 547.925 53.795 ;
        RECT 548.095 52.705 553.440 53.795 ;
        RECT 553.615 52.705 558.960 53.795 ;
        RECT 559.135 52.705 564.480 53.795 ;
        RECT 564.655 52.705 570.000 53.795 ;
        RECT 570.175 52.705 575.520 53.795 ;
        RECT 548.095 52.015 550.675 52.535 ;
        RECT 550.845 52.185 553.440 52.705 ;
        RECT 553.615 52.015 556.195 52.535 ;
        RECT 556.365 52.185 558.960 52.705 ;
        RECT 559.135 52.015 561.715 52.535 ;
        RECT 561.885 52.185 564.480 52.705 ;
        RECT 564.655 52.015 567.235 52.535 ;
        RECT 567.405 52.185 570.000 52.705 ;
        RECT 570.175 52.015 572.755 52.535 ;
        RECT 572.925 52.185 575.520 52.705 ;
        RECT 575.695 52.630 575.985 53.795 ;
        RECT 576.155 52.705 581.500 53.795 ;
        RECT 581.675 52.705 587.020 53.795 ;
        RECT 587.195 52.705 592.540 53.795 ;
        RECT 592.715 52.705 598.060 53.795 ;
        RECT 598.235 52.705 603.580 53.795 ;
        RECT 576.155 52.015 578.735 52.535 ;
        RECT 578.905 52.185 581.500 52.705 ;
        RECT 581.675 52.015 584.255 52.535 ;
        RECT 584.425 52.185 587.020 52.705 ;
        RECT 587.195 52.015 589.775 52.535 ;
        RECT 589.945 52.185 592.540 52.705 ;
        RECT 592.715 52.015 595.295 52.535 ;
        RECT 595.465 52.185 598.060 52.705 ;
        RECT 598.235 52.015 600.815 52.535 ;
        RECT 600.985 52.185 603.580 52.705 ;
        RECT 603.755 52.630 604.045 53.795 ;
        RECT 604.215 52.705 609.560 53.795 ;
        RECT 609.735 52.705 615.080 53.795 ;
        RECT 615.255 52.705 620.600 53.795 ;
        RECT 620.775 52.705 623.365 53.795 ;
        RECT 624.185 53.070 624.515 53.795 ;
        RECT 604.215 52.015 606.795 52.535 ;
        RECT 606.965 52.185 609.560 52.705 ;
        RECT 609.735 52.015 612.315 52.535 ;
        RECT 612.485 52.185 615.080 52.705 ;
        RECT 615.255 52.015 617.835 52.535 ;
        RECT 618.005 52.185 620.600 52.705 ;
        RECT 620.775 52.015 621.985 52.535 ;
        RECT 622.155 52.185 623.365 52.705 ;
        RECT 405.955 51.245 407.165 51.995 ;
        RECT 407.335 51.245 407.625 51.970 ;
        RECT 407.795 51.245 413.140 52.015 ;
        RECT 413.315 51.245 418.660 52.015 ;
        RECT 418.835 51.245 424.180 52.015 ;
        RECT 424.355 51.245 429.700 52.015 ;
        RECT 429.875 51.245 435.220 52.015 ;
        RECT 435.395 51.245 435.685 51.970 ;
        RECT 435.855 51.245 441.200 52.015 ;
        RECT 441.375 51.245 446.720 52.015 ;
        RECT 446.895 51.245 452.240 52.015 ;
        RECT 452.415 51.245 457.760 52.015 ;
        RECT 457.935 51.245 463.280 52.015 ;
        RECT 463.455 51.245 463.745 51.970 ;
        RECT 463.915 51.245 469.260 52.015 ;
        RECT 469.435 51.245 474.780 52.015 ;
        RECT 474.955 51.245 480.300 52.015 ;
        RECT 480.475 51.245 485.820 52.015 ;
        RECT 485.995 51.245 491.340 52.015 ;
        RECT 491.515 51.245 491.805 51.970 ;
        RECT 491.975 51.245 497.320 52.015 ;
        RECT 497.495 51.245 502.840 52.015 ;
        RECT 503.015 51.245 508.360 52.015 ;
        RECT 508.535 51.245 513.880 52.015 ;
        RECT 514.055 51.245 519.400 52.015 ;
        RECT 519.575 51.245 519.865 51.970 ;
        RECT 520.035 51.245 525.380 52.015 ;
        RECT 525.555 51.245 530.900 52.015 ;
        RECT 531.075 51.245 536.420 52.015 ;
        RECT 536.595 51.245 541.940 52.015 ;
        RECT 542.115 51.245 547.460 52.015 ;
        RECT 547.635 51.245 547.925 51.970 ;
        RECT 548.095 51.245 553.440 52.015 ;
        RECT 553.615 51.245 558.960 52.015 ;
        RECT 559.135 51.245 564.480 52.015 ;
        RECT 564.655 51.245 570.000 52.015 ;
        RECT 570.175 51.245 575.520 52.015 ;
        RECT 575.695 51.245 575.985 51.970 ;
        RECT 576.155 51.245 581.500 52.015 ;
        RECT 581.675 51.245 587.020 52.015 ;
        RECT 587.195 51.245 592.540 52.015 ;
        RECT 592.715 51.245 598.060 52.015 ;
        RECT 598.235 51.245 603.580 52.015 ;
        RECT 603.755 51.245 604.045 51.970 ;
        RECT 604.215 51.245 609.560 52.015 ;
        RECT 609.735 51.245 615.080 52.015 ;
        RECT 615.255 51.245 620.600 52.015 ;
        RECT 620.775 51.245 623.365 52.015 ;
        RECT 623.995 51.415 624.515 52.900 ;
        RECT 624.685 52.075 625.205 53.625 ;
        RECT 625.375 52.705 628.885 53.795 ;
        RECT 625.375 52.015 627.025 52.535 ;
        RECT 627.195 52.185 628.885 52.705 ;
        RECT 629.975 52.705 631.185 53.795 ;
        RECT 629.975 52.165 630.495 52.705 ;
        RECT 624.685 51.245 625.025 51.905 ;
        RECT 625.375 51.245 628.885 52.015 ;
        RECT 630.665 51.995 631.185 52.535 ;
        RECT 629.975 51.245 631.185 51.995 ;
        RECT 42.470 51.075 631.270 51.245 ;
        RECT 42.555 50.325 43.765 51.075 ;
        RECT 42.555 49.785 43.075 50.325 ;
        RECT 43.935 50.305 49.280 51.075 ;
        RECT 49.455 50.305 54.800 51.075 ;
        RECT 54.975 50.305 56.645 51.075 ;
        RECT 56.815 50.350 57.105 51.075 ;
        RECT 57.275 50.305 62.620 51.075 ;
        RECT 62.795 50.305 68.140 51.075 ;
        RECT 68.315 50.305 71.825 51.075 ;
        RECT 43.245 49.615 43.765 50.155 ;
        RECT 43.935 49.785 46.515 50.305 ;
        RECT 46.685 49.615 49.280 50.135 ;
        RECT 49.455 49.785 52.035 50.305 ;
        RECT 52.205 49.615 54.800 50.135 ;
        RECT 54.975 49.785 55.725 50.305 ;
        RECT 55.895 49.615 56.645 50.135 ;
        RECT 57.275 49.785 59.855 50.305 ;
        RECT 42.555 48.525 43.765 49.615 ;
        RECT 43.935 48.525 49.280 49.615 ;
        RECT 49.455 48.525 54.800 49.615 ;
        RECT 54.975 48.525 56.645 49.615 ;
        RECT 56.815 48.525 57.105 49.690 ;
        RECT 60.025 49.615 62.620 50.135 ;
        RECT 62.795 49.785 65.375 50.305 ;
        RECT 65.545 49.615 68.140 50.135 ;
        RECT 68.315 49.785 69.965 50.305 ;
        RECT 72.955 50.255 73.185 51.075 ;
        RECT 73.355 50.275 73.685 50.905 ;
        RECT 70.135 49.615 71.825 50.135 ;
        RECT 72.935 49.835 73.265 50.085 ;
        RECT 73.435 49.675 73.685 50.275 ;
        RECT 73.855 50.255 74.065 51.075 ;
        RECT 74.295 50.305 77.805 51.075 ;
        RECT 77.995 50.565 78.235 51.075 ;
        RECT 74.295 49.785 75.945 50.305 ;
        RECT 57.275 48.525 62.620 49.615 ;
        RECT 62.795 48.525 68.140 49.615 ;
        RECT 68.315 48.525 71.825 49.615 ;
        RECT 72.955 48.525 73.185 49.665 ;
        RECT 73.355 48.695 73.685 49.675 ;
        RECT 73.855 48.525 74.065 49.665 ;
        RECT 76.115 49.615 77.805 50.135 ;
        RECT 77.980 49.835 78.235 50.395 ;
        RECT 78.405 50.335 78.735 50.870 ;
        RECT 78.950 50.335 79.120 51.075 ;
        RECT 79.330 50.425 79.660 50.895 ;
        RECT 79.830 50.595 80.000 51.075 ;
        RECT 80.170 50.425 80.500 50.895 ;
        RECT 80.670 50.595 80.840 51.075 ;
        RECT 78.405 49.665 78.585 50.335 ;
        RECT 79.330 50.255 81.025 50.425 ;
        RECT 78.755 49.835 79.130 50.165 ;
        RECT 79.300 49.915 80.510 50.085 ;
        RECT 79.300 49.665 79.505 49.915 ;
        RECT 80.680 49.665 81.025 50.255 ;
        RECT 81.195 50.305 84.705 51.075 ;
        RECT 84.875 50.350 85.165 51.075 ;
        RECT 85.885 50.525 86.055 50.905 ;
        RECT 86.270 50.695 86.600 51.075 ;
        RECT 85.885 50.355 86.600 50.525 ;
        RECT 81.195 49.785 82.845 50.305 ;
        RECT 74.295 48.525 77.805 49.615 ;
        RECT 78.045 49.495 79.505 49.665 ;
        RECT 80.170 49.495 81.025 49.665 ;
        RECT 83.015 49.615 84.705 50.135 ;
        RECT 85.795 49.805 86.150 50.175 ;
        RECT 86.430 50.165 86.600 50.355 ;
        RECT 86.770 50.330 87.025 50.905 ;
        RECT 86.430 49.835 86.685 50.165 ;
        RECT 78.045 48.695 78.405 49.495 ;
        RECT 80.170 49.325 80.500 49.495 ;
        RECT 78.950 48.525 79.120 49.325 ;
        RECT 79.330 49.155 80.500 49.325 ;
        RECT 79.330 48.695 79.660 49.155 ;
        RECT 79.830 48.525 80.000 48.985 ;
        RECT 80.170 48.695 80.500 49.155 ;
        RECT 80.670 48.525 80.840 49.325 ;
        RECT 81.195 48.525 84.705 49.615 ;
        RECT 84.875 48.525 85.165 49.690 ;
        RECT 86.430 49.625 86.600 49.835 ;
        RECT 85.885 49.455 86.600 49.625 ;
        RECT 86.855 49.600 87.025 50.330 ;
        RECT 87.200 50.235 87.460 51.075 ;
        RECT 87.635 50.305 91.145 51.075 ;
        RECT 91.405 50.525 91.575 50.815 ;
        RECT 91.745 50.695 92.075 51.075 ;
        RECT 91.405 50.355 92.070 50.525 ;
        RECT 87.635 49.785 89.285 50.305 ;
        RECT 85.885 48.695 86.055 49.455 ;
        RECT 86.270 48.525 86.600 49.285 ;
        RECT 86.770 48.695 87.025 49.600 ;
        RECT 87.200 48.525 87.460 49.675 ;
        RECT 89.455 49.615 91.145 50.135 ;
        RECT 87.635 48.525 91.145 49.615 ;
        RECT 91.320 49.535 91.670 50.185 ;
        RECT 91.840 49.365 92.070 50.355 ;
        RECT 91.405 49.195 92.070 49.365 ;
        RECT 91.405 48.695 91.575 49.195 ;
        RECT 91.745 48.525 92.075 49.025 ;
        RECT 92.245 48.695 92.470 50.815 ;
        RECT 92.685 50.615 92.935 51.075 ;
        RECT 93.120 50.625 93.450 50.795 ;
        RECT 93.630 50.625 94.380 50.795 ;
        RECT 92.670 49.495 92.950 50.095 ;
        RECT 93.120 49.095 93.290 50.625 ;
        RECT 93.460 50.125 94.040 50.455 ;
        RECT 93.460 49.255 93.700 50.125 ;
        RECT 94.210 49.845 94.380 50.625 ;
        RECT 94.630 50.575 95.000 51.075 ;
        RECT 95.180 50.625 95.640 50.795 ;
        RECT 95.870 50.625 96.540 50.795 ;
        RECT 95.180 50.395 95.350 50.625 ;
        RECT 94.550 50.095 95.350 50.395 ;
        RECT 95.520 50.125 96.070 50.455 ;
        RECT 94.550 50.065 94.720 50.095 ;
        RECT 94.840 49.845 95.010 49.915 ;
        RECT 94.210 49.675 95.010 49.845 ;
        RECT 94.500 49.585 95.010 49.675 ;
        RECT 93.890 49.150 94.330 49.505 ;
        RECT 92.670 48.525 92.935 48.985 ;
        RECT 93.120 48.720 93.355 49.095 ;
        RECT 94.500 48.970 94.670 49.585 ;
        RECT 93.600 48.800 94.670 48.970 ;
        RECT 94.840 48.525 95.010 49.325 ;
        RECT 95.180 49.025 95.350 50.095 ;
        RECT 95.520 49.195 95.710 49.915 ;
        RECT 95.880 49.585 96.070 50.125 ;
        RECT 96.370 50.085 96.540 50.625 ;
        RECT 96.855 50.545 97.025 51.075 ;
        RECT 97.320 50.425 97.680 50.865 ;
        RECT 97.855 50.595 98.025 51.075 ;
        RECT 98.215 50.430 98.550 50.855 ;
        RECT 98.725 50.600 98.895 51.075 ;
        RECT 99.070 50.430 99.405 50.855 ;
        RECT 99.575 50.600 99.745 51.075 ;
        RECT 97.320 50.255 97.820 50.425 ;
        RECT 98.215 50.260 99.885 50.430 ;
        RECT 97.650 50.085 97.820 50.255 ;
        RECT 96.370 49.915 97.460 50.085 ;
        RECT 97.650 49.915 99.470 50.085 ;
        RECT 95.880 49.255 96.200 49.585 ;
        RECT 95.180 48.695 95.430 49.025 ;
        RECT 96.370 48.995 96.540 49.915 ;
        RECT 97.650 49.660 97.820 49.915 ;
        RECT 99.640 49.695 99.885 50.260 ;
        RECT 100.055 50.305 103.565 51.075 ;
        RECT 103.735 50.325 104.945 51.075 ;
        RECT 100.055 49.785 101.705 50.305 ;
        RECT 96.710 49.490 97.820 49.660 ;
        RECT 98.215 49.525 99.885 49.695 ;
        RECT 101.875 49.615 103.565 50.135 ;
        RECT 103.735 49.785 104.255 50.325 ;
        RECT 105.120 50.255 105.395 51.075 ;
        RECT 105.565 50.435 105.895 50.905 ;
        RECT 106.065 50.605 106.235 51.075 ;
        RECT 106.405 50.435 106.735 50.905 ;
        RECT 106.905 50.605 107.075 51.075 ;
        RECT 107.245 50.435 107.575 50.905 ;
        RECT 107.745 50.605 107.915 51.075 ;
        RECT 108.085 50.435 108.415 50.905 ;
        RECT 108.585 50.605 108.870 51.075 ;
        RECT 105.565 50.255 109.085 50.435 ;
        RECT 104.425 49.615 104.945 50.155 ;
        RECT 105.170 49.885 106.830 50.085 ;
        RECT 107.150 49.885 108.515 50.085 ;
        RECT 108.685 49.715 109.085 50.255 ;
        RECT 109.255 50.305 112.765 51.075 ;
        RECT 112.935 50.350 113.225 51.075 ;
        RECT 113.485 50.525 113.655 50.815 ;
        RECT 113.825 50.695 114.155 51.075 ;
        RECT 113.485 50.355 114.150 50.525 ;
        RECT 109.255 49.785 110.905 50.305 ;
        RECT 96.710 49.330 97.570 49.490 ;
        RECT 95.655 48.825 96.540 48.995 ;
        RECT 96.720 48.525 96.935 49.025 ;
        RECT 97.400 48.705 97.570 49.330 ;
        RECT 97.855 48.525 98.035 49.305 ;
        RECT 98.215 48.765 98.550 49.525 ;
        RECT 98.730 48.525 98.900 49.355 ;
        RECT 99.070 48.765 99.400 49.525 ;
        RECT 99.570 48.525 99.740 49.355 ;
        RECT 100.055 48.525 103.565 49.615 ;
        RECT 103.735 48.525 104.945 49.615 ;
        RECT 105.120 49.495 107.155 49.705 ;
        RECT 105.120 48.695 105.395 49.495 ;
        RECT 105.565 48.525 105.895 49.325 ;
        RECT 106.065 48.695 106.235 49.495 ;
        RECT 106.405 48.525 106.655 49.325 ;
        RECT 106.825 48.865 107.155 49.495 ;
        RECT 107.325 49.415 109.085 49.715 ;
        RECT 111.075 49.615 112.765 50.135 ;
        RECT 107.325 49.035 107.495 49.415 ;
        RECT 107.665 48.865 107.995 49.225 ;
        RECT 108.165 49.035 108.335 49.415 ;
        RECT 108.505 48.865 108.920 49.245 ;
        RECT 106.825 48.695 108.920 48.865 ;
        RECT 109.255 48.525 112.765 49.615 ;
        RECT 112.935 48.525 113.225 49.690 ;
        RECT 113.400 49.535 113.750 50.185 ;
        RECT 113.920 49.365 114.150 50.355 ;
        RECT 113.485 49.195 114.150 49.365 ;
        RECT 113.485 48.695 113.655 49.195 ;
        RECT 113.825 48.525 114.155 49.025 ;
        RECT 114.325 48.695 114.550 50.815 ;
        RECT 114.765 50.615 115.015 51.075 ;
        RECT 115.200 50.625 115.530 50.795 ;
        RECT 115.710 50.625 116.460 50.795 ;
        RECT 114.750 49.495 115.030 50.095 ;
        RECT 115.200 49.095 115.370 50.625 ;
        RECT 115.540 50.125 116.120 50.455 ;
        RECT 115.540 49.255 115.780 50.125 ;
        RECT 116.290 49.845 116.460 50.625 ;
        RECT 116.710 50.575 117.080 51.075 ;
        RECT 117.260 50.625 117.720 50.795 ;
        RECT 117.950 50.625 118.620 50.795 ;
        RECT 117.260 50.395 117.430 50.625 ;
        RECT 116.630 50.095 117.430 50.395 ;
        RECT 117.600 50.125 118.150 50.455 ;
        RECT 116.630 50.065 116.800 50.095 ;
        RECT 116.920 49.845 117.090 49.915 ;
        RECT 116.290 49.675 117.090 49.845 ;
        RECT 116.580 49.585 117.090 49.675 ;
        RECT 115.970 49.150 116.410 49.505 ;
        RECT 114.750 48.525 115.015 48.985 ;
        RECT 115.200 48.720 115.435 49.095 ;
        RECT 116.580 48.970 116.750 49.585 ;
        RECT 115.680 48.800 116.750 48.970 ;
        RECT 116.920 48.525 117.090 49.325 ;
        RECT 117.260 49.025 117.430 50.095 ;
        RECT 117.600 49.195 117.790 49.915 ;
        RECT 117.960 49.585 118.150 50.125 ;
        RECT 118.450 50.085 118.620 50.625 ;
        RECT 118.935 50.545 119.105 51.075 ;
        RECT 119.400 50.425 119.760 50.865 ;
        RECT 119.935 50.595 120.105 51.075 ;
        RECT 120.295 50.430 120.630 50.855 ;
        RECT 120.805 50.600 120.975 51.075 ;
        RECT 121.150 50.430 121.485 50.855 ;
        RECT 121.655 50.600 121.825 51.075 ;
        RECT 119.400 50.255 119.900 50.425 ;
        RECT 120.295 50.260 121.965 50.430 ;
        RECT 119.730 50.085 119.900 50.255 ;
        RECT 118.450 49.915 119.540 50.085 ;
        RECT 119.730 49.915 121.550 50.085 ;
        RECT 117.960 49.255 118.280 49.585 ;
        RECT 117.260 48.695 117.510 49.025 ;
        RECT 118.450 48.995 118.620 49.915 ;
        RECT 119.730 49.660 119.900 49.915 ;
        RECT 121.720 49.695 121.965 50.260 ;
        RECT 122.135 50.305 125.645 51.075 ;
        RECT 125.905 50.525 126.075 50.815 ;
        RECT 126.245 50.695 126.575 51.075 ;
        RECT 125.905 50.355 126.570 50.525 ;
        RECT 122.135 49.785 123.785 50.305 ;
        RECT 118.790 49.490 119.900 49.660 ;
        RECT 120.295 49.525 121.965 49.695 ;
        RECT 123.955 49.615 125.645 50.135 ;
        RECT 118.790 49.330 119.650 49.490 ;
        RECT 117.735 48.825 118.620 48.995 ;
        RECT 118.800 48.525 119.015 49.025 ;
        RECT 119.480 48.705 119.650 49.330 ;
        RECT 119.935 48.525 120.115 49.305 ;
        RECT 120.295 48.765 120.630 49.525 ;
        RECT 120.810 48.525 120.980 49.355 ;
        RECT 121.150 48.765 121.480 49.525 ;
        RECT 121.650 48.525 121.820 49.355 ;
        RECT 122.135 48.525 125.645 49.615 ;
        RECT 125.820 49.535 126.170 50.185 ;
        RECT 126.340 49.365 126.570 50.355 ;
        RECT 125.905 49.195 126.570 49.365 ;
        RECT 125.905 48.695 126.075 49.195 ;
        RECT 126.245 48.525 126.575 49.025 ;
        RECT 126.745 48.695 126.970 50.815 ;
        RECT 127.185 50.615 127.435 51.075 ;
        RECT 127.620 50.625 127.950 50.795 ;
        RECT 128.130 50.625 128.880 50.795 ;
        RECT 127.170 49.495 127.450 50.095 ;
        RECT 127.620 49.095 127.790 50.625 ;
        RECT 127.960 50.125 128.540 50.455 ;
        RECT 127.960 49.255 128.200 50.125 ;
        RECT 128.710 49.845 128.880 50.625 ;
        RECT 129.130 50.575 129.500 51.075 ;
        RECT 129.680 50.625 130.140 50.795 ;
        RECT 130.370 50.625 131.040 50.795 ;
        RECT 129.680 50.395 129.850 50.625 ;
        RECT 129.050 50.095 129.850 50.395 ;
        RECT 130.020 50.125 130.570 50.455 ;
        RECT 129.050 50.065 129.220 50.095 ;
        RECT 129.340 49.845 129.510 49.915 ;
        RECT 128.710 49.675 129.510 49.845 ;
        RECT 129.000 49.585 129.510 49.675 ;
        RECT 128.390 49.150 128.830 49.505 ;
        RECT 127.170 48.525 127.435 48.985 ;
        RECT 127.620 48.720 127.855 49.095 ;
        RECT 129.000 48.970 129.170 49.585 ;
        RECT 128.100 48.800 129.170 48.970 ;
        RECT 129.340 48.525 129.510 49.325 ;
        RECT 129.680 49.025 129.850 50.095 ;
        RECT 130.020 49.195 130.210 49.915 ;
        RECT 130.380 49.585 130.570 50.125 ;
        RECT 130.870 50.085 131.040 50.625 ;
        RECT 131.355 50.545 131.525 51.075 ;
        RECT 131.820 50.425 132.180 50.865 ;
        RECT 132.355 50.595 132.525 51.075 ;
        RECT 132.715 50.430 133.050 50.855 ;
        RECT 133.225 50.600 133.395 51.075 ;
        RECT 133.570 50.430 133.905 50.855 ;
        RECT 134.075 50.600 134.245 51.075 ;
        RECT 131.820 50.255 132.320 50.425 ;
        RECT 132.715 50.260 134.385 50.430 ;
        RECT 132.150 50.085 132.320 50.255 ;
        RECT 130.870 49.915 131.960 50.085 ;
        RECT 132.150 49.915 133.970 50.085 ;
        RECT 130.380 49.255 130.700 49.585 ;
        RECT 129.680 48.695 129.930 49.025 ;
        RECT 130.870 48.995 131.040 49.915 ;
        RECT 132.150 49.660 132.320 49.915 ;
        RECT 134.140 49.695 134.385 50.260 ;
        RECT 134.555 50.305 139.900 51.075 ;
        RECT 140.995 50.350 141.285 51.075 ;
        RECT 141.545 50.525 141.715 50.815 ;
        RECT 141.885 50.695 142.215 51.075 ;
        RECT 141.545 50.355 142.210 50.525 ;
        RECT 134.555 49.785 137.135 50.305 ;
        RECT 131.210 49.490 132.320 49.660 ;
        RECT 132.715 49.525 134.385 49.695 ;
        RECT 137.305 49.615 139.900 50.135 ;
        RECT 131.210 49.330 132.070 49.490 ;
        RECT 130.155 48.825 131.040 48.995 ;
        RECT 131.220 48.525 131.435 49.025 ;
        RECT 131.900 48.705 132.070 49.330 ;
        RECT 132.355 48.525 132.535 49.305 ;
        RECT 132.715 48.765 133.050 49.525 ;
        RECT 133.230 48.525 133.400 49.355 ;
        RECT 133.570 48.765 133.900 49.525 ;
        RECT 134.070 48.525 134.240 49.355 ;
        RECT 134.555 48.525 139.900 49.615 ;
        RECT 140.995 48.525 141.285 49.690 ;
        RECT 141.460 49.535 141.810 50.185 ;
        RECT 141.980 49.365 142.210 50.355 ;
        RECT 141.545 49.195 142.210 49.365 ;
        RECT 141.545 48.695 141.715 49.195 ;
        RECT 141.885 48.525 142.215 49.025 ;
        RECT 142.385 48.695 142.610 50.815 ;
        RECT 142.825 50.615 143.075 51.075 ;
        RECT 143.260 50.625 143.590 50.795 ;
        RECT 143.770 50.625 144.520 50.795 ;
        RECT 142.810 49.495 143.090 50.095 ;
        RECT 143.260 49.095 143.430 50.625 ;
        RECT 143.600 50.125 144.180 50.455 ;
        RECT 143.600 49.255 143.840 50.125 ;
        RECT 144.350 49.845 144.520 50.625 ;
        RECT 144.770 50.575 145.140 51.075 ;
        RECT 145.320 50.625 145.780 50.795 ;
        RECT 146.010 50.625 146.680 50.795 ;
        RECT 145.320 50.395 145.490 50.625 ;
        RECT 144.690 50.095 145.490 50.395 ;
        RECT 145.660 50.125 146.210 50.455 ;
        RECT 144.690 50.065 144.860 50.095 ;
        RECT 144.980 49.845 145.150 49.915 ;
        RECT 144.350 49.675 145.150 49.845 ;
        RECT 144.640 49.585 145.150 49.675 ;
        RECT 144.030 49.150 144.470 49.505 ;
        RECT 142.810 48.525 143.075 48.985 ;
        RECT 143.260 48.720 143.495 49.095 ;
        RECT 144.640 48.970 144.810 49.585 ;
        RECT 143.740 48.800 144.810 48.970 ;
        RECT 144.980 48.525 145.150 49.325 ;
        RECT 145.320 49.025 145.490 50.095 ;
        RECT 145.660 49.195 145.850 49.915 ;
        RECT 146.020 49.585 146.210 50.125 ;
        RECT 146.510 50.085 146.680 50.625 ;
        RECT 146.995 50.545 147.165 51.075 ;
        RECT 147.460 50.425 147.820 50.865 ;
        RECT 147.995 50.595 148.165 51.075 ;
        RECT 148.865 50.600 149.035 51.075 ;
        RECT 149.715 50.600 149.885 51.075 ;
        RECT 147.460 50.255 147.960 50.425 ;
        RECT 147.790 50.085 147.960 50.255 ;
        RECT 150.195 50.305 153.705 51.075 ;
        RECT 153.965 50.525 154.135 50.815 ;
        RECT 154.305 50.695 154.635 51.075 ;
        RECT 153.965 50.355 154.630 50.525 ;
        RECT 146.510 49.915 147.600 50.085 ;
        RECT 147.790 49.915 149.610 50.085 ;
        RECT 146.020 49.255 146.340 49.585 ;
        RECT 145.320 48.695 145.570 49.025 ;
        RECT 146.510 48.995 146.680 49.915 ;
        RECT 147.790 49.660 147.960 49.915 ;
        RECT 150.195 49.785 151.845 50.305 ;
        RECT 146.850 49.490 147.960 49.660 ;
        RECT 152.015 49.615 153.705 50.135 ;
        RECT 146.850 49.330 147.710 49.490 ;
        RECT 145.795 48.825 146.680 48.995 ;
        RECT 146.860 48.525 147.075 49.025 ;
        RECT 147.540 48.705 147.710 49.330 ;
        RECT 147.995 48.525 148.175 49.305 ;
        RECT 148.870 48.525 149.040 49.355 ;
        RECT 149.710 48.525 149.880 49.355 ;
        RECT 150.195 48.525 153.705 49.615 ;
        RECT 153.880 49.535 154.230 50.185 ;
        RECT 154.400 49.365 154.630 50.355 ;
        RECT 153.965 49.195 154.630 49.365 ;
        RECT 153.965 48.695 154.135 49.195 ;
        RECT 154.305 48.525 154.635 49.025 ;
        RECT 154.805 48.695 155.030 50.815 ;
        RECT 155.245 50.615 155.495 51.075 ;
        RECT 155.680 50.625 156.010 50.795 ;
        RECT 156.190 50.625 156.940 50.795 ;
        RECT 155.230 49.495 155.510 50.095 ;
        RECT 155.680 49.095 155.850 50.625 ;
        RECT 156.020 50.125 156.600 50.455 ;
        RECT 156.020 49.255 156.260 50.125 ;
        RECT 156.770 49.845 156.940 50.625 ;
        RECT 157.190 50.575 157.560 51.075 ;
        RECT 157.740 50.625 158.200 50.795 ;
        RECT 158.430 50.625 159.100 50.795 ;
        RECT 157.740 50.395 157.910 50.625 ;
        RECT 157.110 50.095 157.910 50.395 ;
        RECT 158.080 50.125 158.630 50.455 ;
        RECT 157.110 50.065 157.280 50.095 ;
        RECT 157.400 49.845 157.570 49.915 ;
        RECT 156.770 49.675 157.570 49.845 ;
        RECT 157.060 49.585 157.570 49.675 ;
        RECT 156.450 49.150 156.890 49.505 ;
        RECT 155.230 48.525 155.495 48.985 ;
        RECT 155.680 48.720 155.915 49.095 ;
        RECT 157.060 48.970 157.230 49.585 ;
        RECT 156.160 48.800 157.230 48.970 ;
        RECT 157.400 48.525 157.570 49.325 ;
        RECT 157.740 49.025 157.910 50.095 ;
        RECT 158.080 49.195 158.270 49.915 ;
        RECT 158.440 49.585 158.630 50.125 ;
        RECT 158.930 50.085 159.100 50.625 ;
        RECT 159.415 50.545 159.585 51.075 ;
        RECT 159.880 50.425 160.240 50.865 ;
        RECT 160.415 50.595 160.585 51.075 ;
        RECT 160.775 50.430 161.110 50.855 ;
        RECT 161.285 50.600 161.455 51.075 ;
        RECT 161.630 50.430 161.965 50.855 ;
        RECT 162.135 50.600 162.305 51.075 ;
        RECT 159.880 50.255 160.380 50.425 ;
        RECT 160.775 50.260 162.445 50.430 ;
        RECT 160.210 50.085 160.380 50.255 ;
        RECT 158.930 49.915 160.020 50.085 ;
        RECT 160.210 49.915 162.030 50.085 ;
        RECT 158.440 49.255 158.760 49.585 ;
        RECT 157.740 48.695 157.990 49.025 ;
        RECT 158.930 48.995 159.100 49.915 ;
        RECT 160.210 49.660 160.380 49.915 ;
        RECT 162.200 49.695 162.445 50.260 ;
        RECT 162.615 50.305 167.960 51.075 ;
        RECT 169.055 50.350 169.345 51.075 ;
        RECT 169.605 50.525 169.775 50.815 ;
        RECT 169.945 50.695 170.275 51.075 ;
        RECT 169.605 50.355 170.270 50.525 ;
        RECT 162.615 49.785 165.195 50.305 ;
        RECT 159.270 49.490 160.380 49.660 ;
        RECT 160.775 49.525 162.445 49.695 ;
        RECT 165.365 49.615 167.960 50.135 ;
        RECT 159.270 49.330 160.130 49.490 ;
        RECT 158.215 48.825 159.100 48.995 ;
        RECT 159.280 48.525 159.495 49.025 ;
        RECT 159.960 48.705 160.130 49.330 ;
        RECT 160.415 48.525 160.595 49.305 ;
        RECT 160.775 48.765 161.110 49.525 ;
        RECT 161.290 48.525 161.460 49.355 ;
        RECT 161.630 48.765 161.960 49.525 ;
        RECT 162.130 48.525 162.300 49.355 ;
        RECT 162.615 48.525 167.960 49.615 ;
        RECT 169.055 48.525 169.345 49.690 ;
        RECT 169.520 49.535 169.870 50.185 ;
        RECT 170.040 49.365 170.270 50.355 ;
        RECT 169.605 49.195 170.270 49.365 ;
        RECT 169.605 48.695 169.775 49.195 ;
        RECT 169.945 48.525 170.275 49.025 ;
        RECT 170.445 48.695 170.670 50.815 ;
        RECT 170.885 50.615 171.135 51.075 ;
        RECT 171.320 50.625 171.650 50.795 ;
        RECT 171.830 50.625 172.580 50.795 ;
        RECT 170.870 49.495 171.150 50.095 ;
        RECT 171.320 49.095 171.490 50.625 ;
        RECT 171.660 50.125 172.240 50.455 ;
        RECT 171.660 49.255 171.900 50.125 ;
        RECT 172.410 49.845 172.580 50.625 ;
        RECT 172.830 50.575 173.200 51.075 ;
        RECT 173.380 50.625 173.840 50.795 ;
        RECT 174.070 50.625 174.740 50.795 ;
        RECT 173.380 50.395 173.550 50.625 ;
        RECT 172.750 50.095 173.550 50.395 ;
        RECT 173.720 50.125 174.270 50.455 ;
        RECT 172.750 50.065 172.920 50.095 ;
        RECT 173.040 49.845 173.210 49.915 ;
        RECT 172.410 49.675 173.210 49.845 ;
        RECT 172.700 49.585 173.210 49.675 ;
        RECT 172.090 49.150 172.530 49.505 ;
        RECT 170.870 48.525 171.135 48.985 ;
        RECT 171.320 48.720 171.555 49.095 ;
        RECT 172.700 48.970 172.870 49.585 ;
        RECT 171.800 48.800 172.870 48.970 ;
        RECT 173.040 48.525 173.210 49.325 ;
        RECT 173.380 49.025 173.550 50.095 ;
        RECT 173.720 49.195 173.910 49.915 ;
        RECT 174.080 49.585 174.270 50.125 ;
        RECT 174.570 50.085 174.740 50.625 ;
        RECT 175.055 50.545 175.225 51.075 ;
        RECT 175.520 50.425 175.880 50.865 ;
        RECT 176.055 50.595 176.225 51.075 ;
        RECT 176.415 50.430 176.750 50.855 ;
        RECT 176.925 50.600 177.095 51.075 ;
        RECT 177.270 50.430 177.605 50.855 ;
        RECT 177.775 50.600 177.945 51.075 ;
        RECT 175.520 50.255 176.020 50.425 ;
        RECT 176.415 50.260 178.085 50.430 ;
        RECT 175.850 50.085 176.020 50.255 ;
        RECT 174.570 49.915 175.660 50.085 ;
        RECT 175.850 49.915 177.670 50.085 ;
        RECT 174.080 49.255 174.400 49.585 ;
        RECT 173.380 48.695 173.630 49.025 ;
        RECT 174.570 48.995 174.740 49.915 ;
        RECT 175.850 49.660 176.020 49.915 ;
        RECT 177.840 49.695 178.085 50.260 ;
        RECT 178.255 50.305 181.765 51.075 ;
        RECT 182.025 50.525 182.195 50.815 ;
        RECT 182.365 50.695 182.695 51.075 ;
        RECT 182.025 50.355 182.690 50.525 ;
        RECT 178.255 49.785 179.905 50.305 ;
        RECT 174.910 49.490 176.020 49.660 ;
        RECT 176.415 49.525 178.085 49.695 ;
        RECT 180.075 49.615 181.765 50.135 ;
        RECT 174.910 49.330 175.770 49.490 ;
        RECT 173.855 48.825 174.740 48.995 ;
        RECT 174.920 48.525 175.135 49.025 ;
        RECT 175.600 48.705 175.770 49.330 ;
        RECT 176.055 48.525 176.235 49.305 ;
        RECT 176.415 48.765 176.750 49.525 ;
        RECT 176.930 48.525 177.100 49.355 ;
        RECT 177.270 48.765 177.600 49.525 ;
        RECT 177.770 48.525 177.940 49.355 ;
        RECT 178.255 48.525 181.765 49.615 ;
        RECT 181.940 49.535 182.290 50.185 ;
        RECT 182.460 49.365 182.690 50.355 ;
        RECT 182.025 49.195 182.690 49.365 ;
        RECT 182.025 48.695 182.195 49.195 ;
        RECT 182.365 48.525 182.695 49.025 ;
        RECT 182.865 48.695 183.090 50.815 ;
        RECT 183.305 50.615 183.555 51.075 ;
        RECT 183.740 50.625 184.070 50.795 ;
        RECT 184.250 50.625 185.000 50.795 ;
        RECT 183.290 49.495 183.570 50.095 ;
        RECT 183.740 49.095 183.910 50.625 ;
        RECT 184.080 50.125 184.660 50.455 ;
        RECT 184.080 49.255 184.320 50.125 ;
        RECT 184.830 49.845 185.000 50.625 ;
        RECT 185.250 50.575 185.620 51.075 ;
        RECT 185.800 50.625 186.260 50.795 ;
        RECT 186.490 50.625 187.160 50.795 ;
        RECT 185.800 50.395 185.970 50.625 ;
        RECT 185.170 50.095 185.970 50.395 ;
        RECT 186.140 50.125 186.690 50.455 ;
        RECT 185.170 50.065 185.340 50.095 ;
        RECT 185.460 49.845 185.630 49.915 ;
        RECT 184.830 49.675 185.630 49.845 ;
        RECT 185.120 49.585 185.630 49.675 ;
        RECT 184.510 49.150 184.950 49.505 ;
        RECT 183.290 48.525 183.555 48.985 ;
        RECT 183.740 48.720 183.975 49.095 ;
        RECT 185.120 48.970 185.290 49.585 ;
        RECT 184.220 48.800 185.290 48.970 ;
        RECT 185.460 48.525 185.630 49.325 ;
        RECT 185.800 49.025 185.970 50.095 ;
        RECT 186.140 49.195 186.330 49.915 ;
        RECT 186.500 49.585 186.690 50.125 ;
        RECT 186.990 50.085 187.160 50.625 ;
        RECT 187.475 50.545 187.645 51.075 ;
        RECT 187.940 50.425 188.300 50.865 ;
        RECT 188.475 50.595 188.645 51.075 ;
        RECT 188.835 50.430 189.170 50.855 ;
        RECT 189.345 50.600 189.515 51.075 ;
        RECT 189.690 50.430 190.025 50.855 ;
        RECT 190.195 50.600 190.365 51.075 ;
        RECT 187.940 50.255 188.440 50.425 ;
        RECT 188.835 50.260 190.505 50.430 ;
        RECT 188.270 50.085 188.440 50.255 ;
        RECT 186.990 49.915 188.080 50.085 ;
        RECT 188.270 49.915 190.090 50.085 ;
        RECT 186.500 49.255 186.820 49.585 ;
        RECT 185.800 48.695 186.050 49.025 ;
        RECT 186.990 48.995 187.160 49.915 ;
        RECT 188.270 49.660 188.440 49.915 ;
        RECT 190.260 49.695 190.505 50.260 ;
        RECT 190.675 50.305 194.185 51.075 ;
        RECT 194.355 50.400 194.615 50.905 ;
        RECT 194.795 50.695 195.125 51.075 ;
        RECT 195.305 50.525 195.475 50.905 ;
        RECT 190.675 49.785 192.325 50.305 ;
        RECT 187.330 49.490 188.440 49.660 ;
        RECT 188.835 49.525 190.505 49.695 ;
        RECT 192.495 49.615 194.185 50.135 ;
        RECT 187.330 49.330 188.190 49.490 ;
        RECT 186.275 48.825 187.160 48.995 ;
        RECT 187.340 48.525 187.555 49.025 ;
        RECT 188.020 48.705 188.190 49.330 ;
        RECT 188.475 48.525 188.655 49.305 ;
        RECT 188.835 48.765 189.170 49.525 ;
        RECT 189.350 48.525 189.520 49.355 ;
        RECT 189.690 48.765 190.020 49.525 ;
        RECT 190.190 48.525 190.360 49.355 ;
        RECT 190.675 48.525 194.185 49.615 ;
        RECT 194.355 49.600 194.525 50.400 ;
        RECT 194.810 50.355 195.475 50.525 ;
        RECT 194.810 50.100 194.980 50.355 ;
        RECT 195.735 50.325 196.945 51.075 ;
        RECT 197.115 50.350 197.405 51.075 ;
        RECT 197.665 50.525 197.835 50.815 ;
        RECT 198.005 50.695 198.335 51.075 ;
        RECT 197.665 50.355 198.330 50.525 ;
        RECT 194.695 49.770 194.980 50.100 ;
        RECT 195.215 49.805 195.545 50.175 ;
        RECT 195.735 49.785 196.255 50.325 ;
        RECT 194.810 49.625 194.980 49.770 ;
        RECT 194.355 48.695 194.625 49.600 ;
        RECT 194.810 49.455 195.475 49.625 ;
        RECT 196.425 49.615 196.945 50.155 ;
        RECT 194.795 48.525 195.125 49.285 ;
        RECT 195.305 48.695 195.475 49.455 ;
        RECT 195.735 48.525 196.945 49.615 ;
        RECT 197.115 48.525 197.405 49.690 ;
        RECT 197.580 49.535 197.930 50.185 ;
        RECT 198.100 49.365 198.330 50.355 ;
        RECT 197.665 49.195 198.330 49.365 ;
        RECT 197.665 48.695 197.835 49.195 ;
        RECT 198.005 48.525 198.335 49.025 ;
        RECT 198.505 48.695 198.730 50.815 ;
        RECT 198.945 50.615 199.195 51.075 ;
        RECT 199.380 50.625 199.710 50.795 ;
        RECT 199.890 50.625 200.640 50.795 ;
        RECT 198.930 49.495 199.210 50.095 ;
        RECT 199.380 49.095 199.550 50.625 ;
        RECT 199.720 50.125 200.300 50.455 ;
        RECT 199.720 49.255 199.960 50.125 ;
        RECT 200.470 49.845 200.640 50.625 ;
        RECT 200.890 50.575 201.260 51.075 ;
        RECT 201.440 50.625 201.900 50.795 ;
        RECT 202.130 50.625 202.800 50.795 ;
        RECT 201.440 50.395 201.610 50.625 ;
        RECT 200.810 50.095 201.610 50.395 ;
        RECT 201.780 50.125 202.330 50.455 ;
        RECT 200.810 50.065 200.980 50.095 ;
        RECT 201.100 49.845 201.270 49.915 ;
        RECT 200.470 49.675 201.270 49.845 ;
        RECT 200.760 49.585 201.270 49.675 ;
        RECT 200.150 49.150 200.590 49.505 ;
        RECT 198.930 48.525 199.195 48.985 ;
        RECT 199.380 48.720 199.615 49.095 ;
        RECT 200.760 48.970 200.930 49.585 ;
        RECT 199.860 48.800 200.930 48.970 ;
        RECT 201.100 48.525 201.270 49.325 ;
        RECT 201.440 49.025 201.610 50.095 ;
        RECT 201.780 49.195 201.970 49.915 ;
        RECT 202.140 49.585 202.330 50.125 ;
        RECT 202.630 50.085 202.800 50.625 ;
        RECT 203.115 50.545 203.285 51.075 ;
        RECT 203.580 50.425 203.940 50.865 ;
        RECT 204.115 50.595 204.285 51.075 ;
        RECT 204.475 50.430 204.810 50.855 ;
        RECT 204.985 50.600 205.155 51.075 ;
        RECT 205.330 50.430 205.665 50.855 ;
        RECT 205.835 50.600 206.005 51.075 ;
        RECT 203.580 50.255 204.080 50.425 ;
        RECT 204.475 50.260 206.145 50.430 ;
        RECT 203.910 50.085 204.080 50.255 ;
        RECT 202.630 49.915 203.720 50.085 ;
        RECT 203.910 49.915 205.730 50.085 ;
        RECT 202.140 49.255 202.460 49.585 ;
        RECT 201.440 48.695 201.690 49.025 ;
        RECT 202.630 48.995 202.800 49.915 ;
        RECT 203.910 49.660 204.080 49.915 ;
        RECT 205.900 49.695 206.145 50.260 ;
        RECT 206.315 50.305 209.825 51.075 ;
        RECT 206.315 49.785 207.965 50.305 ;
        RECT 210.085 50.265 210.255 51.075 ;
        RECT 210.425 50.685 211.595 50.905 ;
        RECT 210.425 50.255 210.675 50.685 ;
        RECT 211.765 50.605 211.935 51.075 ;
        RECT 210.845 50.425 211.180 50.515 ;
        RECT 212.105 50.425 212.435 50.905 ;
        RECT 212.605 50.605 213.295 51.075 ;
        RECT 213.465 50.435 213.795 50.905 ;
        RECT 213.965 50.605 214.135 51.075 ;
        RECT 214.305 50.435 214.635 50.905 ;
        RECT 210.845 50.255 212.435 50.425 ;
        RECT 212.865 50.255 214.635 50.435 ;
        RECT 214.805 50.265 214.975 51.075 ;
        RECT 215.145 50.435 215.475 50.885 ;
        RECT 215.645 50.605 215.815 51.075 ;
        RECT 215.985 50.435 216.315 50.885 ;
        RECT 216.485 50.605 216.655 51.075 ;
        RECT 215.145 50.255 216.830 50.435 ;
        RECT 202.970 49.490 204.080 49.660 ;
        RECT 204.475 49.525 206.145 49.695 ;
        RECT 208.135 49.615 209.825 50.135 ;
        RECT 202.970 49.330 203.830 49.490 ;
        RECT 201.915 48.825 202.800 48.995 ;
        RECT 202.980 48.525 203.195 49.025 ;
        RECT 203.660 48.705 203.830 49.330 ;
        RECT 204.115 48.525 204.295 49.305 ;
        RECT 204.475 48.765 204.810 49.525 ;
        RECT 204.990 48.525 205.160 49.355 ;
        RECT 205.330 48.765 205.660 49.525 ;
        RECT 205.830 48.525 206.000 49.355 ;
        RECT 206.315 48.525 209.825 49.615 ;
        RECT 209.995 49.715 210.485 50.085 ;
        RECT 210.715 49.885 211.255 50.085 ;
        RECT 211.425 49.915 211.805 50.085 ;
        RECT 211.425 49.715 211.595 49.915 ;
        RECT 209.995 49.545 211.595 49.715 ;
        RECT 212.145 49.745 212.355 50.255 ;
        RECT 212.865 50.085 213.055 50.255 ;
        RECT 212.525 49.915 213.055 50.085 ;
        RECT 211.765 49.375 211.975 49.705 ;
        RECT 210.045 49.205 211.975 49.375 ;
        RECT 210.045 48.695 210.295 49.205 ;
        RECT 210.465 48.525 210.715 49.035 ;
        RECT 210.885 48.695 211.135 49.205 ;
        RECT 211.305 48.525 211.555 49.035 ;
        RECT 211.725 48.865 211.975 49.205 ;
        RECT 212.145 49.195 212.530 49.745 ;
        RECT 212.865 49.665 213.055 49.915 ;
        RECT 213.225 49.835 213.555 50.085 ;
        RECT 213.725 49.885 214.345 50.085 ;
        RECT 213.385 49.715 213.555 49.835 ;
        RECT 214.515 49.715 214.875 50.085 ;
        RECT 212.865 49.495 213.215 49.665 ;
        RECT 213.385 49.545 214.875 49.715 ;
        RECT 215.045 49.915 216.350 50.085 ;
        RECT 215.045 49.545 215.370 49.915 ;
        RECT 216.520 49.745 216.830 50.255 ;
        RECT 217.355 50.305 222.700 51.075 ;
        RECT 222.875 50.305 224.545 51.075 ;
        RECT 225.175 50.350 225.465 51.075 ;
        RECT 225.635 50.305 229.145 51.075 ;
        RECT 230.155 50.785 230.490 50.905 ;
        RECT 230.155 50.595 231.415 50.785 ;
        RECT 231.595 50.715 231.925 51.075 ;
        RECT 232.500 50.715 232.830 51.075 ;
        RECT 230.155 50.355 230.490 50.595 ;
        RECT 231.225 50.545 231.415 50.595 ;
        RECT 232.140 50.545 232.330 50.645 ;
        RECT 233.000 50.545 233.190 50.905 ;
        RECT 233.360 50.715 233.690 51.075 ;
        RECT 217.355 49.785 219.935 50.305 ;
        RECT 213.045 49.375 213.215 49.495 ;
        RECT 216.025 49.505 216.830 49.745 ;
        RECT 220.105 49.615 222.700 50.135 ;
        RECT 222.875 49.785 223.625 50.305 ;
        RECT 223.795 49.615 224.545 50.135 ;
        RECT 225.635 49.785 227.285 50.305 ;
        RECT 216.025 49.375 216.275 49.505 ;
        RECT 213.045 49.195 214.175 49.375 ;
        RECT 212.145 49.035 212.395 49.195 ;
        RECT 213.925 49.035 214.175 49.195 ;
        RECT 212.565 48.865 212.815 49.025 ;
        RECT 211.725 48.695 212.815 48.865 ;
        RECT 213.085 48.525 213.335 49.025 ;
        RECT 213.505 48.865 213.755 49.025 ;
        RECT 214.345 48.865 214.595 49.375 ;
        RECT 213.505 48.695 214.595 48.865 ;
        RECT 214.765 48.525 215.015 49.365 ;
        RECT 215.185 49.205 216.275 49.375 ;
        RECT 215.185 48.695 215.435 49.205 ;
        RECT 215.605 48.525 215.855 48.995 ;
        RECT 216.025 48.695 216.275 49.205 ;
        RECT 216.445 48.525 216.695 49.335 ;
        RECT 217.355 48.525 222.700 49.615 ;
        RECT 222.875 48.525 224.545 49.615 ;
        RECT 225.175 48.525 225.465 49.690 ;
        RECT 227.455 49.615 229.145 50.135 ;
        RECT 225.635 48.525 229.145 49.615 ;
        RECT 229.805 49.820 230.565 50.165 ;
        RECT 230.755 49.820 231.045 50.415 ;
        RECT 231.225 50.355 231.970 50.545 ;
        RECT 231.215 49.835 231.590 50.165 ;
        RECT 231.760 50.140 231.970 50.355 ;
        RECT 232.140 50.315 233.745 50.545 ;
        RECT 229.805 48.825 230.055 49.820 ;
        RECT 231.760 49.805 233.295 50.140 ;
        RECT 231.760 49.580 231.970 49.805 ;
        RECT 233.465 49.625 233.745 50.315 ;
        RECT 233.915 50.305 237.425 51.075 ;
        RECT 233.915 49.785 235.565 50.305 ;
        RECT 237.685 50.265 237.855 51.075 ;
        RECT 238.025 50.685 239.195 50.905 ;
        RECT 238.025 50.255 238.275 50.685 ;
        RECT 239.365 50.605 239.535 51.075 ;
        RECT 238.445 50.425 238.780 50.515 ;
        RECT 239.705 50.425 240.035 50.905 ;
        RECT 240.205 50.605 240.895 51.075 ;
        RECT 241.065 50.435 241.395 50.905 ;
        RECT 241.565 50.605 241.735 51.075 ;
        RECT 241.905 50.435 242.235 50.905 ;
        RECT 238.445 50.255 240.035 50.425 ;
        RECT 240.465 50.255 242.235 50.435 ;
        RECT 242.405 50.265 242.575 51.075 ;
        RECT 242.745 50.435 243.075 50.885 ;
        RECT 243.245 50.605 243.415 51.075 ;
        RECT 243.585 50.435 243.915 50.885 ;
        RECT 244.085 50.605 244.255 51.075 ;
        RECT 242.745 50.255 244.430 50.435 ;
        RECT 230.235 49.410 231.970 49.580 ;
        RECT 230.235 48.695 230.415 49.410 ;
        RECT 230.585 48.525 231.035 49.225 ;
        RECT 231.210 48.695 231.390 49.410 ;
        RECT 232.140 49.400 233.745 49.625 ;
        RECT 235.735 49.615 237.425 50.135 ;
        RECT 231.600 48.525 231.930 49.225 ;
        RECT 232.140 49.035 232.330 49.400 ;
        RECT 233.000 49.395 233.745 49.400 ;
        RECT 232.135 48.865 232.330 49.035 ;
        RECT 232.140 48.695 232.330 48.865 ;
        RECT 232.500 48.525 232.830 49.225 ;
        RECT 233.000 48.695 233.190 49.395 ;
        RECT 233.360 48.525 233.690 49.225 ;
        RECT 233.915 48.525 237.425 49.615 ;
        RECT 237.595 49.715 238.085 50.085 ;
        RECT 238.315 49.885 238.855 50.085 ;
        RECT 239.025 49.915 239.405 50.085 ;
        RECT 239.025 49.715 239.195 49.915 ;
        RECT 237.595 49.545 239.195 49.715 ;
        RECT 239.745 49.745 239.955 50.255 ;
        RECT 240.465 50.085 240.655 50.255 ;
        RECT 240.125 49.915 240.655 50.085 ;
        RECT 239.365 49.375 239.575 49.705 ;
        RECT 237.645 49.205 239.575 49.375 ;
        RECT 237.645 48.695 237.895 49.205 ;
        RECT 238.065 48.525 238.315 49.035 ;
        RECT 238.485 48.695 238.735 49.205 ;
        RECT 238.905 48.525 239.155 49.035 ;
        RECT 239.325 48.865 239.575 49.205 ;
        RECT 239.745 49.195 240.130 49.745 ;
        RECT 240.465 49.665 240.655 49.915 ;
        RECT 240.825 49.835 241.155 50.085 ;
        RECT 241.325 49.885 241.945 50.085 ;
        RECT 240.985 49.715 241.155 49.835 ;
        RECT 242.115 49.715 242.475 50.085 ;
        RECT 240.465 49.495 240.815 49.665 ;
        RECT 240.985 49.545 242.475 49.715 ;
        RECT 242.645 49.915 243.950 50.085 ;
        RECT 242.645 49.545 242.970 49.915 ;
        RECT 244.120 49.745 244.430 50.255 ;
        RECT 244.955 50.305 250.300 51.075 ;
        RECT 250.475 50.305 253.065 51.075 ;
        RECT 253.235 50.350 253.525 51.075 ;
        RECT 244.955 49.785 247.535 50.305 ;
        RECT 240.645 49.375 240.815 49.495 ;
        RECT 243.625 49.505 244.430 49.745 ;
        RECT 247.705 49.615 250.300 50.135 ;
        RECT 250.475 49.785 251.685 50.305 ;
        RECT 253.785 50.265 253.955 51.075 ;
        RECT 254.125 50.685 255.295 50.905 ;
        RECT 254.125 50.255 254.375 50.685 ;
        RECT 255.465 50.605 255.635 51.075 ;
        RECT 254.545 50.425 254.880 50.515 ;
        RECT 255.805 50.425 256.135 50.905 ;
        RECT 256.305 50.605 256.995 51.075 ;
        RECT 257.165 50.435 257.495 50.905 ;
        RECT 257.665 50.605 257.835 51.075 ;
        RECT 258.005 50.435 258.335 50.905 ;
        RECT 254.545 50.255 256.135 50.425 ;
        RECT 256.565 50.255 258.335 50.435 ;
        RECT 258.505 50.265 258.675 51.075 ;
        RECT 258.845 50.435 259.175 50.885 ;
        RECT 259.345 50.605 259.515 51.075 ;
        RECT 259.685 50.435 260.015 50.885 ;
        RECT 260.185 50.605 260.355 51.075 ;
        RECT 258.845 50.255 260.530 50.435 ;
        RECT 251.855 49.615 253.065 50.135 ;
        RECT 253.695 49.715 254.185 50.085 ;
        RECT 254.415 49.885 254.955 50.085 ;
        RECT 255.125 49.915 255.505 50.085 ;
        RECT 255.125 49.715 255.295 49.915 ;
        RECT 243.625 49.375 243.875 49.505 ;
        RECT 240.645 49.195 241.775 49.375 ;
        RECT 239.745 49.035 239.995 49.195 ;
        RECT 241.525 49.035 241.775 49.195 ;
        RECT 240.165 48.865 240.415 49.025 ;
        RECT 239.325 48.695 240.415 48.865 ;
        RECT 240.685 48.525 240.935 49.025 ;
        RECT 241.105 48.865 241.355 49.025 ;
        RECT 241.945 48.865 242.195 49.375 ;
        RECT 241.105 48.695 242.195 48.865 ;
        RECT 242.365 48.525 242.615 49.365 ;
        RECT 242.785 49.205 243.875 49.375 ;
        RECT 242.785 48.695 243.035 49.205 ;
        RECT 243.205 48.525 243.455 48.995 ;
        RECT 243.625 48.695 243.875 49.205 ;
        RECT 244.045 48.525 244.295 49.335 ;
        RECT 244.955 48.525 250.300 49.615 ;
        RECT 250.475 48.525 253.065 49.615 ;
        RECT 253.235 48.525 253.525 49.690 ;
        RECT 253.695 49.545 255.295 49.715 ;
        RECT 255.845 49.745 256.055 50.255 ;
        RECT 256.565 50.085 256.755 50.255 ;
        RECT 256.225 49.915 256.755 50.085 ;
        RECT 255.465 49.375 255.675 49.705 ;
        RECT 253.745 49.205 255.675 49.375 ;
        RECT 253.745 48.695 253.995 49.205 ;
        RECT 254.165 48.525 254.415 49.035 ;
        RECT 254.585 48.695 254.835 49.205 ;
        RECT 255.005 48.525 255.255 49.035 ;
        RECT 255.425 48.865 255.675 49.205 ;
        RECT 255.845 49.195 256.230 49.745 ;
        RECT 256.565 49.665 256.755 49.915 ;
        RECT 256.925 49.835 257.255 50.085 ;
        RECT 257.425 49.885 258.045 50.085 ;
        RECT 257.085 49.715 257.255 49.835 ;
        RECT 258.215 49.715 258.575 50.085 ;
        RECT 256.565 49.495 256.915 49.665 ;
        RECT 257.085 49.545 258.575 49.715 ;
        RECT 258.745 49.915 260.050 50.085 ;
        RECT 258.745 49.545 259.070 49.915 ;
        RECT 260.220 49.745 260.530 50.255 ;
        RECT 261.055 50.305 264.565 51.075 ;
        RECT 264.825 50.525 264.995 50.905 ;
        RECT 265.210 50.695 265.540 51.075 ;
        RECT 264.825 50.355 265.540 50.525 ;
        RECT 261.055 49.785 262.705 50.305 ;
        RECT 256.745 49.375 256.915 49.495 ;
        RECT 259.725 49.505 260.530 49.745 ;
        RECT 262.875 49.615 264.565 50.135 ;
        RECT 264.735 49.805 265.090 50.175 ;
        RECT 265.370 50.165 265.540 50.355 ;
        RECT 265.710 50.330 265.965 50.905 ;
        RECT 265.370 49.835 265.625 50.165 ;
        RECT 265.370 49.625 265.540 49.835 ;
        RECT 259.725 49.375 259.975 49.505 ;
        RECT 256.745 49.195 257.875 49.375 ;
        RECT 255.845 49.035 256.095 49.195 ;
        RECT 257.625 49.035 257.875 49.195 ;
        RECT 256.265 48.865 256.515 49.025 ;
        RECT 255.425 48.695 256.515 48.865 ;
        RECT 256.785 48.525 257.035 49.025 ;
        RECT 257.205 48.865 257.455 49.025 ;
        RECT 258.045 48.865 258.295 49.375 ;
        RECT 257.205 48.695 258.295 48.865 ;
        RECT 258.465 48.525 258.715 49.365 ;
        RECT 258.885 49.205 259.975 49.375 ;
        RECT 258.885 48.695 259.135 49.205 ;
        RECT 259.305 48.525 259.555 48.995 ;
        RECT 259.725 48.695 259.975 49.205 ;
        RECT 260.145 48.525 260.395 49.335 ;
        RECT 261.055 48.525 264.565 49.615 ;
        RECT 264.825 49.455 265.540 49.625 ;
        RECT 265.795 49.600 265.965 50.330 ;
        RECT 266.140 50.235 266.400 51.075 ;
        RECT 266.575 50.305 270.085 51.075 ;
        RECT 266.575 49.785 268.225 50.305 ;
        RECT 270.345 50.265 270.515 51.075 ;
        RECT 270.685 50.685 271.855 50.905 ;
        RECT 270.685 50.255 270.935 50.685 ;
        RECT 272.025 50.605 272.195 51.075 ;
        RECT 271.105 50.425 271.440 50.515 ;
        RECT 272.365 50.425 272.695 50.905 ;
        RECT 272.865 50.605 273.555 51.075 ;
        RECT 273.725 50.435 274.055 50.905 ;
        RECT 274.225 50.605 274.395 51.075 ;
        RECT 274.565 50.435 274.895 50.905 ;
        RECT 271.105 50.255 272.695 50.425 ;
        RECT 273.125 50.255 274.895 50.435 ;
        RECT 275.065 50.265 275.235 51.075 ;
        RECT 275.405 50.435 275.735 50.885 ;
        RECT 275.905 50.605 276.075 51.075 ;
        RECT 276.245 50.435 276.575 50.885 ;
        RECT 276.745 50.605 276.915 51.075 ;
        RECT 275.405 50.255 277.090 50.435 ;
        RECT 264.825 48.695 264.995 49.455 ;
        RECT 265.210 48.525 265.540 49.285 ;
        RECT 265.710 48.695 265.965 49.600 ;
        RECT 266.140 48.525 266.400 49.675 ;
        RECT 268.395 49.615 270.085 50.135 ;
        RECT 266.575 48.525 270.085 49.615 ;
        RECT 270.255 49.715 270.745 50.085 ;
        RECT 270.975 49.885 271.515 50.085 ;
        RECT 271.685 49.915 272.065 50.085 ;
        RECT 271.685 49.715 271.855 49.915 ;
        RECT 270.255 49.545 271.855 49.715 ;
        RECT 272.405 49.745 272.615 50.255 ;
        RECT 273.125 50.085 273.315 50.255 ;
        RECT 272.785 49.915 273.315 50.085 ;
        RECT 272.025 49.375 272.235 49.705 ;
        RECT 270.305 49.205 272.235 49.375 ;
        RECT 270.305 48.695 270.555 49.205 ;
        RECT 270.725 48.525 270.975 49.035 ;
        RECT 271.145 48.695 271.395 49.205 ;
        RECT 271.565 48.525 271.815 49.035 ;
        RECT 271.985 48.865 272.235 49.205 ;
        RECT 272.405 49.195 272.790 49.745 ;
        RECT 273.125 49.665 273.315 49.915 ;
        RECT 273.485 49.835 273.815 50.085 ;
        RECT 273.985 49.885 274.605 50.085 ;
        RECT 273.645 49.715 273.815 49.835 ;
        RECT 274.775 49.715 275.135 50.085 ;
        RECT 273.125 49.495 273.475 49.665 ;
        RECT 273.645 49.545 275.135 49.715 ;
        RECT 275.305 49.915 276.610 50.085 ;
        RECT 275.305 49.545 275.630 49.915 ;
        RECT 276.780 49.745 277.090 50.255 ;
        RECT 277.615 50.305 281.125 51.075 ;
        RECT 281.295 50.350 281.585 51.075 ;
        RECT 277.615 49.785 279.265 50.305 ;
        RECT 281.760 50.255 282.035 51.075 ;
        RECT 282.205 50.435 282.535 50.905 ;
        RECT 282.705 50.605 282.875 51.075 ;
        RECT 283.045 50.435 283.375 50.905 ;
        RECT 283.545 50.605 283.715 51.075 ;
        RECT 283.885 50.435 284.215 50.905 ;
        RECT 284.385 50.605 284.555 51.075 ;
        RECT 284.725 50.435 285.055 50.905 ;
        RECT 285.225 50.605 285.510 51.075 ;
        RECT 282.205 50.255 285.725 50.435 ;
        RECT 273.305 49.375 273.475 49.495 ;
        RECT 276.285 49.505 277.090 49.745 ;
        RECT 279.435 49.615 281.125 50.135 ;
        RECT 281.810 49.885 283.470 50.085 ;
        RECT 283.790 49.885 285.155 50.085 ;
        RECT 285.325 49.715 285.725 50.255 ;
        RECT 285.895 50.305 289.405 51.075 ;
        RECT 285.895 49.785 287.545 50.305 ;
        RECT 289.665 50.265 289.835 51.075 ;
        RECT 290.005 50.685 291.175 50.905 ;
        RECT 290.005 50.255 290.255 50.685 ;
        RECT 291.345 50.605 291.515 51.075 ;
        RECT 290.425 50.425 290.760 50.515 ;
        RECT 291.685 50.425 292.015 50.905 ;
        RECT 292.185 50.605 292.875 51.075 ;
        RECT 293.045 50.435 293.375 50.905 ;
        RECT 293.545 50.605 293.715 51.075 ;
        RECT 293.885 50.435 294.215 50.905 ;
        RECT 290.425 50.255 292.015 50.425 ;
        RECT 292.445 50.255 294.215 50.435 ;
        RECT 294.385 50.265 294.555 51.075 ;
        RECT 294.725 50.435 295.055 50.885 ;
        RECT 295.225 50.605 295.395 51.075 ;
        RECT 295.565 50.435 295.895 50.885 ;
        RECT 296.065 50.605 296.235 51.075 ;
        RECT 294.725 50.255 296.410 50.435 ;
        RECT 276.285 49.375 276.535 49.505 ;
        RECT 273.305 49.195 274.435 49.375 ;
        RECT 272.405 49.035 272.655 49.195 ;
        RECT 274.185 49.035 274.435 49.195 ;
        RECT 272.825 48.865 273.075 49.025 ;
        RECT 271.985 48.695 273.075 48.865 ;
        RECT 273.345 48.525 273.595 49.025 ;
        RECT 273.765 48.865 274.015 49.025 ;
        RECT 274.605 48.865 274.855 49.375 ;
        RECT 273.765 48.695 274.855 48.865 ;
        RECT 275.025 48.525 275.275 49.365 ;
        RECT 275.445 49.205 276.535 49.375 ;
        RECT 275.445 48.695 275.695 49.205 ;
        RECT 275.865 48.525 276.115 48.995 ;
        RECT 276.285 48.695 276.535 49.205 ;
        RECT 276.705 48.525 276.955 49.335 ;
        RECT 277.615 48.525 281.125 49.615 ;
        RECT 281.295 48.525 281.585 49.690 ;
        RECT 281.760 49.495 283.795 49.705 ;
        RECT 281.760 48.695 282.035 49.495 ;
        RECT 282.205 48.525 282.535 49.325 ;
        RECT 282.705 48.695 282.875 49.495 ;
        RECT 283.045 48.525 283.295 49.325 ;
        RECT 283.465 48.865 283.795 49.495 ;
        RECT 283.965 49.415 285.725 49.715 ;
        RECT 287.715 49.615 289.405 50.135 ;
        RECT 283.965 49.035 284.135 49.415 ;
        RECT 284.305 48.865 284.635 49.225 ;
        RECT 284.805 49.035 284.975 49.415 ;
        RECT 285.145 48.865 285.560 49.245 ;
        RECT 283.465 48.695 285.560 48.865 ;
        RECT 285.895 48.525 289.405 49.615 ;
        RECT 289.575 49.715 290.065 50.085 ;
        RECT 290.295 49.885 290.835 50.085 ;
        RECT 291.005 49.915 291.385 50.085 ;
        RECT 291.005 49.715 291.175 49.915 ;
        RECT 289.575 49.545 291.175 49.715 ;
        RECT 291.725 49.745 291.935 50.255 ;
        RECT 292.445 50.085 292.635 50.255 ;
        RECT 296.075 50.225 296.410 50.255 ;
        RECT 292.105 49.915 292.635 50.085 ;
        RECT 291.345 49.375 291.555 49.705 ;
        RECT 289.625 49.205 291.555 49.375 ;
        RECT 289.625 48.695 289.875 49.205 ;
        RECT 290.045 48.525 290.295 49.035 ;
        RECT 290.465 48.695 290.715 49.205 ;
        RECT 290.885 48.525 291.135 49.035 ;
        RECT 291.305 48.865 291.555 49.205 ;
        RECT 291.725 49.195 292.110 49.745 ;
        RECT 292.445 49.665 292.635 49.915 ;
        RECT 292.805 49.835 293.135 50.085 ;
        RECT 293.305 49.885 293.925 50.085 ;
        RECT 292.965 49.715 293.135 49.835 ;
        RECT 294.095 49.715 294.455 50.085 ;
        RECT 292.445 49.495 292.795 49.665 ;
        RECT 292.965 49.545 294.455 49.715 ;
        RECT 294.625 49.915 295.930 50.085 ;
        RECT 294.625 49.545 294.950 49.915 ;
        RECT 296.100 49.745 296.410 50.225 ;
        RECT 296.935 50.305 300.445 51.075 ;
        RECT 296.935 49.785 298.585 50.305 ;
        RECT 300.620 50.255 300.895 51.075 ;
        RECT 301.065 50.435 301.395 50.905 ;
        RECT 301.565 50.605 301.735 51.075 ;
        RECT 301.905 50.435 302.235 50.905 ;
        RECT 302.405 50.605 302.575 51.075 ;
        RECT 302.745 50.435 303.075 50.905 ;
        RECT 303.245 50.605 303.415 51.075 ;
        RECT 303.585 50.435 303.915 50.905 ;
        RECT 304.085 50.605 304.370 51.075 ;
        RECT 301.065 50.255 304.585 50.435 ;
        RECT 292.625 49.375 292.795 49.495 ;
        RECT 295.605 49.505 296.410 49.745 ;
        RECT 298.755 49.615 300.445 50.135 ;
        RECT 300.670 49.885 302.330 50.085 ;
        RECT 302.650 49.885 304.015 50.085 ;
        RECT 304.185 49.715 304.585 50.255 ;
        RECT 304.755 50.305 308.265 51.075 ;
        RECT 309.355 50.350 309.645 51.075 ;
        RECT 309.815 50.305 313.325 51.075 ;
        RECT 304.755 49.785 306.405 50.305 ;
        RECT 295.605 49.375 295.855 49.505 ;
        RECT 292.625 49.195 293.755 49.375 ;
        RECT 291.725 49.035 291.975 49.195 ;
        RECT 293.505 49.035 293.755 49.195 ;
        RECT 292.145 48.865 292.395 49.025 ;
        RECT 291.305 48.695 292.395 48.865 ;
        RECT 292.665 48.525 292.915 49.025 ;
        RECT 293.085 48.865 293.335 49.025 ;
        RECT 293.925 48.865 294.175 49.375 ;
        RECT 293.085 48.695 294.175 48.865 ;
        RECT 294.345 48.525 294.595 49.365 ;
        RECT 294.765 49.205 295.855 49.375 ;
        RECT 294.765 48.695 295.015 49.205 ;
        RECT 295.185 48.525 295.435 48.995 ;
        RECT 295.605 48.695 295.855 49.205 ;
        RECT 296.025 48.525 296.275 49.335 ;
        RECT 296.935 48.525 300.445 49.615 ;
        RECT 300.620 49.495 302.655 49.705 ;
        RECT 300.620 48.695 300.895 49.495 ;
        RECT 301.065 48.525 301.395 49.325 ;
        RECT 301.565 48.695 301.735 49.495 ;
        RECT 301.905 48.525 302.155 49.325 ;
        RECT 302.325 48.865 302.655 49.495 ;
        RECT 302.825 49.415 304.585 49.715 ;
        RECT 306.575 49.615 308.265 50.135 ;
        RECT 309.815 49.785 311.465 50.305 ;
        RECT 314.420 50.255 314.695 51.075 ;
        RECT 314.865 50.435 315.195 50.905 ;
        RECT 315.365 50.605 315.535 51.075 ;
        RECT 315.705 50.435 316.035 50.905 ;
        RECT 316.205 50.605 316.375 51.075 ;
        RECT 316.545 50.435 316.875 50.905 ;
        RECT 317.045 50.605 317.215 51.075 ;
        RECT 317.385 50.435 317.715 50.905 ;
        RECT 317.885 50.605 318.170 51.075 ;
        RECT 314.865 50.255 318.385 50.435 ;
        RECT 302.825 49.035 302.995 49.415 ;
        RECT 303.165 48.865 303.495 49.225 ;
        RECT 303.665 49.035 303.835 49.415 ;
        RECT 304.005 48.865 304.420 49.245 ;
        RECT 302.325 48.695 304.420 48.865 ;
        RECT 304.755 48.525 308.265 49.615 ;
        RECT 309.355 48.525 309.645 49.690 ;
        RECT 311.635 49.615 313.325 50.135 ;
        RECT 314.470 49.885 316.130 50.085 ;
        RECT 316.450 49.885 317.815 50.085 ;
        RECT 317.985 49.715 318.385 50.255 ;
        RECT 318.555 50.305 322.065 51.075 ;
        RECT 318.555 49.785 320.205 50.305 ;
        RECT 323.245 50.265 323.415 51.075 ;
        RECT 323.585 50.685 324.755 50.905 ;
        RECT 323.585 50.255 323.835 50.685 ;
        RECT 324.925 50.605 325.095 51.075 ;
        RECT 324.005 50.425 324.340 50.515 ;
        RECT 325.265 50.425 325.595 50.905 ;
        RECT 325.765 50.605 326.455 51.075 ;
        RECT 326.625 50.435 326.955 50.905 ;
        RECT 327.125 50.605 327.295 51.075 ;
        RECT 327.465 50.435 327.795 50.905 ;
        RECT 324.005 50.255 325.595 50.425 ;
        RECT 326.025 50.255 327.795 50.435 ;
        RECT 327.965 50.265 328.135 51.075 ;
        RECT 328.305 50.435 328.635 50.885 ;
        RECT 328.805 50.605 328.975 51.075 ;
        RECT 329.145 50.435 329.475 50.885 ;
        RECT 329.645 50.605 329.815 51.075 ;
        RECT 328.305 50.255 329.990 50.435 ;
        RECT 309.815 48.525 313.325 49.615 ;
        RECT 314.420 49.495 316.455 49.705 ;
        RECT 314.420 48.695 314.695 49.495 ;
        RECT 314.865 48.525 315.195 49.325 ;
        RECT 315.365 48.695 315.535 49.495 ;
        RECT 315.705 48.525 315.955 49.325 ;
        RECT 316.125 48.865 316.455 49.495 ;
        RECT 316.625 49.415 318.385 49.715 ;
        RECT 320.375 49.615 322.065 50.135 ;
        RECT 316.625 49.035 316.795 49.415 ;
        RECT 316.965 48.865 317.295 49.225 ;
        RECT 317.465 49.035 317.635 49.415 ;
        RECT 317.805 48.865 318.220 49.245 ;
        RECT 316.125 48.695 318.220 48.865 ;
        RECT 318.555 48.525 322.065 49.615 ;
        RECT 323.155 49.715 323.645 50.085 ;
        RECT 323.875 49.885 324.415 50.085 ;
        RECT 324.585 49.915 324.965 50.085 ;
        RECT 324.585 49.715 324.755 49.915 ;
        RECT 323.155 49.545 324.755 49.715 ;
        RECT 325.305 49.745 325.515 50.255 ;
        RECT 326.025 50.085 326.215 50.255 ;
        RECT 329.655 50.225 329.990 50.255 ;
        RECT 325.685 49.915 326.215 50.085 ;
        RECT 324.925 49.375 325.135 49.705 ;
        RECT 323.205 49.205 325.135 49.375 ;
        RECT 323.205 48.695 323.455 49.205 ;
        RECT 323.625 48.525 323.875 49.035 ;
        RECT 324.045 48.695 324.295 49.205 ;
        RECT 324.465 48.525 324.715 49.035 ;
        RECT 324.885 48.865 325.135 49.205 ;
        RECT 325.305 49.195 325.690 49.745 ;
        RECT 326.025 49.665 326.215 49.915 ;
        RECT 326.385 49.835 326.715 50.085 ;
        RECT 326.885 49.885 327.505 50.085 ;
        RECT 326.545 49.715 326.715 49.835 ;
        RECT 327.675 49.715 328.035 50.085 ;
        RECT 326.025 49.495 326.375 49.665 ;
        RECT 326.545 49.545 328.035 49.715 ;
        RECT 328.205 49.915 329.510 50.085 ;
        RECT 328.205 49.545 328.530 49.915 ;
        RECT 329.680 49.745 329.990 50.225 ;
        RECT 330.515 50.305 335.860 51.075 ;
        RECT 336.035 50.325 337.245 51.075 ;
        RECT 337.415 50.350 337.705 51.075 ;
        RECT 337.965 50.525 338.135 50.905 ;
        RECT 338.350 50.695 338.680 51.075 ;
        RECT 337.965 50.355 338.680 50.525 ;
        RECT 330.515 49.785 333.095 50.305 ;
        RECT 326.205 49.375 326.375 49.495 ;
        RECT 329.185 49.505 329.990 49.745 ;
        RECT 333.265 49.615 335.860 50.135 ;
        RECT 336.035 49.785 336.555 50.325 ;
        RECT 336.725 49.615 337.245 50.155 ;
        RECT 337.875 49.805 338.230 50.175 ;
        RECT 338.510 50.165 338.680 50.355 ;
        RECT 339.280 50.235 339.540 51.075 ;
        RECT 339.715 50.305 343.225 51.075 ;
        RECT 338.510 49.835 338.765 50.165 ;
        RECT 329.185 49.375 329.435 49.505 ;
        RECT 326.205 49.195 327.335 49.375 ;
        RECT 325.305 49.035 325.555 49.195 ;
        RECT 327.085 49.035 327.335 49.195 ;
        RECT 325.725 48.865 325.975 49.025 ;
        RECT 324.885 48.695 325.975 48.865 ;
        RECT 326.245 48.525 326.495 49.025 ;
        RECT 326.665 48.865 326.915 49.025 ;
        RECT 327.505 48.865 327.755 49.375 ;
        RECT 326.665 48.695 327.755 48.865 ;
        RECT 327.925 48.525 328.175 49.365 ;
        RECT 328.345 49.205 329.435 49.375 ;
        RECT 328.345 48.695 328.595 49.205 ;
        RECT 328.765 48.525 329.015 48.995 ;
        RECT 329.185 48.695 329.435 49.205 ;
        RECT 329.605 48.525 329.855 49.335 ;
        RECT 330.515 48.525 335.860 49.615 ;
        RECT 336.035 48.525 337.245 49.615 ;
        RECT 337.415 48.525 337.705 49.690 ;
        RECT 338.510 49.625 338.680 49.835 ;
        RECT 339.715 49.785 341.365 50.305 ;
        RECT 343.485 50.265 343.655 51.075 ;
        RECT 343.825 50.685 344.995 50.905 ;
        RECT 343.825 50.255 344.075 50.685 ;
        RECT 345.165 50.605 345.335 51.075 ;
        RECT 344.245 50.425 344.580 50.515 ;
        RECT 345.505 50.425 345.835 50.905 ;
        RECT 346.005 50.605 346.695 51.075 ;
        RECT 346.865 50.435 347.195 50.905 ;
        RECT 347.365 50.605 347.535 51.075 ;
        RECT 347.705 50.435 348.035 50.905 ;
        RECT 344.245 50.255 345.835 50.425 ;
        RECT 346.265 50.255 348.035 50.435 ;
        RECT 348.205 50.265 348.375 51.075 ;
        RECT 348.545 50.435 348.875 50.885 ;
        RECT 349.045 50.605 349.215 51.075 ;
        RECT 349.385 50.435 349.715 50.885 ;
        RECT 349.885 50.605 350.055 51.075 ;
        RECT 348.545 50.255 350.230 50.435 ;
        RECT 337.965 49.455 338.680 49.625 ;
        RECT 337.965 48.695 338.135 49.455 ;
        RECT 338.350 48.525 338.680 49.285 ;
        RECT 339.280 48.525 339.540 49.675 ;
        RECT 341.535 49.615 343.225 50.135 ;
        RECT 339.715 48.525 343.225 49.615 ;
        RECT 343.395 49.715 343.885 50.085 ;
        RECT 344.115 49.885 344.655 50.085 ;
        RECT 344.825 49.915 345.205 50.085 ;
        RECT 344.825 49.715 344.995 49.915 ;
        RECT 343.395 49.545 344.995 49.715 ;
        RECT 345.545 49.745 345.755 50.255 ;
        RECT 346.265 50.085 346.455 50.255 ;
        RECT 345.925 49.915 346.455 50.085 ;
        RECT 345.165 49.375 345.375 49.705 ;
        RECT 343.445 49.205 345.375 49.375 ;
        RECT 343.445 48.695 343.695 49.205 ;
        RECT 343.865 48.525 344.115 49.035 ;
        RECT 344.285 48.695 344.535 49.205 ;
        RECT 344.705 48.525 344.955 49.035 ;
        RECT 345.125 48.865 345.375 49.205 ;
        RECT 345.545 49.195 345.930 49.745 ;
        RECT 346.265 49.665 346.455 49.915 ;
        RECT 346.625 49.835 346.955 50.085 ;
        RECT 347.125 49.885 347.745 50.085 ;
        RECT 346.785 49.715 346.955 49.835 ;
        RECT 347.915 49.715 348.275 50.085 ;
        RECT 346.265 49.495 346.615 49.665 ;
        RECT 346.785 49.545 348.275 49.715 ;
        RECT 348.445 49.915 349.750 50.085 ;
        RECT 348.445 49.545 348.770 49.915 ;
        RECT 349.920 49.745 350.230 50.255 ;
        RECT 350.755 50.305 354.265 51.075 ;
        RECT 350.755 49.785 352.405 50.305 ;
        RECT 354.440 50.255 354.715 51.075 ;
        RECT 354.885 50.435 355.215 50.905 ;
        RECT 355.385 50.605 355.555 51.075 ;
        RECT 355.725 50.435 356.055 50.905 ;
        RECT 356.225 50.605 356.395 51.075 ;
        RECT 356.565 50.435 356.895 50.905 ;
        RECT 357.065 50.605 357.235 51.075 ;
        RECT 357.405 50.435 357.735 50.905 ;
        RECT 357.905 50.605 358.190 51.075 ;
        RECT 354.885 50.255 358.405 50.435 ;
        RECT 346.445 49.375 346.615 49.495 ;
        RECT 349.425 49.505 350.230 49.745 ;
        RECT 352.575 49.615 354.265 50.135 ;
        RECT 354.490 49.885 356.150 50.085 ;
        RECT 356.470 49.885 357.835 50.085 ;
        RECT 358.005 49.715 358.405 50.255 ;
        RECT 358.575 50.305 363.920 51.075 ;
        RECT 364.095 50.325 365.305 51.075 ;
        RECT 365.475 50.350 365.765 51.075 ;
        RECT 358.575 49.785 361.155 50.305 ;
        RECT 349.425 49.375 349.675 49.505 ;
        RECT 346.445 49.195 347.575 49.375 ;
        RECT 345.545 49.035 345.795 49.195 ;
        RECT 347.325 49.035 347.575 49.195 ;
        RECT 345.965 48.865 346.215 49.025 ;
        RECT 345.125 48.695 346.215 48.865 ;
        RECT 346.485 48.525 346.735 49.025 ;
        RECT 346.905 48.865 347.155 49.025 ;
        RECT 347.745 48.865 347.995 49.375 ;
        RECT 346.905 48.695 347.995 48.865 ;
        RECT 348.165 48.525 348.415 49.365 ;
        RECT 348.585 49.205 349.675 49.375 ;
        RECT 348.585 48.695 348.835 49.205 ;
        RECT 349.005 48.525 349.255 48.995 ;
        RECT 349.425 48.695 349.675 49.205 ;
        RECT 349.845 48.525 350.095 49.335 ;
        RECT 350.755 48.525 354.265 49.615 ;
        RECT 354.440 49.495 356.475 49.705 ;
        RECT 354.440 48.695 354.715 49.495 ;
        RECT 354.885 48.525 355.215 49.325 ;
        RECT 355.385 48.695 355.555 49.495 ;
        RECT 355.725 48.525 355.975 49.325 ;
        RECT 356.145 48.865 356.475 49.495 ;
        RECT 356.645 49.415 358.405 49.715 ;
        RECT 361.325 49.615 363.920 50.135 ;
        RECT 364.095 49.785 364.615 50.325 ;
        RECT 365.940 50.255 366.215 51.075 ;
        RECT 366.385 50.435 366.715 50.905 ;
        RECT 366.885 50.605 367.055 51.075 ;
        RECT 367.225 50.435 367.555 50.905 ;
        RECT 367.725 50.605 367.895 51.075 ;
        RECT 368.065 50.435 368.395 50.905 ;
        RECT 368.565 50.605 368.735 51.075 ;
        RECT 368.905 50.435 369.235 50.905 ;
        RECT 369.405 50.605 369.690 51.075 ;
        RECT 366.385 50.255 369.905 50.435 ;
        RECT 364.785 49.615 365.305 50.155 ;
        RECT 365.990 49.885 367.650 50.085 ;
        RECT 367.970 49.885 369.335 50.085 ;
        RECT 369.505 49.715 369.905 50.255 ;
        RECT 370.075 50.305 373.585 51.075 ;
        RECT 370.075 49.785 371.725 50.305 ;
        RECT 373.760 50.255 374.035 51.075 ;
        RECT 374.205 50.435 374.535 50.905 ;
        RECT 374.705 50.605 374.875 51.075 ;
        RECT 375.045 50.435 375.375 50.905 ;
        RECT 375.545 50.605 375.715 51.075 ;
        RECT 375.885 50.435 376.215 50.905 ;
        RECT 376.385 50.605 376.555 51.075 ;
        RECT 376.725 50.435 377.055 50.905 ;
        RECT 377.225 50.605 377.510 51.075 ;
        RECT 374.205 50.255 377.725 50.435 ;
        RECT 356.645 49.035 356.815 49.415 ;
        RECT 356.985 48.865 357.315 49.225 ;
        RECT 357.485 49.035 357.655 49.415 ;
        RECT 357.825 48.865 358.240 49.245 ;
        RECT 356.145 48.695 358.240 48.865 ;
        RECT 358.575 48.525 363.920 49.615 ;
        RECT 364.095 48.525 365.305 49.615 ;
        RECT 365.475 48.525 365.765 49.690 ;
        RECT 365.940 49.495 367.975 49.705 ;
        RECT 365.940 48.695 366.215 49.495 ;
        RECT 366.385 48.525 366.715 49.325 ;
        RECT 366.885 48.695 367.055 49.495 ;
        RECT 367.225 48.525 367.475 49.325 ;
        RECT 367.645 48.865 367.975 49.495 ;
        RECT 368.145 49.415 369.905 49.715 ;
        RECT 371.895 49.615 373.585 50.135 ;
        RECT 373.810 49.885 375.470 50.085 ;
        RECT 375.790 49.885 377.155 50.085 ;
        RECT 377.325 49.715 377.725 50.255 ;
        RECT 377.895 50.305 381.405 51.075 ;
        RECT 377.895 49.785 379.545 50.305 ;
        RECT 368.145 49.035 368.315 49.415 ;
        RECT 368.485 48.865 368.815 49.225 ;
        RECT 368.985 49.035 369.155 49.415 ;
        RECT 369.325 48.865 369.740 49.245 ;
        RECT 367.645 48.695 369.740 48.865 ;
        RECT 370.075 48.525 373.585 49.615 ;
        RECT 373.760 49.495 375.795 49.705 ;
        RECT 373.760 48.695 374.035 49.495 ;
        RECT 374.205 48.525 374.535 49.325 ;
        RECT 374.705 48.695 374.875 49.495 ;
        RECT 375.045 48.525 375.295 49.325 ;
        RECT 375.465 48.865 375.795 49.495 ;
        RECT 375.965 49.415 377.725 49.715 ;
        RECT 379.715 49.615 381.405 50.135 ;
        RECT 375.965 49.035 376.135 49.415 ;
        RECT 376.305 48.865 376.635 49.225 ;
        RECT 376.805 49.035 376.975 49.415 ;
        RECT 377.145 48.865 377.560 49.245 ;
        RECT 375.465 48.695 377.560 48.865 ;
        RECT 377.895 48.525 381.405 49.615 ;
        RECT 381.575 49.420 382.095 50.905 ;
        RECT 382.265 50.415 382.605 51.075 ;
        RECT 382.955 50.305 386.465 51.075 ;
        RECT 381.765 48.525 382.095 49.250 ;
        RECT 382.265 48.695 382.785 50.245 ;
        RECT 382.955 49.785 384.605 50.305 ;
        RECT 384.775 49.615 386.465 50.135 ;
        RECT 382.955 48.525 386.465 49.615 ;
        RECT 386.635 49.420 387.155 50.905 ;
        RECT 387.325 50.415 387.665 51.075 ;
        RECT 388.015 50.305 393.360 51.075 ;
        RECT 393.535 50.350 393.825 51.075 ;
        RECT 386.825 48.525 387.155 49.250 ;
        RECT 387.325 48.695 387.845 50.245 ;
        RECT 388.015 49.785 390.595 50.305 ;
        RECT 390.765 49.615 393.360 50.135 ;
        RECT 388.015 48.525 393.360 49.615 ;
        RECT 393.535 48.525 393.825 49.690 ;
        RECT 393.995 49.420 394.515 50.905 ;
        RECT 394.685 50.415 395.025 51.075 ;
        RECT 395.375 50.305 398.885 51.075 ;
        RECT 394.185 48.525 394.515 49.250 ;
        RECT 394.685 48.695 395.205 50.245 ;
        RECT 395.375 49.785 397.025 50.305 ;
        RECT 397.195 49.615 398.885 50.135 ;
        RECT 395.375 48.525 398.885 49.615 ;
        RECT 399.055 49.420 399.575 50.905 ;
        RECT 399.745 50.415 400.085 51.075 ;
        RECT 400.435 50.305 403.945 51.075 ;
        RECT 399.245 48.525 399.575 49.250 ;
        RECT 399.745 48.695 400.265 50.245 ;
        RECT 400.435 49.785 402.085 50.305 ;
        RECT 402.255 49.615 403.945 50.135 ;
        RECT 400.435 48.525 403.945 49.615 ;
        RECT 404.115 49.420 404.635 50.905 ;
        RECT 404.805 50.415 405.145 51.075 ;
        RECT 405.495 50.305 410.840 51.075 ;
        RECT 411.015 50.305 412.685 51.075 ;
        RECT 404.305 48.525 404.635 49.250 ;
        RECT 404.805 48.695 405.325 50.245 ;
        RECT 405.495 49.785 408.075 50.305 ;
        RECT 408.245 49.615 410.840 50.135 ;
        RECT 411.015 49.785 411.765 50.305 ;
        RECT 411.935 49.615 412.685 50.135 ;
        RECT 405.495 48.525 410.840 49.615 ;
        RECT 411.015 48.525 412.685 49.615 ;
        RECT 413.315 49.420 413.835 50.905 ;
        RECT 414.005 50.415 414.345 51.075 ;
        RECT 414.695 50.305 420.040 51.075 ;
        RECT 420.215 50.325 421.425 51.075 ;
        RECT 421.595 50.350 421.885 51.075 ;
        RECT 413.505 48.525 413.835 49.250 ;
        RECT 414.005 48.695 414.525 50.245 ;
        RECT 414.695 49.785 417.275 50.305 ;
        RECT 417.445 49.615 420.040 50.135 ;
        RECT 420.215 49.785 420.735 50.325 ;
        RECT 422.055 50.305 427.400 51.075 ;
        RECT 420.905 49.615 421.425 50.155 ;
        RECT 422.055 49.785 424.635 50.305 ;
        RECT 414.695 48.525 420.040 49.615 ;
        RECT 420.215 48.525 421.425 49.615 ;
        RECT 421.595 48.525 421.885 49.690 ;
        RECT 424.805 49.615 427.400 50.135 ;
        RECT 422.055 48.525 427.400 49.615 ;
        RECT 428.035 49.420 428.555 50.905 ;
        RECT 428.725 50.415 429.065 51.075 ;
        RECT 429.415 50.305 434.760 51.075 ;
        RECT 428.225 48.525 428.555 49.250 ;
        RECT 428.725 48.695 429.245 50.245 ;
        RECT 429.415 49.785 431.995 50.305 ;
        RECT 432.165 49.615 434.760 50.135 ;
        RECT 429.415 48.525 434.760 49.615 ;
        RECT 435.395 49.420 435.915 50.905 ;
        RECT 436.085 50.415 436.425 51.075 ;
        RECT 436.775 50.305 442.120 51.075 ;
        RECT 442.295 50.305 447.640 51.075 ;
        RECT 447.815 50.305 449.485 51.075 ;
        RECT 449.655 50.350 449.945 51.075 ;
        RECT 435.585 48.525 435.915 49.250 ;
        RECT 436.085 48.695 436.605 50.245 ;
        RECT 436.775 49.785 439.355 50.305 ;
        RECT 439.525 49.615 442.120 50.135 ;
        RECT 442.295 49.785 444.875 50.305 ;
        RECT 445.045 49.615 447.640 50.135 ;
        RECT 447.815 49.785 448.565 50.305 ;
        RECT 448.735 49.615 449.485 50.135 ;
        RECT 436.775 48.525 442.120 49.615 ;
        RECT 442.295 48.525 447.640 49.615 ;
        RECT 447.815 48.525 449.485 49.615 ;
        RECT 449.655 48.525 449.945 49.690 ;
        RECT 450.115 49.420 450.635 50.905 ;
        RECT 450.805 50.415 451.145 51.075 ;
        RECT 451.495 50.305 456.840 51.075 ;
        RECT 450.305 48.525 450.635 49.250 ;
        RECT 450.805 48.695 451.325 50.245 ;
        RECT 451.495 49.785 454.075 50.305 ;
        RECT 454.245 49.615 456.840 50.135 ;
        RECT 451.495 48.525 456.840 49.615 ;
        RECT 457.475 49.420 457.995 50.905 ;
        RECT 458.165 50.415 458.505 51.075 ;
        RECT 458.855 50.305 464.200 51.075 ;
        RECT 464.375 50.305 467.885 51.075 ;
        RECT 457.665 48.525 457.995 49.250 ;
        RECT 458.165 48.695 458.685 50.245 ;
        RECT 458.855 49.785 461.435 50.305 ;
        RECT 461.605 49.615 464.200 50.135 ;
        RECT 464.375 49.785 466.025 50.305 ;
        RECT 466.195 49.615 467.885 50.135 ;
        RECT 458.855 48.525 464.200 49.615 ;
        RECT 464.375 48.525 467.885 49.615 ;
        RECT 468.515 49.420 469.035 50.905 ;
        RECT 469.205 50.415 469.545 51.075 ;
        RECT 469.895 50.305 475.240 51.075 ;
        RECT 475.415 50.305 477.085 51.075 ;
        RECT 477.715 50.350 478.005 51.075 ;
        RECT 478.175 50.325 479.385 51.075 ;
        RECT 468.705 48.525 469.035 49.250 ;
        RECT 469.205 48.695 469.725 50.245 ;
        RECT 469.895 49.785 472.475 50.305 ;
        RECT 472.645 49.615 475.240 50.135 ;
        RECT 475.415 49.785 476.165 50.305 ;
        RECT 476.335 49.615 477.085 50.135 ;
        RECT 478.175 49.785 478.695 50.325 ;
        RECT 469.895 48.525 475.240 49.615 ;
        RECT 475.415 48.525 477.085 49.615 ;
        RECT 477.715 48.525 478.005 49.690 ;
        RECT 478.865 49.615 479.385 50.155 ;
        RECT 478.175 48.525 479.385 49.615 ;
        RECT 479.555 49.420 480.075 50.905 ;
        RECT 480.245 50.415 480.585 51.075 ;
        RECT 480.935 50.305 486.280 51.075 ;
        RECT 479.745 48.525 480.075 49.250 ;
        RECT 480.245 48.695 480.765 50.245 ;
        RECT 480.935 49.785 483.515 50.305 ;
        RECT 483.685 49.615 486.280 50.135 ;
        RECT 480.935 48.525 486.280 49.615 ;
        RECT 486.915 49.420 487.435 50.905 ;
        RECT 487.605 50.415 487.945 51.075 ;
        RECT 488.295 50.305 493.640 51.075 ;
        RECT 493.815 50.305 499.160 51.075 ;
        RECT 499.335 50.305 504.680 51.075 ;
        RECT 505.775 50.350 506.065 51.075 ;
        RECT 506.235 50.305 511.580 51.075 ;
        RECT 487.105 48.525 487.435 49.250 ;
        RECT 487.605 48.695 488.125 50.245 ;
        RECT 488.295 49.785 490.875 50.305 ;
        RECT 491.045 49.615 493.640 50.135 ;
        RECT 493.815 49.785 496.395 50.305 ;
        RECT 496.565 49.615 499.160 50.135 ;
        RECT 499.335 49.785 501.915 50.305 ;
        RECT 502.085 49.615 504.680 50.135 ;
        RECT 506.235 49.785 508.815 50.305 ;
        RECT 488.295 48.525 493.640 49.615 ;
        RECT 493.815 48.525 499.160 49.615 ;
        RECT 499.335 48.525 504.680 49.615 ;
        RECT 505.775 48.525 506.065 49.690 ;
        RECT 508.985 49.615 511.580 50.135 ;
        RECT 506.235 48.525 511.580 49.615 ;
        RECT 512.675 49.420 513.195 50.905 ;
        RECT 513.365 50.415 513.705 51.075 ;
        RECT 514.055 50.305 519.400 51.075 ;
        RECT 512.865 48.525 513.195 49.250 ;
        RECT 513.365 48.695 513.885 50.245 ;
        RECT 514.055 49.785 516.635 50.305 ;
        RECT 516.805 49.615 519.400 50.135 ;
        RECT 514.055 48.525 519.400 49.615 ;
        RECT 520.035 49.420 520.555 50.905 ;
        RECT 520.725 50.415 521.065 51.075 ;
        RECT 521.415 50.305 526.760 51.075 ;
        RECT 526.935 50.305 532.280 51.075 ;
        RECT 532.455 50.325 533.665 51.075 ;
        RECT 533.835 50.350 534.125 51.075 ;
        RECT 520.225 48.525 520.555 49.250 ;
        RECT 520.725 48.695 521.245 50.245 ;
        RECT 521.415 49.785 523.995 50.305 ;
        RECT 524.165 49.615 526.760 50.135 ;
        RECT 526.935 49.785 529.515 50.305 ;
        RECT 529.685 49.615 532.280 50.135 ;
        RECT 532.455 49.785 532.975 50.325 ;
        RECT 533.145 49.615 533.665 50.155 ;
        RECT 521.415 48.525 526.760 49.615 ;
        RECT 526.935 48.525 532.280 49.615 ;
        RECT 532.455 48.525 533.665 49.615 ;
        RECT 533.835 48.525 534.125 49.690 ;
        RECT 534.755 49.420 535.275 50.905 ;
        RECT 535.445 50.415 535.785 51.075 ;
        RECT 536.135 50.305 541.480 51.075 ;
        RECT 534.945 48.525 535.275 49.250 ;
        RECT 535.445 48.695 535.965 50.245 ;
        RECT 536.135 49.785 538.715 50.305 ;
        RECT 538.885 49.615 541.480 50.135 ;
        RECT 536.135 48.525 541.480 49.615 ;
        RECT 542.115 49.420 542.635 50.905 ;
        RECT 542.805 50.415 543.145 51.075 ;
        RECT 543.495 50.305 548.840 51.075 ;
        RECT 549.015 50.305 552.525 51.075 ;
        RECT 542.305 48.525 542.635 49.250 ;
        RECT 542.805 48.695 543.325 50.245 ;
        RECT 543.495 49.785 546.075 50.305 ;
        RECT 546.245 49.615 548.840 50.135 ;
        RECT 549.015 49.785 550.665 50.305 ;
        RECT 550.835 49.615 552.525 50.135 ;
        RECT 543.495 48.525 548.840 49.615 ;
        RECT 549.015 48.525 552.525 49.615 ;
        RECT 553.155 49.420 553.675 50.905 ;
        RECT 553.845 50.415 554.185 51.075 ;
        RECT 554.535 50.305 559.880 51.075 ;
        RECT 560.055 50.305 561.725 51.075 ;
        RECT 561.895 50.350 562.185 51.075 ;
        RECT 562.355 50.325 563.565 51.075 ;
        RECT 553.345 48.525 553.675 49.250 ;
        RECT 553.845 48.695 554.365 50.245 ;
        RECT 554.535 49.785 557.115 50.305 ;
        RECT 557.285 49.615 559.880 50.135 ;
        RECT 560.055 49.785 560.805 50.305 ;
        RECT 560.975 49.615 561.725 50.135 ;
        RECT 562.355 49.785 562.875 50.325 ;
        RECT 554.535 48.525 559.880 49.615 ;
        RECT 560.055 48.525 561.725 49.615 ;
        RECT 561.895 48.525 562.185 49.690 ;
        RECT 563.045 49.615 563.565 50.155 ;
        RECT 562.355 48.525 563.565 49.615 ;
        RECT 563.735 49.420 564.255 50.905 ;
        RECT 564.425 50.415 564.765 51.075 ;
        RECT 565.115 50.305 570.460 51.075 ;
        RECT 563.925 48.525 564.255 49.250 ;
        RECT 564.425 48.695 564.945 50.245 ;
        RECT 565.115 49.785 567.695 50.305 ;
        RECT 567.865 49.615 570.460 50.135 ;
        RECT 565.115 48.525 570.460 49.615 ;
        RECT 571.095 49.420 571.615 50.905 ;
        RECT 571.785 50.415 572.125 51.075 ;
        RECT 572.475 50.305 577.820 51.075 ;
        RECT 577.995 50.305 583.340 51.075 ;
        RECT 583.515 50.305 588.860 51.075 ;
        RECT 589.955 50.350 590.245 51.075 ;
        RECT 590.415 50.305 595.760 51.075 ;
        RECT 571.285 48.525 571.615 49.250 ;
        RECT 571.785 48.695 572.305 50.245 ;
        RECT 572.475 49.785 575.055 50.305 ;
        RECT 575.225 49.615 577.820 50.135 ;
        RECT 577.995 49.785 580.575 50.305 ;
        RECT 580.745 49.615 583.340 50.135 ;
        RECT 583.515 49.785 586.095 50.305 ;
        RECT 586.265 49.615 588.860 50.135 ;
        RECT 590.415 49.785 592.995 50.305 ;
        RECT 572.475 48.525 577.820 49.615 ;
        RECT 577.995 48.525 583.340 49.615 ;
        RECT 583.515 48.525 588.860 49.615 ;
        RECT 589.955 48.525 590.245 49.690 ;
        RECT 593.165 49.615 595.760 50.135 ;
        RECT 590.415 48.525 595.760 49.615 ;
        RECT 596.855 49.420 597.375 50.905 ;
        RECT 597.545 50.415 597.885 51.075 ;
        RECT 598.235 50.305 603.580 51.075 ;
        RECT 597.045 48.525 597.375 49.250 ;
        RECT 597.545 48.695 598.065 50.245 ;
        RECT 598.235 49.785 600.815 50.305 ;
        RECT 600.985 49.615 603.580 50.135 ;
        RECT 598.235 48.525 603.580 49.615 ;
        RECT 604.215 49.420 604.735 50.905 ;
        RECT 604.905 50.415 605.245 51.075 ;
        RECT 605.595 50.305 610.940 51.075 ;
        RECT 611.115 50.305 616.460 51.075 ;
        RECT 616.635 50.325 617.845 51.075 ;
        RECT 618.015 50.350 618.305 51.075 ;
        RECT 605.595 49.785 608.175 50.305 ;
        RECT 608.345 49.615 610.940 50.135 ;
        RECT 611.115 49.785 613.695 50.305 ;
        RECT 613.865 49.615 616.460 50.135 ;
        RECT 616.635 49.785 617.155 50.325 ;
        RECT 617.325 49.615 617.845 50.155 ;
        RECT 604.405 48.525 604.735 49.250 ;
        RECT 605.595 48.525 610.940 49.615 ;
        RECT 611.115 48.525 616.460 49.615 ;
        RECT 616.635 48.525 617.845 49.615 ;
        RECT 618.015 48.525 618.305 49.690 ;
        RECT 618.935 49.420 619.455 50.905 ;
        RECT 619.625 50.415 619.965 51.075 ;
        RECT 620.315 50.305 623.825 51.075 ;
        RECT 619.125 48.525 619.455 49.250 ;
        RECT 619.625 48.695 620.145 50.245 ;
        RECT 620.315 49.785 621.965 50.305 ;
        RECT 622.135 49.615 623.825 50.135 ;
        RECT 620.315 48.525 623.825 49.615 ;
        RECT 623.995 49.420 624.515 50.905 ;
        RECT 624.685 50.415 625.025 51.075 ;
        RECT 625.375 50.305 628.885 51.075 ;
        RECT 629.975 50.325 631.185 51.075 ;
        RECT 624.185 48.525 624.515 49.250 ;
        RECT 624.685 48.695 625.205 50.245 ;
        RECT 625.375 49.785 627.025 50.305 ;
        RECT 627.195 49.615 628.885 50.135 ;
        RECT 625.375 48.525 628.885 49.615 ;
        RECT 629.975 49.615 630.495 50.155 ;
        RECT 630.665 49.785 631.185 50.325 ;
        RECT 629.975 48.525 631.185 49.615 ;
        RECT 42.470 48.355 631.270 48.525 ;
        RECT 42.555 47.265 43.765 48.355 ;
        RECT 43.935 47.265 49.280 48.355 ;
        RECT 49.455 47.265 54.800 48.355 ;
        RECT 54.975 47.265 60.320 48.355 ;
        RECT 60.495 47.265 65.840 48.355 ;
        RECT 66.015 47.265 69.525 48.355 ;
        RECT 42.555 46.555 43.075 47.095 ;
        RECT 43.245 46.725 43.765 47.265 ;
        RECT 43.935 46.575 46.515 47.095 ;
        RECT 46.685 46.745 49.280 47.265 ;
        RECT 49.455 46.575 52.035 47.095 ;
        RECT 52.205 46.745 54.800 47.265 ;
        RECT 54.975 46.575 57.555 47.095 ;
        RECT 57.725 46.745 60.320 47.265 ;
        RECT 60.495 46.575 63.075 47.095 ;
        RECT 63.245 46.745 65.840 47.265 ;
        RECT 66.015 46.575 67.665 47.095 ;
        RECT 67.835 46.745 69.525 47.265 ;
        RECT 70.615 47.190 70.905 48.355 ;
        RECT 71.075 47.265 72.285 48.355 ;
        RECT 42.555 45.805 43.765 46.555 ;
        RECT 43.935 45.805 49.280 46.575 ;
        RECT 49.455 45.805 54.800 46.575 ;
        RECT 54.975 45.805 60.320 46.575 ;
        RECT 60.495 45.805 65.840 46.575 ;
        RECT 66.015 45.805 69.525 46.575 ;
        RECT 71.075 46.555 71.595 47.095 ;
        RECT 71.765 46.725 72.285 47.265 ;
        RECT 72.495 47.215 72.725 48.355 ;
        RECT 72.895 47.205 73.225 48.185 ;
        RECT 73.395 47.215 73.605 48.355 ;
        RECT 73.835 47.265 77.345 48.355 ;
        RECT 77.525 47.600 77.855 48.355 ;
        RECT 78.035 47.470 78.215 48.185 ;
        RECT 78.420 47.655 78.750 48.355 ;
        RECT 78.960 47.480 79.150 48.185 ;
        RECT 79.320 47.655 79.650 48.355 ;
        RECT 79.820 47.485 80.010 48.185 ;
        RECT 80.180 47.655 80.510 48.355 ;
        RECT 79.820 47.480 80.565 47.485 ;
        RECT 72.475 46.795 72.805 47.045 ;
        RECT 70.615 45.805 70.905 46.530 ;
        RECT 71.075 45.805 72.285 46.555 ;
        RECT 72.495 45.805 72.725 46.625 ;
        RECT 72.975 46.605 73.225 47.205 ;
        RECT 72.895 45.975 73.225 46.605 ;
        RECT 73.395 45.805 73.605 46.625 ;
        RECT 73.835 46.575 75.485 47.095 ;
        RECT 75.655 46.745 77.345 47.265 ;
        RECT 77.555 46.715 77.865 47.335 ;
        RECT 78.035 47.300 78.790 47.470 ;
        RECT 78.580 47.075 78.790 47.300 ;
        RECT 78.960 47.255 80.565 47.480 ;
        RECT 80.735 47.265 84.245 48.355 ;
        RECT 78.035 46.715 78.410 47.045 ;
        RECT 78.580 46.740 80.115 47.075 ;
        RECT 73.835 45.805 77.345 46.575 ;
        RECT 78.580 46.525 78.790 46.740 ;
        RECT 80.285 46.565 80.565 47.255 ;
        RECT 77.525 46.335 78.790 46.525 ;
        RECT 78.960 46.335 80.565 46.565 ;
        RECT 80.735 46.575 82.385 47.095 ;
        RECT 82.555 46.745 84.245 47.265 ;
        RECT 85.425 47.425 85.595 48.185 ;
        RECT 85.810 47.595 86.140 48.355 ;
        RECT 85.425 47.255 86.140 47.425 ;
        RECT 86.310 47.280 86.565 48.185 ;
        RECT 85.335 46.705 85.690 47.075 ;
        RECT 85.970 47.045 86.140 47.255 ;
        RECT 85.970 46.715 86.225 47.045 ;
        RECT 77.525 45.975 77.855 46.335 ;
        RECT 78.960 46.235 79.150 46.335 ;
        RECT 78.385 45.805 78.715 46.165 ;
        RECT 79.320 45.805 79.650 46.165 ;
        RECT 79.820 45.975 80.010 46.335 ;
        RECT 80.180 45.805 80.510 46.165 ;
        RECT 80.735 45.805 84.245 46.575 ;
        RECT 85.970 46.525 86.140 46.715 ;
        RECT 86.395 46.550 86.565 47.280 ;
        RECT 86.740 47.205 87.000 48.355 ;
        RECT 87.175 47.265 90.685 48.355 ;
        RECT 85.425 46.355 86.140 46.525 ;
        RECT 85.425 45.975 85.595 46.355 ;
        RECT 85.810 45.805 86.140 46.185 ;
        RECT 86.310 45.975 86.565 46.550 ;
        RECT 86.740 45.805 87.000 46.645 ;
        RECT 87.175 46.575 88.825 47.095 ;
        RECT 88.995 46.745 90.685 47.265 ;
        RECT 90.860 47.385 91.135 48.185 ;
        RECT 91.305 47.555 91.635 48.355 ;
        RECT 91.805 47.385 91.975 48.185 ;
        RECT 92.145 47.555 92.395 48.355 ;
        RECT 92.565 48.015 94.660 48.185 ;
        RECT 92.565 47.385 92.895 48.015 ;
        RECT 90.860 47.175 92.895 47.385 ;
        RECT 93.065 47.465 93.235 47.845 ;
        RECT 93.405 47.655 93.735 48.015 ;
        RECT 93.905 47.465 94.075 47.845 ;
        RECT 94.245 47.635 94.660 48.015 ;
        RECT 93.065 47.165 94.825 47.465 ;
        RECT 94.995 47.265 98.505 48.355 ;
        RECT 90.910 46.795 92.570 46.995 ;
        RECT 92.890 46.795 94.255 46.995 ;
        RECT 94.425 46.625 94.825 47.165 ;
        RECT 87.175 45.805 90.685 46.575 ;
        RECT 90.860 45.805 91.135 46.625 ;
        RECT 91.305 46.445 94.825 46.625 ;
        RECT 94.995 46.575 96.645 47.095 ;
        RECT 96.815 46.745 98.505 47.265 ;
        RECT 98.675 47.190 98.965 48.355 ;
        RECT 99.135 47.265 102.645 48.355 ;
        RECT 99.135 46.575 100.785 47.095 ;
        RECT 100.955 46.745 102.645 47.265 ;
        RECT 103.280 47.385 103.555 48.185 ;
        RECT 103.725 47.555 104.055 48.355 ;
        RECT 104.225 47.385 104.395 48.185 ;
        RECT 104.565 47.555 104.815 48.355 ;
        RECT 104.985 48.015 107.080 48.185 ;
        RECT 104.985 47.385 105.315 48.015 ;
        RECT 103.280 47.175 105.315 47.385 ;
        RECT 105.485 47.465 105.655 47.845 ;
        RECT 105.825 47.655 106.155 48.015 ;
        RECT 106.325 47.465 106.495 47.845 ;
        RECT 106.665 47.635 107.080 48.015 ;
        RECT 105.485 47.165 107.245 47.465 ;
        RECT 107.415 47.265 110.925 48.355 ;
        RECT 103.330 46.795 104.990 46.995 ;
        RECT 105.310 46.795 106.675 46.995 ;
        RECT 106.845 46.625 107.245 47.165 ;
        RECT 91.305 45.975 91.635 46.445 ;
        RECT 91.805 45.805 91.975 46.275 ;
        RECT 92.145 45.975 92.475 46.445 ;
        RECT 92.645 45.805 92.815 46.275 ;
        RECT 92.985 45.975 93.315 46.445 ;
        RECT 93.485 45.805 93.655 46.275 ;
        RECT 93.825 45.975 94.155 46.445 ;
        RECT 94.325 45.805 94.610 46.275 ;
        RECT 94.995 45.805 98.505 46.575 ;
        RECT 98.675 45.805 98.965 46.530 ;
        RECT 99.135 45.805 102.645 46.575 ;
        RECT 103.280 45.805 103.555 46.625 ;
        RECT 103.725 46.445 107.245 46.625 ;
        RECT 107.415 46.575 109.065 47.095 ;
        RECT 109.235 46.745 110.925 47.265 ;
        RECT 111.100 47.385 111.375 48.185 ;
        RECT 111.545 47.555 111.875 48.355 ;
        RECT 112.045 47.385 112.215 48.185 ;
        RECT 112.385 47.555 112.635 48.355 ;
        RECT 112.805 48.015 114.900 48.185 ;
        RECT 112.805 47.385 113.135 48.015 ;
        RECT 111.100 47.175 113.135 47.385 ;
        RECT 113.305 47.465 113.475 47.845 ;
        RECT 113.645 47.655 113.975 48.015 ;
        RECT 114.145 47.465 114.315 47.845 ;
        RECT 114.485 47.635 114.900 48.015 ;
        RECT 113.305 47.165 115.065 47.465 ;
        RECT 115.235 47.265 118.745 48.355 ;
        RECT 111.150 46.795 112.810 46.995 ;
        RECT 113.130 46.795 114.495 46.995 ;
        RECT 114.665 46.625 115.065 47.165 ;
        RECT 103.725 45.975 104.055 46.445 ;
        RECT 104.225 45.805 104.395 46.275 ;
        RECT 104.565 45.975 104.895 46.445 ;
        RECT 105.065 45.805 105.235 46.275 ;
        RECT 105.405 45.975 105.735 46.445 ;
        RECT 105.905 45.805 106.075 46.275 ;
        RECT 106.245 45.975 106.575 46.445 ;
        RECT 106.745 45.805 107.030 46.275 ;
        RECT 107.415 45.805 110.925 46.575 ;
        RECT 111.100 45.805 111.375 46.625 ;
        RECT 111.545 46.445 115.065 46.625 ;
        RECT 115.235 46.575 116.885 47.095 ;
        RECT 117.055 46.745 118.745 47.265 ;
        RECT 118.945 47.385 119.280 48.170 ;
        RECT 118.945 47.215 119.540 47.385 ;
        RECT 111.545 45.975 111.875 46.445 ;
        RECT 112.045 45.805 112.215 46.275 ;
        RECT 112.385 45.975 112.715 46.445 ;
        RECT 112.885 45.805 113.055 46.275 ;
        RECT 113.225 45.975 113.555 46.445 ;
        RECT 113.725 45.805 113.895 46.275 ;
        RECT 114.065 45.975 114.395 46.445 ;
        RECT 114.565 45.805 114.850 46.275 ;
        RECT 115.235 45.805 118.745 46.575 ;
        RECT 118.915 46.475 119.200 47.045 ;
        RECT 119.370 46.545 119.540 47.215 ;
        RECT 119.710 47.340 120.060 48.095 ;
        RECT 120.230 47.505 120.550 48.095 ;
        RECT 120.835 47.515 121.085 48.355 ;
        RECT 119.710 46.715 119.880 47.340 ;
        RECT 120.230 47.170 120.440 47.505 ;
        RECT 121.310 47.345 121.560 48.185 ;
        RECT 121.730 47.515 121.980 48.355 ;
        RECT 122.150 47.345 122.400 48.185 ;
        RECT 122.570 47.515 122.820 48.355 ;
        RECT 120.110 46.715 120.440 47.170 ;
        RECT 120.670 47.165 121.105 47.335 ;
        RECT 121.310 47.175 122.885 47.345 ;
        RECT 123.055 47.265 126.565 48.355 ;
        RECT 120.670 46.715 120.840 47.165 ;
        RECT 121.010 46.795 122.470 46.965 ;
        RECT 121.010 46.545 121.180 46.795 ;
        RECT 122.640 46.625 122.885 47.175 ;
        RECT 119.370 46.375 121.180 46.545 ;
        RECT 121.350 46.445 122.885 46.625 ;
        RECT 123.055 46.575 124.705 47.095 ;
        RECT 124.875 46.745 126.565 47.265 ;
        RECT 126.735 47.190 127.025 48.355 ;
        RECT 127.745 47.685 127.915 48.185 ;
        RECT 128.085 47.855 128.415 48.355 ;
        RECT 127.745 47.515 128.410 47.685 ;
        RECT 127.660 46.695 128.010 47.345 ;
        RECT 118.950 45.805 119.200 46.305 ;
        RECT 119.530 46.025 119.700 46.375 ;
        RECT 119.900 45.805 120.230 46.205 ;
        RECT 120.400 46.025 120.570 46.375 ;
        RECT 120.790 45.805 121.170 46.205 ;
        RECT 121.350 45.975 121.600 46.445 ;
        RECT 121.770 45.805 121.940 46.275 ;
        RECT 122.110 45.975 122.440 46.445 ;
        RECT 122.610 45.805 122.780 46.275 ;
        RECT 123.055 45.805 126.565 46.575 ;
        RECT 126.735 45.805 127.025 46.530 ;
        RECT 128.180 46.525 128.410 47.515 ;
        RECT 127.745 46.355 128.410 46.525 ;
        RECT 127.745 46.065 127.915 46.355 ;
        RECT 128.085 45.805 128.415 46.185 ;
        RECT 128.585 46.065 128.810 48.185 ;
        RECT 129.010 47.895 129.275 48.355 ;
        RECT 129.460 47.785 129.695 48.160 ;
        RECT 129.940 47.910 131.010 48.080 ;
        RECT 129.010 46.785 129.290 47.385 ;
        RECT 129.025 45.805 129.275 46.265 ;
        RECT 129.460 46.255 129.630 47.785 ;
        RECT 129.800 46.755 130.040 47.625 ;
        RECT 130.230 47.375 130.670 47.730 ;
        RECT 130.840 47.295 131.010 47.910 ;
        RECT 131.180 47.555 131.350 48.355 ;
        RECT 131.520 47.855 131.770 48.185 ;
        RECT 131.995 47.885 132.880 48.055 ;
        RECT 130.840 47.205 131.350 47.295 ;
        RECT 130.550 47.035 131.350 47.205 ;
        RECT 129.800 46.425 130.380 46.755 ;
        RECT 130.550 46.255 130.720 47.035 ;
        RECT 131.180 46.965 131.350 47.035 ;
        RECT 130.890 46.785 131.060 46.815 ;
        RECT 131.520 46.785 131.690 47.855 ;
        RECT 131.860 46.965 132.050 47.685 ;
        RECT 132.220 47.295 132.540 47.625 ;
        RECT 130.890 46.485 131.690 46.785 ;
        RECT 132.220 46.755 132.410 47.295 ;
        RECT 129.460 46.085 129.790 46.255 ;
        RECT 129.970 46.085 130.720 46.255 ;
        RECT 130.970 45.805 131.340 46.305 ;
        RECT 131.520 46.255 131.690 46.485 ;
        RECT 131.860 46.425 132.410 46.755 ;
        RECT 132.710 46.965 132.880 47.885 ;
        RECT 133.060 47.855 133.275 48.355 ;
        RECT 133.740 47.550 133.910 48.175 ;
        RECT 134.195 47.575 134.375 48.355 ;
        RECT 133.050 47.390 133.910 47.550 ;
        RECT 133.050 47.220 134.160 47.390 ;
        RECT 133.990 46.965 134.160 47.220 ;
        RECT 134.555 47.355 134.890 48.115 ;
        RECT 135.070 47.525 135.240 48.355 ;
        RECT 135.410 47.355 135.740 48.115 ;
        RECT 135.910 47.525 136.080 48.355 ;
        RECT 134.555 47.185 136.225 47.355 ;
        RECT 136.395 47.265 141.740 48.355 ;
        RECT 141.915 47.265 143.585 48.355 ;
        RECT 143.805 47.675 144.055 48.185 ;
        RECT 144.225 47.845 144.475 48.355 ;
        RECT 144.645 47.675 144.895 48.185 ;
        RECT 145.065 47.845 145.315 48.355 ;
        RECT 145.485 48.015 146.575 48.185 ;
        RECT 145.485 47.675 145.735 48.015 ;
        RECT 146.325 47.855 146.575 48.015 ;
        RECT 146.845 47.855 147.095 48.355 ;
        RECT 147.265 48.015 148.355 48.185 ;
        RECT 147.265 47.855 147.515 48.015 ;
        RECT 143.805 47.505 145.735 47.675 ;
        RECT 132.710 46.795 133.800 46.965 ;
        RECT 133.990 46.795 135.810 46.965 ;
        RECT 132.710 46.255 132.880 46.795 ;
        RECT 133.990 46.625 134.160 46.795 ;
        RECT 133.660 46.455 134.160 46.625 ;
        RECT 135.980 46.620 136.225 47.185 ;
        RECT 131.520 46.085 131.980 46.255 ;
        RECT 132.210 46.085 132.880 46.255 ;
        RECT 133.195 45.805 133.365 46.335 ;
        RECT 133.660 46.015 134.020 46.455 ;
        RECT 134.555 46.450 136.225 46.620 ;
        RECT 136.395 46.575 138.975 47.095 ;
        RECT 139.145 46.745 141.740 47.265 ;
        RECT 141.915 46.575 142.665 47.095 ;
        RECT 142.835 46.745 143.585 47.265 ;
        RECT 143.755 47.165 145.355 47.335 ;
        RECT 145.525 47.175 145.735 47.505 ;
        RECT 145.905 47.685 146.155 47.845 ;
        RECT 147.685 47.685 147.935 47.845 ;
        RECT 143.755 46.795 144.245 47.165 ;
        RECT 145.185 46.995 145.355 47.165 ;
        RECT 145.905 47.135 146.290 47.685 ;
        RECT 146.805 47.505 147.935 47.685 ;
        RECT 148.105 47.505 148.355 48.015 ;
        RECT 148.525 47.515 148.775 48.355 ;
        RECT 148.945 47.675 149.195 48.185 ;
        RECT 149.365 47.885 149.615 48.355 ;
        RECT 149.785 47.675 150.035 48.185 ;
        RECT 148.945 47.505 150.035 47.675 ;
        RECT 150.205 47.545 150.455 48.355 ;
        RECT 146.805 47.385 146.975 47.505 ;
        RECT 146.625 47.215 146.975 47.385 ;
        RECT 149.785 47.375 150.035 47.505 ;
        RECT 144.475 46.795 145.015 46.995 ;
        RECT 145.185 46.965 145.365 46.995 ;
        RECT 145.185 46.795 145.565 46.965 ;
        RECT 145.905 46.625 146.115 47.135 ;
        RECT 146.625 46.965 146.815 47.215 ;
        RECT 147.145 47.165 148.635 47.335 ;
        RECT 147.145 47.045 147.315 47.165 ;
        RECT 146.285 46.795 146.815 46.965 ;
        RECT 146.985 46.795 147.315 47.045 ;
        RECT 147.485 46.795 148.105 46.995 ;
        RECT 148.275 46.795 148.635 47.165 ;
        RECT 148.805 46.965 149.130 47.335 ;
        RECT 149.785 47.135 150.590 47.375 ;
        RECT 151.115 47.265 154.625 48.355 ;
        RECT 148.805 46.795 150.110 46.965 ;
        RECT 146.625 46.625 146.815 46.795 ;
        RECT 150.280 46.625 150.590 47.135 ;
        RECT 134.195 45.805 134.365 46.285 ;
        RECT 134.555 46.025 134.890 46.450 ;
        RECT 135.065 45.805 135.235 46.280 ;
        RECT 135.410 46.025 135.745 46.450 ;
        RECT 135.915 45.805 136.085 46.280 ;
        RECT 136.395 45.805 141.740 46.575 ;
        RECT 141.915 45.805 143.585 46.575 ;
        RECT 143.845 45.805 144.015 46.615 ;
        RECT 144.185 46.195 144.435 46.625 ;
        RECT 144.605 46.455 146.195 46.625 ;
        RECT 144.605 46.365 144.940 46.455 ;
        RECT 144.185 45.975 145.355 46.195 ;
        RECT 145.525 45.805 145.695 46.275 ;
        RECT 145.865 45.975 146.195 46.455 ;
        RECT 146.625 46.445 148.395 46.625 ;
        RECT 146.365 45.805 147.055 46.275 ;
        RECT 147.225 45.975 147.555 46.445 ;
        RECT 147.725 45.805 147.895 46.275 ;
        RECT 148.065 45.975 148.395 46.445 ;
        RECT 148.565 45.805 148.735 46.615 ;
        RECT 148.905 46.445 150.590 46.625 ;
        RECT 151.115 46.575 152.765 47.095 ;
        RECT 152.935 46.745 154.625 47.265 ;
        RECT 154.795 47.190 155.085 48.355 ;
        RECT 155.345 47.685 155.515 48.185 ;
        RECT 155.685 47.855 156.015 48.355 ;
        RECT 155.345 47.515 156.010 47.685 ;
        RECT 155.260 46.695 155.610 47.345 ;
        RECT 148.905 45.995 149.235 46.445 ;
        RECT 149.405 45.805 149.575 46.275 ;
        RECT 149.745 45.995 150.075 46.445 ;
        RECT 150.245 45.805 150.415 46.275 ;
        RECT 151.115 45.805 154.625 46.575 ;
        RECT 154.795 45.805 155.085 46.530 ;
        RECT 155.780 46.525 156.010 47.515 ;
        RECT 155.345 46.355 156.010 46.525 ;
        RECT 155.345 46.065 155.515 46.355 ;
        RECT 155.685 45.805 156.015 46.185 ;
        RECT 156.185 46.065 156.410 48.185 ;
        RECT 156.610 47.895 156.875 48.355 ;
        RECT 157.060 47.785 157.295 48.160 ;
        RECT 157.540 47.910 158.610 48.080 ;
        RECT 156.610 46.785 156.890 47.385 ;
        RECT 156.625 45.805 156.875 46.265 ;
        RECT 157.060 46.255 157.230 47.785 ;
        RECT 157.400 46.755 157.640 47.625 ;
        RECT 157.830 47.375 158.270 47.730 ;
        RECT 158.440 47.295 158.610 47.910 ;
        RECT 158.780 47.555 158.950 48.355 ;
        RECT 159.120 47.855 159.370 48.185 ;
        RECT 159.595 47.885 160.480 48.055 ;
        RECT 158.440 47.205 158.950 47.295 ;
        RECT 158.150 47.035 158.950 47.205 ;
        RECT 157.400 46.425 157.980 46.755 ;
        RECT 158.150 46.255 158.320 47.035 ;
        RECT 158.780 46.965 158.950 47.035 ;
        RECT 158.490 46.785 158.660 46.815 ;
        RECT 159.120 46.785 159.290 47.855 ;
        RECT 159.460 46.965 159.650 47.685 ;
        RECT 159.820 47.295 160.140 47.625 ;
        RECT 158.490 46.485 159.290 46.785 ;
        RECT 159.820 46.755 160.010 47.295 ;
        RECT 157.060 46.085 157.390 46.255 ;
        RECT 157.570 46.085 158.320 46.255 ;
        RECT 158.570 45.805 158.940 46.305 ;
        RECT 159.120 46.255 159.290 46.485 ;
        RECT 159.460 46.425 160.010 46.755 ;
        RECT 160.310 46.965 160.480 47.885 ;
        RECT 160.660 47.855 160.875 48.355 ;
        RECT 161.340 47.550 161.510 48.175 ;
        RECT 161.795 47.575 161.975 48.355 ;
        RECT 160.650 47.390 161.510 47.550 ;
        RECT 160.650 47.220 161.760 47.390 ;
        RECT 161.590 46.965 161.760 47.220 ;
        RECT 162.155 47.355 162.490 48.115 ;
        RECT 162.670 47.525 162.840 48.355 ;
        RECT 163.010 47.355 163.340 48.115 ;
        RECT 163.510 47.525 163.680 48.355 ;
        RECT 162.155 47.185 163.825 47.355 ;
        RECT 163.995 47.265 167.505 48.355 ;
        RECT 167.675 47.265 168.885 48.355 ;
        RECT 169.145 47.685 169.315 48.185 ;
        RECT 169.485 47.855 169.815 48.355 ;
        RECT 169.145 47.515 169.810 47.685 ;
        RECT 160.310 46.795 161.400 46.965 ;
        RECT 161.590 46.795 163.410 46.965 ;
        RECT 160.310 46.255 160.480 46.795 ;
        RECT 161.590 46.625 161.760 46.795 ;
        RECT 161.260 46.455 161.760 46.625 ;
        RECT 163.580 46.620 163.825 47.185 ;
        RECT 159.120 46.085 159.580 46.255 ;
        RECT 159.810 46.085 160.480 46.255 ;
        RECT 160.795 45.805 160.965 46.335 ;
        RECT 161.260 46.015 161.620 46.455 ;
        RECT 162.155 46.450 163.825 46.620 ;
        RECT 163.995 46.575 165.645 47.095 ;
        RECT 165.815 46.745 167.505 47.265 ;
        RECT 161.795 45.805 161.965 46.285 ;
        RECT 162.155 46.025 162.490 46.450 ;
        RECT 162.665 45.805 162.835 46.280 ;
        RECT 163.010 46.025 163.345 46.450 ;
        RECT 163.515 45.805 163.685 46.280 ;
        RECT 163.995 45.805 167.505 46.575 ;
        RECT 167.675 46.555 168.195 47.095 ;
        RECT 168.365 46.725 168.885 47.265 ;
        RECT 169.060 46.695 169.410 47.345 ;
        RECT 167.675 45.805 168.885 46.555 ;
        RECT 169.580 46.525 169.810 47.515 ;
        RECT 169.145 46.355 169.810 46.525 ;
        RECT 169.145 46.065 169.315 46.355 ;
        RECT 169.485 45.805 169.815 46.185 ;
        RECT 169.985 46.065 170.210 48.185 ;
        RECT 170.410 47.895 170.675 48.355 ;
        RECT 170.860 47.785 171.095 48.160 ;
        RECT 171.340 47.910 172.410 48.080 ;
        RECT 170.410 46.785 170.690 47.385 ;
        RECT 170.425 45.805 170.675 46.265 ;
        RECT 170.860 46.255 171.030 47.785 ;
        RECT 171.200 46.755 171.440 47.625 ;
        RECT 171.630 47.375 172.070 47.730 ;
        RECT 172.240 47.295 172.410 47.910 ;
        RECT 172.580 47.555 172.750 48.355 ;
        RECT 172.920 47.855 173.170 48.185 ;
        RECT 173.395 47.885 174.280 48.055 ;
        RECT 172.240 47.205 172.750 47.295 ;
        RECT 171.950 47.035 172.750 47.205 ;
        RECT 171.200 46.425 171.780 46.755 ;
        RECT 171.950 46.255 172.120 47.035 ;
        RECT 172.580 46.965 172.750 47.035 ;
        RECT 172.290 46.785 172.460 46.815 ;
        RECT 172.920 46.785 173.090 47.855 ;
        RECT 173.260 46.965 173.450 47.685 ;
        RECT 173.620 47.295 173.940 47.625 ;
        RECT 172.290 46.485 173.090 46.785 ;
        RECT 173.620 46.755 173.810 47.295 ;
        RECT 170.860 46.085 171.190 46.255 ;
        RECT 171.370 46.085 172.120 46.255 ;
        RECT 172.370 45.805 172.740 46.305 ;
        RECT 172.920 46.255 173.090 46.485 ;
        RECT 173.260 46.425 173.810 46.755 ;
        RECT 174.110 46.965 174.280 47.885 ;
        RECT 174.460 47.855 174.675 48.355 ;
        RECT 175.140 47.550 175.310 48.175 ;
        RECT 175.595 47.575 175.775 48.355 ;
        RECT 174.450 47.390 175.310 47.550 ;
        RECT 176.470 47.525 176.640 48.355 ;
        RECT 177.310 47.525 177.480 48.355 ;
        RECT 174.450 47.220 175.560 47.390 ;
        RECT 177.795 47.265 181.305 48.355 ;
        RECT 181.475 47.265 182.685 48.355 ;
        RECT 175.390 46.965 175.560 47.220 ;
        RECT 174.110 46.795 175.200 46.965 ;
        RECT 175.390 46.795 177.210 46.965 ;
        RECT 174.110 46.255 174.280 46.795 ;
        RECT 175.390 46.625 175.560 46.795 ;
        RECT 175.060 46.455 175.560 46.625 ;
        RECT 177.795 46.575 179.445 47.095 ;
        RECT 179.615 46.745 181.305 47.265 ;
        RECT 172.920 46.085 173.380 46.255 ;
        RECT 173.610 46.085 174.280 46.255 ;
        RECT 174.595 45.805 174.765 46.335 ;
        RECT 175.060 46.015 175.420 46.455 ;
        RECT 175.595 45.805 175.765 46.285 ;
        RECT 176.465 45.805 176.635 46.280 ;
        RECT 177.315 45.805 177.485 46.280 ;
        RECT 177.795 45.805 181.305 46.575 ;
        RECT 181.475 46.555 181.995 47.095 ;
        RECT 182.165 46.725 182.685 47.265 ;
        RECT 182.855 47.190 183.145 48.355 ;
        RECT 183.315 47.265 184.525 48.355 ;
        RECT 184.785 47.685 184.955 48.185 ;
        RECT 185.125 47.855 185.455 48.355 ;
        RECT 184.785 47.515 185.450 47.685 ;
        RECT 183.315 46.555 183.835 47.095 ;
        RECT 184.005 46.725 184.525 47.265 ;
        RECT 184.700 46.695 185.050 47.345 ;
        RECT 181.475 45.805 182.685 46.555 ;
        RECT 182.855 45.805 183.145 46.530 ;
        RECT 183.315 45.805 184.525 46.555 ;
        RECT 185.220 46.525 185.450 47.515 ;
        RECT 184.785 46.355 185.450 46.525 ;
        RECT 184.785 46.065 184.955 46.355 ;
        RECT 185.125 45.805 185.455 46.185 ;
        RECT 185.625 46.065 185.850 48.185 ;
        RECT 186.050 47.895 186.315 48.355 ;
        RECT 186.500 47.785 186.735 48.160 ;
        RECT 186.980 47.910 188.050 48.080 ;
        RECT 186.050 46.785 186.330 47.385 ;
        RECT 186.065 45.805 186.315 46.265 ;
        RECT 186.500 46.255 186.670 47.785 ;
        RECT 186.840 46.755 187.080 47.625 ;
        RECT 187.270 47.375 187.710 47.730 ;
        RECT 187.880 47.295 188.050 47.910 ;
        RECT 188.220 47.555 188.390 48.355 ;
        RECT 188.560 47.855 188.810 48.185 ;
        RECT 189.035 47.885 189.920 48.055 ;
        RECT 187.880 47.205 188.390 47.295 ;
        RECT 187.590 47.035 188.390 47.205 ;
        RECT 186.840 46.425 187.420 46.755 ;
        RECT 187.590 46.255 187.760 47.035 ;
        RECT 188.220 46.965 188.390 47.035 ;
        RECT 187.930 46.785 188.100 46.815 ;
        RECT 188.560 46.785 188.730 47.855 ;
        RECT 188.900 46.965 189.090 47.685 ;
        RECT 189.260 47.295 189.580 47.625 ;
        RECT 187.930 46.485 188.730 46.785 ;
        RECT 189.260 46.755 189.450 47.295 ;
        RECT 186.500 46.085 186.830 46.255 ;
        RECT 187.010 46.085 187.760 46.255 ;
        RECT 188.010 45.805 188.380 46.305 ;
        RECT 188.560 46.255 188.730 46.485 ;
        RECT 188.900 46.425 189.450 46.755 ;
        RECT 189.750 46.965 189.920 47.885 ;
        RECT 190.100 47.855 190.315 48.355 ;
        RECT 190.780 47.550 190.950 48.175 ;
        RECT 191.235 47.575 191.415 48.355 ;
        RECT 190.090 47.390 190.950 47.550 ;
        RECT 190.090 47.220 191.200 47.390 ;
        RECT 191.030 46.965 191.200 47.220 ;
        RECT 191.595 47.355 191.930 48.115 ;
        RECT 192.110 47.525 192.280 48.355 ;
        RECT 192.450 47.355 192.780 48.115 ;
        RECT 192.950 47.525 193.120 48.355 ;
        RECT 191.595 47.185 193.265 47.355 ;
        RECT 193.435 47.265 196.945 48.355 ;
        RECT 197.205 47.685 197.375 48.185 ;
        RECT 197.545 47.855 197.875 48.355 ;
        RECT 197.205 47.515 197.870 47.685 ;
        RECT 189.750 46.795 190.840 46.965 ;
        RECT 191.030 46.795 192.850 46.965 ;
        RECT 189.750 46.255 189.920 46.795 ;
        RECT 191.030 46.625 191.200 46.795 ;
        RECT 190.700 46.455 191.200 46.625 ;
        RECT 193.020 46.620 193.265 47.185 ;
        RECT 188.560 46.085 189.020 46.255 ;
        RECT 189.250 46.085 189.920 46.255 ;
        RECT 190.235 45.805 190.405 46.335 ;
        RECT 190.700 46.015 191.060 46.455 ;
        RECT 191.595 46.450 193.265 46.620 ;
        RECT 193.435 46.575 195.085 47.095 ;
        RECT 195.255 46.745 196.945 47.265 ;
        RECT 197.120 46.695 197.470 47.345 ;
        RECT 191.235 45.805 191.405 46.285 ;
        RECT 191.595 46.025 191.930 46.450 ;
        RECT 192.105 45.805 192.275 46.280 ;
        RECT 192.450 46.025 192.785 46.450 ;
        RECT 192.955 45.805 193.125 46.280 ;
        RECT 193.435 45.805 196.945 46.575 ;
        RECT 197.640 46.525 197.870 47.515 ;
        RECT 197.205 46.355 197.870 46.525 ;
        RECT 197.205 46.065 197.375 46.355 ;
        RECT 197.545 45.805 197.875 46.185 ;
        RECT 198.045 46.065 198.270 48.185 ;
        RECT 198.470 47.895 198.735 48.355 ;
        RECT 198.920 47.785 199.155 48.160 ;
        RECT 199.400 47.910 200.470 48.080 ;
        RECT 198.470 46.785 198.750 47.385 ;
        RECT 198.485 45.805 198.735 46.265 ;
        RECT 198.920 46.255 199.090 47.785 ;
        RECT 199.260 46.755 199.500 47.625 ;
        RECT 199.690 47.375 200.130 47.730 ;
        RECT 200.300 47.295 200.470 47.910 ;
        RECT 200.640 47.555 200.810 48.355 ;
        RECT 200.980 47.855 201.230 48.185 ;
        RECT 201.455 47.885 202.340 48.055 ;
        RECT 200.300 47.205 200.810 47.295 ;
        RECT 200.010 47.035 200.810 47.205 ;
        RECT 199.260 46.425 199.840 46.755 ;
        RECT 200.010 46.255 200.180 47.035 ;
        RECT 200.640 46.965 200.810 47.035 ;
        RECT 200.350 46.785 200.520 46.815 ;
        RECT 200.980 46.785 201.150 47.855 ;
        RECT 201.320 46.965 201.510 47.685 ;
        RECT 201.680 47.295 202.000 47.625 ;
        RECT 200.350 46.485 201.150 46.785 ;
        RECT 201.680 46.755 201.870 47.295 ;
        RECT 198.920 46.085 199.250 46.255 ;
        RECT 199.430 46.085 200.180 46.255 ;
        RECT 200.430 45.805 200.800 46.305 ;
        RECT 200.980 46.255 201.150 46.485 ;
        RECT 201.320 46.425 201.870 46.755 ;
        RECT 202.170 46.965 202.340 47.885 ;
        RECT 202.520 47.855 202.735 48.355 ;
        RECT 203.200 47.550 203.370 48.175 ;
        RECT 203.655 47.575 203.835 48.355 ;
        RECT 202.510 47.390 203.370 47.550 ;
        RECT 202.510 47.220 203.620 47.390 ;
        RECT 203.450 46.965 203.620 47.220 ;
        RECT 204.015 47.355 204.350 48.115 ;
        RECT 204.530 47.525 204.700 48.355 ;
        RECT 204.870 47.355 205.200 48.115 ;
        RECT 205.370 47.525 205.540 48.355 ;
        RECT 204.015 47.185 205.685 47.355 ;
        RECT 205.855 47.265 209.365 48.355 ;
        RECT 209.535 47.265 210.745 48.355 ;
        RECT 202.170 46.795 203.260 46.965 ;
        RECT 203.450 46.795 205.270 46.965 ;
        RECT 202.170 46.255 202.340 46.795 ;
        RECT 203.450 46.625 203.620 46.795 ;
        RECT 203.120 46.455 203.620 46.625 ;
        RECT 205.440 46.620 205.685 47.185 ;
        RECT 200.980 46.085 201.440 46.255 ;
        RECT 201.670 46.085 202.340 46.255 ;
        RECT 202.655 45.805 202.825 46.335 ;
        RECT 203.120 46.015 203.480 46.455 ;
        RECT 204.015 46.450 205.685 46.620 ;
        RECT 205.855 46.575 207.505 47.095 ;
        RECT 207.675 46.745 209.365 47.265 ;
        RECT 203.655 45.805 203.825 46.285 ;
        RECT 204.015 46.025 204.350 46.450 ;
        RECT 204.525 45.805 204.695 46.280 ;
        RECT 204.870 46.025 205.205 46.450 ;
        RECT 205.375 45.805 205.545 46.280 ;
        RECT 205.855 45.805 209.365 46.575 ;
        RECT 209.535 46.555 210.055 47.095 ;
        RECT 210.225 46.725 210.745 47.265 ;
        RECT 210.915 47.190 211.205 48.355 ;
        RECT 211.405 47.385 211.740 48.170 ;
        RECT 211.405 47.215 212.000 47.385 ;
        RECT 209.535 45.805 210.745 46.555 ;
        RECT 210.915 45.805 211.205 46.530 ;
        RECT 211.375 46.475 211.660 47.045 ;
        RECT 211.830 46.545 212.000 47.215 ;
        RECT 212.170 47.340 212.520 48.095 ;
        RECT 212.690 47.505 213.010 48.095 ;
        RECT 213.295 47.515 213.545 48.355 ;
        RECT 212.170 46.715 212.340 47.340 ;
        RECT 212.690 47.170 212.900 47.505 ;
        RECT 213.770 47.345 214.020 48.185 ;
        RECT 214.190 47.515 214.440 48.355 ;
        RECT 214.610 47.345 214.860 48.185 ;
        RECT 215.030 47.515 215.280 48.355 ;
        RECT 212.570 46.715 212.900 47.170 ;
        RECT 213.130 47.165 213.565 47.335 ;
        RECT 213.770 47.175 215.345 47.345 ;
        RECT 215.515 47.265 219.025 48.355 ;
        RECT 213.130 46.715 213.300 47.165 ;
        RECT 213.470 46.795 214.930 46.965 ;
        RECT 213.470 46.545 213.640 46.795 ;
        RECT 215.100 46.625 215.345 47.175 ;
        RECT 211.830 46.375 213.640 46.545 ;
        RECT 213.810 46.445 215.345 46.625 ;
        RECT 215.515 46.575 217.165 47.095 ;
        RECT 217.335 46.745 219.025 47.265 ;
        RECT 219.225 47.060 219.475 48.055 ;
        RECT 219.655 47.470 219.835 48.185 ;
        RECT 220.005 47.655 220.455 48.355 ;
        RECT 220.630 47.470 220.810 48.185 ;
        RECT 221.020 47.655 221.350 48.355 ;
        RECT 221.560 47.480 221.750 48.185 ;
        RECT 221.920 47.655 222.250 48.355 ;
        RECT 222.420 47.485 222.610 48.185 ;
        RECT 222.780 47.655 223.110 48.355 ;
        RECT 222.420 47.480 223.165 47.485 ;
        RECT 219.655 47.300 221.390 47.470 ;
        RECT 221.180 47.075 221.390 47.300 ;
        RECT 221.560 47.255 223.165 47.480 ;
        RECT 223.335 47.265 228.680 48.355 ;
        RECT 228.855 47.265 230.525 48.355 ;
        RECT 219.225 46.715 219.985 47.060 ;
        RECT 211.410 45.805 211.660 46.305 ;
        RECT 211.990 46.025 212.160 46.375 ;
        RECT 212.360 45.805 212.690 46.205 ;
        RECT 212.860 46.025 213.030 46.375 ;
        RECT 213.250 45.805 213.630 46.205 ;
        RECT 213.810 45.975 214.060 46.445 ;
        RECT 214.230 45.805 214.400 46.275 ;
        RECT 214.570 45.975 214.900 46.445 ;
        RECT 215.070 45.805 215.240 46.275 ;
        RECT 215.515 45.805 219.025 46.575 ;
        RECT 219.575 46.285 219.910 46.525 ;
        RECT 220.175 46.465 220.465 47.060 ;
        RECT 220.635 46.715 221.010 47.045 ;
        RECT 221.180 46.740 222.715 47.075 ;
        RECT 221.180 46.525 221.390 46.740 ;
        RECT 222.885 46.565 223.165 47.255 ;
        RECT 220.645 46.335 221.390 46.525 ;
        RECT 221.560 46.335 223.165 46.565 ;
        RECT 223.335 46.575 225.915 47.095 ;
        RECT 226.085 46.745 228.680 47.265 ;
        RECT 228.855 46.575 229.605 47.095 ;
        RECT 229.775 46.745 230.525 47.265 ;
        RECT 230.725 47.385 231.060 48.170 ;
        RECT 230.725 47.215 231.320 47.385 ;
        RECT 220.645 46.285 220.835 46.335 ;
        RECT 219.575 46.095 220.835 46.285 ;
        RECT 221.560 46.235 221.750 46.335 ;
        RECT 219.575 45.975 219.910 46.095 ;
        RECT 221.015 45.805 221.345 46.165 ;
        RECT 221.920 45.805 222.250 46.165 ;
        RECT 222.420 45.975 222.610 46.335 ;
        RECT 222.780 45.805 223.110 46.165 ;
        RECT 223.335 45.805 228.680 46.575 ;
        RECT 228.855 45.805 230.525 46.575 ;
        RECT 230.695 46.475 230.980 47.045 ;
        RECT 231.150 46.545 231.320 47.215 ;
        RECT 231.490 47.340 231.840 48.095 ;
        RECT 232.010 47.505 232.330 48.095 ;
        RECT 232.615 47.515 232.865 48.355 ;
        RECT 231.490 46.715 231.660 47.340 ;
        RECT 232.010 47.170 232.220 47.505 ;
        RECT 233.090 47.345 233.340 48.185 ;
        RECT 233.510 47.515 233.760 48.355 ;
        RECT 233.930 47.345 234.180 48.185 ;
        RECT 234.350 47.515 234.600 48.355 ;
        RECT 231.890 46.715 232.220 47.170 ;
        RECT 232.450 47.165 232.885 47.335 ;
        RECT 233.090 47.175 234.665 47.345 ;
        RECT 234.835 47.265 238.345 48.355 ;
        RECT 232.450 46.715 232.620 47.165 ;
        RECT 232.790 46.795 234.250 46.965 ;
        RECT 232.790 46.545 232.960 46.795 ;
        RECT 234.420 46.625 234.665 47.175 ;
        RECT 231.150 46.375 232.960 46.545 ;
        RECT 233.130 46.445 234.665 46.625 ;
        RECT 234.835 46.575 236.485 47.095 ;
        RECT 236.655 46.745 238.345 47.265 ;
        RECT 238.975 47.190 239.265 48.355 ;
        RECT 239.485 47.675 239.735 48.185 ;
        RECT 239.905 47.845 240.155 48.355 ;
        RECT 240.325 47.675 240.575 48.185 ;
        RECT 240.745 47.845 240.995 48.355 ;
        RECT 241.165 48.015 242.255 48.185 ;
        RECT 241.165 47.675 241.415 48.015 ;
        RECT 242.005 47.855 242.255 48.015 ;
        RECT 242.525 47.855 242.775 48.355 ;
        RECT 242.945 48.015 244.035 48.185 ;
        RECT 242.945 47.855 243.195 48.015 ;
        RECT 239.485 47.505 241.415 47.675 ;
        RECT 239.435 47.165 241.035 47.335 ;
        RECT 241.205 47.175 241.415 47.505 ;
        RECT 241.585 47.685 241.835 47.845 ;
        RECT 243.365 47.685 243.615 47.845 ;
        RECT 239.435 46.795 239.925 47.165 ;
        RECT 240.155 46.795 240.695 46.995 ;
        RECT 240.865 46.965 241.035 47.165 ;
        RECT 241.585 47.135 241.970 47.685 ;
        RECT 242.485 47.505 243.615 47.685 ;
        RECT 243.785 47.505 244.035 48.015 ;
        RECT 244.205 47.515 244.455 48.355 ;
        RECT 244.625 47.675 244.875 48.185 ;
        RECT 245.045 47.885 245.295 48.355 ;
        RECT 245.465 47.675 245.715 48.185 ;
        RECT 244.625 47.505 245.715 47.675 ;
        RECT 245.885 47.545 246.135 48.355 ;
        RECT 242.485 47.385 242.655 47.505 ;
        RECT 242.305 47.215 242.655 47.385 ;
        RECT 245.465 47.375 245.715 47.505 ;
        RECT 240.865 46.795 241.245 46.965 ;
        RECT 241.585 46.625 241.795 47.135 ;
        RECT 242.305 46.965 242.495 47.215 ;
        RECT 242.825 47.165 244.315 47.335 ;
        RECT 242.825 47.045 242.995 47.165 ;
        RECT 241.965 46.795 242.495 46.965 ;
        RECT 242.665 46.795 242.995 47.045 ;
        RECT 243.165 46.795 243.785 46.995 ;
        RECT 243.955 46.795 244.315 47.165 ;
        RECT 244.485 46.965 244.810 47.335 ;
        RECT 245.465 47.135 246.270 47.375 ;
        RECT 246.795 47.265 250.305 48.355 ;
        RECT 244.485 46.795 245.790 46.965 ;
        RECT 242.305 46.625 242.495 46.795 ;
        RECT 245.960 46.625 246.270 47.135 ;
        RECT 230.730 45.805 230.980 46.305 ;
        RECT 231.310 46.025 231.480 46.375 ;
        RECT 231.680 45.805 232.010 46.205 ;
        RECT 232.180 46.025 232.350 46.375 ;
        RECT 232.570 45.805 232.950 46.205 ;
        RECT 233.130 45.975 233.380 46.445 ;
        RECT 233.550 45.805 233.720 46.275 ;
        RECT 233.890 45.975 234.220 46.445 ;
        RECT 234.390 45.805 234.560 46.275 ;
        RECT 234.835 45.805 238.345 46.575 ;
        RECT 238.975 45.805 239.265 46.530 ;
        RECT 239.525 45.805 239.695 46.615 ;
        RECT 239.865 46.195 240.115 46.625 ;
        RECT 240.285 46.455 241.875 46.625 ;
        RECT 240.285 46.365 240.620 46.455 ;
        RECT 239.865 45.975 241.035 46.195 ;
        RECT 241.205 45.805 241.375 46.275 ;
        RECT 241.545 45.975 241.875 46.455 ;
        RECT 242.305 46.445 244.075 46.625 ;
        RECT 242.045 45.805 242.735 46.275 ;
        RECT 242.905 45.975 243.235 46.445 ;
        RECT 243.405 45.805 243.575 46.275 ;
        RECT 243.745 45.975 244.075 46.445 ;
        RECT 244.245 45.805 244.415 46.615 ;
        RECT 244.585 46.445 246.270 46.625 ;
        RECT 246.795 46.575 248.445 47.095 ;
        RECT 248.615 46.745 250.305 47.265 ;
        RECT 250.505 47.385 250.840 48.170 ;
        RECT 251.270 47.675 251.620 48.095 ;
        RECT 251.225 47.505 251.620 47.675 ;
        RECT 250.505 47.215 251.100 47.385 ;
        RECT 244.585 45.995 244.915 46.445 ;
        RECT 245.085 45.805 245.255 46.275 ;
        RECT 245.425 45.995 245.755 46.445 ;
        RECT 245.925 45.805 246.095 46.275 ;
        RECT 246.795 45.805 250.305 46.575 ;
        RECT 250.475 46.475 250.760 47.045 ;
        RECT 250.930 46.545 251.100 47.215 ;
        RECT 251.270 47.340 251.620 47.505 ;
        RECT 251.790 47.505 252.110 48.095 ;
        RECT 252.395 47.515 252.645 48.355 ;
        RECT 252.870 48.015 253.120 48.185 ;
        RECT 252.835 47.845 253.120 48.015 ;
        RECT 251.270 46.715 251.440 47.340 ;
        RECT 251.790 47.170 252.000 47.505 ;
        RECT 252.870 47.345 253.120 47.845 ;
        RECT 253.290 47.515 253.540 48.355 ;
        RECT 253.710 47.345 253.960 48.185 ;
        RECT 254.130 47.515 254.380 48.355 ;
        RECT 251.670 46.715 252.000 47.170 ;
        RECT 252.230 47.165 252.665 47.335 ;
        RECT 252.870 47.175 254.445 47.345 ;
        RECT 254.615 47.265 258.125 48.355 ;
        RECT 252.230 46.715 252.400 47.165 ;
        RECT 252.570 46.795 254.030 46.965 ;
        RECT 252.570 46.545 252.740 46.795 ;
        RECT 254.200 46.625 254.445 47.175 ;
        RECT 250.930 46.375 252.740 46.545 ;
        RECT 252.910 46.445 254.445 46.625 ;
        RECT 254.615 46.575 256.265 47.095 ;
        RECT 256.435 46.745 258.125 47.265 ;
        RECT 258.365 47.385 258.725 48.185 ;
        RECT 259.270 47.555 259.440 48.355 ;
        RECT 259.650 47.725 259.980 48.185 ;
        RECT 260.150 47.895 260.320 48.355 ;
        RECT 260.490 47.725 260.820 48.185 ;
        RECT 259.650 47.555 260.820 47.725 ;
        RECT 260.990 47.555 261.160 48.355 ;
        RECT 260.490 47.385 260.820 47.555 ;
        RECT 258.365 47.215 259.825 47.385 ;
        RECT 260.490 47.215 261.345 47.385 ;
        RECT 261.515 47.265 266.860 48.355 ;
        RECT 250.510 45.805 250.760 46.305 ;
        RECT 251.090 46.025 251.260 46.375 ;
        RECT 251.460 45.805 251.790 46.205 ;
        RECT 251.960 46.025 252.130 46.375 ;
        RECT 252.350 45.805 252.730 46.205 ;
        RECT 252.910 45.975 253.160 46.445 ;
        RECT 253.330 45.805 253.500 46.275 ;
        RECT 253.670 45.975 254.000 46.445 ;
        RECT 254.170 45.805 254.340 46.275 ;
        RECT 254.615 45.805 258.125 46.575 ;
        RECT 258.300 46.485 258.555 47.045 ;
        RECT 258.725 46.545 258.905 47.215 ;
        RECT 259.075 46.715 259.450 47.045 ;
        RECT 259.620 46.965 259.825 47.215 ;
        RECT 259.620 46.795 260.830 46.965 ;
        RECT 261.000 46.625 261.345 47.215 ;
        RECT 258.315 45.805 258.555 46.315 ;
        RECT 258.725 46.010 259.055 46.545 ;
        RECT 259.270 45.805 259.440 46.545 ;
        RECT 259.650 46.455 261.345 46.625 ;
        RECT 261.515 46.575 264.095 47.095 ;
        RECT 264.265 46.745 266.860 47.265 ;
        RECT 267.035 47.190 267.325 48.355 ;
        RECT 267.585 47.425 267.755 48.185 ;
        RECT 267.970 47.595 268.300 48.355 ;
        RECT 267.585 47.255 268.300 47.425 ;
        RECT 268.470 47.280 268.725 48.185 ;
        RECT 267.495 46.705 267.850 47.075 ;
        RECT 268.130 47.045 268.300 47.255 ;
        RECT 268.130 46.715 268.385 47.045 ;
        RECT 259.650 45.985 259.980 46.455 ;
        RECT 260.150 45.805 260.320 46.285 ;
        RECT 260.490 45.985 260.820 46.455 ;
        RECT 260.990 45.805 261.160 46.285 ;
        RECT 261.515 45.805 266.860 46.575 ;
        RECT 267.035 45.805 267.325 46.530 ;
        RECT 268.130 46.525 268.300 46.715 ;
        RECT 268.555 46.550 268.725 47.280 ;
        RECT 268.900 47.205 269.160 48.355 ;
        RECT 269.335 47.265 272.845 48.355 ;
        RECT 267.585 46.355 268.300 46.525 ;
        RECT 267.585 45.975 267.755 46.355 ;
        RECT 267.970 45.805 268.300 46.185 ;
        RECT 268.470 45.975 268.725 46.550 ;
        RECT 268.900 45.805 269.160 46.645 ;
        RECT 269.335 46.575 270.985 47.095 ;
        RECT 271.155 46.745 272.845 47.265 ;
        RECT 273.020 47.385 273.295 48.185 ;
        RECT 273.465 47.555 273.795 48.355 ;
        RECT 273.965 47.385 274.135 48.185 ;
        RECT 274.305 47.555 274.555 48.355 ;
        RECT 274.725 48.015 276.820 48.185 ;
        RECT 274.725 47.385 275.055 48.015 ;
        RECT 273.020 47.175 275.055 47.385 ;
        RECT 275.225 47.465 275.395 47.845 ;
        RECT 275.565 47.655 275.895 48.015 ;
        RECT 276.065 47.465 276.235 47.845 ;
        RECT 276.405 47.635 276.820 48.015 ;
        RECT 275.225 47.165 276.985 47.465 ;
        RECT 277.155 47.265 282.500 48.355 ;
        RECT 282.675 47.265 283.885 48.355 ;
        RECT 273.070 46.795 274.730 46.995 ;
        RECT 275.050 46.795 276.415 46.995 ;
        RECT 276.585 46.625 276.985 47.165 ;
        RECT 269.335 45.805 272.845 46.575 ;
        RECT 273.020 45.805 273.295 46.625 ;
        RECT 273.465 46.445 276.985 46.625 ;
        RECT 277.155 46.575 279.735 47.095 ;
        RECT 279.905 46.745 282.500 47.265 ;
        RECT 273.465 45.975 273.795 46.445 ;
        RECT 273.965 45.805 274.135 46.275 ;
        RECT 274.305 45.975 274.635 46.445 ;
        RECT 274.805 45.805 274.975 46.275 ;
        RECT 275.145 45.975 275.475 46.445 ;
        RECT 275.645 45.805 275.815 46.275 ;
        RECT 275.985 45.975 276.315 46.445 ;
        RECT 276.485 45.805 276.770 46.275 ;
        RECT 277.155 45.805 282.500 46.575 ;
        RECT 282.675 46.555 283.195 47.095 ;
        RECT 283.365 46.725 283.885 47.265 ;
        RECT 282.675 45.805 283.885 46.555 ;
        RECT 284.055 45.975 284.805 48.185 ;
        RECT 285.110 47.545 285.360 48.355 ;
        RECT 285.530 47.335 285.780 48.185 ;
        RECT 285.950 47.515 286.200 48.355 ;
        RECT 286.370 47.335 286.620 48.185 ;
        RECT 286.790 47.845 287.560 48.355 ;
        RECT 287.730 48.015 288.820 48.185 ;
        RECT 287.730 47.845 287.980 48.015 ;
        RECT 288.570 47.845 288.820 48.015 ;
        RECT 288.990 47.845 289.320 48.355 ;
        RECT 289.490 48.015 290.580 48.185 ;
        RECT 289.490 47.845 289.740 48.015 ;
        RECT 288.150 47.675 288.400 47.845 ;
        RECT 289.910 47.675 290.160 47.845 ;
        RECT 284.975 47.165 286.620 47.335 ;
        RECT 286.790 47.505 290.160 47.675 ;
        RECT 290.330 47.505 290.580 48.015 ;
        RECT 284.975 46.625 285.260 47.165 ;
        RECT 286.790 46.995 287.120 47.505 ;
        RECT 285.430 46.795 287.120 46.995 ;
        RECT 287.310 47.165 289.070 47.335 ;
        RECT 287.310 46.795 287.845 47.165 ;
        RECT 288.015 46.795 288.570 46.995 ;
        RECT 288.740 46.795 289.070 47.165 ;
        RECT 289.240 47.165 290.625 47.335 ;
        RECT 290.795 47.175 291.000 48.355 ;
        RECT 291.415 47.265 294.925 48.355 ;
        RECT 289.240 46.795 289.570 47.165 ;
        RECT 290.455 46.995 290.625 47.165 ;
        RECT 289.790 46.795 290.285 46.995 ;
        RECT 290.455 46.795 291.245 46.995 ;
        RECT 286.830 46.625 287.120 46.795 ;
        RECT 284.975 46.445 286.660 46.625 ;
        RECT 286.830 46.455 288.860 46.625 ;
        RECT 285.150 45.805 285.320 46.275 ;
        RECT 285.490 45.985 285.820 46.445 ;
        RECT 285.990 45.805 286.160 46.275 ;
        RECT 286.330 45.975 286.660 46.445 ;
        RECT 287.305 46.365 288.860 46.455 ;
        RECT 289.030 46.455 291.040 46.625 ;
        RECT 286.830 45.805 287.000 46.275 ;
        RECT 289.030 46.195 289.360 46.455 ;
        RECT 289.870 46.445 291.040 46.455 ;
        RECT 287.270 45.975 289.360 46.195 ;
        RECT 289.530 45.805 289.700 46.275 ;
        RECT 289.870 45.975 290.200 46.445 ;
        RECT 290.370 45.805 290.540 46.275 ;
        RECT 290.710 45.975 291.040 46.445 ;
        RECT 291.415 46.575 293.065 47.095 ;
        RECT 293.235 46.745 294.925 47.265 ;
        RECT 295.095 47.190 295.385 48.355 ;
        RECT 295.560 47.385 295.835 48.185 ;
        RECT 296.005 47.555 296.335 48.355 ;
        RECT 296.505 47.385 296.675 48.185 ;
        RECT 296.845 47.555 297.095 48.355 ;
        RECT 297.265 48.015 299.360 48.185 ;
        RECT 297.265 47.385 297.595 48.015 ;
        RECT 295.560 47.175 297.595 47.385 ;
        RECT 297.765 47.465 297.935 47.845 ;
        RECT 298.105 47.655 298.435 48.015 ;
        RECT 298.605 47.465 298.775 47.845 ;
        RECT 298.945 47.635 299.360 48.015 ;
        RECT 297.765 47.165 299.525 47.465 ;
        RECT 299.695 47.265 303.205 48.355 ;
        RECT 297.590 46.795 298.955 46.995 ;
        RECT 299.125 46.625 299.525 47.165 ;
        RECT 291.415 45.805 294.925 46.575 ;
        RECT 295.095 45.805 295.385 46.530 ;
        RECT 295.560 45.805 295.835 46.625 ;
        RECT 296.005 46.445 299.525 46.625 ;
        RECT 299.695 46.575 301.345 47.095 ;
        RECT 301.515 46.745 303.205 47.265 ;
        RECT 303.380 47.385 303.655 48.185 ;
        RECT 303.825 47.555 304.155 48.355 ;
        RECT 304.325 47.385 304.495 48.185 ;
        RECT 304.665 47.555 304.915 48.355 ;
        RECT 305.085 48.015 307.180 48.185 ;
        RECT 305.085 47.385 305.415 48.015 ;
        RECT 303.380 47.175 305.415 47.385 ;
        RECT 305.585 47.465 305.755 47.845 ;
        RECT 305.925 47.655 306.255 48.015 ;
        RECT 306.425 47.465 306.595 47.845 ;
        RECT 306.765 47.635 307.180 48.015 ;
        RECT 305.585 47.165 307.345 47.465 ;
        RECT 307.515 47.265 311.025 48.355 ;
        RECT 303.430 46.795 305.090 46.995 ;
        RECT 305.410 46.795 306.775 46.995 ;
        RECT 306.945 46.625 307.345 47.165 ;
        RECT 296.005 45.975 296.335 46.445 ;
        RECT 296.505 45.805 296.675 46.275 ;
        RECT 296.845 45.975 297.175 46.445 ;
        RECT 297.345 45.805 297.515 46.275 ;
        RECT 297.685 45.975 298.015 46.445 ;
        RECT 298.185 45.805 298.355 46.275 ;
        RECT 298.525 45.975 298.855 46.445 ;
        RECT 299.025 45.805 299.310 46.275 ;
        RECT 299.695 45.805 303.205 46.575 ;
        RECT 303.380 45.805 303.655 46.625 ;
        RECT 303.825 46.445 307.345 46.625 ;
        RECT 307.515 46.575 309.165 47.095 ;
        RECT 309.335 46.745 311.025 47.265 ;
        RECT 311.200 47.385 311.475 48.185 ;
        RECT 311.645 47.555 311.975 48.355 ;
        RECT 312.145 47.385 312.315 48.185 ;
        RECT 312.485 47.555 312.735 48.355 ;
        RECT 312.905 48.015 315.000 48.185 ;
        RECT 312.905 47.385 313.235 48.015 ;
        RECT 311.200 47.175 313.235 47.385 ;
        RECT 313.405 47.465 313.575 47.845 ;
        RECT 313.745 47.655 314.075 48.015 ;
        RECT 314.245 47.465 314.415 47.845 ;
        RECT 314.585 47.635 315.000 48.015 ;
        RECT 313.405 47.165 315.165 47.465 ;
        RECT 315.335 47.265 320.680 48.355 ;
        RECT 320.855 47.265 322.525 48.355 ;
        RECT 311.250 46.795 312.910 46.995 ;
        RECT 313.230 46.795 314.595 46.995 ;
        RECT 314.765 46.625 315.165 47.165 ;
        RECT 303.825 45.975 304.155 46.445 ;
        RECT 304.325 45.805 304.495 46.275 ;
        RECT 304.665 45.975 304.995 46.445 ;
        RECT 305.165 45.805 305.335 46.275 ;
        RECT 305.505 45.975 305.835 46.445 ;
        RECT 306.005 45.805 306.175 46.275 ;
        RECT 306.345 45.975 306.675 46.445 ;
        RECT 306.845 45.805 307.130 46.275 ;
        RECT 307.515 45.805 311.025 46.575 ;
        RECT 311.200 45.805 311.475 46.625 ;
        RECT 311.645 46.445 315.165 46.625 ;
        RECT 315.335 46.575 317.915 47.095 ;
        RECT 318.085 46.745 320.680 47.265 ;
        RECT 320.855 46.575 321.605 47.095 ;
        RECT 321.775 46.745 322.525 47.265 ;
        RECT 323.155 47.190 323.445 48.355 ;
        RECT 323.620 47.385 323.895 48.185 ;
        RECT 324.065 47.555 324.395 48.355 ;
        RECT 324.565 47.385 324.735 48.185 ;
        RECT 324.905 47.555 325.155 48.355 ;
        RECT 325.325 48.015 327.420 48.185 ;
        RECT 325.325 47.385 325.655 48.015 ;
        RECT 323.620 47.175 325.655 47.385 ;
        RECT 325.825 47.465 325.995 47.845 ;
        RECT 326.165 47.655 326.495 48.015 ;
        RECT 326.665 47.465 326.835 47.845 ;
        RECT 327.005 47.635 327.420 48.015 ;
        RECT 325.825 47.165 327.585 47.465 ;
        RECT 327.755 47.265 331.265 48.355 ;
        RECT 323.670 46.795 325.330 46.995 ;
        RECT 325.650 46.795 327.015 46.995 ;
        RECT 327.185 46.625 327.585 47.165 ;
        RECT 311.645 45.975 311.975 46.445 ;
        RECT 312.145 45.805 312.315 46.275 ;
        RECT 312.485 45.975 312.815 46.445 ;
        RECT 312.985 45.805 313.155 46.275 ;
        RECT 313.325 45.975 313.655 46.445 ;
        RECT 313.825 45.805 313.995 46.275 ;
        RECT 314.165 45.975 314.495 46.445 ;
        RECT 314.665 45.805 314.950 46.275 ;
        RECT 315.335 45.805 320.680 46.575 ;
        RECT 320.855 45.805 322.525 46.575 ;
        RECT 323.155 45.805 323.445 46.530 ;
        RECT 323.620 45.805 323.895 46.625 ;
        RECT 324.065 46.445 327.585 46.625 ;
        RECT 327.755 46.575 329.405 47.095 ;
        RECT 329.575 46.745 331.265 47.265 ;
        RECT 331.440 47.385 331.715 48.185 ;
        RECT 331.885 47.555 332.215 48.355 ;
        RECT 332.385 47.385 332.555 48.185 ;
        RECT 332.725 47.555 332.975 48.355 ;
        RECT 333.145 48.015 335.240 48.185 ;
        RECT 333.145 47.385 333.475 48.015 ;
        RECT 331.440 47.175 333.475 47.385 ;
        RECT 333.645 47.465 333.815 47.845 ;
        RECT 333.985 47.655 334.315 48.015 ;
        RECT 334.485 47.465 334.655 47.845 ;
        RECT 334.825 47.635 335.240 48.015 ;
        RECT 333.645 47.165 335.405 47.465 ;
        RECT 335.575 47.265 339.085 48.355 ;
        RECT 331.490 46.795 333.150 46.995 ;
        RECT 333.470 46.795 334.835 46.995 ;
        RECT 335.005 46.625 335.405 47.165 ;
        RECT 324.065 45.975 324.395 46.445 ;
        RECT 324.565 45.805 324.735 46.275 ;
        RECT 324.905 45.975 325.235 46.445 ;
        RECT 325.405 45.805 325.575 46.275 ;
        RECT 325.745 45.975 326.075 46.445 ;
        RECT 326.245 45.805 326.415 46.275 ;
        RECT 326.585 45.975 326.915 46.445 ;
        RECT 327.085 45.805 327.370 46.275 ;
        RECT 327.755 45.805 331.265 46.575 ;
        RECT 331.440 45.805 331.715 46.625 ;
        RECT 331.885 46.445 335.405 46.625 ;
        RECT 335.575 46.575 337.225 47.095 ;
        RECT 337.395 46.745 339.085 47.265 ;
        RECT 339.260 47.385 339.535 48.185 ;
        RECT 339.705 47.555 340.035 48.355 ;
        RECT 340.205 47.385 340.375 48.185 ;
        RECT 340.545 47.555 340.795 48.355 ;
        RECT 340.965 48.015 343.060 48.185 ;
        RECT 340.965 47.385 341.295 48.015 ;
        RECT 339.260 47.175 341.295 47.385 ;
        RECT 341.465 47.465 341.635 47.845 ;
        RECT 341.805 47.655 342.135 48.015 ;
        RECT 342.305 47.465 342.475 47.845 ;
        RECT 342.645 47.635 343.060 48.015 ;
        RECT 341.465 47.165 343.225 47.465 ;
        RECT 343.395 47.265 348.740 48.355 ;
        RECT 348.915 47.265 350.585 48.355 ;
        RECT 339.310 46.795 340.970 46.995 ;
        RECT 341.290 46.795 342.655 46.995 ;
        RECT 342.825 46.625 343.225 47.165 ;
        RECT 331.885 45.975 332.215 46.445 ;
        RECT 332.385 45.805 332.555 46.275 ;
        RECT 332.725 45.975 333.055 46.445 ;
        RECT 333.225 45.805 333.395 46.275 ;
        RECT 333.565 45.975 333.895 46.445 ;
        RECT 334.065 45.805 334.235 46.275 ;
        RECT 334.405 45.975 334.735 46.445 ;
        RECT 334.905 45.805 335.190 46.275 ;
        RECT 335.575 45.805 339.085 46.575 ;
        RECT 339.260 45.805 339.535 46.625 ;
        RECT 339.705 46.445 343.225 46.625 ;
        RECT 343.395 46.575 345.975 47.095 ;
        RECT 346.145 46.745 348.740 47.265 ;
        RECT 348.915 46.575 349.665 47.095 ;
        RECT 349.835 46.745 350.585 47.265 ;
        RECT 351.215 47.190 351.505 48.355 ;
        RECT 351.680 47.385 351.955 48.185 ;
        RECT 352.125 47.555 352.455 48.355 ;
        RECT 352.625 47.385 352.795 48.185 ;
        RECT 352.965 47.555 353.215 48.355 ;
        RECT 353.385 48.015 355.480 48.185 ;
        RECT 353.385 47.385 353.715 48.015 ;
        RECT 351.680 47.175 353.715 47.385 ;
        RECT 353.885 47.465 354.055 47.845 ;
        RECT 354.225 47.655 354.555 48.015 ;
        RECT 354.725 47.465 354.895 47.845 ;
        RECT 355.065 47.635 355.480 48.015 ;
        RECT 353.885 47.165 355.645 47.465 ;
        RECT 355.815 47.265 359.325 48.355 ;
        RECT 351.730 46.795 353.390 46.995 ;
        RECT 353.710 46.795 355.075 46.995 ;
        RECT 355.245 46.625 355.645 47.165 ;
        RECT 339.705 45.975 340.035 46.445 ;
        RECT 340.205 45.805 340.375 46.275 ;
        RECT 340.545 45.975 340.875 46.445 ;
        RECT 341.045 45.805 341.215 46.275 ;
        RECT 341.385 45.975 341.715 46.445 ;
        RECT 341.885 45.805 342.055 46.275 ;
        RECT 342.225 45.975 342.555 46.445 ;
        RECT 342.725 45.805 343.010 46.275 ;
        RECT 343.395 45.805 348.740 46.575 ;
        RECT 348.915 45.805 350.585 46.575 ;
        RECT 351.215 45.805 351.505 46.530 ;
        RECT 351.680 45.805 351.955 46.625 ;
        RECT 352.125 46.445 355.645 46.625 ;
        RECT 355.815 46.575 357.465 47.095 ;
        RECT 357.635 46.745 359.325 47.265 ;
        RECT 359.500 47.385 359.775 48.185 ;
        RECT 359.945 47.555 360.275 48.355 ;
        RECT 360.445 47.385 360.615 48.185 ;
        RECT 360.785 47.555 361.035 48.355 ;
        RECT 361.205 48.015 363.300 48.185 ;
        RECT 361.205 47.385 361.535 48.015 ;
        RECT 359.500 47.175 361.535 47.385 ;
        RECT 361.705 47.465 361.875 47.845 ;
        RECT 362.045 47.655 362.375 48.015 ;
        RECT 362.545 47.465 362.715 47.845 ;
        RECT 362.885 47.635 363.300 48.015 ;
        RECT 361.705 47.165 363.465 47.465 ;
        RECT 363.635 47.265 367.145 48.355 ;
        RECT 359.550 46.795 361.210 46.995 ;
        RECT 361.530 46.795 362.895 46.995 ;
        RECT 363.065 46.625 363.465 47.165 ;
        RECT 352.125 45.975 352.455 46.445 ;
        RECT 352.625 45.805 352.795 46.275 ;
        RECT 352.965 45.975 353.295 46.445 ;
        RECT 353.465 45.805 353.635 46.275 ;
        RECT 353.805 45.975 354.135 46.445 ;
        RECT 354.305 45.805 354.475 46.275 ;
        RECT 354.645 45.975 354.975 46.445 ;
        RECT 355.145 45.805 355.430 46.275 ;
        RECT 355.815 45.805 359.325 46.575 ;
        RECT 359.500 45.805 359.775 46.625 ;
        RECT 359.945 46.445 363.465 46.625 ;
        RECT 363.635 46.575 365.285 47.095 ;
        RECT 365.455 46.745 367.145 47.265 ;
        RECT 367.320 47.385 367.595 48.185 ;
        RECT 367.765 47.555 368.095 48.355 ;
        RECT 368.265 47.385 368.435 48.185 ;
        RECT 368.605 47.555 368.855 48.355 ;
        RECT 369.025 48.015 371.120 48.185 ;
        RECT 369.025 47.385 369.355 48.015 ;
        RECT 367.320 47.175 369.355 47.385 ;
        RECT 369.525 47.465 369.695 47.845 ;
        RECT 369.865 47.655 370.195 48.015 ;
        RECT 370.365 47.465 370.535 47.845 ;
        RECT 370.705 47.635 371.120 48.015 ;
        RECT 369.525 47.165 371.285 47.465 ;
        RECT 371.455 47.265 376.800 48.355 ;
        RECT 376.975 47.265 378.645 48.355 ;
        RECT 367.370 46.795 369.030 46.995 ;
        RECT 369.350 46.795 370.715 46.995 ;
        RECT 370.885 46.625 371.285 47.165 ;
        RECT 359.945 45.975 360.275 46.445 ;
        RECT 360.445 45.805 360.615 46.275 ;
        RECT 360.785 45.975 361.115 46.445 ;
        RECT 361.285 45.805 361.455 46.275 ;
        RECT 361.625 45.975 361.955 46.445 ;
        RECT 362.125 45.805 362.295 46.275 ;
        RECT 362.465 45.975 362.795 46.445 ;
        RECT 362.965 45.805 363.250 46.275 ;
        RECT 363.635 45.805 367.145 46.575 ;
        RECT 367.320 45.805 367.595 46.625 ;
        RECT 367.765 46.445 371.285 46.625 ;
        RECT 371.455 46.575 374.035 47.095 ;
        RECT 374.205 46.745 376.800 47.265 ;
        RECT 376.975 46.575 377.725 47.095 ;
        RECT 377.895 46.745 378.645 47.265 ;
        RECT 379.275 47.190 379.565 48.355 ;
        RECT 379.925 47.630 380.255 48.355 ;
        RECT 367.765 45.975 368.095 46.445 ;
        RECT 368.265 45.805 368.435 46.275 ;
        RECT 368.605 45.975 368.935 46.445 ;
        RECT 369.105 45.805 369.275 46.275 ;
        RECT 369.445 45.975 369.775 46.445 ;
        RECT 369.945 45.805 370.115 46.275 ;
        RECT 370.285 45.975 370.615 46.445 ;
        RECT 370.785 45.805 371.070 46.275 ;
        RECT 371.455 45.805 376.800 46.575 ;
        RECT 376.975 45.805 378.645 46.575 ;
        RECT 379.275 45.805 379.565 46.530 ;
        RECT 379.735 45.975 380.255 47.460 ;
        RECT 381.115 47.265 384.625 48.355 ;
        RECT 384.985 47.630 385.315 48.355 ;
        RECT 381.115 46.575 382.765 47.095 ;
        RECT 382.935 46.745 384.625 47.265 ;
        RECT 380.425 45.805 380.765 46.465 ;
        RECT 381.115 45.805 384.625 46.575 ;
        RECT 384.795 45.975 385.315 47.460 ;
        RECT 385.485 46.635 386.005 48.185 ;
        RECT 386.175 47.265 389.685 48.355 ;
        RECT 390.045 47.630 390.375 48.355 ;
        RECT 386.175 46.575 387.825 47.095 ;
        RECT 387.995 46.745 389.685 47.265 ;
        RECT 385.485 45.805 385.825 46.465 ;
        RECT 386.175 45.805 389.685 46.575 ;
        RECT 389.855 45.975 390.375 47.460 ;
        RECT 390.545 46.635 391.065 48.185 ;
        RECT 391.235 47.265 394.745 48.355 ;
        RECT 395.105 47.630 395.435 48.355 ;
        RECT 391.235 46.575 392.885 47.095 ;
        RECT 393.055 46.745 394.745 47.265 ;
        RECT 390.545 45.805 390.885 46.465 ;
        RECT 391.235 45.805 394.745 46.575 ;
        RECT 394.915 45.975 395.435 47.460 ;
        RECT 396.295 47.265 399.805 48.355 ;
        RECT 400.165 47.630 400.495 48.355 ;
        RECT 396.295 46.575 397.945 47.095 ;
        RECT 398.115 46.745 399.805 47.265 ;
        RECT 395.605 45.805 395.945 46.465 ;
        RECT 396.295 45.805 399.805 46.575 ;
        RECT 399.975 45.975 400.495 47.460 ;
        RECT 400.665 46.635 401.185 48.185 ;
        RECT 401.355 47.265 406.700 48.355 ;
        RECT 401.355 46.575 403.935 47.095 ;
        RECT 404.105 46.745 406.700 47.265 ;
        RECT 407.335 47.190 407.625 48.355 ;
        RECT 407.985 47.630 408.315 48.355 ;
        RECT 400.665 45.805 401.005 46.465 ;
        RECT 401.355 45.805 406.700 46.575 ;
        RECT 407.335 45.805 407.625 46.530 ;
        RECT 407.795 45.975 408.315 47.460 ;
        RECT 408.485 46.635 409.005 48.185 ;
        RECT 409.175 47.265 412.685 48.355 ;
        RECT 413.045 47.630 413.375 48.355 ;
        RECT 409.175 46.575 410.825 47.095 ;
        RECT 410.995 46.745 412.685 47.265 ;
        RECT 408.485 45.805 408.825 46.465 ;
        RECT 409.175 45.805 412.685 46.575 ;
        RECT 412.855 45.975 413.375 47.460 ;
        RECT 413.545 46.635 414.065 48.185 ;
        RECT 414.235 47.265 417.745 48.355 ;
        RECT 418.105 47.630 418.435 48.355 ;
        RECT 414.235 46.575 415.885 47.095 ;
        RECT 416.055 46.745 417.745 47.265 ;
        RECT 413.545 45.805 413.885 46.465 ;
        RECT 414.235 45.805 417.745 46.575 ;
        RECT 417.915 45.975 418.435 47.460 ;
        RECT 418.605 46.635 419.125 48.185 ;
        RECT 419.295 47.265 422.805 48.355 ;
        RECT 423.165 47.630 423.495 48.355 ;
        RECT 419.295 46.575 420.945 47.095 ;
        RECT 421.115 46.745 422.805 47.265 ;
        RECT 418.605 45.805 418.945 46.465 ;
        RECT 419.295 45.805 422.805 46.575 ;
        RECT 422.975 45.975 423.495 47.460 ;
        RECT 423.665 46.635 424.185 48.185 ;
        RECT 424.355 47.265 427.865 48.355 ;
        RECT 428.225 47.630 428.555 48.355 ;
        RECT 424.355 46.575 426.005 47.095 ;
        RECT 426.175 46.745 427.865 47.265 ;
        RECT 423.665 45.805 424.005 46.465 ;
        RECT 424.355 45.805 427.865 46.575 ;
        RECT 428.035 45.975 428.555 47.460 ;
        RECT 428.725 46.635 429.245 48.185 ;
        RECT 429.415 47.265 434.760 48.355 ;
        RECT 429.415 46.575 431.995 47.095 ;
        RECT 432.165 46.745 434.760 47.265 ;
        RECT 435.395 47.190 435.685 48.355 ;
        RECT 436.045 47.630 436.375 48.355 ;
        RECT 428.725 45.805 429.065 46.465 ;
        RECT 429.415 45.805 434.760 46.575 ;
        RECT 435.395 45.805 435.685 46.530 ;
        RECT 435.855 45.975 436.375 47.460 ;
        RECT 437.235 47.265 440.745 48.355 ;
        RECT 441.105 47.630 441.435 48.355 ;
        RECT 437.235 46.575 438.885 47.095 ;
        RECT 439.055 46.745 440.745 47.265 ;
        RECT 436.545 45.805 436.885 46.465 ;
        RECT 437.235 45.805 440.745 46.575 ;
        RECT 440.915 45.975 441.435 47.460 ;
        RECT 441.605 46.635 442.125 48.185 ;
        RECT 442.295 47.265 445.805 48.355 ;
        RECT 446.165 47.630 446.495 48.355 ;
        RECT 442.295 46.575 443.945 47.095 ;
        RECT 444.115 46.745 445.805 47.265 ;
        RECT 441.605 45.805 441.945 46.465 ;
        RECT 442.295 45.805 445.805 46.575 ;
        RECT 445.975 45.975 446.495 47.460 ;
        RECT 446.665 46.635 447.185 48.185 ;
        RECT 447.355 47.265 450.865 48.355 ;
        RECT 451.225 47.630 451.555 48.355 ;
        RECT 447.355 46.575 449.005 47.095 ;
        RECT 449.175 46.745 450.865 47.265 ;
        RECT 446.665 45.805 447.005 46.465 ;
        RECT 447.355 45.805 450.865 46.575 ;
        RECT 451.035 45.975 451.555 47.460 ;
        RECT 451.725 46.635 452.245 48.185 ;
        RECT 452.415 47.265 455.925 48.355 ;
        RECT 456.285 47.630 456.615 48.355 ;
        RECT 452.415 46.575 454.065 47.095 ;
        RECT 454.235 46.745 455.925 47.265 ;
        RECT 451.725 45.805 452.065 46.465 ;
        RECT 452.415 45.805 455.925 46.575 ;
        RECT 456.095 45.975 456.615 47.460 ;
        RECT 456.785 46.635 457.305 48.185 ;
        RECT 457.475 47.265 462.820 48.355 ;
        RECT 457.475 46.575 460.055 47.095 ;
        RECT 460.225 46.745 462.820 47.265 ;
        RECT 463.455 47.190 463.745 48.355 ;
        RECT 464.105 47.630 464.435 48.355 ;
        RECT 456.785 45.805 457.125 46.465 ;
        RECT 457.475 45.805 462.820 46.575 ;
        RECT 463.455 45.805 463.745 46.530 ;
        RECT 463.915 45.975 464.435 47.460 ;
        RECT 465.295 47.265 468.805 48.355 ;
        RECT 469.165 47.630 469.495 48.355 ;
        RECT 465.295 46.575 466.945 47.095 ;
        RECT 467.115 46.745 468.805 47.265 ;
        RECT 464.605 45.805 464.945 46.465 ;
        RECT 465.295 45.805 468.805 46.575 ;
        RECT 468.975 45.975 469.495 47.460 ;
        RECT 469.665 46.635 470.185 48.185 ;
        RECT 470.355 47.265 473.865 48.355 ;
        RECT 474.225 47.630 474.555 48.355 ;
        RECT 470.355 46.575 472.005 47.095 ;
        RECT 472.175 46.745 473.865 47.265 ;
        RECT 469.665 45.805 470.005 46.465 ;
        RECT 470.355 45.805 473.865 46.575 ;
        RECT 474.035 45.975 474.555 47.460 ;
        RECT 474.725 46.635 475.245 48.185 ;
        RECT 475.415 47.265 478.925 48.355 ;
        RECT 479.285 47.630 479.615 48.355 ;
        RECT 475.415 46.575 477.065 47.095 ;
        RECT 477.235 46.745 478.925 47.265 ;
        RECT 474.725 45.805 475.065 46.465 ;
        RECT 475.415 45.805 478.925 46.575 ;
        RECT 479.095 45.975 479.615 47.460 ;
        RECT 479.785 46.635 480.305 48.185 ;
        RECT 480.475 47.265 483.985 48.355 ;
        RECT 484.345 47.630 484.675 48.355 ;
        RECT 480.475 46.575 482.125 47.095 ;
        RECT 482.295 46.745 483.985 47.265 ;
        RECT 479.785 45.805 480.125 46.465 ;
        RECT 480.475 45.805 483.985 46.575 ;
        RECT 484.155 45.975 484.675 47.460 ;
        RECT 484.845 46.635 485.365 48.185 ;
        RECT 485.535 47.265 490.880 48.355 ;
        RECT 485.535 46.575 488.115 47.095 ;
        RECT 488.285 46.745 490.880 47.265 ;
        RECT 491.515 47.190 491.805 48.355 ;
        RECT 492.165 47.630 492.495 48.355 ;
        RECT 484.845 45.805 485.185 46.465 ;
        RECT 485.535 45.805 490.880 46.575 ;
        RECT 491.515 45.805 491.805 46.530 ;
        RECT 491.975 45.975 492.495 47.460 ;
        RECT 492.665 46.635 493.185 48.185 ;
        RECT 493.355 47.265 496.865 48.355 ;
        RECT 497.225 47.630 497.555 48.355 ;
        RECT 493.355 46.575 495.005 47.095 ;
        RECT 495.175 46.745 496.865 47.265 ;
        RECT 492.665 45.805 493.005 46.465 ;
        RECT 493.355 45.805 496.865 46.575 ;
        RECT 497.035 45.975 497.555 47.460 ;
        RECT 497.725 46.635 498.245 48.185 ;
        RECT 498.415 47.265 501.925 48.355 ;
        RECT 502.285 47.630 502.615 48.355 ;
        RECT 498.415 46.575 500.065 47.095 ;
        RECT 500.235 46.745 501.925 47.265 ;
        RECT 497.725 45.805 498.065 46.465 ;
        RECT 498.415 45.805 501.925 46.575 ;
        RECT 502.095 45.975 502.615 47.460 ;
        RECT 502.785 46.635 503.305 48.185 ;
        RECT 503.475 47.265 506.985 48.355 ;
        RECT 507.345 47.630 507.675 48.355 ;
        RECT 503.475 46.575 505.125 47.095 ;
        RECT 505.295 46.745 506.985 47.265 ;
        RECT 502.785 45.805 503.125 46.465 ;
        RECT 503.475 45.805 506.985 46.575 ;
        RECT 507.155 45.975 507.675 47.460 ;
        RECT 507.845 46.635 508.365 48.185 ;
        RECT 508.535 47.265 512.045 48.355 ;
        RECT 512.405 47.630 512.735 48.355 ;
        RECT 508.535 46.575 510.185 47.095 ;
        RECT 510.355 46.745 512.045 47.265 ;
        RECT 507.845 45.805 508.185 46.465 ;
        RECT 508.535 45.805 512.045 46.575 ;
        RECT 512.215 45.975 512.735 47.460 ;
        RECT 513.595 47.265 518.940 48.355 ;
        RECT 513.595 46.575 516.175 47.095 ;
        RECT 516.345 46.745 518.940 47.265 ;
        RECT 519.575 47.190 519.865 48.355 ;
        RECT 520.225 47.630 520.555 48.355 ;
        RECT 512.905 45.805 513.245 46.465 ;
        RECT 513.595 45.805 518.940 46.575 ;
        RECT 519.575 45.805 519.865 46.530 ;
        RECT 520.035 45.975 520.555 47.460 ;
        RECT 520.725 46.635 521.245 48.185 ;
        RECT 521.415 47.265 524.925 48.355 ;
        RECT 525.285 47.630 525.615 48.355 ;
        RECT 521.415 46.575 523.065 47.095 ;
        RECT 523.235 46.745 524.925 47.265 ;
        RECT 520.725 45.805 521.065 46.465 ;
        RECT 521.415 45.805 524.925 46.575 ;
        RECT 525.095 45.975 525.615 47.460 ;
        RECT 525.785 46.635 526.305 48.185 ;
        RECT 526.475 47.265 529.985 48.355 ;
        RECT 530.345 47.630 530.675 48.355 ;
        RECT 526.475 46.575 528.125 47.095 ;
        RECT 528.295 46.745 529.985 47.265 ;
        RECT 525.785 45.805 526.125 46.465 ;
        RECT 526.475 45.805 529.985 46.575 ;
        RECT 530.155 45.975 530.675 47.460 ;
        RECT 530.845 46.635 531.365 48.185 ;
        RECT 531.535 47.265 535.045 48.355 ;
        RECT 535.405 47.630 535.735 48.355 ;
        RECT 531.535 46.575 533.185 47.095 ;
        RECT 533.355 46.745 535.045 47.265 ;
        RECT 530.845 45.805 531.185 46.465 ;
        RECT 531.535 45.805 535.045 46.575 ;
        RECT 535.215 45.975 535.735 47.460 ;
        RECT 535.905 46.635 536.425 48.185 ;
        RECT 536.595 47.265 540.105 48.355 ;
        RECT 540.465 47.630 540.795 48.355 ;
        RECT 536.595 46.575 538.245 47.095 ;
        RECT 538.415 46.745 540.105 47.265 ;
        RECT 535.905 45.805 536.245 46.465 ;
        RECT 536.595 45.805 540.105 46.575 ;
        RECT 540.275 45.975 540.795 47.460 ;
        RECT 540.965 46.635 541.485 48.185 ;
        RECT 541.655 47.265 547.000 48.355 ;
        RECT 541.655 46.575 544.235 47.095 ;
        RECT 544.405 46.745 547.000 47.265 ;
        RECT 547.635 47.190 547.925 48.355 ;
        RECT 548.285 47.630 548.615 48.355 ;
        RECT 540.965 45.805 541.305 46.465 ;
        RECT 541.655 45.805 547.000 46.575 ;
        RECT 547.635 45.805 547.925 46.530 ;
        RECT 548.095 45.975 548.615 47.460 ;
        RECT 548.785 46.635 549.305 48.185 ;
        RECT 549.475 47.265 552.985 48.355 ;
        RECT 553.345 47.630 553.675 48.355 ;
        RECT 549.475 46.575 551.125 47.095 ;
        RECT 551.295 46.745 552.985 47.265 ;
        RECT 548.785 45.805 549.125 46.465 ;
        RECT 549.475 45.805 552.985 46.575 ;
        RECT 553.155 45.975 553.675 47.460 ;
        RECT 553.845 46.635 554.365 48.185 ;
        RECT 554.535 47.265 558.045 48.355 ;
        RECT 558.405 47.630 558.735 48.355 ;
        RECT 554.535 46.575 556.185 47.095 ;
        RECT 556.355 46.745 558.045 47.265 ;
        RECT 553.845 45.805 554.185 46.465 ;
        RECT 554.535 45.805 558.045 46.575 ;
        RECT 558.215 45.975 558.735 47.460 ;
        RECT 558.905 46.635 559.425 48.185 ;
        RECT 559.595 47.265 563.105 48.355 ;
        RECT 563.465 47.630 563.795 48.355 ;
        RECT 559.595 46.575 561.245 47.095 ;
        RECT 561.415 46.745 563.105 47.265 ;
        RECT 558.905 45.805 559.245 46.465 ;
        RECT 559.595 45.805 563.105 46.575 ;
        RECT 563.275 45.975 563.795 47.460 ;
        RECT 563.965 46.635 564.485 48.185 ;
        RECT 564.655 47.265 568.165 48.355 ;
        RECT 568.525 47.630 568.855 48.355 ;
        RECT 564.655 46.575 566.305 47.095 ;
        RECT 566.475 46.745 568.165 47.265 ;
        RECT 563.965 45.805 564.305 46.465 ;
        RECT 564.655 45.805 568.165 46.575 ;
        RECT 568.335 45.975 568.855 47.460 ;
        RECT 569.025 46.635 569.545 48.185 ;
        RECT 569.715 47.265 575.060 48.355 ;
        RECT 569.715 46.575 572.295 47.095 ;
        RECT 572.465 46.745 575.060 47.265 ;
        RECT 575.695 47.190 575.985 48.355 ;
        RECT 576.345 47.630 576.675 48.355 ;
        RECT 569.025 45.805 569.365 46.465 ;
        RECT 569.715 45.805 575.060 46.575 ;
        RECT 575.695 45.805 575.985 46.530 ;
        RECT 576.155 45.975 576.675 47.460 ;
        RECT 576.845 46.635 577.365 48.185 ;
        RECT 577.535 47.265 581.045 48.355 ;
        RECT 581.405 47.630 581.735 48.355 ;
        RECT 577.535 46.575 579.185 47.095 ;
        RECT 579.355 46.745 581.045 47.265 ;
        RECT 576.845 45.805 577.185 46.465 ;
        RECT 577.535 45.805 581.045 46.575 ;
        RECT 581.215 45.975 581.735 47.460 ;
        RECT 581.905 46.635 582.425 48.185 ;
        RECT 582.595 47.265 586.105 48.355 ;
        RECT 586.465 47.630 586.795 48.355 ;
        RECT 582.595 46.575 584.245 47.095 ;
        RECT 584.415 46.745 586.105 47.265 ;
        RECT 581.905 45.805 582.245 46.465 ;
        RECT 582.595 45.805 586.105 46.575 ;
        RECT 586.275 45.975 586.795 47.460 ;
        RECT 586.965 46.635 587.485 48.185 ;
        RECT 587.655 47.265 591.165 48.355 ;
        RECT 591.525 47.630 591.855 48.355 ;
        RECT 587.655 46.575 589.305 47.095 ;
        RECT 589.475 46.745 591.165 47.265 ;
        RECT 586.965 45.805 587.305 46.465 ;
        RECT 587.655 45.805 591.165 46.575 ;
        RECT 591.335 45.975 591.855 47.460 ;
        RECT 592.025 46.635 592.545 48.185 ;
        RECT 592.715 47.265 596.225 48.355 ;
        RECT 596.585 47.630 596.915 48.355 ;
        RECT 592.715 46.575 594.365 47.095 ;
        RECT 594.535 46.745 596.225 47.265 ;
        RECT 592.025 45.805 592.365 46.465 ;
        RECT 592.715 45.805 596.225 46.575 ;
        RECT 596.395 45.975 596.915 47.460 ;
        RECT 597.085 46.635 597.605 48.185 ;
        RECT 597.775 47.265 603.120 48.355 ;
        RECT 597.775 46.575 600.355 47.095 ;
        RECT 600.525 46.745 603.120 47.265 ;
        RECT 603.755 47.190 604.045 48.355 ;
        RECT 604.405 47.630 604.735 48.355 ;
        RECT 597.085 45.805 597.425 46.465 ;
        RECT 597.775 45.805 603.120 46.575 ;
        RECT 603.755 45.805 604.045 46.530 ;
        RECT 604.215 45.975 604.735 47.460 ;
        RECT 604.905 46.635 605.425 48.185 ;
        RECT 605.595 47.265 609.105 48.355 ;
        RECT 609.465 47.630 609.795 48.355 ;
        RECT 605.595 46.575 607.245 47.095 ;
        RECT 607.415 46.745 609.105 47.265 ;
        RECT 604.905 45.805 605.245 46.465 ;
        RECT 605.595 45.805 609.105 46.575 ;
        RECT 609.275 45.975 609.795 47.460 ;
        RECT 609.965 46.635 610.485 48.185 ;
        RECT 610.655 47.265 614.165 48.355 ;
        RECT 614.525 47.630 614.855 48.355 ;
        RECT 610.655 46.575 612.305 47.095 ;
        RECT 612.475 46.745 614.165 47.265 ;
        RECT 609.965 45.805 610.305 46.465 ;
        RECT 610.655 45.805 614.165 46.575 ;
        RECT 614.335 45.975 614.855 47.460 ;
        RECT 615.025 46.635 615.545 48.185 ;
        RECT 615.715 47.265 619.225 48.355 ;
        RECT 619.585 47.630 619.915 48.355 ;
        RECT 615.715 46.575 617.365 47.095 ;
        RECT 617.535 46.745 619.225 47.265 ;
        RECT 615.025 45.805 615.365 46.465 ;
        RECT 615.715 45.805 619.225 46.575 ;
        RECT 619.395 45.975 619.915 47.460 ;
        RECT 620.085 46.635 620.605 48.185 ;
        RECT 620.775 47.265 624.285 48.355 ;
        RECT 624.645 47.630 624.975 48.355 ;
        RECT 620.775 46.575 622.425 47.095 ;
        RECT 622.595 46.745 624.285 47.265 ;
        RECT 620.085 45.805 620.425 46.465 ;
        RECT 620.775 45.805 624.285 46.575 ;
        RECT 624.455 45.975 624.975 47.460 ;
        RECT 625.145 46.635 625.665 48.185 ;
        RECT 625.835 47.265 629.345 48.355 ;
        RECT 625.835 46.575 627.485 47.095 ;
        RECT 627.655 46.745 629.345 47.265 ;
        RECT 629.975 47.265 631.185 48.355 ;
        RECT 629.975 46.725 630.495 47.265 ;
        RECT 625.145 45.805 625.485 46.465 ;
        RECT 625.835 45.805 629.345 46.575 ;
        RECT 630.665 46.555 631.185 47.095 ;
        RECT 629.975 45.805 631.185 46.555 ;
        RECT 42.470 45.635 631.270 45.805 ;
        RECT 42.555 44.885 43.765 45.635 ;
        RECT 42.555 44.345 43.075 44.885 ;
        RECT 43.935 44.865 49.280 45.635 ;
        RECT 49.455 44.865 54.800 45.635 ;
        RECT 54.975 44.865 56.645 45.635 ;
        RECT 56.815 44.910 57.105 45.635 ;
        RECT 57.275 44.865 62.620 45.635 ;
        RECT 62.795 44.865 68.140 45.635 ;
        RECT 68.315 44.865 70.905 45.635 ;
        RECT 71.075 44.910 71.365 45.635 ;
        RECT 71.535 44.865 76.880 45.635 ;
        RECT 77.055 44.885 78.265 45.635 ;
        RECT 78.455 45.125 78.695 45.635 ;
        RECT 43.245 44.175 43.765 44.715 ;
        RECT 43.935 44.345 46.515 44.865 ;
        RECT 46.685 44.175 49.280 44.695 ;
        RECT 49.455 44.345 52.035 44.865 ;
        RECT 52.205 44.175 54.800 44.695 ;
        RECT 54.975 44.345 55.725 44.865 ;
        RECT 55.895 44.175 56.645 44.695 ;
        RECT 57.275 44.345 59.855 44.865 ;
        RECT 42.555 43.085 43.765 44.175 ;
        RECT 43.935 43.085 49.280 44.175 ;
        RECT 49.455 43.085 54.800 44.175 ;
        RECT 54.975 43.085 56.645 44.175 ;
        RECT 56.815 43.085 57.105 44.250 ;
        RECT 60.025 44.175 62.620 44.695 ;
        RECT 62.795 44.345 65.375 44.865 ;
        RECT 65.545 44.175 68.140 44.695 ;
        RECT 68.315 44.345 69.525 44.865 ;
        RECT 69.695 44.175 70.905 44.695 ;
        RECT 71.535 44.345 74.115 44.865 ;
        RECT 57.275 43.085 62.620 44.175 ;
        RECT 62.795 43.085 68.140 44.175 ;
        RECT 68.315 43.085 70.905 44.175 ;
        RECT 71.075 43.085 71.365 44.250 ;
        RECT 74.285 44.175 76.880 44.695 ;
        RECT 77.055 44.345 77.575 44.885 ;
        RECT 77.745 44.175 78.265 44.715 ;
        RECT 78.440 44.395 78.695 44.955 ;
        RECT 78.865 44.895 79.195 45.430 ;
        RECT 79.410 44.895 79.580 45.635 ;
        RECT 79.790 44.985 80.120 45.455 ;
        RECT 80.290 45.155 80.460 45.635 ;
        RECT 80.630 44.985 80.960 45.455 ;
        RECT 81.130 45.155 81.300 45.635 ;
        RECT 78.865 44.225 79.045 44.895 ;
        RECT 79.790 44.815 81.485 44.985 ;
        RECT 79.215 44.395 79.590 44.725 ;
        RECT 79.760 44.475 80.970 44.645 ;
        RECT 79.760 44.225 79.965 44.475 ;
        RECT 81.140 44.225 81.485 44.815 ;
        RECT 81.655 44.865 85.165 45.635 ;
        RECT 85.335 44.910 85.625 45.635 ;
        RECT 81.655 44.345 83.305 44.865 ;
        RECT 86.755 44.815 86.985 45.635 ;
        RECT 87.155 44.835 87.485 45.465 ;
        RECT 71.535 43.085 76.880 44.175 ;
        RECT 77.055 43.085 78.265 44.175 ;
        RECT 78.505 44.055 79.965 44.225 ;
        RECT 80.630 44.055 81.485 44.225 ;
        RECT 83.475 44.175 85.165 44.695 ;
        RECT 86.735 44.395 87.065 44.645 ;
        RECT 78.505 43.255 78.865 44.055 ;
        RECT 80.630 43.885 80.960 44.055 ;
        RECT 79.410 43.085 79.580 43.885 ;
        RECT 79.790 43.715 80.960 43.885 ;
        RECT 79.790 43.255 80.120 43.715 ;
        RECT 80.290 43.085 80.460 43.545 ;
        RECT 80.630 43.255 80.960 43.715 ;
        RECT 81.130 43.085 81.300 43.885 ;
        RECT 81.655 43.085 85.165 44.175 ;
        RECT 85.335 43.085 85.625 44.250 ;
        RECT 87.235 44.235 87.485 44.835 ;
        RECT 87.655 44.815 87.865 45.635 ;
        RECT 88.095 44.865 91.605 45.635 ;
        RECT 88.095 44.345 89.745 44.865 ;
        RECT 91.780 44.815 92.055 45.635 ;
        RECT 92.225 44.995 92.555 45.465 ;
        RECT 92.725 45.165 92.895 45.635 ;
        RECT 93.065 44.995 93.395 45.465 ;
        RECT 93.565 45.165 93.735 45.635 ;
        RECT 93.905 44.995 94.235 45.465 ;
        RECT 94.405 45.165 94.575 45.635 ;
        RECT 94.745 44.995 95.075 45.465 ;
        RECT 95.245 45.165 95.530 45.635 ;
        RECT 92.225 44.815 95.745 44.995 ;
        RECT 86.755 43.085 86.985 44.225 ;
        RECT 87.155 43.255 87.485 44.235 ;
        RECT 87.655 43.085 87.865 44.225 ;
        RECT 89.915 44.175 91.605 44.695 ;
        RECT 93.810 44.445 95.175 44.645 ;
        RECT 95.345 44.275 95.745 44.815 ;
        RECT 95.915 44.865 99.425 45.635 ;
        RECT 99.595 44.910 99.885 45.635 ;
        RECT 100.605 45.085 100.775 45.465 ;
        RECT 100.990 45.255 101.320 45.635 ;
        RECT 100.605 44.915 101.320 45.085 ;
        RECT 95.915 44.345 97.565 44.865 ;
        RECT 88.095 43.085 91.605 44.175 ;
        RECT 91.780 44.055 93.815 44.265 ;
        RECT 91.780 43.255 92.055 44.055 ;
        RECT 92.225 43.085 92.555 43.885 ;
        RECT 92.725 43.255 92.895 44.055 ;
        RECT 93.065 43.085 93.315 43.885 ;
        RECT 93.485 43.425 93.815 44.055 ;
        RECT 93.985 43.975 95.745 44.275 ;
        RECT 97.735 44.175 99.425 44.695 ;
        RECT 100.515 44.365 100.870 44.735 ;
        RECT 101.150 44.725 101.320 44.915 ;
        RECT 101.490 44.890 101.745 45.465 ;
        RECT 101.150 44.395 101.405 44.725 ;
        RECT 93.985 43.595 94.155 43.975 ;
        RECT 94.325 43.425 94.655 43.785 ;
        RECT 94.825 43.595 94.995 43.975 ;
        RECT 95.165 43.425 95.580 43.805 ;
        RECT 93.485 43.255 95.580 43.425 ;
        RECT 95.915 43.085 99.425 44.175 ;
        RECT 99.595 43.085 99.885 44.250 ;
        RECT 101.150 44.185 101.320 44.395 ;
        RECT 100.605 44.015 101.320 44.185 ;
        RECT 101.575 44.160 101.745 44.890 ;
        RECT 101.920 44.795 102.180 45.635 ;
        RECT 102.355 44.865 105.865 45.635 ;
        RECT 106.070 45.135 106.320 45.635 ;
        RECT 106.650 45.065 106.820 45.415 ;
        RECT 107.020 45.235 107.350 45.635 ;
        RECT 107.520 45.065 107.690 45.415 ;
        RECT 107.910 45.235 108.290 45.635 ;
        RECT 102.355 44.345 104.005 44.865 ;
        RECT 100.605 43.255 100.775 44.015 ;
        RECT 100.990 43.085 101.320 43.845 ;
        RECT 101.490 43.255 101.745 44.160 ;
        RECT 101.920 43.085 102.180 44.235 ;
        RECT 104.175 44.175 105.865 44.695 ;
        RECT 106.035 44.395 106.320 44.965 ;
        RECT 106.490 44.895 108.300 45.065 ;
        RECT 106.490 44.225 106.660 44.895 ;
        RECT 102.355 43.085 105.865 44.175 ;
        RECT 106.065 44.055 106.660 44.225 ;
        RECT 106.830 44.100 107.000 44.725 ;
        RECT 107.230 44.270 107.560 44.725 ;
        RECT 106.065 43.270 106.400 44.055 ;
        RECT 106.830 43.595 107.180 44.100 ;
        RECT 106.785 43.425 107.180 43.595 ;
        RECT 106.830 43.345 107.180 43.425 ;
        RECT 107.350 43.935 107.560 44.270 ;
        RECT 107.790 44.275 107.960 44.725 ;
        RECT 108.130 44.645 108.300 44.895 ;
        RECT 108.470 44.995 108.720 45.465 ;
        RECT 108.890 45.165 109.060 45.635 ;
        RECT 109.230 44.995 109.560 45.465 ;
        RECT 109.730 45.165 109.900 45.635 ;
        RECT 108.470 44.815 110.005 44.995 ;
        RECT 108.130 44.475 109.590 44.645 ;
        RECT 107.790 44.105 108.225 44.275 ;
        RECT 109.760 44.265 110.005 44.815 ;
        RECT 110.175 44.865 113.685 45.635 ;
        RECT 113.855 44.910 114.145 45.635 ;
        RECT 115.270 45.135 115.520 45.635 ;
        RECT 115.850 45.065 116.020 45.415 ;
        RECT 116.220 45.235 116.550 45.635 ;
        RECT 116.720 45.065 116.890 45.415 ;
        RECT 117.110 45.235 117.490 45.635 ;
        RECT 110.175 44.345 111.825 44.865 ;
        RECT 108.430 44.095 110.005 44.265 ;
        RECT 111.995 44.175 113.685 44.695 ;
        RECT 115.235 44.395 115.520 44.965 ;
        RECT 115.690 44.895 117.500 45.065 ;
        RECT 107.350 43.345 107.670 43.935 ;
        RECT 107.955 43.085 108.205 43.925 ;
        RECT 108.430 43.255 108.680 44.095 ;
        RECT 108.850 43.085 109.100 43.925 ;
        RECT 109.270 43.255 109.520 44.095 ;
        RECT 109.690 43.085 109.940 43.925 ;
        RECT 110.175 43.085 113.685 44.175 ;
        RECT 113.855 43.085 114.145 44.250 ;
        RECT 115.690 44.225 115.860 44.895 ;
        RECT 115.265 44.055 115.860 44.225 ;
        RECT 116.030 44.100 116.200 44.725 ;
        RECT 116.430 44.270 116.760 44.725 ;
        RECT 115.265 43.270 115.600 44.055 ;
        RECT 116.030 43.935 116.380 44.100 ;
        RECT 115.985 43.765 116.380 43.935 ;
        RECT 116.030 43.345 116.380 43.765 ;
        RECT 116.550 43.935 116.760 44.270 ;
        RECT 116.990 44.275 117.160 44.725 ;
        RECT 117.330 44.645 117.500 44.895 ;
        RECT 117.670 44.995 117.920 45.465 ;
        RECT 118.090 45.165 118.260 45.635 ;
        RECT 118.430 44.995 118.760 45.465 ;
        RECT 118.930 45.165 119.100 45.635 ;
        RECT 117.670 44.815 119.205 44.995 ;
        RECT 117.330 44.475 118.790 44.645 ;
        RECT 116.990 44.105 117.425 44.275 ;
        RECT 118.960 44.265 119.205 44.815 ;
        RECT 119.375 44.865 122.885 45.635 ;
        RECT 119.375 44.345 121.025 44.865 ;
        RECT 123.095 44.815 123.325 45.635 ;
        RECT 123.495 44.835 123.825 45.465 ;
        RECT 117.630 44.095 119.205 44.265 ;
        RECT 121.195 44.175 122.885 44.695 ;
        RECT 123.075 44.395 123.405 44.645 ;
        RECT 123.575 44.235 123.825 44.835 ;
        RECT 123.995 44.815 124.205 45.635 ;
        RECT 124.435 44.865 127.945 45.635 ;
        RECT 128.115 44.910 128.405 45.635 ;
        RECT 128.610 45.135 128.860 45.635 ;
        RECT 129.190 45.065 129.360 45.415 ;
        RECT 129.560 45.235 129.890 45.635 ;
        RECT 130.060 45.065 130.230 45.415 ;
        RECT 130.450 45.235 130.830 45.635 ;
        RECT 124.435 44.345 126.085 44.865 ;
        RECT 116.550 43.345 116.870 43.935 ;
        RECT 117.155 43.085 117.405 43.925 ;
        RECT 117.630 43.255 117.880 44.095 ;
        RECT 118.050 43.085 118.300 43.925 ;
        RECT 118.470 43.255 118.720 44.095 ;
        RECT 118.890 43.085 119.140 43.925 ;
        RECT 119.375 43.085 122.885 44.175 ;
        RECT 123.095 43.085 123.325 44.225 ;
        RECT 123.495 43.255 123.825 44.235 ;
        RECT 123.995 43.085 124.205 44.225 ;
        RECT 126.255 44.175 127.945 44.695 ;
        RECT 128.575 44.395 128.860 44.965 ;
        RECT 129.030 44.895 130.840 45.065 ;
        RECT 124.435 43.085 127.945 44.175 ;
        RECT 128.115 43.085 128.405 44.250 ;
        RECT 129.030 44.225 129.200 44.895 ;
        RECT 128.605 44.055 129.200 44.225 ;
        RECT 129.370 44.100 129.540 44.725 ;
        RECT 129.770 44.270 130.100 44.725 ;
        RECT 128.605 43.270 128.940 44.055 ;
        RECT 129.370 43.345 129.720 44.100 ;
        RECT 129.890 43.935 130.100 44.270 ;
        RECT 130.330 44.275 130.500 44.725 ;
        RECT 130.670 44.645 130.840 44.895 ;
        RECT 131.010 44.995 131.260 45.465 ;
        RECT 131.430 45.165 131.600 45.635 ;
        RECT 131.770 44.995 132.100 45.465 ;
        RECT 132.270 45.165 132.440 45.635 ;
        RECT 131.010 44.815 132.545 44.995 ;
        RECT 130.670 44.475 132.130 44.645 ;
        RECT 130.330 44.105 130.765 44.275 ;
        RECT 132.300 44.265 132.545 44.815 ;
        RECT 132.715 44.865 136.225 45.635 ;
        RECT 136.945 45.085 137.115 45.465 ;
        RECT 137.330 45.255 137.660 45.635 ;
        RECT 136.945 44.915 137.660 45.085 ;
        RECT 132.715 44.345 134.365 44.865 ;
        RECT 130.970 44.095 132.545 44.265 ;
        RECT 134.535 44.175 136.225 44.695 ;
        RECT 136.855 44.365 137.210 44.735 ;
        RECT 137.490 44.725 137.660 44.915 ;
        RECT 137.830 44.890 138.085 45.465 ;
        RECT 137.490 44.395 137.745 44.725 ;
        RECT 137.490 44.185 137.660 44.395 ;
        RECT 129.890 43.345 130.210 43.935 ;
        RECT 130.495 43.085 130.745 43.925 ;
        RECT 130.970 43.255 131.220 44.095 ;
        RECT 131.390 43.085 131.640 43.925 ;
        RECT 131.810 43.255 132.060 44.095 ;
        RECT 132.230 43.085 132.480 43.925 ;
        RECT 132.715 43.085 136.225 44.175 ;
        RECT 136.945 44.015 137.660 44.185 ;
        RECT 137.915 44.160 138.085 44.890 ;
        RECT 138.260 44.795 138.520 45.635 ;
        RECT 138.695 44.865 142.205 45.635 ;
        RECT 142.375 44.910 142.665 45.635 ;
        RECT 143.385 45.085 143.555 45.465 ;
        RECT 143.770 45.255 144.100 45.635 ;
        RECT 143.385 44.915 144.100 45.085 ;
        RECT 138.695 44.345 140.345 44.865 ;
        RECT 136.945 43.255 137.115 44.015 ;
        RECT 137.330 43.085 137.660 43.845 ;
        RECT 137.830 43.255 138.085 44.160 ;
        RECT 138.260 43.085 138.520 44.235 ;
        RECT 140.515 44.175 142.205 44.695 ;
        RECT 143.295 44.365 143.650 44.735 ;
        RECT 143.930 44.725 144.100 44.915 ;
        RECT 144.270 44.890 144.525 45.465 ;
        RECT 143.930 44.395 144.185 44.725 ;
        RECT 138.695 43.085 142.205 44.175 ;
        RECT 142.375 43.085 142.665 44.250 ;
        RECT 143.930 44.185 144.100 44.395 ;
        RECT 143.385 44.015 144.100 44.185 ;
        RECT 144.355 44.160 144.525 44.890 ;
        RECT 144.700 44.795 144.960 45.635 ;
        RECT 145.135 44.865 148.645 45.635 ;
        RECT 145.135 44.345 146.785 44.865 ;
        RECT 148.820 44.815 149.095 45.635 ;
        RECT 149.265 44.995 149.595 45.465 ;
        RECT 149.765 45.165 149.935 45.635 ;
        RECT 150.105 44.995 150.435 45.465 ;
        RECT 150.605 45.165 150.775 45.635 ;
        RECT 150.945 44.995 151.275 45.465 ;
        RECT 151.445 45.165 151.615 45.635 ;
        RECT 151.785 44.995 152.115 45.465 ;
        RECT 152.285 45.165 152.570 45.635 ;
        RECT 149.265 44.815 152.785 44.995 ;
        RECT 143.385 43.255 143.555 44.015 ;
        RECT 143.770 43.085 144.100 43.845 ;
        RECT 144.270 43.255 144.525 44.160 ;
        RECT 144.700 43.085 144.960 44.235 ;
        RECT 146.955 44.175 148.645 44.695 ;
        RECT 148.870 44.445 150.530 44.645 ;
        RECT 150.850 44.445 152.215 44.645 ;
        RECT 152.385 44.275 152.785 44.815 ;
        RECT 152.955 44.865 156.465 45.635 ;
        RECT 156.635 44.910 156.925 45.635 ;
        RECT 157.185 45.085 157.355 45.375 ;
        RECT 157.525 45.255 157.855 45.635 ;
        RECT 157.185 44.915 157.850 45.085 ;
        RECT 152.955 44.345 154.605 44.865 ;
        RECT 145.135 43.085 148.645 44.175 ;
        RECT 148.820 44.055 150.855 44.265 ;
        RECT 148.820 43.255 149.095 44.055 ;
        RECT 149.265 43.085 149.595 43.885 ;
        RECT 149.765 43.255 149.935 44.055 ;
        RECT 150.105 43.085 150.355 43.885 ;
        RECT 150.525 43.425 150.855 44.055 ;
        RECT 151.025 43.975 152.785 44.275 ;
        RECT 154.775 44.175 156.465 44.695 ;
        RECT 151.025 43.595 151.195 43.975 ;
        RECT 151.365 43.425 151.695 43.785 ;
        RECT 151.865 43.595 152.035 43.975 ;
        RECT 152.205 43.425 152.620 43.805 ;
        RECT 150.525 43.255 152.620 43.425 ;
        RECT 152.955 43.085 156.465 44.175 ;
        RECT 156.635 43.085 156.925 44.250 ;
        RECT 157.100 44.095 157.450 44.745 ;
        RECT 157.620 43.925 157.850 44.915 ;
        RECT 157.185 43.755 157.850 43.925 ;
        RECT 157.185 43.255 157.355 43.755 ;
        RECT 157.525 43.085 157.855 43.585 ;
        RECT 158.025 43.255 158.250 45.375 ;
        RECT 158.465 45.175 158.715 45.635 ;
        RECT 158.900 45.185 159.230 45.355 ;
        RECT 159.410 45.185 160.160 45.355 ;
        RECT 158.450 44.055 158.730 44.655 ;
        RECT 158.900 43.655 159.070 45.185 ;
        RECT 159.240 44.685 159.820 45.015 ;
        RECT 159.240 43.815 159.480 44.685 ;
        RECT 159.990 44.405 160.160 45.185 ;
        RECT 160.410 45.135 160.780 45.635 ;
        RECT 160.960 45.185 161.420 45.355 ;
        RECT 161.650 45.185 162.320 45.355 ;
        RECT 160.960 44.955 161.130 45.185 ;
        RECT 160.330 44.655 161.130 44.955 ;
        RECT 161.300 44.685 161.850 45.015 ;
        RECT 160.330 44.625 160.500 44.655 ;
        RECT 160.620 44.405 160.790 44.475 ;
        RECT 159.990 44.235 160.790 44.405 ;
        RECT 160.280 44.145 160.790 44.235 ;
        RECT 159.670 43.710 160.110 44.065 ;
        RECT 158.450 43.085 158.715 43.545 ;
        RECT 158.900 43.280 159.135 43.655 ;
        RECT 160.280 43.530 160.450 44.145 ;
        RECT 159.380 43.360 160.450 43.530 ;
        RECT 160.620 43.085 160.790 43.885 ;
        RECT 160.960 43.585 161.130 44.655 ;
        RECT 161.300 43.755 161.490 44.475 ;
        RECT 161.660 44.145 161.850 44.685 ;
        RECT 162.150 44.645 162.320 45.185 ;
        RECT 162.635 45.105 162.805 45.635 ;
        RECT 163.100 44.985 163.460 45.425 ;
        RECT 163.635 45.155 163.805 45.635 ;
        RECT 163.995 44.990 164.330 45.415 ;
        RECT 164.505 45.160 164.675 45.635 ;
        RECT 164.850 44.990 165.185 45.415 ;
        RECT 165.355 45.160 165.525 45.635 ;
        RECT 163.100 44.815 163.600 44.985 ;
        RECT 163.995 44.820 165.665 44.990 ;
        RECT 163.430 44.645 163.600 44.815 ;
        RECT 162.150 44.475 163.240 44.645 ;
        RECT 163.430 44.475 165.250 44.645 ;
        RECT 161.660 43.815 161.980 44.145 ;
        RECT 160.960 43.255 161.210 43.585 ;
        RECT 162.150 43.555 162.320 44.475 ;
        RECT 163.430 44.220 163.600 44.475 ;
        RECT 165.420 44.255 165.665 44.820 ;
        RECT 165.835 44.865 169.345 45.635 ;
        RECT 169.515 44.885 170.725 45.635 ;
        RECT 170.895 44.910 171.185 45.635 ;
        RECT 165.835 44.345 167.485 44.865 ;
        RECT 162.490 44.050 163.600 44.220 ;
        RECT 163.995 44.085 165.665 44.255 ;
        RECT 167.655 44.175 169.345 44.695 ;
        RECT 169.515 44.345 170.035 44.885 ;
        RECT 171.355 44.865 173.025 45.635 ;
        RECT 170.205 44.175 170.725 44.715 ;
        RECT 171.355 44.345 172.105 44.865 ;
        RECT 173.745 44.825 173.915 45.635 ;
        RECT 174.085 45.245 175.255 45.465 ;
        RECT 174.085 44.815 174.335 45.245 ;
        RECT 175.425 45.165 175.595 45.635 ;
        RECT 174.505 44.985 174.840 45.075 ;
        RECT 175.765 44.985 176.095 45.465 ;
        RECT 176.265 45.165 176.955 45.635 ;
        RECT 177.125 44.995 177.455 45.465 ;
        RECT 177.625 45.165 177.795 45.635 ;
        RECT 177.965 44.995 178.295 45.465 ;
        RECT 174.505 44.815 176.095 44.985 ;
        RECT 176.525 44.815 178.295 44.995 ;
        RECT 178.465 44.825 178.635 45.635 ;
        RECT 178.805 44.995 179.135 45.445 ;
        RECT 179.305 45.165 179.475 45.635 ;
        RECT 179.645 44.995 179.975 45.445 ;
        RECT 180.145 45.165 180.315 45.635 ;
        RECT 178.805 44.815 180.490 44.995 ;
        RECT 162.490 43.890 163.350 44.050 ;
        RECT 161.435 43.385 162.320 43.555 ;
        RECT 162.500 43.085 162.715 43.585 ;
        RECT 163.180 43.265 163.350 43.890 ;
        RECT 163.635 43.085 163.815 43.865 ;
        RECT 163.995 43.325 164.330 44.085 ;
        RECT 164.510 43.085 164.680 43.915 ;
        RECT 164.850 43.325 165.180 44.085 ;
        RECT 165.350 43.085 165.520 43.915 ;
        RECT 165.835 43.085 169.345 44.175 ;
        RECT 169.515 43.085 170.725 44.175 ;
        RECT 170.895 43.085 171.185 44.250 ;
        RECT 172.275 44.175 173.025 44.695 ;
        RECT 171.355 43.085 173.025 44.175 ;
        RECT 173.655 44.275 174.145 44.645 ;
        RECT 174.375 44.445 174.915 44.645 ;
        RECT 175.085 44.475 175.465 44.645 ;
        RECT 175.085 44.275 175.255 44.475 ;
        RECT 173.655 44.105 175.255 44.275 ;
        RECT 175.805 44.305 176.015 44.815 ;
        RECT 176.525 44.645 176.715 44.815 ;
        RECT 176.185 44.475 176.715 44.645 ;
        RECT 175.425 43.935 175.635 44.265 ;
        RECT 173.705 43.765 175.635 43.935 ;
        RECT 173.705 43.255 173.955 43.765 ;
        RECT 174.125 43.085 174.375 43.595 ;
        RECT 174.545 43.255 174.795 43.765 ;
        RECT 174.965 43.085 175.215 43.595 ;
        RECT 175.385 43.425 175.635 43.765 ;
        RECT 175.805 43.755 176.190 44.305 ;
        RECT 176.525 44.225 176.715 44.475 ;
        RECT 176.885 44.395 177.215 44.645 ;
        RECT 177.385 44.445 178.005 44.645 ;
        RECT 177.045 44.275 177.215 44.395 ;
        RECT 178.175 44.275 178.535 44.645 ;
        RECT 176.525 44.055 176.875 44.225 ;
        RECT 177.045 44.105 178.535 44.275 ;
        RECT 178.705 44.475 180.010 44.645 ;
        RECT 178.705 44.105 179.030 44.475 ;
        RECT 180.180 44.305 180.490 44.815 ;
        RECT 181.015 44.865 184.525 45.635 ;
        RECT 185.155 44.910 185.445 45.635 ;
        RECT 186.165 45.085 186.335 45.375 ;
        RECT 186.505 45.255 186.835 45.635 ;
        RECT 186.165 44.915 186.830 45.085 ;
        RECT 181.015 44.345 182.665 44.865 ;
        RECT 176.705 43.935 176.875 44.055 ;
        RECT 179.685 44.065 180.490 44.305 ;
        RECT 182.835 44.175 184.525 44.695 ;
        RECT 179.685 43.935 179.935 44.065 ;
        RECT 176.705 43.755 177.835 43.935 ;
        RECT 175.805 43.595 176.055 43.755 ;
        RECT 177.585 43.595 177.835 43.755 ;
        RECT 176.225 43.425 176.475 43.585 ;
        RECT 175.385 43.255 176.475 43.425 ;
        RECT 176.745 43.085 176.995 43.585 ;
        RECT 177.165 43.425 177.415 43.585 ;
        RECT 178.005 43.425 178.255 43.935 ;
        RECT 177.165 43.255 178.255 43.425 ;
        RECT 178.425 43.085 178.675 43.925 ;
        RECT 178.845 43.765 179.935 43.935 ;
        RECT 178.845 43.255 179.095 43.765 ;
        RECT 179.265 43.085 179.515 43.555 ;
        RECT 179.685 43.255 179.935 43.765 ;
        RECT 180.105 43.085 180.355 43.895 ;
        RECT 181.015 43.085 184.525 44.175 ;
        RECT 185.155 43.085 185.445 44.250 ;
        RECT 186.080 44.095 186.430 44.745 ;
        RECT 186.600 43.925 186.830 44.915 ;
        RECT 186.165 43.755 186.830 43.925 ;
        RECT 186.165 43.255 186.335 43.755 ;
        RECT 186.505 43.085 186.835 43.585 ;
        RECT 187.005 43.255 187.230 45.375 ;
        RECT 187.445 45.175 187.695 45.635 ;
        RECT 187.880 45.185 188.210 45.355 ;
        RECT 188.390 45.185 189.140 45.355 ;
        RECT 187.430 44.055 187.710 44.655 ;
        RECT 187.880 43.655 188.050 45.185 ;
        RECT 188.220 44.685 188.800 45.015 ;
        RECT 188.220 43.815 188.460 44.685 ;
        RECT 188.970 44.405 189.140 45.185 ;
        RECT 189.390 45.135 189.760 45.635 ;
        RECT 189.940 45.185 190.400 45.355 ;
        RECT 190.630 45.185 191.300 45.355 ;
        RECT 189.940 44.955 190.110 45.185 ;
        RECT 189.310 44.655 190.110 44.955 ;
        RECT 190.280 44.685 190.830 45.015 ;
        RECT 189.310 44.625 189.480 44.655 ;
        RECT 189.600 44.405 189.770 44.475 ;
        RECT 188.970 44.235 189.770 44.405 ;
        RECT 189.260 44.145 189.770 44.235 ;
        RECT 188.650 43.710 189.090 44.065 ;
        RECT 187.430 43.085 187.695 43.545 ;
        RECT 187.880 43.280 188.115 43.655 ;
        RECT 189.260 43.530 189.430 44.145 ;
        RECT 188.360 43.360 189.430 43.530 ;
        RECT 189.600 43.085 189.770 43.885 ;
        RECT 189.940 43.585 190.110 44.655 ;
        RECT 190.280 43.755 190.470 44.475 ;
        RECT 190.640 44.145 190.830 44.685 ;
        RECT 191.130 44.645 191.300 45.185 ;
        RECT 191.615 45.105 191.785 45.635 ;
        RECT 192.080 44.985 192.440 45.425 ;
        RECT 192.615 45.155 192.785 45.635 ;
        RECT 192.975 44.990 193.310 45.415 ;
        RECT 193.485 45.160 193.655 45.635 ;
        RECT 193.830 44.990 194.165 45.415 ;
        RECT 194.335 45.160 194.505 45.635 ;
        RECT 192.080 44.815 192.580 44.985 ;
        RECT 192.975 44.820 194.645 44.990 ;
        RECT 192.410 44.645 192.580 44.815 ;
        RECT 191.130 44.475 192.220 44.645 ;
        RECT 192.410 44.475 194.230 44.645 ;
        RECT 190.640 43.815 190.960 44.145 ;
        RECT 189.940 43.255 190.190 43.585 ;
        RECT 191.130 43.555 191.300 44.475 ;
        RECT 192.410 44.220 192.580 44.475 ;
        RECT 194.400 44.255 194.645 44.820 ;
        RECT 194.815 44.865 198.325 45.635 ;
        RECT 199.415 44.910 199.705 45.635 ;
        RECT 199.875 44.865 203.385 45.635 ;
        RECT 204.035 45.275 204.375 45.635 ;
        RECT 204.905 45.275 205.235 45.635 ;
        RECT 205.840 45.275 206.615 45.635 ;
        RECT 206.805 45.105 206.975 45.465 ;
        RECT 207.185 45.275 207.515 45.635 ;
        RECT 204.075 44.935 205.665 45.105 ;
        RECT 205.965 45.050 206.975 45.105 ;
        RECT 208.015 45.050 208.295 45.315 ;
        RECT 205.965 44.935 208.295 45.050 ;
        RECT 194.815 44.345 196.465 44.865 ;
        RECT 191.470 44.050 192.580 44.220 ;
        RECT 192.975 44.085 194.645 44.255 ;
        RECT 196.635 44.175 198.325 44.695 ;
        RECT 199.875 44.345 201.525 44.865 ;
        RECT 191.470 43.890 192.330 44.050 ;
        RECT 190.415 43.385 191.300 43.555 ;
        RECT 191.480 43.085 191.695 43.585 ;
        RECT 192.160 43.265 192.330 43.890 ;
        RECT 192.615 43.085 192.795 43.865 ;
        RECT 192.975 43.325 193.310 44.085 ;
        RECT 193.490 43.085 193.660 43.915 ;
        RECT 193.830 43.325 194.160 44.085 ;
        RECT 194.330 43.085 194.500 43.915 ;
        RECT 194.815 43.085 198.325 44.175 ;
        RECT 199.415 43.085 199.705 44.250 ;
        RECT 201.695 44.175 203.385 44.695 ;
        RECT 199.875 43.085 203.385 44.175 ;
        RECT 204.075 44.135 204.560 44.935 ;
        RECT 205.965 44.725 206.135 44.935 ;
        RECT 206.805 44.880 208.295 44.935 ;
        RECT 204.730 44.395 206.135 44.725 ;
        RECT 204.075 43.965 205.665 44.135 ;
        RECT 204.045 43.085 204.375 43.785 ;
        RECT 204.555 43.535 204.725 43.965 ;
        RECT 204.905 43.085 205.235 43.785 ;
        RECT 205.415 43.535 205.665 43.965 ;
        RECT 205.845 43.085 206.095 44.205 ;
        RECT 206.325 44.195 206.635 44.725 ;
        RECT 206.385 43.425 206.555 44.025 ;
        RECT 206.805 43.595 206.975 44.880 ;
        RECT 208.875 44.835 209.155 45.635 ;
        RECT 209.535 44.865 213.045 45.635 ;
        RECT 213.675 44.910 213.965 45.635 ;
        RECT 214.515 45.345 214.850 45.465 ;
        RECT 214.515 45.155 215.775 45.345 ;
        RECT 215.955 45.275 216.285 45.635 ;
        RECT 216.860 45.275 217.190 45.635 ;
        RECT 214.515 44.915 214.850 45.155 ;
        RECT 215.585 45.105 215.775 45.155 ;
        RECT 216.500 45.105 216.690 45.205 ;
        RECT 217.360 45.105 217.550 45.465 ;
        RECT 217.720 45.275 218.050 45.635 ;
        RECT 207.355 44.445 207.750 44.710 ;
        RECT 207.920 44.445 208.445 44.710 ;
        RECT 207.215 43.870 207.395 44.275 ;
        RECT 207.575 44.210 207.750 44.445 ;
        RECT 208.615 44.430 209.030 44.665 ;
        RECT 208.615 44.210 208.865 44.430 ;
        RECT 209.535 44.345 211.185 44.865 ;
        RECT 207.575 44.040 208.865 44.210 ;
        RECT 209.035 43.870 209.290 44.260 ;
        RECT 211.355 44.175 213.045 44.695 ;
        RECT 214.165 44.380 214.925 44.725 ;
        RECT 215.115 44.380 215.405 44.975 ;
        RECT 215.585 44.915 216.330 45.105 ;
        RECT 215.575 44.395 215.950 44.725 ;
        RECT 216.120 44.700 216.330 44.915 ;
        RECT 216.500 44.875 218.105 45.105 ;
        RECT 207.215 43.700 209.290 43.870 ;
        RECT 207.215 43.425 207.395 43.700 ;
        RECT 206.385 43.255 207.395 43.425 ;
        RECT 207.565 43.085 207.895 43.445 ;
        RECT 208.065 43.255 208.235 43.700 ;
        RECT 208.405 43.085 208.735 43.445 ;
        RECT 208.960 43.325 209.290 43.700 ;
        RECT 209.535 43.085 213.045 44.175 ;
        RECT 213.675 43.085 213.965 44.250 ;
        RECT 214.165 43.385 214.415 44.380 ;
        RECT 216.120 44.365 217.655 44.700 ;
        RECT 216.120 44.140 216.330 44.365 ;
        RECT 217.825 44.185 218.105 44.875 ;
        RECT 218.275 44.865 221.785 45.635 ;
        RECT 222.045 45.085 222.215 45.465 ;
        RECT 222.430 45.255 222.760 45.635 ;
        RECT 222.045 44.915 222.760 45.085 ;
        RECT 218.275 44.345 219.925 44.865 ;
        RECT 214.595 43.970 216.330 44.140 ;
        RECT 214.595 43.255 214.775 43.970 ;
        RECT 214.945 43.085 215.395 43.785 ;
        RECT 215.570 43.255 215.750 43.970 ;
        RECT 216.500 43.960 218.105 44.185 ;
        RECT 220.095 44.175 221.785 44.695 ;
        RECT 221.955 44.365 222.310 44.735 ;
        RECT 222.590 44.725 222.760 44.915 ;
        RECT 222.930 44.890 223.185 45.465 ;
        RECT 222.590 44.395 222.845 44.725 ;
        RECT 222.590 44.185 222.760 44.395 ;
        RECT 215.960 43.085 216.290 43.785 ;
        RECT 216.500 43.255 216.690 43.960 ;
        RECT 217.360 43.955 218.105 43.960 ;
        RECT 216.860 43.085 217.190 43.785 ;
        RECT 217.360 43.255 217.550 43.955 ;
        RECT 217.720 43.085 218.050 43.785 ;
        RECT 218.275 43.085 221.785 44.175 ;
        RECT 222.045 44.015 222.760 44.185 ;
        RECT 223.015 44.160 223.185 44.890 ;
        RECT 223.360 44.795 223.620 45.635 ;
        RECT 223.795 44.865 227.305 45.635 ;
        RECT 227.935 44.910 228.225 45.635 ;
        RECT 228.395 44.995 228.735 45.465 ;
        RECT 228.905 45.165 229.075 45.635 ;
        RECT 229.245 44.995 229.575 45.465 ;
        RECT 229.745 45.165 230.445 45.635 ;
        RECT 223.795 44.345 225.445 44.865 ;
        RECT 228.395 44.815 230.400 44.995 ;
        RECT 230.615 44.985 230.945 45.455 ;
        RECT 231.115 45.165 231.285 45.635 ;
        RECT 231.455 44.985 231.785 45.455 ;
        RECT 231.955 45.165 232.125 45.635 ;
        RECT 230.615 44.815 232.365 44.985 ;
        RECT 222.045 43.255 222.215 44.015 ;
        RECT 222.430 43.085 222.760 43.845 ;
        RECT 222.930 43.255 223.185 44.160 ;
        RECT 223.360 43.085 223.620 44.235 ;
        RECT 225.615 44.175 227.305 44.695 ;
        RECT 230.180 44.645 230.400 44.815 ;
        RECT 228.395 44.395 228.735 44.645 ;
        RECT 228.905 44.395 229.365 44.645 ;
        RECT 229.535 44.395 230.010 44.645 ;
        RECT 230.180 44.475 231.905 44.645 ;
        RECT 223.795 43.085 227.305 44.175 ;
        RECT 227.935 43.085 228.225 44.250 ;
        RECT 228.395 43.425 228.735 44.225 ;
        RECT 228.905 43.670 229.140 44.395 ;
        RECT 230.180 44.225 230.400 44.475 ;
        RECT 230.755 44.265 230.925 44.275 ;
        RECT 232.075 44.265 232.365 44.815 ;
        RECT 232.535 44.865 236.045 45.635 ;
        RECT 236.305 45.085 236.475 45.465 ;
        RECT 236.690 45.255 237.020 45.635 ;
        RECT 236.305 44.915 237.020 45.085 ;
        RECT 232.535 44.345 234.185 44.865 ;
        RECT 229.310 44.055 230.400 44.225 ;
        RECT 230.655 44.095 232.365 44.265 ;
        RECT 234.355 44.175 236.045 44.695 ;
        RECT 236.215 44.365 236.570 44.735 ;
        RECT 236.850 44.725 237.020 44.915 ;
        RECT 237.190 44.890 237.445 45.465 ;
        RECT 236.850 44.395 237.105 44.725 ;
        RECT 236.850 44.185 237.020 44.395 ;
        RECT 229.310 43.425 229.575 44.055 ;
        RECT 228.395 43.255 229.575 43.425 ;
        RECT 229.745 43.085 230.445 43.885 ;
        RECT 230.655 43.255 230.905 44.095 ;
        RECT 231.075 43.085 231.325 43.925 ;
        RECT 231.495 43.255 231.745 44.095 ;
        RECT 231.915 43.085 232.165 43.925 ;
        RECT 232.535 43.085 236.045 44.175 ;
        RECT 236.305 44.015 237.020 44.185 ;
        RECT 237.275 44.160 237.445 44.890 ;
        RECT 237.620 44.795 237.880 45.635 ;
        RECT 238.055 44.865 241.565 45.635 ;
        RECT 242.195 44.910 242.485 45.635 ;
        RECT 242.675 45.125 242.915 45.635 ;
        RECT 238.055 44.345 239.705 44.865 ;
        RECT 236.305 43.255 236.475 44.015 ;
        RECT 236.690 43.085 237.020 43.845 ;
        RECT 237.190 43.255 237.445 44.160 ;
        RECT 237.620 43.085 237.880 44.235 ;
        RECT 239.875 44.175 241.565 44.695 ;
        RECT 242.660 44.395 242.915 44.955 ;
        RECT 243.085 44.895 243.415 45.430 ;
        RECT 243.630 44.895 243.800 45.635 ;
        RECT 244.010 44.985 244.340 45.455 ;
        RECT 244.510 45.155 244.680 45.635 ;
        RECT 244.850 44.985 245.180 45.455 ;
        RECT 245.350 45.155 245.520 45.635 ;
        RECT 238.055 43.085 241.565 44.175 ;
        RECT 242.195 43.085 242.485 44.250 ;
        RECT 243.085 44.225 243.265 44.895 ;
        RECT 244.010 44.815 245.705 44.985 ;
        RECT 243.435 44.395 243.810 44.725 ;
        RECT 243.980 44.475 245.190 44.645 ;
        RECT 243.980 44.225 244.185 44.475 ;
        RECT 245.360 44.225 245.705 44.815 ;
        RECT 245.875 44.865 249.385 45.635 ;
        RECT 249.575 45.125 249.815 45.635 ;
        RECT 245.875 44.345 247.525 44.865 ;
        RECT 242.725 44.055 244.185 44.225 ;
        RECT 244.850 44.055 245.705 44.225 ;
        RECT 247.695 44.175 249.385 44.695 ;
        RECT 249.560 44.395 249.815 44.955 ;
        RECT 249.985 44.895 250.315 45.430 ;
        RECT 250.530 44.895 250.700 45.635 ;
        RECT 250.910 44.985 251.240 45.455 ;
        RECT 251.410 45.155 251.580 45.635 ;
        RECT 251.750 44.985 252.080 45.455 ;
        RECT 252.250 45.155 252.420 45.635 ;
        RECT 249.985 44.225 250.165 44.895 ;
        RECT 250.910 44.815 252.605 44.985 ;
        RECT 250.335 44.395 250.710 44.725 ;
        RECT 250.880 44.475 252.090 44.645 ;
        RECT 250.880 44.225 251.085 44.475 ;
        RECT 252.260 44.225 252.605 44.815 ;
        RECT 252.775 44.865 256.285 45.635 ;
        RECT 256.455 44.910 256.745 45.635 ;
        RECT 256.935 45.125 257.175 45.635 ;
        RECT 252.775 44.345 254.425 44.865 ;
        RECT 242.725 43.255 243.085 44.055 ;
        RECT 244.850 43.885 245.180 44.055 ;
        RECT 243.630 43.085 243.800 43.885 ;
        RECT 244.010 43.715 245.180 43.885 ;
        RECT 244.010 43.255 244.340 43.715 ;
        RECT 244.510 43.085 244.680 43.545 ;
        RECT 244.850 43.255 245.180 43.715 ;
        RECT 245.350 43.085 245.520 43.885 ;
        RECT 245.875 43.085 249.385 44.175 ;
        RECT 249.625 44.055 251.085 44.225 ;
        RECT 251.750 44.055 252.605 44.225 ;
        RECT 254.595 44.175 256.285 44.695 ;
        RECT 256.920 44.395 257.175 44.955 ;
        RECT 257.345 44.895 257.675 45.430 ;
        RECT 257.890 44.895 258.060 45.635 ;
        RECT 258.270 44.985 258.600 45.455 ;
        RECT 258.770 45.155 258.940 45.635 ;
        RECT 259.110 44.985 259.440 45.455 ;
        RECT 259.610 45.155 259.780 45.635 ;
        RECT 249.625 43.255 249.985 44.055 ;
        RECT 251.750 43.885 252.080 44.055 ;
        RECT 250.530 43.085 250.700 43.885 ;
        RECT 250.910 43.715 252.080 43.885 ;
        RECT 250.910 43.255 251.240 43.715 ;
        RECT 251.410 43.085 251.580 43.545 ;
        RECT 251.750 43.255 252.080 43.715 ;
        RECT 252.250 43.085 252.420 43.885 ;
        RECT 252.775 43.085 256.285 44.175 ;
        RECT 256.455 43.085 256.745 44.250 ;
        RECT 257.345 44.225 257.525 44.895 ;
        RECT 258.270 44.815 259.965 44.985 ;
        RECT 257.695 44.395 258.070 44.725 ;
        RECT 258.240 44.475 259.450 44.645 ;
        RECT 258.240 44.225 258.445 44.475 ;
        RECT 259.620 44.225 259.965 44.815 ;
        RECT 260.135 44.865 263.645 45.635 ;
        RECT 263.905 45.085 264.075 45.465 ;
        RECT 264.290 45.255 264.620 45.635 ;
        RECT 263.905 44.915 264.620 45.085 ;
        RECT 260.135 44.345 261.785 44.865 ;
        RECT 256.985 44.055 258.445 44.225 ;
        RECT 259.110 44.055 259.965 44.225 ;
        RECT 261.955 44.175 263.645 44.695 ;
        RECT 263.815 44.365 264.170 44.735 ;
        RECT 264.450 44.725 264.620 44.915 ;
        RECT 264.790 44.890 265.045 45.465 ;
        RECT 264.450 44.395 264.705 44.725 ;
        RECT 264.450 44.185 264.620 44.395 ;
        RECT 256.985 43.255 257.345 44.055 ;
        RECT 259.110 43.885 259.440 44.055 ;
        RECT 257.890 43.085 258.060 43.885 ;
        RECT 258.270 43.715 259.440 43.885 ;
        RECT 258.270 43.255 258.600 43.715 ;
        RECT 258.770 43.085 258.940 43.545 ;
        RECT 259.110 43.255 259.440 43.715 ;
        RECT 259.610 43.085 259.780 43.885 ;
        RECT 260.135 43.085 263.645 44.175 ;
        RECT 263.905 44.015 264.620 44.185 ;
        RECT 264.875 44.160 265.045 44.890 ;
        RECT 265.220 44.795 265.480 45.635 ;
        RECT 265.655 44.865 269.165 45.635 ;
        RECT 269.335 44.885 270.545 45.635 ;
        RECT 270.715 44.910 271.005 45.635 ;
        RECT 271.265 45.085 271.435 45.465 ;
        RECT 271.650 45.255 271.980 45.635 ;
        RECT 271.265 44.915 271.980 45.085 ;
        RECT 265.655 44.345 267.305 44.865 ;
        RECT 263.905 43.255 264.075 44.015 ;
        RECT 264.290 43.085 264.620 43.845 ;
        RECT 264.790 43.255 265.045 44.160 ;
        RECT 265.220 43.085 265.480 44.235 ;
        RECT 267.475 44.175 269.165 44.695 ;
        RECT 269.335 44.345 269.855 44.885 ;
        RECT 270.025 44.175 270.545 44.715 ;
        RECT 271.175 44.365 271.530 44.735 ;
        RECT 271.810 44.725 271.980 44.915 ;
        RECT 272.150 44.890 272.405 45.465 ;
        RECT 271.810 44.395 272.065 44.725 ;
        RECT 265.655 43.085 269.165 44.175 ;
        RECT 269.335 43.085 270.545 44.175 ;
        RECT 270.715 43.085 271.005 44.250 ;
        RECT 271.810 44.185 271.980 44.395 ;
        RECT 271.265 44.015 271.980 44.185 ;
        RECT 272.235 44.160 272.405 44.890 ;
        RECT 272.580 44.795 272.840 45.635 ;
        RECT 273.015 44.865 276.525 45.635 ;
        RECT 273.015 44.345 274.665 44.865 ;
        RECT 276.700 44.815 276.975 45.635 ;
        RECT 277.145 44.995 277.475 45.465 ;
        RECT 277.645 45.165 277.815 45.635 ;
        RECT 277.985 44.995 278.315 45.465 ;
        RECT 278.485 45.165 278.655 45.635 ;
        RECT 278.825 44.995 279.155 45.465 ;
        RECT 279.325 45.165 279.495 45.635 ;
        RECT 279.665 44.995 279.995 45.465 ;
        RECT 280.165 45.165 280.450 45.635 ;
        RECT 277.145 44.815 280.665 44.995 ;
        RECT 271.265 43.255 271.435 44.015 ;
        RECT 271.650 43.085 271.980 43.845 ;
        RECT 272.150 43.255 272.405 44.160 ;
        RECT 272.580 43.085 272.840 44.235 ;
        RECT 274.835 44.175 276.525 44.695 ;
        RECT 276.750 44.445 278.410 44.645 ;
        RECT 278.730 44.445 280.095 44.645 ;
        RECT 280.265 44.275 280.665 44.815 ;
        RECT 280.835 44.865 284.345 45.635 ;
        RECT 284.975 44.910 285.265 45.635 ;
        RECT 280.835 44.345 282.485 44.865 ;
        RECT 285.440 44.815 285.715 45.635 ;
        RECT 285.885 44.995 286.215 45.465 ;
        RECT 286.385 45.165 286.555 45.635 ;
        RECT 286.725 44.995 287.055 45.465 ;
        RECT 287.225 45.165 287.395 45.635 ;
        RECT 287.565 44.995 287.895 45.465 ;
        RECT 288.065 45.165 288.235 45.635 ;
        RECT 288.405 44.995 288.735 45.465 ;
        RECT 288.905 45.165 289.190 45.635 ;
        RECT 285.885 44.815 289.405 44.995 ;
        RECT 273.015 43.085 276.525 44.175 ;
        RECT 276.700 44.055 278.735 44.265 ;
        RECT 276.700 43.255 276.975 44.055 ;
        RECT 277.145 43.085 277.475 43.885 ;
        RECT 277.645 43.255 277.815 44.055 ;
        RECT 277.985 43.085 278.235 43.885 ;
        RECT 278.405 43.425 278.735 44.055 ;
        RECT 278.905 43.975 280.665 44.275 ;
        RECT 282.655 44.175 284.345 44.695 ;
        RECT 285.490 44.445 287.150 44.645 ;
        RECT 287.470 44.445 288.835 44.645 ;
        RECT 289.005 44.275 289.405 44.815 ;
        RECT 289.575 44.865 293.085 45.635 ;
        RECT 293.345 45.085 293.515 45.465 ;
        RECT 293.730 45.255 294.060 45.635 ;
        RECT 293.345 44.915 294.060 45.085 ;
        RECT 289.575 44.345 291.225 44.865 ;
        RECT 278.905 43.595 279.075 43.975 ;
        RECT 279.245 43.425 279.575 43.785 ;
        RECT 279.745 43.595 279.915 43.975 ;
        RECT 280.085 43.425 280.500 43.805 ;
        RECT 278.405 43.255 280.500 43.425 ;
        RECT 280.835 43.085 284.345 44.175 ;
        RECT 284.975 43.085 285.265 44.250 ;
        RECT 285.440 44.055 287.475 44.265 ;
        RECT 285.440 43.255 285.715 44.055 ;
        RECT 285.885 43.085 286.215 43.885 ;
        RECT 286.385 43.255 286.555 44.055 ;
        RECT 286.725 43.085 286.975 43.885 ;
        RECT 287.145 43.425 287.475 44.055 ;
        RECT 287.645 43.975 289.405 44.275 ;
        RECT 291.395 44.175 293.085 44.695 ;
        RECT 293.255 44.365 293.610 44.735 ;
        RECT 293.890 44.725 294.060 44.915 ;
        RECT 294.230 44.890 294.485 45.465 ;
        RECT 293.890 44.395 294.145 44.725 ;
        RECT 293.890 44.185 294.060 44.395 ;
        RECT 287.645 43.595 287.815 43.975 ;
        RECT 287.985 43.425 288.315 43.785 ;
        RECT 288.485 43.595 288.655 43.975 ;
        RECT 288.825 43.425 289.240 43.805 ;
        RECT 287.145 43.255 289.240 43.425 ;
        RECT 289.575 43.085 293.085 44.175 ;
        RECT 293.345 44.015 294.060 44.185 ;
        RECT 294.315 44.160 294.485 44.890 ;
        RECT 294.660 44.795 294.920 45.635 ;
        RECT 295.095 44.865 298.605 45.635 ;
        RECT 299.235 44.910 299.525 45.635 ;
        RECT 295.095 44.345 296.745 44.865 ;
        RECT 299.700 44.815 299.975 45.635 ;
        RECT 300.145 44.995 300.475 45.465 ;
        RECT 300.645 45.165 300.815 45.635 ;
        RECT 300.985 44.995 301.315 45.465 ;
        RECT 301.485 45.165 301.655 45.635 ;
        RECT 301.825 44.995 302.155 45.465 ;
        RECT 302.325 45.165 302.495 45.635 ;
        RECT 302.665 44.995 302.995 45.465 ;
        RECT 303.165 45.165 303.450 45.635 ;
        RECT 300.145 44.815 303.665 44.995 ;
        RECT 293.345 43.255 293.515 44.015 ;
        RECT 293.730 43.085 294.060 43.845 ;
        RECT 294.230 43.255 294.485 44.160 ;
        RECT 294.660 43.085 294.920 44.235 ;
        RECT 296.915 44.175 298.605 44.695 ;
        RECT 299.750 44.445 301.410 44.645 ;
        RECT 301.730 44.445 303.095 44.645 ;
        RECT 303.265 44.275 303.665 44.815 ;
        RECT 303.835 44.865 307.345 45.635 ;
        RECT 307.605 45.085 307.775 45.465 ;
        RECT 307.990 45.255 308.320 45.635 ;
        RECT 307.605 44.915 308.320 45.085 ;
        RECT 303.835 44.345 305.485 44.865 ;
        RECT 295.095 43.085 298.605 44.175 ;
        RECT 299.235 43.085 299.525 44.250 ;
        RECT 299.700 44.055 301.735 44.265 ;
        RECT 299.700 43.255 299.975 44.055 ;
        RECT 300.145 43.085 300.475 43.885 ;
        RECT 300.645 43.255 300.815 44.055 ;
        RECT 300.985 43.085 301.235 43.885 ;
        RECT 301.405 43.425 301.735 44.055 ;
        RECT 301.905 43.975 303.665 44.275 ;
        RECT 305.655 44.175 307.345 44.695 ;
        RECT 307.515 44.365 307.870 44.735 ;
        RECT 308.150 44.725 308.320 44.915 ;
        RECT 308.490 44.890 308.745 45.465 ;
        RECT 308.150 44.395 308.405 44.725 ;
        RECT 308.150 44.185 308.320 44.395 ;
        RECT 301.905 43.595 302.075 43.975 ;
        RECT 302.245 43.425 302.575 43.785 ;
        RECT 302.745 43.595 302.915 43.975 ;
        RECT 303.085 43.425 303.500 43.805 ;
        RECT 301.405 43.255 303.500 43.425 ;
        RECT 303.835 43.085 307.345 44.175 ;
        RECT 307.605 44.015 308.320 44.185 ;
        RECT 308.575 44.160 308.745 44.890 ;
        RECT 308.920 44.795 309.180 45.635 ;
        RECT 309.355 44.865 312.865 45.635 ;
        RECT 313.495 44.910 313.785 45.635 ;
        RECT 309.355 44.345 311.005 44.865 ;
        RECT 313.960 44.815 314.235 45.635 ;
        RECT 314.405 44.995 314.735 45.465 ;
        RECT 314.905 45.165 315.075 45.635 ;
        RECT 315.245 44.995 315.575 45.465 ;
        RECT 315.745 45.165 315.915 45.635 ;
        RECT 316.085 44.995 316.415 45.465 ;
        RECT 316.585 45.165 316.755 45.635 ;
        RECT 316.925 44.995 317.255 45.465 ;
        RECT 317.425 45.165 317.710 45.635 ;
        RECT 314.405 44.815 317.925 44.995 ;
        RECT 307.605 43.255 307.775 44.015 ;
        RECT 307.990 43.085 308.320 43.845 ;
        RECT 308.490 43.255 308.745 44.160 ;
        RECT 308.920 43.085 309.180 44.235 ;
        RECT 311.175 44.175 312.865 44.695 ;
        RECT 314.010 44.445 315.670 44.645 ;
        RECT 315.990 44.445 317.355 44.645 ;
        RECT 317.525 44.275 317.925 44.815 ;
        RECT 318.095 44.865 321.605 45.635 ;
        RECT 321.865 45.085 322.035 45.465 ;
        RECT 322.250 45.255 322.580 45.635 ;
        RECT 321.865 44.915 322.580 45.085 ;
        RECT 318.095 44.345 319.745 44.865 ;
        RECT 309.355 43.085 312.865 44.175 ;
        RECT 313.495 43.085 313.785 44.250 ;
        RECT 313.960 44.055 315.995 44.265 ;
        RECT 313.960 43.255 314.235 44.055 ;
        RECT 314.405 43.085 314.735 43.885 ;
        RECT 314.905 43.255 315.075 44.055 ;
        RECT 315.245 43.085 315.495 43.885 ;
        RECT 315.665 43.425 315.995 44.055 ;
        RECT 316.165 43.975 317.925 44.275 ;
        RECT 319.915 44.175 321.605 44.695 ;
        RECT 321.775 44.365 322.130 44.735 ;
        RECT 322.410 44.725 322.580 44.915 ;
        RECT 322.750 44.890 323.005 45.465 ;
        RECT 322.410 44.395 322.665 44.725 ;
        RECT 322.410 44.185 322.580 44.395 ;
        RECT 316.165 43.595 316.335 43.975 ;
        RECT 316.505 43.425 316.835 43.785 ;
        RECT 317.005 43.595 317.175 43.975 ;
        RECT 317.345 43.425 317.760 43.805 ;
        RECT 315.665 43.255 317.760 43.425 ;
        RECT 318.095 43.085 321.605 44.175 ;
        RECT 321.865 44.015 322.580 44.185 ;
        RECT 322.835 44.160 323.005 44.890 ;
        RECT 323.180 44.795 323.440 45.635 ;
        RECT 323.615 44.865 327.125 45.635 ;
        RECT 327.755 44.910 328.045 45.635 ;
        RECT 323.615 44.345 325.265 44.865 ;
        RECT 328.220 44.815 328.495 45.635 ;
        RECT 328.665 44.995 328.995 45.465 ;
        RECT 329.165 45.165 329.335 45.635 ;
        RECT 329.505 44.995 329.835 45.465 ;
        RECT 330.005 45.165 330.175 45.635 ;
        RECT 330.345 44.995 330.675 45.465 ;
        RECT 330.845 45.165 331.015 45.635 ;
        RECT 331.185 44.995 331.515 45.465 ;
        RECT 331.685 45.165 331.970 45.635 ;
        RECT 328.665 44.815 332.185 44.995 ;
        RECT 321.865 43.255 322.035 44.015 ;
        RECT 322.250 43.085 322.580 43.845 ;
        RECT 322.750 43.255 323.005 44.160 ;
        RECT 323.180 43.085 323.440 44.235 ;
        RECT 325.435 44.175 327.125 44.695 ;
        RECT 328.270 44.445 329.930 44.645 ;
        RECT 330.250 44.445 331.615 44.645 ;
        RECT 331.785 44.275 332.185 44.815 ;
        RECT 332.355 44.865 335.865 45.635 ;
        RECT 336.125 45.085 336.295 45.465 ;
        RECT 336.510 45.255 336.840 45.635 ;
        RECT 336.125 44.915 336.840 45.085 ;
        RECT 332.355 44.345 334.005 44.865 ;
        RECT 323.615 43.085 327.125 44.175 ;
        RECT 327.755 43.085 328.045 44.250 ;
        RECT 328.220 44.055 330.255 44.265 ;
        RECT 328.220 43.255 328.495 44.055 ;
        RECT 328.665 43.085 328.995 43.885 ;
        RECT 329.165 43.255 329.335 44.055 ;
        RECT 329.505 43.085 329.755 43.885 ;
        RECT 329.925 43.425 330.255 44.055 ;
        RECT 330.425 43.975 332.185 44.275 ;
        RECT 334.175 44.175 335.865 44.695 ;
        RECT 336.035 44.365 336.390 44.735 ;
        RECT 336.670 44.725 336.840 44.915 ;
        RECT 337.010 44.890 337.265 45.465 ;
        RECT 336.670 44.395 336.925 44.725 ;
        RECT 336.670 44.185 336.840 44.395 ;
        RECT 330.425 43.595 330.595 43.975 ;
        RECT 330.765 43.425 331.095 43.785 ;
        RECT 331.265 43.595 331.435 43.975 ;
        RECT 331.605 43.425 332.020 43.805 ;
        RECT 329.925 43.255 332.020 43.425 ;
        RECT 332.355 43.085 335.865 44.175 ;
        RECT 336.125 44.015 336.840 44.185 ;
        RECT 337.095 44.160 337.265 44.890 ;
        RECT 337.440 44.795 337.700 45.635 ;
        RECT 337.875 44.865 341.385 45.635 ;
        RECT 342.015 44.910 342.305 45.635 ;
        RECT 342.475 44.865 344.145 45.635 ;
        RECT 337.875 44.345 339.525 44.865 ;
        RECT 336.125 43.255 336.295 44.015 ;
        RECT 336.510 43.085 336.840 43.845 ;
        RECT 337.010 43.255 337.265 44.160 ;
        RECT 337.440 43.085 337.700 44.235 ;
        RECT 339.695 44.175 341.385 44.695 ;
        RECT 342.475 44.345 343.225 44.865 ;
        RECT 337.875 43.085 341.385 44.175 ;
        RECT 342.015 43.085 342.305 44.250 ;
        RECT 343.395 44.175 344.145 44.695 ;
        RECT 342.475 43.085 344.145 44.175 ;
        RECT 344.775 43.255 345.525 45.465 ;
        RECT 345.870 45.165 346.040 45.635 ;
        RECT 346.210 44.995 346.540 45.455 ;
        RECT 346.710 45.165 346.880 45.635 ;
        RECT 347.050 44.995 347.380 45.465 ;
        RECT 347.550 45.165 347.720 45.635 ;
        RECT 347.990 45.245 350.080 45.465 ;
        RECT 345.695 44.815 347.380 44.995 ;
        RECT 348.025 44.985 349.580 45.075 ;
        RECT 347.550 44.815 349.580 44.985 ;
        RECT 349.750 44.985 350.080 45.245 ;
        RECT 350.250 45.165 350.420 45.635 ;
        RECT 350.590 44.995 350.920 45.465 ;
        RECT 351.090 45.165 351.260 45.635 ;
        RECT 351.430 44.995 351.760 45.465 ;
        RECT 350.590 44.985 351.760 44.995 ;
        RECT 349.750 44.815 351.760 44.985 ;
        RECT 352.135 44.865 355.645 45.635 ;
        RECT 356.275 44.910 356.565 45.635 ;
        RECT 345.695 44.275 345.980 44.815 ;
        RECT 347.550 44.645 347.840 44.815 ;
        RECT 346.150 44.445 347.840 44.645 ;
        RECT 345.695 44.105 347.340 44.275 ;
        RECT 345.830 43.085 346.080 43.895 ;
        RECT 346.250 43.255 346.500 44.105 ;
        RECT 346.670 43.085 346.920 43.925 ;
        RECT 347.090 43.255 347.340 44.105 ;
        RECT 347.510 43.935 347.840 44.445 ;
        RECT 348.030 44.275 348.565 44.645 ;
        RECT 348.735 44.445 349.290 44.645 ;
        RECT 349.460 44.275 349.790 44.645 ;
        RECT 348.030 44.105 349.790 44.275 ;
        RECT 349.960 44.275 350.290 44.645 ;
        RECT 350.510 44.445 351.005 44.645 ;
        RECT 351.175 44.445 351.965 44.645 ;
        RECT 351.175 44.275 351.345 44.445 ;
        RECT 352.135 44.345 353.785 44.865 ;
        RECT 356.740 44.815 357.015 45.635 ;
        RECT 357.185 44.995 357.515 45.465 ;
        RECT 357.685 45.165 357.855 45.635 ;
        RECT 358.025 44.995 358.355 45.465 ;
        RECT 358.525 45.165 358.695 45.635 ;
        RECT 358.865 44.995 359.195 45.465 ;
        RECT 359.365 45.165 359.535 45.635 ;
        RECT 359.705 44.995 360.035 45.465 ;
        RECT 360.205 45.165 360.490 45.635 ;
        RECT 357.185 44.815 360.705 44.995 ;
        RECT 349.960 44.105 351.345 44.275 ;
        RECT 347.510 43.765 350.880 43.935 ;
        RECT 348.870 43.595 349.120 43.765 ;
        RECT 350.630 43.595 350.880 43.765 ;
        RECT 347.510 43.085 348.280 43.595 ;
        RECT 348.450 43.425 348.700 43.595 ;
        RECT 349.290 43.425 349.540 43.595 ;
        RECT 348.450 43.255 349.540 43.425 ;
        RECT 349.710 43.085 350.040 43.595 ;
        RECT 350.210 43.425 350.460 43.595 ;
        RECT 351.050 43.425 351.300 43.935 ;
        RECT 350.210 43.255 351.300 43.425 ;
        RECT 351.515 43.085 351.720 44.265 ;
        RECT 353.955 44.175 355.645 44.695 ;
        RECT 356.790 44.445 358.450 44.645 ;
        RECT 358.770 44.445 360.135 44.645 ;
        RECT 360.305 44.275 360.705 44.815 ;
        RECT 360.875 44.865 364.385 45.635 ;
        RECT 360.875 44.345 362.525 44.865 ;
        RECT 364.595 44.815 364.825 45.635 ;
        RECT 364.995 44.835 365.325 45.465 ;
        RECT 352.135 43.085 355.645 44.175 ;
        RECT 356.275 43.085 356.565 44.250 ;
        RECT 356.740 44.055 358.775 44.265 ;
        RECT 356.740 43.255 357.015 44.055 ;
        RECT 357.185 43.085 357.515 43.885 ;
        RECT 357.685 43.255 357.855 44.055 ;
        RECT 358.025 43.085 358.275 43.885 ;
        RECT 358.445 43.425 358.775 44.055 ;
        RECT 358.945 43.975 360.705 44.275 ;
        RECT 362.695 44.175 364.385 44.695 ;
        RECT 364.575 44.395 364.905 44.645 ;
        RECT 365.075 44.235 365.325 44.835 ;
        RECT 365.495 44.815 365.705 45.635 ;
        RECT 365.935 44.865 369.445 45.635 ;
        RECT 370.535 44.910 370.825 45.635 ;
        RECT 365.935 44.345 367.585 44.865 ;
        RECT 371.000 44.815 371.275 45.635 ;
        RECT 371.445 44.995 371.775 45.465 ;
        RECT 371.945 45.165 372.115 45.635 ;
        RECT 372.285 44.995 372.615 45.465 ;
        RECT 372.785 45.165 372.955 45.635 ;
        RECT 373.125 44.995 373.455 45.465 ;
        RECT 373.625 45.165 373.795 45.635 ;
        RECT 373.965 44.995 374.295 45.465 ;
        RECT 374.465 45.165 374.750 45.635 ;
        RECT 371.445 44.815 374.965 44.995 ;
        RECT 358.945 43.595 359.115 43.975 ;
        RECT 359.285 43.425 359.615 43.785 ;
        RECT 359.785 43.595 359.955 43.975 ;
        RECT 360.125 43.425 360.540 43.805 ;
        RECT 358.445 43.255 360.540 43.425 ;
        RECT 360.875 43.085 364.385 44.175 ;
        RECT 364.595 43.085 364.825 44.225 ;
        RECT 364.995 43.255 365.325 44.235 ;
        RECT 365.495 43.085 365.705 44.225 ;
        RECT 367.755 44.175 369.445 44.695 ;
        RECT 371.050 44.445 372.710 44.645 ;
        RECT 373.030 44.445 374.395 44.645 ;
        RECT 374.565 44.275 374.965 44.815 ;
        RECT 375.135 44.865 378.645 45.635 ;
        RECT 375.135 44.345 376.785 44.865 ;
        RECT 365.935 43.085 369.445 44.175 ;
        RECT 370.535 43.085 370.825 44.250 ;
        RECT 371.000 44.055 373.035 44.265 ;
        RECT 371.000 43.255 371.275 44.055 ;
        RECT 371.445 43.085 371.775 43.885 ;
        RECT 371.945 43.255 372.115 44.055 ;
        RECT 372.285 43.085 372.535 43.885 ;
        RECT 372.705 43.425 373.035 44.055 ;
        RECT 373.205 43.975 374.965 44.275 ;
        RECT 376.955 44.175 378.645 44.695 ;
        RECT 373.205 43.595 373.375 43.975 ;
        RECT 373.545 43.425 373.875 43.785 ;
        RECT 374.045 43.595 374.215 43.975 ;
        RECT 374.385 43.425 374.800 43.805 ;
        RECT 372.705 43.255 374.800 43.425 ;
        RECT 375.135 43.085 378.645 44.175 ;
        RECT 378.815 43.980 379.335 45.465 ;
        RECT 379.505 44.975 379.845 45.635 ;
        RECT 380.195 44.865 383.705 45.635 ;
        RECT 384.795 44.910 385.085 45.635 ;
        RECT 379.005 43.085 379.335 43.810 ;
        RECT 379.505 43.255 380.025 44.805 ;
        RECT 380.195 44.345 381.845 44.865 ;
        RECT 382.015 44.175 383.705 44.695 ;
        RECT 380.195 43.085 383.705 44.175 ;
        RECT 384.795 43.085 385.085 44.250 ;
        RECT 385.255 43.980 385.775 45.465 ;
        RECT 385.945 44.975 386.285 45.635 ;
        RECT 386.635 44.865 390.145 45.635 ;
        RECT 385.445 43.085 385.775 43.810 ;
        RECT 385.945 43.255 386.465 44.805 ;
        RECT 386.635 44.345 388.285 44.865 ;
        RECT 388.455 44.175 390.145 44.695 ;
        RECT 386.635 43.085 390.145 44.175 ;
        RECT 390.315 43.980 390.835 45.465 ;
        RECT 391.005 44.975 391.345 45.635 ;
        RECT 391.695 44.865 397.040 45.635 ;
        RECT 397.215 44.865 398.885 45.635 ;
        RECT 399.055 44.910 399.345 45.635 ;
        RECT 399.515 44.865 404.860 45.635 ;
        RECT 405.035 44.865 410.380 45.635 ;
        RECT 410.555 44.865 413.145 45.635 ;
        RECT 413.315 44.910 413.605 45.635 ;
        RECT 413.775 44.865 419.120 45.635 ;
        RECT 419.295 44.865 424.640 45.635 ;
        RECT 424.815 44.865 427.405 45.635 ;
        RECT 427.575 44.910 427.865 45.635 ;
        RECT 428.035 44.865 433.380 45.635 ;
        RECT 433.555 44.865 438.900 45.635 ;
        RECT 439.075 44.865 441.665 45.635 ;
        RECT 441.835 44.910 442.125 45.635 ;
        RECT 442.295 44.865 447.640 45.635 ;
        RECT 447.815 44.865 453.160 45.635 ;
        RECT 453.335 44.865 455.925 45.635 ;
        RECT 456.095 44.910 456.385 45.635 ;
        RECT 456.555 44.865 461.900 45.635 ;
        RECT 462.075 44.865 467.420 45.635 ;
        RECT 467.595 44.865 470.185 45.635 ;
        RECT 470.355 44.910 470.645 45.635 ;
        RECT 470.815 44.865 476.160 45.635 ;
        RECT 476.335 44.865 481.680 45.635 ;
        RECT 481.855 44.865 484.445 45.635 ;
        RECT 484.615 44.910 484.905 45.635 ;
        RECT 485.075 44.865 490.420 45.635 ;
        RECT 490.595 44.865 495.940 45.635 ;
        RECT 496.115 44.865 498.705 45.635 ;
        RECT 498.875 44.910 499.165 45.635 ;
        RECT 499.335 44.865 501.005 45.635 ;
        RECT 390.505 43.085 390.835 43.810 ;
        RECT 391.005 43.255 391.525 44.805 ;
        RECT 391.695 44.345 394.275 44.865 ;
        RECT 394.445 44.175 397.040 44.695 ;
        RECT 397.215 44.345 397.965 44.865 ;
        RECT 398.135 44.175 398.885 44.695 ;
        RECT 399.515 44.345 402.095 44.865 ;
        RECT 391.695 43.085 397.040 44.175 ;
        RECT 397.215 43.085 398.885 44.175 ;
        RECT 399.055 43.085 399.345 44.250 ;
        RECT 402.265 44.175 404.860 44.695 ;
        RECT 405.035 44.345 407.615 44.865 ;
        RECT 407.785 44.175 410.380 44.695 ;
        RECT 410.555 44.345 411.765 44.865 ;
        RECT 411.935 44.175 413.145 44.695 ;
        RECT 413.775 44.345 416.355 44.865 ;
        RECT 399.515 43.085 404.860 44.175 ;
        RECT 405.035 43.085 410.380 44.175 ;
        RECT 410.555 43.085 413.145 44.175 ;
        RECT 413.315 43.085 413.605 44.250 ;
        RECT 416.525 44.175 419.120 44.695 ;
        RECT 419.295 44.345 421.875 44.865 ;
        RECT 422.045 44.175 424.640 44.695 ;
        RECT 424.815 44.345 426.025 44.865 ;
        RECT 426.195 44.175 427.405 44.695 ;
        RECT 428.035 44.345 430.615 44.865 ;
        RECT 413.775 43.085 419.120 44.175 ;
        RECT 419.295 43.085 424.640 44.175 ;
        RECT 424.815 43.085 427.405 44.175 ;
        RECT 427.575 43.085 427.865 44.250 ;
        RECT 430.785 44.175 433.380 44.695 ;
        RECT 433.555 44.345 436.135 44.865 ;
        RECT 436.305 44.175 438.900 44.695 ;
        RECT 439.075 44.345 440.285 44.865 ;
        RECT 440.455 44.175 441.665 44.695 ;
        RECT 442.295 44.345 444.875 44.865 ;
        RECT 428.035 43.085 433.380 44.175 ;
        RECT 433.555 43.085 438.900 44.175 ;
        RECT 439.075 43.085 441.665 44.175 ;
        RECT 441.835 43.085 442.125 44.250 ;
        RECT 445.045 44.175 447.640 44.695 ;
        RECT 447.815 44.345 450.395 44.865 ;
        RECT 450.565 44.175 453.160 44.695 ;
        RECT 453.335 44.345 454.545 44.865 ;
        RECT 454.715 44.175 455.925 44.695 ;
        RECT 456.555 44.345 459.135 44.865 ;
        RECT 442.295 43.085 447.640 44.175 ;
        RECT 447.815 43.085 453.160 44.175 ;
        RECT 453.335 43.085 455.925 44.175 ;
        RECT 456.095 43.085 456.385 44.250 ;
        RECT 459.305 44.175 461.900 44.695 ;
        RECT 462.075 44.345 464.655 44.865 ;
        RECT 464.825 44.175 467.420 44.695 ;
        RECT 467.595 44.345 468.805 44.865 ;
        RECT 468.975 44.175 470.185 44.695 ;
        RECT 470.815 44.345 473.395 44.865 ;
        RECT 456.555 43.085 461.900 44.175 ;
        RECT 462.075 43.085 467.420 44.175 ;
        RECT 467.595 43.085 470.185 44.175 ;
        RECT 470.355 43.085 470.645 44.250 ;
        RECT 473.565 44.175 476.160 44.695 ;
        RECT 476.335 44.345 478.915 44.865 ;
        RECT 479.085 44.175 481.680 44.695 ;
        RECT 481.855 44.345 483.065 44.865 ;
        RECT 483.235 44.175 484.445 44.695 ;
        RECT 485.075 44.345 487.655 44.865 ;
        RECT 470.815 43.085 476.160 44.175 ;
        RECT 476.335 43.085 481.680 44.175 ;
        RECT 481.855 43.085 484.445 44.175 ;
        RECT 484.615 43.085 484.905 44.250 ;
        RECT 487.825 44.175 490.420 44.695 ;
        RECT 490.595 44.345 493.175 44.865 ;
        RECT 493.345 44.175 495.940 44.695 ;
        RECT 496.115 44.345 497.325 44.865 ;
        RECT 497.495 44.175 498.705 44.695 ;
        RECT 499.335 44.345 500.085 44.865 ;
        RECT 485.075 43.085 490.420 44.175 ;
        RECT 490.595 43.085 495.940 44.175 ;
        RECT 496.115 43.085 498.705 44.175 ;
        RECT 498.875 43.085 499.165 44.250 ;
        RECT 500.255 44.175 501.005 44.695 ;
        RECT 499.335 43.085 501.005 44.175 ;
        RECT 501.635 43.980 502.155 45.465 ;
        RECT 502.325 44.975 502.665 45.635 ;
        RECT 503.015 44.865 508.360 45.635 ;
        RECT 508.535 44.865 512.045 45.635 ;
        RECT 513.135 44.910 513.425 45.635 ;
        RECT 513.595 44.865 518.940 45.635 ;
        RECT 519.115 44.865 524.460 45.635 ;
        RECT 524.635 44.865 527.225 45.635 ;
        RECT 527.395 44.910 527.685 45.635 ;
        RECT 527.855 44.865 533.200 45.635 ;
        RECT 533.375 44.865 538.720 45.635 ;
        RECT 538.895 44.865 541.485 45.635 ;
        RECT 541.655 44.910 541.945 45.635 ;
        RECT 542.115 44.865 547.460 45.635 ;
        RECT 547.635 44.865 552.980 45.635 ;
        RECT 553.155 44.865 555.745 45.635 ;
        RECT 555.915 44.910 556.205 45.635 ;
        RECT 556.375 44.865 561.720 45.635 ;
        RECT 561.895 44.865 567.240 45.635 ;
        RECT 567.415 44.865 570.005 45.635 ;
        RECT 570.175 44.910 570.465 45.635 ;
        RECT 570.635 44.865 575.980 45.635 ;
        RECT 576.155 44.865 581.500 45.635 ;
        RECT 581.675 44.865 584.265 45.635 ;
        RECT 584.435 44.910 584.725 45.635 ;
        RECT 501.825 43.085 502.155 43.810 ;
        RECT 502.325 43.255 502.845 44.805 ;
        RECT 503.015 44.345 505.595 44.865 ;
        RECT 505.765 44.175 508.360 44.695 ;
        RECT 508.535 44.345 510.185 44.865 ;
        RECT 510.355 44.175 512.045 44.695 ;
        RECT 513.595 44.345 516.175 44.865 ;
        RECT 503.015 43.085 508.360 44.175 ;
        RECT 508.535 43.085 512.045 44.175 ;
        RECT 513.135 43.085 513.425 44.250 ;
        RECT 516.345 44.175 518.940 44.695 ;
        RECT 519.115 44.345 521.695 44.865 ;
        RECT 521.865 44.175 524.460 44.695 ;
        RECT 524.635 44.345 525.845 44.865 ;
        RECT 526.015 44.175 527.225 44.695 ;
        RECT 527.855 44.345 530.435 44.865 ;
        RECT 513.595 43.085 518.940 44.175 ;
        RECT 519.115 43.085 524.460 44.175 ;
        RECT 524.635 43.085 527.225 44.175 ;
        RECT 527.395 43.085 527.685 44.250 ;
        RECT 530.605 44.175 533.200 44.695 ;
        RECT 533.375 44.345 535.955 44.865 ;
        RECT 536.125 44.175 538.720 44.695 ;
        RECT 538.895 44.345 540.105 44.865 ;
        RECT 540.275 44.175 541.485 44.695 ;
        RECT 542.115 44.345 544.695 44.865 ;
        RECT 527.855 43.085 533.200 44.175 ;
        RECT 533.375 43.085 538.720 44.175 ;
        RECT 538.895 43.085 541.485 44.175 ;
        RECT 541.655 43.085 541.945 44.250 ;
        RECT 544.865 44.175 547.460 44.695 ;
        RECT 547.635 44.345 550.215 44.865 ;
        RECT 550.385 44.175 552.980 44.695 ;
        RECT 553.155 44.345 554.365 44.865 ;
        RECT 554.535 44.175 555.745 44.695 ;
        RECT 556.375 44.345 558.955 44.865 ;
        RECT 542.115 43.085 547.460 44.175 ;
        RECT 547.635 43.085 552.980 44.175 ;
        RECT 553.155 43.085 555.745 44.175 ;
        RECT 555.915 43.085 556.205 44.250 ;
        RECT 559.125 44.175 561.720 44.695 ;
        RECT 561.895 44.345 564.475 44.865 ;
        RECT 564.645 44.175 567.240 44.695 ;
        RECT 567.415 44.345 568.625 44.865 ;
        RECT 568.795 44.175 570.005 44.695 ;
        RECT 570.635 44.345 573.215 44.865 ;
        RECT 556.375 43.085 561.720 44.175 ;
        RECT 561.895 43.085 567.240 44.175 ;
        RECT 567.415 43.085 570.005 44.175 ;
        RECT 570.175 43.085 570.465 44.250 ;
        RECT 573.385 44.175 575.980 44.695 ;
        RECT 576.155 44.345 578.735 44.865 ;
        RECT 578.905 44.175 581.500 44.695 ;
        RECT 581.675 44.345 582.885 44.865 ;
        RECT 583.055 44.175 584.265 44.695 ;
        RECT 570.635 43.085 575.980 44.175 ;
        RECT 576.155 43.085 581.500 44.175 ;
        RECT 581.675 43.085 584.265 44.175 ;
        RECT 584.435 43.085 584.725 44.250 ;
        RECT 585.815 43.980 586.335 45.465 ;
        RECT 586.505 44.975 586.845 45.635 ;
        RECT 587.195 44.865 592.540 45.635 ;
        RECT 592.715 44.865 598.060 45.635 ;
        RECT 598.695 44.910 598.985 45.635 ;
        RECT 599.155 44.865 604.500 45.635 ;
        RECT 604.675 44.865 610.020 45.635 ;
        RECT 610.195 44.865 612.785 45.635 ;
        RECT 612.955 44.910 613.245 45.635 ;
        RECT 613.415 44.865 618.760 45.635 ;
        RECT 618.935 44.865 621.525 45.635 ;
        RECT 586.005 43.085 586.335 43.810 ;
        RECT 586.505 43.255 587.025 44.805 ;
        RECT 587.195 44.345 589.775 44.865 ;
        RECT 589.945 44.175 592.540 44.695 ;
        RECT 592.715 44.345 595.295 44.865 ;
        RECT 595.465 44.175 598.060 44.695 ;
        RECT 599.155 44.345 601.735 44.865 ;
        RECT 587.195 43.085 592.540 44.175 ;
        RECT 592.715 43.085 598.060 44.175 ;
        RECT 598.695 43.085 598.985 44.250 ;
        RECT 601.905 44.175 604.500 44.695 ;
        RECT 604.675 44.345 607.255 44.865 ;
        RECT 607.425 44.175 610.020 44.695 ;
        RECT 610.195 44.345 611.405 44.865 ;
        RECT 611.575 44.175 612.785 44.695 ;
        RECT 613.415 44.345 615.995 44.865 ;
        RECT 599.155 43.085 604.500 44.175 ;
        RECT 604.675 43.085 610.020 44.175 ;
        RECT 610.195 43.085 612.785 44.175 ;
        RECT 612.955 43.085 613.245 44.250 ;
        RECT 616.165 44.175 618.760 44.695 ;
        RECT 618.935 44.345 620.145 44.865 ;
        RECT 620.315 44.175 621.525 44.695 ;
        RECT 613.415 43.085 618.760 44.175 ;
        RECT 618.935 43.085 621.525 44.175 ;
        RECT 622.155 43.980 622.675 45.465 ;
        RECT 622.845 44.975 623.185 45.635 ;
        RECT 623.535 44.865 627.045 45.635 ;
        RECT 627.215 44.910 627.505 45.635 ;
        RECT 627.675 44.865 629.345 45.635 ;
        RECT 629.975 44.885 631.185 45.635 ;
        RECT 623.535 44.345 625.185 44.865 ;
        RECT 625.355 44.175 627.045 44.695 ;
        RECT 627.675 44.345 628.425 44.865 ;
        RECT 622.345 43.085 622.675 43.810 ;
        RECT 623.535 43.085 627.045 44.175 ;
        RECT 627.215 43.085 627.505 44.250 ;
        RECT 628.595 44.175 629.345 44.695 ;
        RECT 627.675 43.085 629.345 44.175 ;
        RECT 629.975 44.175 630.495 44.715 ;
        RECT 630.665 44.345 631.185 44.885 ;
        RECT 629.975 43.085 631.185 44.175 ;
        RECT 42.470 42.915 631.270 43.085 ;
        RECT 155.775 40.705 155.945 42.235 ;
        RECT 163.135 39.685 163.305 41.895 ;
        RECT 175.095 38.665 175.265 41.895 ;
        RECT 215.115 39.005 215.285 42.575 ;
        RECT 221.555 39.345 221.725 42.575 ;
        RECT 223.855 41.725 224.485 41.895 ;
        RECT 224.775 41.215 224.945 42.235 ;
        RECT 223.395 41.045 224.945 41.215 ;
        RECT 258.355 39.685 258.525 40.875 ;
      LAYER L1M1_PR_C ;
        RECT 42.615 53.795 42.785 53.965 ;
        RECT 43.075 53.795 43.245 53.965 ;
        RECT 43.535 53.795 43.705 53.965 ;
        RECT 43.995 53.795 44.165 53.965 ;
        RECT 44.455 53.795 44.625 53.965 ;
        RECT 44.915 53.795 45.085 53.965 ;
        RECT 45.375 53.795 45.545 53.965 ;
        RECT 45.835 53.795 46.005 53.965 ;
        RECT 46.295 53.795 46.465 53.965 ;
        RECT 46.755 53.795 46.925 53.965 ;
        RECT 47.215 53.795 47.385 53.965 ;
        RECT 47.675 53.795 47.845 53.965 ;
        RECT 48.135 53.795 48.305 53.965 ;
        RECT 48.595 53.795 48.765 53.965 ;
        RECT 49.055 53.795 49.225 53.965 ;
        RECT 49.515 53.795 49.685 53.965 ;
        RECT 49.975 53.795 50.145 53.965 ;
        RECT 50.435 53.795 50.605 53.965 ;
        RECT 50.895 53.795 51.065 53.965 ;
        RECT 51.355 53.795 51.525 53.965 ;
        RECT 51.815 53.795 51.985 53.965 ;
        RECT 52.275 53.795 52.445 53.965 ;
        RECT 52.735 53.795 52.905 53.965 ;
        RECT 53.195 53.795 53.365 53.965 ;
        RECT 53.655 53.795 53.825 53.965 ;
        RECT 54.115 53.795 54.285 53.965 ;
        RECT 54.575 53.795 54.745 53.965 ;
        RECT 55.035 53.795 55.205 53.965 ;
        RECT 55.495 53.795 55.665 53.965 ;
        RECT 55.955 53.795 56.125 53.965 ;
        RECT 56.415 53.795 56.585 53.965 ;
        RECT 56.875 53.795 57.045 53.965 ;
        RECT 57.335 53.795 57.505 53.965 ;
        RECT 57.795 53.795 57.965 53.965 ;
        RECT 58.255 53.795 58.425 53.965 ;
        RECT 58.715 53.795 58.885 53.965 ;
        RECT 59.175 53.795 59.345 53.965 ;
        RECT 59.635 53.795 59.805 53.965 ;
        RECT 60.095 53.795 60.265 53.965 ;
        RECT 60.555 53.795 60.725 53.965 ;
        RECT 61.015 53.795 61.185 53.965 ;
        RECT 61.475 53.795 61.645 53.965 ;
        RECT 61.935 53.795 62.105 53.965 ;
        RECT 62.395 53.795 62.565 53.965 ;
        RECT 62.855 53.795 63.025 53.965 ;
        RECT 63.315 53.795 63.485 53.965 ;
        RECT 63.775 53.795 63.945 53.965 ;
        RECT 64.235 53.795 64.405 53.965 ;
        RECT 64.695 53.795 64.865 53.965 ;
        RECT 65.155 53.795 65.325 53.965 ;
        RECT 65.615 53.795 65.785 53.965 ;
        RECT 66.075 53.795 66.245 53.965 ;
        RECT 66.535 53.795 66.705 53.965 ;
        RECT 66.995 53.795 67.165 53.965 ;
        RECT 67.455 53.795 67.625 53.965 ;
        RECT 67.915 53.795 68.085 53.965 ;
        RECT 68.375 53.795 68.545 53.965 ;
        RECT 68.835 53.795 69.005 53.965 ;
        RECT 69.295 53.795 69.465 53.965 ;
        RECT 69.755 53.795 69.925 53.965 ;
        RECT 70.215 53.795 70.385 53.965 ;
        RECT 70.675 53.795 70.845 53.965 ;
        RECT 71.135 53.795 71.305 53.965 ;
        RECT 71.595 53.795 71.765 53.965 ;
        RECT 72.055 53.795 72.225 53.965 ;
        RECT 72.515 53.795 72.685 53.965 ;
        RECT 72.975 53.795 73.145 53.965 ;
        RECT 73.435 53.795 73.605 53.965 ;
        RECT 73.895 53.795 74.065 53.965 ;
        RECT 74.355 53.795 74.525 53.965 ;
        RECT 74.815 53.795 74.985 53.965 ;
        RECT 75.275 53.795 75.445 53.965 ;
        RECT 75.735 53.795 75.905 53.965 ;
        RECT 76.195 53.795 76.365 53.965 ;
        RECT 76.655 53.795 76.825 53.965 ;
        RECT 77.115 53.795 77.285 53.965 ;
        RECT 77.575 53.795 77.745 53.965 ;
        RECT 78.035 53.795 78.205 53.965 ;
        RECT 78.495 53.795 78.665 53.965 ;
        RECT 78.955 53.795 79.125 53.965 ;
        RECT 79.415 53.795 79.585 53.965 ;
        RECT 79.875 53.795 80.045 53.965 ;
        RECT 80.335 53.795 80.505 53.965 ;
        RECT 80.795 53.795 80.965 53.965 ;
        RECT 81.255 53.795 81.425 53.965 ;
        RECT 81.715 53.795 81.885 53.965 ;
        RECT 82.175 53.795 82.345 53.965 ;
        RECT 82.635 53.795 82.805 53.965 ;
        RECT 83.095 53.795 83.265 53.965 ;
        RECT 83.555 53.795 83.725 53.965 ;
        RECT 84.015 53.795 84.185 53.965 ;
        RECT 84.475 53.795 84.645 53.965 ;
        RECT 84.935 53.795 85.105 53.965 ;
        RECT 85.395 53.795 85.565 53.965 ;
        RECT 85.855 53.795 86.025 53.965 ;
        RECT 86.315 53.795 86.485 53.965 ;
        RECT 86.775 53.795 86.945 53.965 ;
        RECT 87.235 53.795 87.405 53.965 ;
        RECT 87.695 53.795 87.865 53.965 ;
        RECT 88.155 53.795 88.325 53.965 ;
        RECT 88.615 53.795 88.785 53.965 ;
        RECT 89.075 53.795 89.245 53.965 ;
        RECT 89.535 53.795 89.705 53.965 ;
        RECT 89.995 53.795 90.165 53.965 ;
        RECT 90.455 53.795 90.625 53.965 ;
        RECT 90.915 53.795 91.085 53.965 ;
        RECT 91.375 53.795 91.545 53.965 ;
        RECT 91.835 53.795 92.005 53.965 ;
        RECT 92.295 53.795 92.465 53.965 ;
        RECT 92.755 53.795 92.925 53.965 ;
        RECT 93.215 53.795 93.385 53.965 ;
        RECT 93.675 53.795 93.845 53.965 ;
        RECT 94.135 53.795 94.305 53.965 ;
        RECT 94.595 53.795 94.765 53.965 ;
        RECT 95.055 53.795 95.225 53.965 ;
        RECT 95.515 53.795 95.685 53.965 ;
        RECT 95.975 53.795 96.145 53.965 ;
        RECT 96.435 53.795 96.605 53.965 ;
        RECT 96.895 53.795 97.065 53.965 ;
        RECT 97.355 53.795 97.525 53.965 ;
        RECT 97.815 53.795 97.985 53.965 ;
        RECT 98.275 53.795 98.445 53.965 ;
        RECT 98.735 53.795 98.905 53.965 ;
        RECT 99.195 53.795 99.365 53.965 ;
        RECT 99.655 53.795 99.825 53.965 ;
        RECT 100.115 53.795 100.285 53.965 ;
        RECT 100.575 53.795 100.745 53.965 ;
        RECT 101.035 53.795 101.205 53.965 ;
        RECT 101.495 53.795 101.665 53.965 ;
        RECT 101.955 53.795 102.125 53.965 ;
        RECT 102.415 53.795 102.585 53.965 ;
        RECT 102.875 53.795 103.045 53.965 ;
        RECT 103.335 53.795 103.505 53.965 ;
        RECT 103.795 53.795 103.965 53.965 ;
        RECT 104.255 53.795 104.425 53.965 ;
        RECT 104.715 53.795 104.885 53.965 ;
        RECT 105.175 53.795 105.345 53.965 ;
        RECT 105.635 53.795 105.805 53.965 ;
        RECT 106.095 53.795 106.265 53.965 ;
        RECT 106.555 53.795 106.725 53.965 ;
        RECT 107.015 53.795 107.185 53.965 ;
        RECT 107.475 53.795 107.645 53.965 ;
        RECT 107.935 53.795 108.105 53.965 ;
        RECT 108.395 53.795 108.565 53.965 ;
        RECT 108.855 53.795 109.025 53.965 ;
        RECT 109.315 53.795 109.485 53.965 ;
        RECT 109.775 53.795 109.945 53.965 ;
        RECT 110.235 53.795 110.405 53.965 ;
        RECT 110.695 53.795 110.865 53.965 ;
        RECT 111.155 53.795 111.325 53.965 ;
        RECT 111.615 53.795 111.785 53.965 ;
        RECT 112.075 53.795 112.245 53.965 ;
        RECT 112.535 53.795 112.705 53.965 ;
        RECT 112.995 53.795 113.165 53.965 ;
        RECT 113.455 53.795 113.625 53.965 ;
        RECT 113.915 53.795 114.085 53.965 ;
        RECT 114.375 53.795 114.545 53.965 ;
        RECT 114.835 53.795 115.005 53.965 ;
        RECT 115.295 53.795 115.465 53.965 ;
        RECT 115.755 53.795 115.925 53.965 ;
        RECT 116.215 53.795 116.385 53.965 ;
        RECT 116.675 53.795 116.845 53.965 ;
        RECT 117.135 53.795 117.305 53.965 ;
        RECT 117.595 53.795 117.765 53.965 ;
        RECT 118.055 53.795 118.225 53.965 ;
        RECT 118.515 53.795 118.685 53.965 ;
        RECT 118.975 53.795 119.145 53.965 ;
        RECT 119.435 53.795 119.605 53.965 ;
        RECT 119.895 53.795 120.065 53.965 ;
        RECT 120.355 53.795 120.525 53.965 ;
        RECT 120.815 53.795 120.985 53.965 ;
        RECT 121.275 53.795 121.445 53.965 ;
        RECT 121.735 53.795 121.905 53.965 ;
        RECT 122.195 53.795 122.365 53.965 ;
        RECT 122.655 53.795 122.825 53.965 ;
        RECT 123.115 53.795 123.285 53.965 ;
        RECT 123.575 53.795 123.745 53.965 ;
        RECT 124.035 53.795 124.205 53.965 ;
        RECT 124.495 53.795 124.665 53.965 ;
        RECT 124.955 53.795 125.125 53.965 ;
        RECT 125.415 53.795 125.585 53.965 ;
        RECT 125.875 53.795 126.045 53.965 ;
        RECT 126.335 53.795 126.505 53.965 ;
        RECT 126.795 53.795 126.965 53.965 ;
        RECT 127.255 53.795 127.425 53.965 ;
        RECT 127.715 53.795 127.885 53.965 ;
        RECT 128.175 53.795 128.345 53.965 ;
        RECT 128.635 53.795 128.805 53.965 ;
        RECT 129.095 53.795 129.265 53.965 ;
        RECT 129.555 53.795 129.725 53.965 ;
        RECT 130.015 53.795 130.185 53.965 ;
        RECT 130.475 53.795 130.645 53.965 ;
        RECT 130.935 53.795 131.105 53.965 ;
        RECT 131.395 53.795 131.565 53.965 ;
        RECT 131.855 53.795 132.025 53.965 ;
        RECT 132.315 53.795 132.485 53.965 ;
        RECT 132.775 53.795 132.945 53.965 ;
        RECT 133.235 53.795 133.405 53.965 ;
        RECT 133.695 53.795 133.865 53.965 ;
        RECT 134.155 53.795 134.325 53.965 ;
        RECT 134.615 53.795 134.785 53.965 ;
        RECT 135.075 53.795 135.245 53.965 ;
        RECT 135.535 53.795 135.705 53.965 ;
        RECT 135.995 53.795 136.165 53.965 ;
        RECT 136.455 53.795 136.625 53.965 ;
        RECT 136.915 53.795 137.085 53.965 ;
        RECT 137.375 53.795 137.545 53.965 ;
        RECT 137.835 53.795 138.005 53.965 ;
        RECT 138.295 53.795 138.465 53.965 ;
        RECT 138.755 53.795 138.925 53.965 ;
        RECT 139.215 53.795 139.385 53.965 ;
        RECT 139.675 53.795 139.845 53.965 ;
        RECT 140.135 53.795 140.305 53.965 ;
        RECT 140.595 53.795 140.765 53.965 ;
        RECT 141.055 53.795 141.225 53.965 ;
        RECT 141.515 53.795 141.685 53.965 ;
        RECT 141.975 53.795 142.145 53.965 ;
        RECT 142.435 53.795 142.605 53.965 ;
        RECT 142.895 53.795 143.065 53.965 ;
        RECT 143.355 53.795 143.525 53.965 ;
        RECT 143.815 53.795 143.985 53.965 ;
        RECT 144.275 53.795 144.445 53.965 ;
        RECT 144.735 53.795 144.905 53.965 ;
        RECT 145.195 53.795 145.365 53.965 ;
        RECT 145.655 53.795 145.825 53.965 ;
        RECT 146.115 53.795 146.285 53.965 ;
        RECT 146.575 53.795 146.745 53.965 ;
        RECT 147.035 53.795 147.205 53.965 ;
        RECT 147.495 53.795 147.665 53.965 ;
        RECT 147.955 53.795 148.125 53.965 ;
        RECT 148.415 53.795 148.585 53.965 ;
        RECT 148.875 53.795 149.045 53.965 ;
        RECT 149.335 53.795 149.505 53.965 ;
        RECT 149.795 53.795 149.965 53.965 ;
        RECT 150.255 53.795 150.425 53.965 ;
        RECT 150.715 53.795 150.885 53.965 ;
        RECT 151.175 53.795 151.345 53.965 ;
        RECT 151.635 53.795 151.805 53.965 ;
        RECT 152.095 53.795 152.265 53.965 ;
        RECT 152.555 53.795 152.725 53.965 ;
        RECT 153.015 53.795 153.185 53.965 ;
        RECT 153.475 53.795 153.645 53.965 ;
        RECT 153.935 53.795 154.105 53.965 ;
        RECT 154.395 53.795 154.565 53.965 ;
        RECT 154.855 53.795 155.025 53.965 ;
        RECT 155.315 53.795 155.485 53.965 ;
        RECT 155.775 53.795 155.945 53.965 ;
        RECT 156.235 53.795 156.405 53.965 ;
        RECT 156.695 53.795 156.865 53.965 ;
        RECT 157.155 53.795 157.325 53.965 ;
        RECT 157.615 53.795 157.785 53.965 ;
        RECT 158.075 53.795 158.245 53.965 ;
        RECT 158.535 53.795 158.705 53.965 ;
        RECT 158.995 53.795 159.165 53.965 ;
        RECT 159.455 53.795 159.625 53.965 ;
        RECT 159.915 53.795 160.085 53.965 ;
        RECT 160.375 53.795 160.545 53.965 ;
        RECT 160.835 53.795 161.005 53.965 ;
        RECT 161.295 53.795 161.465 53.965 ;
        RECT 161.755 53.795 161.925 53.965 ;
        RECT 162.215 53.795 162.385 53.965 ;
        RECT 162.675 53.795 162.845 53.965 ;
        RECT 163.135 53.795 163.305 53.965 ;
        RECT 163.595 53.795 163.765 53.965 ;
        RECT 164.055 53.795 164.225 53.965 ;
        RECT 164.515 53.795 164.685 53.965 ;
        RECT 164.975 53.795 165.145 53.965 ;
        RECT 165.435 53.795 165.605 53.965 ;
        RECT 165.895 53.795 166.065 53.965 ;
        RECT 166.355 53.795 166.525 53.965 ;
        RECT 166.815 53.795 166.985 53.965 ;
        RECT 167.275 53.795 167.445 53.965 ;
        RECT 167.735 53.795 167.905 53.965 ;
        RECT 168.195 53.795 168.365 53.965 ;
        RECT 168.655 53.795 168.825 53.965 ;
        RECT 169.115 53.795 169.285 53.965 ;
        RECT 169.575 53.795 169.745 53.965 ;
        RECT 170.035 53.795 170.205 53.965 ;
        RECT 170.495 53.795 170.665 53.965 ;
        RECT 170.955 53.795 171.125 53.965 ;
        RECT 171.415 53.795 171.585 53.965 ;
        RECT 171.875 53.795 172.045 53.965 ;
        RECT 172.335 53.795 172.505 53.965 ;
        RECT 172.795 53.795 172.965 53.965 ;
        RECT 173.255 53.795 173.425 53.965 ;
        RECT 173.715 53.795 173.885 53.965 ;
        RECT 174.175 53.795 174.345 53.965 ;
        RECT 174.635 53.795 174.805 53.965 ;
        RECT 175.095 53.795 175.265 53.965 ;
        RECT 175.555 53.795 175.725 53.965 ;
        RECT 176.015 53.795 176.185 53.965 ;
        RECT 176.475 53.795 176.645 53.965 ;
        RECT 176.935 53.795 177.105 53.965 ;
        RECT 177.395 53.795 177.565 53.965 ;
        RECT 177.855 53.795 178.025 53.965 ;
        RECT 178.315 53.795 178.485 53.965 ;
        RECT 178.775 53.795 178.945 53.965 ;
        RECT 179.235 53.795 179.405 53.965 ;
        RECT 179.695 53.795 179.865 53.965 ;
        RECT 180.155 53.795 180.325 53.965 ;
        RECT 180.615 53.795 180.785 53.965 ;
        RECT 181.075 53.795 181.245 53.965 ;
        RECT 181.535 53.795 181.705 53.965 ;
        RECT 181.995 53.795 182.165 53.965 ;
        RECT 182.455 53.795 182.625 53.965 ;
        RECT 182.915 53.795 183.085 53.965 ;
        RECT 183.375 53.795 183.545 53.965 ;
        RECT 183.835 53.795 184.005 53.965 ;
        RECT 184.295 53.795 184.465 53.965 ;
        RECT 184.755 53.795 184.925 53.965 ;
        RECT 185.215 53.795 185.385 53.965 ;
        RECT 185.675 53.795 185.845 53.965 ;
        RECT 186.135 53.795 186.305 53.965 ;
        RECT 186.595 53.795 186.765 53.965 ;
        RECT 187.055 53.795 187.225 53.965 ;
        RECT 187.515 53.795 187.685 53.965 ;
        RECT 187.975 53.795 188.145 53.965 ;
        RECT 188.435 53.795 188.605 53.965 ;
        RECT 188.895 53.795 189.065 53.965 ;
        RECT 189.355 53.795 189.525 53.965 ;
        RECT 189.815 53.795 189.985 53.965 ;
        RECT 190.275 53.795 190.445 53.965 ;
        RECT 190.735 53.795 190.905 53.965 ;
        RECT 191.195 53.795 191.365 53.965 ;
        RECT 191.655 53.795 191.825 53.965 ;
        RECT 192.115 53.795 192.285 53.965 ;
        RECT 192.575 53.795 192.745 53.965 ;
        RECT 193.035 53.795 193.205 53.965 ;
        RECT 193.495 53.795 193.665 53.965 ;
        RECT 193.955 53.795 194.125 53.965 ;
        RECT 194.415 53.795 194.585 53.965 ;
        RECT 194.875 53.795 195.045 53.965 ;
        RECT 195.335 53.795 195.505 53.965 ;
        RECT 195.795 53.795 195.965 53.965 ;
        RECT 196.255 53.795 196.425 53.965 ;
        RECT 196.715 53.795 196.885 53.965 ;
        RECT 197.175 53.795 197.345 53.965 ;
        RECT 197.635 53.795 197.805 53.965 ;
        RECT 198.095 53.795 198.265 53.965 ;
        RECT 198.555 53.795 198.725 53.965 ;
        RECT 199.015 53.795 199.185 53.965 ;
        RECT 199.475 53.795 199.645 53.965 ;
        RECT 199.935 53.795 200.105 53.965 ;
        RECT 200.395 53.795 200.565 53.965 ;
        RECT 200.855 53.795 201.025 53.965 ;
        RECT 201.315 53.795 201.485 53.965 ;
        RECT 201.775 53.795 201.945 53.965 ;
        RECT 202.235 53.795 202.405 53.965 ;
        RECT 202.695 53.795 202.865 53.965 ;
        RECT 203.155 53.795 203.325 53.965 ;
        RECT 203.615 53.795 203.785 53.965 ;
        RECT 204.075 53.795 204.245 53.965 ;
        RECT 204.535 53.795 204.705 53.965 ;
        RECT 204.995 53.795 205.165 53.965 ;
        RECT 205.455 53.795 205.625 53.965 ;
        RECT 205.915 53.795 206.085 53.965 ;
        RECT 206.375 53.795 206.545 53.965 ;
        RECT 206.835 53.795 207.005 53.965 ;
        RECT 207.295 53.795 207.465 53.965 ;
        RECT 207.755 53.795 207.925 53.965 ;
        RECT 208.215 53.795 208.385 53.965 ;
        RECT 208.675 53.795 208.845 53.965 ;
        RECT 209.135 53.795 209.305 53.965 ;
        RECT 209.595 53.795 209.765 53.965 ;
        RECT 210.055 53.795 210.225 53.965 ;
        RECT 210.515 53.795 210.685 53.965 ;
        RECT 210.975 53.795 211.145 53.965 ;
        RECT 211.435 53.795 211.605 53.965 ;
        RECT 211.895 53.795 212.065 53.965 ;
        RECT 212.355 53.795 212.525 53.965 ;
        RECT 212.815 53.795 212.985 53.965 ;
        RECT 213.275 53.795 213.445 53.965 ;
        RECT 213.735 53.795 213.905 53.965 ;
        RECT 214.195 53.795 214.365 53.965 ;
        RECT 214.655 53.795 214.825 53.965 ;
        RECT 215.115 53.795 215.285 53.965 ;
        RECT 215.575 53.795 215.745 53.965 ;
        RECT 216.035 53.795 216.205 53.965 ;
        RECT 216.495 53.795 216.665 53.965 ;
        RECT 216.955 53.795 217.125 53.965 ;
        RECT 217.415 53.795 217.585 53.965 ;
        RECT 217.875 53.795 218.045 53.965 ;
        RECT 218.335 53.795 218.505 53.965 ;
        RECT 218.795 53.795 218.965 53.965 ;
        RECT 219.255 53.795 219.425 53.965 ;
        RECT 219.715 53.795 219.885 53.965 ;
        RECT 220.175 53.795 220.345 53.965 ;
        RECT 220.635 53.795 220.805 53.965 ;
        RECT 221.095 53.795 221.265 53.965 ;
        RECT 221.555 53.795 221.725 53.965 ;
        RECT 222.015 53.795 222.185 53.965 ;
        RECT 222.475 53.795 222.645 53.965 ;
        RECT 222.935 53.795 223.105 53.965 ;
        RECT 223.395 53.795 223.565 53.965 ;
        RECT 223.855 53.795 224.025 53.965 ;
        RECT 224.315 53.795 224.485 53.965 ;
        RECT 224.775 53.795 224.945 53.965 ;
        RECT 225.235 53.795 225.405 53.965 ;
        RECT 225.695 53.795 225.865 53.965 ;
        RECT 226.155 53.795 226.325 53.965 ;
        RECT 226.615 53.795 226.785 53.965 ;
        RECT 227.075 53.795 227.245 53.965 ;
        RECT 227.535 53.795 227.705 53.965 ;
        RECT 227.995 53.795 228.165 53.965 ;
        RECT 228.455 53.795 228.625 53.965 ;
        RECT 228.915 53.795 229.085 53.965 ;
        RECT 229.375 53.795 229.545 53.965 ;
        RECT 229.835 53.795 230.005 53.965 ;
        RECT 230.295 53.795 230.465 53.965 ;
        RECT 230.755 53.795 230.925 53.965 ;
        RECT 231.215 53.795 231.385 53.965 ;
        RECT 231.675 53.795 231.845 53.965 ;
        RECT 232.135 53.795 232.305 53.965 ;
        RECT 232.595 53.795 232.765 53.965 ;
        RECT 233.055 53.795 233.225 53.965 ;
        RECT 233.515 53.795 233.685 53.965 ;
        RECT 233.975 53.795 234.145 53.965 ;
        RECT 234.435 53.795 234.605 53.965 ;
        RECT 234.895 53.795 235.065 53.965 ;
        RECT 235.355 53.795 235.525 53.965 ;
        RECT 235.815 53.795 235.985 53.965 ;
        RECT 236.275 53.795 236.445 53.965 ;
        RECT 236.735 53.795 236.905 53.965 ;
        RECT 237.195 53.795 237.365 53.965 ;
        RECT 237.655 53.795 237.825 53.965 ;
        RECT 238.115 53.795 238.285 53.965 ;
        RECT 238.575 53.795 238.745 53.965 ;
        RECT 239.035 53.795 239.205 53.965 ;
        RECT 239.495 53.795 239.665 53.965 ;
        RECT 239.955 53.795 240.125 53.965 ;
        RECT 240.415 53.795 240.585 53.965 ;
        RECT 240.875 53.795 241.045 53.965 ;
        RECT 241.335 53.795 241.505 53.965 ;
        RECT 241.795 53.795 241.965 53.965 ;
        RECT 242.255 53.795 242.425 53.965 ;
        RECT 242.715 53.795 242.885 53.965 ;
        RECT 243.175 53.795 243.345 53.965 ;
        RECT 243.635 53.795 243.805 53.965 ;
        RECT 244.095 53.795 244.265 53.965 ;
        RECT 244.555 53.795 244.725 53.965 ;
        RECT 245.015 53.795 245.185 53.965 ;
        RECT 245.475 53.795 245.645 53.965 ;
        RECT 245.935 53.795 246.105 53.965 ;
        RECT 246.395 53.795 246.565 53.965 ;
        RECT 246.855 53.795 247.025 53.965 ;
        RECT 247.315 53.795 247.485 53.965 ;
        RECT 247.775 53.795 247.945 53.965 ;
        RECT 248.235 53.795 248.405 53.965 ;
        RECT 248.695 53.795 248.865 53.965 ;
        RECT 249.155 53.795 249.325 53.965 ;
        RECT 249.615 53.795 249.785 53.965 ;
        RECT 250.075 53.795 250.245 53.965 ;
        RECT 250.535 53.795 250.705 53.965 ;
        RECT 250.995 53.795 251.165 53.965 ;
        RECT 251.455 53.795 251.625 53.965 ;
        RECT 251.915 53.795 252.085 53.965 ;
        RECT 252.375 53.795 252.545 53.965 ;
        RECT 252.835 53.795 253.005 53.965 ;
        RECT 253.295 53.795 253.465 53.965 ;
        RECT 253.755 53.795 253.925 53.965 ;
        RECT 254.215 53.795 254.385 53.965 ;
        RECT 254.675 53.795 254.845 53.965 ;
        RECT 255.135 53.795 255.305 53.965 ;
        RECT 255.595 53.795 255.765 53.965 ;
        RECT 256.055 53.795 256.225 53.965 ;
        RECT 256.515 53.795 256.685 53.965 ;
        RECT 256.975 53.795 257.145 53.965 ;
        RECT 257.435 53.795 257.605 53.965 ;
        RECT 257.895 53.795 258.065 53.965 ;
        RECT 258.355 53.795 258.525 53.965 ;
        RECT 258.815 53.795 258.985 53.965 ;
        RECT 259.275 53.795 259.445 53.965 ;
        RECT 259.735 53.795 259.905 53.965 ;
        RECT 260.195 53.795 260.365 53.965 ;
        RECT 260.655 53.795 260.825 53.965 ;
        RECT 261.115 53.795 261.285 53.965 ;
        RECT 261.575 53.795 261.745 53.965 ;
        RECT 262.035 53.795 262.205 53.965 ;
        RECT 262.495 53.795 262.665 53.965 ;
        RECT 262.955 53.795 263.125 53.965 ;
        RECT 263.415 53.795 263.585 53.965 ;
        RECT 263.875 53.795 264.045 53.965 ;
        RECT 264.335 53.795 264.505 53.965 ;
        RECT 264.795 53.795 264.965 53.965 ;
        RECT 265.255 53.795 265.425 53.965 ;
        RECT 265.715 53.795 265.885 53.965 ;
        RECT 266.175 53.795 266.345 53.965 ;
        RECT 266.635 53.795 266.805 53.965 ;
        RECT 267.095 53.795 267.265 53.965 ;
        RECT 267.555 53.795 267.725 53.965 ;
        RECT 268.015 53.795 268.185 53.965 ;
        RECT 268.475 53.795 268.645 53.965 ;
        RECT 268.935 53.795 269.105 53.965 ;
        RECT 269.395 53.795 269.565 53.965 ;
        RECT 269.855 53.795 270.025 53.965 ;
        RECT 270.315 53.795 270.485 53.965 ;
        RECT 270.775 53.795 270.945 53.965 ;
        RECT 271.235 53.795 271.405 53.965 ;
        RECT 271.695 53.795 271.865 53.965 ;
        RECT 272.155 53.795 272.325 53.965 ;
        RECT 272.615 53.795 272.785 53.965 ;
        RECT 273.075 53.795 273.245 53.965 ;
        RECT 273.535 53.795 273.705 53.965 ;
        RECT 273.995 53.795 274.165 53.965 ;
        RECT 274.455 53.795 274.625 53.965 ;
        RECT 274.915 53.795 275.085 53.965 ;
        RECT 275.375 53.795 275.545 53.965 ;
        RECT 275.835 53.795 276.005 53.965 ;
        RECT 276.295 53.795 276.465 53.965 ;
        RECT 276.755 53.795 276.925 53.965 ;
        RECT 277.215 53.795 277.385 53.965 ;
        RECT 277.675 53.795 277.845 53.965 ;
        RECT 278.135 53.795 278.305 53.965 ;
        RECT 278.595 53.795 278.765 53.965 ;
        RECT 279.055 53.795 279.225 53.965 ;
        RECT 279.515 53.795 279.685 53.965 ;
        RECT 279.975 53.795 280.145 53.965 ;
        RECT 280.435 53.795 280.605 53.965 ;
        RECT 280.895 53.795 281.065 53.965 ;
        RECT 281.355 53.795 281.525 53.965 ;
        RECT 281.815 53.795 281.985 53.965 ;
        RECT 282.275 53.795 282.445 53.965 ;
        RECT 282.735 53.795 282.905 53.965 ;
        RECT 283.195 53.795 283.365 53.965 ;
        RECT 283.655 53.795 283.825 53.965 ;
        RECT 284.115 53.795 284.285 53.965 ;
        RECT 284.575 53.795 284.745 53.965 ;
        RECT 285.035 53.795 285.205 53.965 ;
        RECT 285.495 53.795 285.665 53.965 ;
        RECT 285.955 53.795 286.125 53.965 ;
        RECT 286.415 53.795 286.585 53.965 ;
        RECT 286.875 53.795 287.045 53.965 ;
        RECT 287.335 53.795 287.505 53.965 ;
        RECT 287.795 53.795 287.965 53.965 ;
        RECT 288.255 53.795 288.425 53.965 ;
        RECT 288.715 53.795 288.885 53.965 ;
        RECT 289.175 53.795 289.345 53.965 ;
        RECT 289.635 53.795 289.805 53.965 ;
        RECT 290.095 53.795 290.265 53.965 ;
        RECT 290.555 53.795 290.725 53.965 ;
        RECT 291.015 53.795 291.185 53.965 ;
        RECT 291.475 53.795 291.645 53.965 ;
        RECT 291.935 53.795 292.105 53.965 ;
        RECT 292.395 53.795 292.565 53.965 ;
        RECT 292.855 53.795 293.025 53.965 ;
        RECT 293.315 53.795 293.485 53.965 ;
        RECT 293.775 53.795 293.945 53.965 ;
        RECT 294.235 53.795 294.405 53.965 ;
        RECT 294.695 53.795 294.865 53.965 ;
        RECT 295.155 53.795 295.325 53.965 ;
        RECT 295.615 53.795 295.785 53.965 ;
        RECT 296.075 53.795 296.245 53.965 ;
        RECT 296.535 53.795 296.705 53.965 ;
        RECT 296.995 53.795 297.165 53.965 ;
        RECT 297.455 53.795 297.625 53.965 ;
        RECT 297.915 53.795 298.085 53.965 ;
        RECT 298.375 53.795 298.545 53.965 ;
        RECT 298.835 53.795 299.005 53.965 ;
        RECT 299.295 53.795 299.465 53.965 ;
        RECT 299.755 53.795 299.925 53.965 ;
        RECT 300.215 53.795 300.385 53.965 ;
        RECT 300.675 53.795 300.845 53.965 ;
        RECT 301.135 53.795 301.305 53.965 ;
        RECT 301.595 53.795 301.765 53.965 ;
        RECT 302.055 53.795 302.225 53.965 ;
        RECT 302.515 53.795 302.685 53.965 ;
        RECT 302.975 53.795 303.145 53.965 ;
        RECT 303.435 53.795 303.605 53.965 ;
        RECT 303.895 53.795 304.065 53.965 ;
        RECT 304.355 53.795 304.525 53.965 ;
        RECT 304.815 53.795 304.985 53.965 ;
        RECT 305.275 53.795 305.445 53.965 ;
        RECT 305.735 53.795 305.905 53.965 ;
        RECT 306.195 53.795 306.365 53.965 ;
        RECT 306.655 53.795 306.825 53.965 ;
        RECT 307.115 53.795 307.285 53.965 ;
        RECT 307.575 53.795 307.745 53.965 ;
        RECT 308.035 53.795 308.205 53.965 ;
        RECT 308.495 53.795 308.665 53.965 ;
        RECT 308.955 53.795 309.125 53.965 ;
        RECT 309.415 53.795 309.585 53.965 ;
        RECT 309.875 53.795 310.045 53.965 ;
        RECT 310.335 53.795 310.505 53.965 ;
        RECT 310.795 53.795 310.965 53.965 ;
        RECT 311.255 53.795 311.425 53.965 ;
        RECT 311.715 53.795 311.885 53.965 ;
        RECT 312.175 53.795 312.345 53.965 ;
        RECT 312.635 53.795 312.805 53.965 ;
        RECT 313.095 53.795 313.265 53.965 ;
        RECT 313.555 53.795 313.725 53.965 ;
        RECT 314.015 53.795 314.185 53.965 ;
        RECT 314.475 53.795 314.645 53.965 ;
        RECT 314.935 53.795 315.105 53.965 ;
        RECT 315.395 53.795 315.565 53.965 ;
        RECT 315.855 53.795 316.025 53.965 ;
        RECT 316.315 53.795 316.485 53.965 ;
        RECT 316.775 53.795 316.945 53.965 ;
        RECT 317.235 53.795 317.405 53.965 ;
        RECT 317.695 53.795 317.865 53.965 ;
        RECT 318.155 53.795 318.325 53.965 ;
        RECT 318.615 53.795 318.785 53.965 ;
        RECT 319.075 53.795 319.245 53.965 ;
        RECT 319.535 53.795 319.705 53.965 ;
        RECT 319.995 53.795 320.165 53.965 ;
        RECT 320.455 53.795 320.625 53.965 ;
        RECT 320.915 53.795 321.085 53.965 ;
        RECT 321.375 53.795 321.545 53.965 ;
        RECT 321.835 53.795 322.005 53.965 ;
        RECT 322.295 53.795 322.465 53.965 ;
        RECT 322.755 53.795 322.925 53.965 ;
        RECT 323.215 53.795 323.385 53.965 ;
        RECT 323.675 53.795 323.845 53.965 ;
        RECT 324.135 53.795 324.305 53.965 ;
        RECT 324.595 53.795 324.765 53.965 ;
        RECT 325.055 53.795 325.225 53.965 ;
        RECT 325.515 53.795 325.685 53.965 ;
        RECT 325.975 53.795 326.145 53.965 ;
        RECT 326.435 53.795 326.605 53.965 ;
        RECT 326.895 53.795 327.065 53.965 ;
        RECT 327.355 53.795 327.525 53.965 ;
        RECT 327.815 53.795 327.985 53.965 ;
        RECT 328.275 53.795 328.445 53.965 ;
        RECT 328.735 53.795 328.905 53.965 ;
        RECT 329.195 53.795 329.365 53.965 ;
        RECT 329.655 53.795 329.825 53.965 ;
        RECT 330.115 53.795 330.285 53.965 ;
        RECT 330.575 53.795 330.745 53.965 ;
        RECT 331.035 53.795 331.205 53.965 ;
        RECT 331.495 53.795 331.665 53.965 ;
        RECT 331.955 53.795 332.125 53.965 ;
        RECT 332.415 53.795 332.585 53.965 ;
        RECT 332.875 53.795 333.045 53.965 ;
        RECT 333.335 53.795 333.505 53.965 ;
        RECT 333.795 53.795 333.965 53.965 ;
        RECT 334.255 53.795 334.425 53.965 ;
        RECT 334.715 53.795 334.885 53.965 ;
        RECT 335.175 53.795 335.345 53.965 ;
        RECT 335.635 53.795 335.805 53.965 ;
        RECT 336.095 53.795 336.265 53.965 ;
        RECT 336.555 53.795 336.725 53.965 ;
        RECT 337.015 53.795 337.185 53.965 ;
        RECT 337.475 53.795 337.645 53.965 ;
        RECT 337.935 53.795 338.105 53.965 ;
        RECT 338.395 53.795 338.565 53.965 ;
        RECT 338.855 53.795 339.025 53.965 ;
        RECT 339.315 53.795 339.485 53.965 ;
        RECT 339.775 53.795 339.945 53.965 ;
        RECT 340.235 53.795 340.405 53.965 ;
        RECT 340.695 53.795 340.865 53.965 ;
        RECT 341.155 53.795 341.325 53.965 ;
        RECT 341.615 53.795 341.785 53.965 ;
        RECT 342.075 53.795 342.245 53.965 ;
        RECT 342.535 53.795 342.705 53.965 ;
        RECT 342.995 53.795 343.165 53.965 ;
        RECT 343.455 53.795 343.625 53.965 ;
        RECT 343.915 53.795 344.085 53.965 ;
        RECT 344.375 53.795 344.545 53.965 ;
        RECT 344.835 53.795 345.005 53.965 ;
        RECT 345.295 53.795 345.465 53.965 ;
        RECT 345.755 53.795 345.925 53.965 ;
        RECT 346.215 53.795 346.385 53.965 ;
        RECT 346.675 53.795 346.845 53.965 ;
        RECT 347.135 53.795 347.305 53.965 ;
        RECT 347.595 53.795 347.765 53.965 ;
        RECT 348.055 53.795 348.225 53.965 ;
        RECT 348.515 53.795 348.685 53.965 ;
        RECT 348.975 53.795 349.145 53.965 ;
        RECT 349.435 53.795 349.605 53.965 ;
        RECT 349.895 53.795 350.065 53.965 ;
        RECT 350.355 53.795 350.525 53.965 ;
        RECT 350.815 53.795 350.985 53.965 ;
        RECT 351.275 53.795 351.445 53.965 ;
        RECT 351.735 53.795 351.905 53.965 ;
        RECT 352.195 53.795 352.365 53.965 ;
        RECT 352.655 53.795 352.825 53.965 ;
        RECT 353.115 53.795 353.285 53.965 ;
        RECT 353.575 53.795 353.745 53.965 ;
        RECT 354.035 53.795 354.205 53.965 ;
        RECT 354.495 53.795 354.665 53.965 ;
        RECT 354.955 53.795 355.125 53.965 ;
        RECT 355.415 53.795 355.585 53.965 ;
        RECT 355.875 53.795 356.045 53.965 ;
        RECT 356.335 53.795 356.505 53.965 ;
        RECT 356.795 53.795 356.965 53.965 ;
        RECT 357.255 53.795 357.425 53.965 ;
        RECT 357.715 53.795 357.885 53.965 ;
        RECT 358.175 53.795 358.345 53.965 ;
        RECT 358.635 53.795 358.805 53.965 ;
        RECT 359.095 53.795 359.265 53.965 ;
        RECT 359.555 53.795 359.725 53.965 ;
        RECT 360.015 53.795 360.185 53.965 ;
        RECT 360.475 53.795 360.645 53.965 ;
        RECT 360.935 53.795 361.105 53.965 ;
        RECT 361.395 53.795 361.565 53.965 ;
        RECT 361.855 53.795 362.025 53.965 ;
        RECT 362.315 53.795 362.485 53.965 ;
        RECT 362.775 53.795 362.945 53.965 ;
        RECT 363.235 53.795 363.405 53.965 ;
        RECT 363.695 53.795 363.865 53.965 ;
        RECT 364.155 53.795 364.325 53.965 ;
        RECT 364.615 53.795 364.785 53.965 ;
        RECT 365.075 53.795 365.245 53.965 ;
        RECT 365.535 53.795 365.705 53.965 ;
        RECT 365.995 53.795 366.165 53.965 ;
        RECT 366.455 53.795 366.625 53.965 ;
        RECT 366.915 53.795 367.085 53.965 ;
        RECT 367.375 53.795 367.545 53.965 ;
        RECT 367.835 53.795 368.005 53.965 ;
        RECT 368.295 53.795 368.465 53.965 ;
        RECT 368.755 53.795 368.925 53.965 ;
        RECT 369.215 53.795 369.385 53.965 ;
        RECT 369.675 53.795 369.845 53.965 ;
        RECT 370.135 53.795 370.305 53.965 ;
        RECT 370.595 53.795 370.765 53.965 ;
        RECT 371.055 53.795 371.225 53.965 ;
        RECT 371.515 53.795 371.685 53.965 ;
        RECT 371.975 53.795 372.145 53.965 ;
        RECT 372.435 53.795 372.605 53.965 ;
        RECT 372.895 53.795 373.065 53.965 ;
        RECT 373.355 53.795 373.525 53.965 ;
        RECT 373.815 53.795 373.985 53.965 ;
        RECT 374.275 53.795 374.445 53.965 ;
        RECT 374.735 53.795 374.905 53.965 ;
        RECT 375.195 53.795 375.365 53.965 ;
        RECT 375.655 53.795 375.825 53.965 ;
        RECT 376.115 53.795 376.285 53.965 ;
        RECT 376.575 53.795 376.745 53.965 ;
        RECT 377.035 53.795 377.205 53.965 ;
        RECT 377.495 53.795 377.665 53.965 ;
        RECT 377.955 53.795 378.125 53.965 ;
        RECT 378.415 53.795 378.585 53.965 ;
        RECT 378.875 53.795 379.045 53.965 ;
        RECT 379.335 53.795 379.505 53.965 ;
        RECT 379.795 53.795 379.965 53.965 ;
        RECT 380.255 53.795 380.425 53.965 ;
        RECT 380.715 53.795 380.885 53.965 ;
        RECT 381.175 53.795 381.345 53.965 ;
        RECT 381.635 53.795 381.805 53.965 ;
        RECT 382.095 53.795 382.265 53.965 ;
        RECT 382.555 53.795 382.725 53.965 ;
        RECT 383.015 53.795 383.185 53.965 ;
        RECT 383.475 53.795 383.645 53.965 ;
        RECT 383.935 53.795 384.105 53.965 ;
        RECT 384.395 53.795 384.565 53.965 ;
        RECT 384.855 53.795 385.025 53.965 ;
        RECT 385.315 53.795 385.485 53.965 ;
        RECT 385.775 53.795 385.945 53.965 ;
        RECT 386.235 53.795 386.405 53.965 ;
        RECT 386.695 53.795 386.865 53.965 ;
        RECT 387.155 53.795 387.325 53.965 ;
        RECT 387.615 53.795 387.785 53.965 ;
        RECT 388.075 53.795 388.245 53.965 ;
        RECT 388.535 53.795 388.705 53.965 ;
        RECT 388.995 53.795 389.165 53.965 ;
        RECT 389.455 53.795 389.625 53.965 ;
        RECT 389.915 53.795 390.085 53.965 ;
        RECT 390.375 53.795 390.545 53.965 ;
        RECT 390.835 53.795 391.005 53.965 ;
        RECT 391.295 53.795 391.465 53.965 ;
        RECT 391.755 53.795 391.925 53.965 ;
        RECT 392.215 53.795 392.385 53.965 ;
        RECT 392.675 53.795 392.845 53.965 ;
        RECT 393.135 53.795 393.305 53.965 ;
        RECT 393.595 53.795 393.765 53.965 ;
        RECT 394.055 53.795 394.225 53.965 ;
        RECT 394.515 53.795 394.685 53.965 ;
        RECT 394.975 53.795 395.145 53.965 ;
        RECT 395.435 53.795 395.605 53.965 ;
        RECT 395.895 53.795 396.065 53.965 ;
        RECT 396.355 53.795 396.525 53.965 ;
        RECT 396.815 53.795 396.985 53.965 ;
        RECT 397.275 53.795 397.445 53.965 ;
        RECT 397.735 53.795 397.905 53.965 ;
        RECT 398.195 53.795 398.365 53.965 ;
        RECT 398.655 53.795 398.825 53.965 ;
        RECT 399.115 53.795 399.285 53.965 ;
        RECT 399.575 53.795 399.745 53.965 ;
        RECT 400.035 53.795 400.205 53.965 ;
        RECT 400.495 53.795 400.665 53.965 ;
        RECT 400.955 53.795 401.125 53.965 ;
        RECT 401.415 53.795 401.585 53.965 ;
        RECT 401.875 53.795 402.045 53.965 ;
        RECT 402.335 53.795 402.505 53.965 ;
        RECT 402.795 53.795 402.965 53.965 ;
        RECT 403.255 53.795 403.425 53.965 ;
        RECT 403.715 53.795 403.885 53.965 ;
        RECT 404.175 53.795 404.345 53.965 ;
        RECT 404.635 53.795 404.805 53.965 ;
        RECT 405.095 53.795 405.265 53.965 ;
        RECT 405.555 53.795 405.725 53.965 ;
        RECT 406.015 53.795 406.185 53.965 ;
        RECT 406.475 53.795 406.645 53.965 ;
        RECT 406.935 53.795 407.105 53.965 ;
        RECT 407.395 53.795 407.565 53.965 ;
        RECT 407.855 53.795 408.025 53.965 ;
        RECT 408.315 53.795 408.485 53.965 ;
        RECT 408.775 53.795 408.945 53.965 ;
        RECT 409.235 53.795 409.405 53.965 ;
        RECT 409.695 53.795 409.865 53.965 ;
        RECT 410.155 53.795 410.325 53.965 ;
        RECT 410.615 53.795 410.785 53.965 ;
        RECT 411.075 53.795 411.245 53.965 ;
        RECT 411.535 53.795 411.705 53.965 ;
        RECT 411.995 53.795 412.165 53.965 ;
        RECT 412.455 53.795 412.625 53.965 ;
        RECT 412.915 53.795 413.085 53.965 ;
        RECT 413.375 53.795 413.545 53.965 ;
        RECT 413.835 53.795 414.005 53.965 ;
        RECT 414.295 53.795 414.465 53.965 ;
        RECT 414.755 53.795 414.925 53.965 ;
        RECT 415.215 53.795 415.385 53.965 ;
        RECT 415.675 53.795 415.845 53.965 ;
        RECT 416.135 53.795 416.305 53.965 ;
        RECT 416.595 53.795 416.765 53.965 ;
        RECT 417.055 53.795 417.225 53.965 ;
        RECT 417.515 53.795 417.685 53.965 ;
        RECT 417.975 53.795 418.145 53.965 ;
        RECT 418.435 53.795 418.605 53.965 ;
        RECT 418.895 53.795 419.065 53.965 ;
        RECT 419.355 53.795 419.525 53.965 ;
        RECT 419.815 53.795 419.985 53.965 ;
        RECT 420.275 53.795 420.445 53.965 ;
        RECT 420.735 53.795 420.905 53.965 ;
        RECT 421.195 53.795 421.365 53.965 ;
        RECT 421.655 53.795 421.825 53.965 ;
        RECT 422.115 53.795 422.285 53.965 ;
        RECT 422.575 53.795 422.745 53.965 ;
        RECT 423.035 53.795 423.205 53.965 ;
        RECT 423.495 53.795 423.665 53.965 ;
        RECT 423.955 53.795 424.125 53.965 ;
        RECT 424.415 53.795 424.585 53.965 ;
        RECT 424.875 53.795 425.045 53.965 ;
        RECT 425.335 53.795 425.505 53.965 ;
        RECT 425.795 53.795 425.965 53.965 ;
        RECT 426.255 53.795 426.425 53.965 ;
        RECT 426.715 53.795 426.885 53.965 ;
        RECT 427.175 53.795 427.345 53.965 ;
        RECT 427.635 53.795 427.805 53.965 ;
        RECT 428.095 53.795 428.265 53.965 ;
        RECT 428.555 53.795 428.725 53.965 ;
        RECT 429.015 53.795 429.185 53.965 ;
        RECT 429.475 53.795 429.645 53.965 ;
        RECT 429.935 53.795 430.105 53.965 ;
        RECT 430.395 53.795 430.565 53.965 ;
        RECT 430.855 53.795 431.025 53.965 ;
        RECT 431.315 53.795 431.485 53.965 ;
        RECT 431.775 53.795 431.945 53.965 ;
        RECT 432.235 53.795 432.405 53.965 ;
        RECT 432.695 53.795 432.865 53.965 ;
        RECT 433.155 53.795 433.325 53.965 ;
        RECT 433.615 53.795 433.785 53.965 ;
        RECT 434.075 53.795 434.245 53.965 ;
        RECT 434.535 53.795 434.705 53.965 ;
        RECT 434.995 53.795 435.165 53.965 ;
        RECT 435.455 53.795 435.625 53.965 ;
        RECT 435.915 53.795 436.085 53.965 ;
        RECT 436.375 53.795 436.545 53.965 ;
        RECT 436.835 53.795 437.005 53.965 ;
        RECT 437.295 53.795 437.465 53.965 ;
        RECT 437.755 53.795 437.925 53.965 ;
        RECT 438.215 53.795 438.385 53.965 ;
        RECT 438.675 53.795 438.845 53.965 ;
        RECT 439.135 53.795 439.305 53.965 ;
        RECT 439.595 53.795 439.765 53.965 ;
        RECT 440.055 53.795 440.225 53.965 ;
        RECT 440.515 53.795 440.685 53.965 ;
        RECT 440.975 53.795 441.145 53.965 ;
        RECT 441.435 53.795 441.605 53.965 ;
        RECT 441.895 53.795 442.065 53.965 ;
        RECT 442.355 53.795 442.525 53.965 ;
        RECT 442.815 53.795 442.985 53.965 ;
        RECT 443.275 53.795 443.445 53.965 ;
        RECT 443.735 53.795 443.905 53.965 ;
        RECT 444.195 53.795 444.365 53.965 ;
        RECT 444.655 53.795 444.825 53.965 ;
        RECT 445.115 53.795 445.285 53.965 ;
        RECT 445.575 53.795 445.745 53.965 ;
        RECT 446.035 53.795 446.205 53.965 ;
        RECT 446.495 53.795 446.665 53.965 ;
        RECT 446.955 53.795 447.125 53.965 ;
        RECT 447.415 53.795 447.585 53.965 ;
        RECT 447.875 53.795 448.045 53.965 ;
        RECT 448.335 53.795 448.505 53.965 ;
        RECT 448.795 53.795 448.965 53.965 ;
        RECT 449.255 53.795 449.425 53.965 ;
        RECT 449.715 53.795 449.885 53.965 ;
        RECT 450.175 53.795 450.345 53.965 ;
        RECT 450.635 53.795 450.805 53.965 ;
        RECT 451.095 53.795 451.265 53.965 ;
        RECT 451.555 53.795 451.725 53.965 ;
        RECT 452.015 53.795 452.185 53.965 ;
        RECT 452.475 53.795 452.645 53.965 ;
        RECT 452.935 53.795 453.105 53.965 ;
        RECT 453.395 53.795 453.565 53.965 ;
        RECT 453.855 53.795 454.025 53.965 ;
        RECT 454.315 53.795 454.485 53.965 ;
        RECT 454.775 53.795 454.945 53.965 ;
        RECT 455.235 53.795 455.405 53.965 ;
        RECT 455.695 53.795 455.865 53.965 ;
        RECT 456.155 53.795 456.325 53.965 ;
        RECT 456.615 53.795 456.785 53.965 ;
        RECT 457.075 53.795 457.245 53.965 ;
        RECT 457.535 53.795 457.705 53.965 ;
        RECT 457.995 53.795 458.165 53.965 ;
        RECT 458.455 53.795 458.625 53.965 ;
        RECT 458.915 53.795 459.085 53.965 ;
        RECT 459.375 53.795 459.545 53.965 ;
        RECT 459.835 53.795 460.005 53.965 ;
        RECT 460.295 53.795 460.465 53.965 ;
        RECT 460.755 53.795 460.925 53.965 ;
        RECT 461.215 53.795 461.385 53.965 ;
        RECT 461.675 53.795 461.845 53.965 ;
        RECT 462.135 53.795 462.305 53.965 ;
        RECT 462.595 53.795 462.765 53.965 ;
        RECT 463.055 53.795 463.225 53.965 ;
        RECT 463.515 53.795 463.685 53.965 ;
        RECT 463.975 53.795 464.145 53.965 ;
        RECT 464.435 53.795 464.605 53.965 ;
        RECT 464.895 53.795 465.065 53.965 ;
        RECT 465.355 53.795 465.525 53.965 ;
        RECT 465.815 53.795 465.985 53.965 ;
        RECT 466.275 53.795 466.445 53.965 ;
        RECT 466.735 53.795 466.905 53.965 ;
        RECT 467.195 53.795 467.365 53.965 ;
        RECT 467.655 53.795 467.825 53.965 ;
        RECT 468.115 53.795 468.285 53.965 ;
        RECT 468.575 53.795 468.745 53.965 ;
        RECT 469.035 53.795 469.205 53.965 ;
        RECT 469.495 53.795 469.665 53.965 ;
        RECT 469.955 53.795 470.125 53.965 ;
        RECT 470.415 53.795 470.585 53.965 ;
        RECT 470.875 53.795 471.045 53.965 ;
        RECT 471.335 53.795 471.505 53.965 ;
        RECT 471.795 53.795 471.965 53.965 ;
        RECT 472.255 53.795 472.425 53.965 ;
        RECT 472.715 53.795 472.885 53.965 ;
        RECT 473.175 53.795 473.345 53.965 ;
        RECT 473.635 53.795 473.805 53.965 ;
        RECT 474.095 53.795 474.265 53.965 ;
        RECT 474.555 53.795 474.725 53.965 ;
        RECT 475.015 53.795 475.185 53.965 ;
        RECT 475.475 53.795 475.645 53.965 ;
        RECT 475.935 53.795 476.105 53.965 ;
        RECT 476.395 53.795 476.565 53.965 ;
        RECT 476.855 53.795 477.025 53.965 ;
        RECT 477.315 53.795 477.485 53.965 ;
        RECT 477.775 53.795 477.945 53.965 ;
        RECT 478.235 53.795 478.405 53.965 ;
        RECT 478.695 53.795 478.865 53.965 ;
        RECT 479.155 53.795 479.325 53.965 ;
        RECT 479.615 53.795 479.785 53.965 ;
        RECT 480.075 53.795 480.245 53.965 ;
        RECT 480.535 53.795 480.705 53.965 ;
        RECT 480.995 53.795 481.165 53.965 ;
        RECT 481.455 53.795 481.625 53.965 ;
        RECT 481.915 53.795 482.085 53.965 ;
        RECT 482.375 53.795 482.545 53.965 ;
        RECT 482.835 53.795 483.005 53.965 ;
        RECT 483.295 53.795 483.465 53.965 ;
        RECT 483.755 53.795 483.925 53.965 ;
        RECT 484.215 53.795 484.385 53.965 ;
        RECT 484.675 53.795 484.845 53.965 ;
        RECT 485.135 53.795 485.305 53.965 ;
        RECT 485.595 53.795 485.765 53.965 ;
        RECT 486.055 53.795 486.225 53.965 ;
        RECT 486.515 53.795 486.685 53.965 ;
        RECT 486.975 53.795 487.145 53.965 ;
        RECT 487.435 53.795 487.605 53.965 ;
        RECT 487.895 53.795 488.065 53.965 ;
        RECT 488.355 53.795 488.525 53.965 ;
        RECT 488.815 53.795 488.985 53.965 ;
        RECT 489.275 53.795 489.445 53.965 ;
        RECT 489.735 53.795 489.905 53.965 ;
        RECT 490.195 53.795 490.365 53.965 ;
        RECT 490.655 53.795 490.825 53.965 ;
        RECT 491.115 53.795 491.285 53.965 ;
        RECT 491.575 53.795 491.745 53.965 ;
        RECT 492.035 53.795 492.205 53.965 ;
        RECT 492.495 53.795 492.665 53.965 ;
        RECT 492.955 53.795 493.125 53.965 ;
        RECT 493.415 53.795 493.585 53.965 ;
        RECT 493.875 53.795 494.045 53.965 ;
        RECT 494.335 53.795 494.505 53.965 ;
        RECT 494.795 53.795 494.965 53.965 ;
        RECT 495.255 53.795 495.425 53.965 ;
        RECT 495.715 53.795 495.885 53.965 ;
        RECT 496.175 53.795 496.345 53.965 ;
        RECT 496.635 53.795 496.805 53.965 ;
        RECT 497.095 53.795 497.265 53.965 ;
        RECT 497.555 53.795 497.725 53.965 ;
        RECT 498.015 53.795 498.185 53.965 ;
        RECT 498.475 53.795 498.645 53.965 ;
        RECT 498.935 53.795 499.105 53.965 ;
        RECT 499.395 53.795 499.565 53.965 ;
        RECT 499.855 53.795 500.025 53.965 ;
        RECT 500.315 53.795 500.485 53.965 ;
        RECT 500.775 53.795 500.945 53.965 ;
        RECT 501.235 53.795 501.405 53.965 ;
        RECT 501.695 53.795 501.865 53.965 ;
        RECT 502.155 53.795 502.325 53.965 ;
        RECT 502.615 53.795 502.785 53.965 ;
        RECT 503.075 53.795 503.245 53.965 ;
        RECT 503.535 53.795 503.705 53.965 ;
        RECT 503.995 53.795 504.165 53.965 ;
        RECT 504.455 53.795 504.625 53.965 ;
        RECT 504.915 53.795 505.085 53.965 ;
        RECT 505.375 53.795 505.545 53.965 ;
        RECT 505.835 53.795 506.005 53.965 ;
        RECT 506.295 53.795 506.465 53.965 ;
        RECT 506.755 53.795 506.925 53.965 ;
        RECT 507.215 53.795 507.385 53.965 ;
        RECT 507.675 53.795 507.845 53.965 ;
        RECT 508.135 53.795 508.305 53.965 ;
        RECT 508.595 53.795 508.765 53.965 ;
        RECT 509.055 53.795 509.225 53.965 ;
        RECT 509.515 53.795 509.685 53.965 ;
        RECT 509.975 53.795 510.145 53.965 ;
        RECT 510.435 53.795 510.605 53.965 ;
        RECT 510.895 53.795 511.065 53.965 ;
        RECT 511.355 53.795 511.525 53.965 ;
        RECT 511.815 53.795 511.985 53.965 ;
        RECT 512.275 53.795 512.445 53.965 ;
        RECT 512.735 53.795 512.905 53.965 ;
        RECT 513.195 53.795 513.365 53.965 ;
        RECT 513.655 53.795 513.825 53.965 ;
        RECT 514.115 53.795 514.285 53.965 ;
        RECT 514.575 53.795 514.745 53.965 ;
        RECT 515.035 53.795 515.205 53.965 ;
        RECT 515.495 53.795 515.665 53.965 ;
        RECT 515.955 53.795 516.125 53.965 ;
        RECT 516.415 53.795 516.585 53.965 ;
        RECT 516.875 53.795 517.045 53.965 ;
        RECT 517.335 53.795 517.505 53.965 ;
        RECT 517.795 53.795 517.965 53.965 ;
        RECT 518.255 53.795 518.425 53.965 ;
        RECT 518.715 53.795 518.885 53.965 ;
        RECT 519.175 53.795 519.345 53.965 ;
        RECT 519.635 53.795 519.805 53.965 ;
        RECT 520.095 53.795 520.265 53.965 ;
        RECT 520.555 53.795 520.725 53.965 ;
        RECT 521.015 53.795 521.185 53.965 ;
        RECT 521.475 53.795 521.645 53.965 ;
        RECT 521.935 53.795 522.105 53.965 ;
        RECT 522.395 53.795 522.565 53.965 ;
        RECT 522.855 53.795 523.025 53.965 ;
        RECT 523.315 53.795 523.485 53.965 ;
        RECT 523.775 53.795 523.945 53.965 ;
        RECT 524.235 53.795 524.405 53.965 ;
        RECT 524.695 53.795 524.865 53.965 ;
        RECT 525.155 53.795 525.325 53.965 ;
        RECT 525.615 53.795 525.785 53.965 ;
        RECT 526.075 53.795 526.245 53.965 ;
        RECT 526.535 53.795 526.705 53.965 ;
        RECT 526.995 53.795 527.165 53.965 ;
        RECT 527.455 53.795 527.625 53.965 ;
        RECT 527.915 53.795 528.085 53.965 ;
        RECT 528.375 53.795 528.545 53.965 ;
        RECT 528.835 53.795 529.005 53.965 ;
        RECT 529.295 53.795 529.465 53.965 ;
        RECT 529.755 53.795 529.925 53.965 ;
        RECT 530.215 53.795 530.385 53.965 ;
        RECT 530.675 53.795 530.845 53.965 ;
        RECT 531.135 53.795 531.305 53.965 ;
        RECT 531.595 53.795 531.765 53.965 ;
        RECT 532.055 53.795 532.225 53.965 ;
        RECT 532.515 53.795 532.685 53.965 ;
        RECT 532.975 53.795 533.145 53.965 ;
        RECT 533.435 53.795 533.605 53.965 ;
        RECT 533.895 53.795 534.065 53.965 ;
        RECT 534.355 53.795 534.525 53.965 ;
        RECT 534.815 53.795 534.985 53.965 ;
        RECT 535.275 53.795 535.445 53.965 ;
        RECT 535.735 53.795 535.905 53.965 ;
        RECT 536.195 53.795 536.365 53.965 ;
        RECT 536.655 53.795 536.825 53.965 ;
        RECT 537.115 53.795 537.285 53.965 ;
        RECT 537.575 53.795 537.745 53.965 ;
        RECT 538.035 53.795 538.205 53.965 ;
        RECT 538.495 53.795 538.665 53.965 ;
        RECT 538.955 53.795 539.125 53.965 ;
        RECT 539.415 53.795 539.585 53.965 ;
        RECT 539.875 53.795 540.045 53.965 ;
        RECT 540.335 53.795 540.505 53.965 ;
        RECT 540.795 53.795 540.965 53.965 ;
        RECT 541.255 53.795 541.425 53.965 ;
        RECT 541.715 53.795 541.885 53.965 ;
        RECT 542.175 53.795 542.345 53.965 ;
        RECT 542.635 53.795 542.805 53.965 ;
        RECT 543.095 53.795 543.265 53.965 ;
        RECT 543.555 53.795 543.725 53.965 ;
        RECT 544.015 53.795 544.185 53.965 ;
        RECT 544.475 53.795 544.645 53.965 ;
        RECT 544.935 53.795 545.105 53.965 ;
        RECT 545.395 53.795 545.565 53.965 ;
        RECT 545.855 53.795 546.025 53.965 ;
        RECT 546.315 53.795 546.485 53.965 ;
        RECT 546.775 53.795 546.945 53.965 ;
        RECT 547.235 53.795 547.405 53.965 ;
        RECT 547.695 53.795 547.865 53.965 ;
        RECT 548.155 53.795 548.325 53.965 ;
        RECT 548.615 53.795 548.785 53.965 ;
        RECT 549.075 53.795 549.245 53.965 ;
        RECT 549.535 53.795 549.705 53.965 ;
        RECT 549.995 53.795 550.165 53.965 ;
        RECT 550.455 53.795 550.625 53.965 ;
        RECT 550.915 53.795 551.085 53.965 ;
        RECT 551.375 53.795 551.545 53.965 ;
        RECT 551.835 53.795 552.005 53.965 ;
        RECT 552.295 53.795 552.465 53.965 ;
        RECT 552.755 53.795 552.925 53.965 ;
        RECT 553.215 53.795 553.385 53.965 ;
        RECT 553.675 53.795 553.845 53.965 ;
        RECT 554.135 53.795 554.305 53.965 ;
        RECT 554.595 53.795 554.765 53.965 ;
        RECT 555.055 53.795 555.225 53.965 ;
        RECT 555.515 53.795 555.685 53.965 ;
        RECT 555.975 53.795 556.145 53.965 ;
        RECT 556.435 53.795 556.605 53.965 ;
        RECT 556.895 53.795 557.065 53.965 ;
        RECT 557.355 53.795 557.525 53.965 ;
        RECT 557.815 53.795 557.985 53.965 ;
        RECT 558.275 53.795 558.445 53.965 ;
        RECT 558.735 53.795 558.905 53.965 ;
        RECT 559.195 53.795 559.365 53.965 ;
        RECT 559.655 53.795 559.825 53.965 ;
        RECT 560.115 53.795 560.285 53.965 ;
        RECT 560.575 53.795 560.745 53.965 ;
        RECT 561.035 53.795 561.205 53.965 ;
        RECT 561.495 53.795 561.665 53.965 ;
        RECT 561.955 53.795 562.125 53.965 ;
        RECT 562.415 53.795 562.585 53.965 ;
        RECT 562.875 53.795 563.045 53.965 ;
        RECT 563.335 53.795 563.505 53.965 ;
        RECT 563.795 53.795 563.965 53.965 ;
        RECT 564.255 53.795 564.425 53.965 ;
        RECT 564.715 53.795 564.885 53.965 ;
        RECT 565.175 53.795 565.345 53.965 ;
        RECT 565.635 53.795 565.805 53.965 ;
        RECT 566.095 53.795 566.265 53.965 ;
        RECT 566.555 53.795 566.725 53.965 ;
        RECT 567.015 53.795 567.185 53.965 ;
        RECT 567.475 53.795 567.645 53.965 ;
        RECT 567.935 53.795 568.105 53.965 ;
        RECT 568.395 53.795 568.565 53.965 ;
        RECT 568.855 53.795 569.025 53.965 ;
        RECT 569.315 53.795 569.485 53.965 ;
        RECT 569.775 53.795 569.945 53.965 ;
        RECT 570.235 53.795 570.405 53.965 ;
        RECT 570.695 53.795 570.865 53.965 ;
        RECT 571.155 53.795 571.325 53.965 ;
        RECT 571.615 53.795 571.785 53.965 ;
        RECT 572.075 53.795 572.245 53.965 ;
        RECT 572.535 53.795 572.705 53.965 ;
        RECT 572.995 53.795 573.165 53.965 ;
        RECT 573.455 53.795 573.625 53.965 ;
        RECT 573.915 53.795 574.085 53.965 ;
        RECT 574.375 53.795 574.545 53.965 ;
        RECT 574.835 53.795 575.005 53.965 ;
        RECT 575.295 53.795 575.465 53.965 ;
        RECT 575.755 53.795 575.925 53.965 ;
        RECT 576.215 53.795 576.385 53.965 ;
        RECT 576.675 53.795 576.845 53.965 ;
        RECT 577.135 53.795 577.305 53.965 ;
        RECT 577.595 53.795 577.765 53.965 ;
        RECT 578.055 53.795 578.225 53.965 ;
        RECT 578.515 53.795 578.685 53.965 ;
        RECT 578.975 53.795 579.145 53.965 ;
        RECT 579.435 53.795 579.605 53.965 ;
        RECT 579.895 53.795 580.065 53.965 ;
        RECT 580.355 53.795 580.525 53.965 ;
        RECT 580.815 53.795 580.985 53.965 ;
        RECT 581.275 53.795 581.445 53.965 ;
        RECT 581.735 53.795 581.905 53.965 ;
        RECT 582.195 53.795 582.365 53.965 ;
        RECT 582.655 53.795 582.825 53.965 ;
        RECT 583.115 53.795 583.285 53.965 ;
        RECT 583.575 53.795 583.745 53.965 ;
        RECT 584.035 53.795 584.205 53.965 ;
        RECT 584.495 53.795 584.665 53.965 ;
        RECT 584.955 53.795 585.125 53.965 ;
        RECT 585.415 53.795 585.585 53.965 ;
        RECT 585.875 53.795 586.045 53.965 ;
        RECT 586.335 53.795 586.505 53.965 ;
        RECT 586.795 53.795 586.965 53.965 ;
        RECT 587.255 53.795 587.425 53.965 ;
        RECT 587.715 53.795 587.885 53.965 ;
        RECT 588.175 53.795 588.345 53.965 ;
        RECT 588.635 53.795 588.805 53.965 ;
        RECT 589.095 53.795 589.265 53.965 ;
        RECT 589.555 53.795 589.725 53.965 ;
        RECT 590.015 53.795 590.185 53.965 ;
        RECT 590.475 53.795 590.645 53.965 ;
        RECT 590.935 53.795 591.105 53.965 ;
        RECT 591.395 53.795 591.565 53.965 ;
        RECT 591.855 53.795 592.025 53.965 ;
        RECT 592.315 53.795 592.485 53.965 ;
        RECT 592.775 53.795 592.945 53.965 ;
        RECT 593.235 53.795 593.405 53.965 ;
        RECT 593.695 53.795 593.865 53.965 ;
        RECT 594.155 53.795 594.325 53.965 ;
        RECT 594.615 53.795 594.785 53.965 ;
        RECT 595.075 53.795 595.245 53.965 ;
        RECT 595.535 53.795 595.705 53.965 ;
        RECT 595.995 53.795 596.165 53.965 ;
        RECT 596.455 53.795 596.625 53.965 ;
        RECT 596.915 53.795 597.085 53.965 ;
        RECT 597.375 53.795 597.545 53.965 ;
        RECT 597.835 53.795 598.005 53.965 ;
        RECT 598.295 53.795 598.465 53.965 ;
        RECT 598.755 53.795 598.925 53.965 ;
        RECT 599.215 53.795 599.385 53.965 ;
        RECT 599.675 53.795 599.845 53.965 ;
        RECT 600.135 53.795 600.305 53.965 ;
        RECT 600.595 53.795 600.765 53.965 ;
        RECT 601.055 53.795 601.225 53.965 ;
        RECT 601.515 53.795 601.685 53.965 ;
        RECT 601.975 53.795 602.145 53.965 ;
        RECT 602.435 53.795 602.605 53.965 ;
        RECT 602.895 53.795 603.065 53.965 ;
        RECT 603.355 53.795 603.525 53.965 ;
        RECT 603.815 53.795 603.985 53.965 ;
        RECT 604.275 53.795 604.445 53.965 ;
        RECT 604.735 53.795 604.905 53.965 ;
        RECT 605.195 53.795 605.365 53.965 ;
        RECT 605.655 53.795 605.825 53.965 ;
        RECT 606.115 53.795 606.285 53.965 ;
        RECT 606.575 53.795 606.745 53.965 ;
        RECT 607.035 53.795 607.205 53.965 ;
        RECT 607.495 53.795 607.665 53.965 ;
        RECT 607.955 53.795 608.125 53.965 ;
        RECT 608.415 53.795 608.585 53.965 ;
        RECT 608.875 53.795 609.045 53.965 ;
        RECT 609.335 53.795 609.505 53.965 ;
        RECT 609.795 53.795 609.965 53.965 ;
        RECT 610.255 53.795 610.425 53.965 ;
        RECT 610.715 53.795 610.885 53.965 ;
        RECT 611.175 53.795 611.345 53.965 ;
        RECT 611.635 53.795 611.805 53.965 ;
        RECT 612.095 53.795 612.265 53.965 ;
        RECT 612.555 53.795 612.725 53.965 ;
        RECT 613.015 53.795 613.185 53.965 ;
        RECT 613.475 53.795 613.645 53.965 ;
        RECT 613.935 53.795 614.105 53.965 ;
        RECT 614.395 53.795 614.565 53.965 ;
        RECT 614.855 53.795 615.025 53.965 ;
        RECT 615.315 53.795 615.485 53.965 ;
        RECT 615.775 53.795 615.945 53.965 ;
        RECT 616.235 53.795 616.405 53.965 ;
        RECT 616.695 53.795 616.865 53.965 ;
        RECT 617.155 53.795 617.325 53.965 ;
        RECT 617.615 53.795 617.785 53.965 ;
        RECT 618.075 53.795 618.245 53.965 ;
        RECT 618.535 53.795 618.705 53.965 ;
        RECT 618.995 53.795 619.165 53.965 ;
        RECT 619.455 53.795 619.625 53.965 ;
        RECT 619.915 53.795 620.085 53.965 ;
        RECT 620.375 53.795 620.545 53.965 ;
        RECT 620.835 53.795 621.005 53.965 ;
        RECT 621.295 53.795 621.465 53.965 ;
        RECT 621.755 53.795 621.925 53.965 ;
        RECT 622.215 53.795 622.385 53.965 ;
        RECT 622.675 53.795 622.845 53.965 ;
        RECT 623.135 53.795 623.305 53.965 ;
        RECT 623.595 53.795 623.765 53.965 ;
        RECT 624.055 53.795 624.225 53.965 ;
        RECT 624.515 53.795 624.685 53.965 ;
        RECT 624.975 53.795 625.145 53.965 ;
        RECT 625.435 53.795 625.605 53.965 ;
        RECT 625.895 53.795 626.065 53.965 ;
        RECT 626.355 53.795 626.525 53.965 ;
        RECT 626.815 53.795 626.985 53.965 ;
        RECT 627.275 53.795 627.445 53.965 ;
        RECT 627.735 53.795 627.905 53.965 ;
        RECT 628.195 53.795 628.365 53.965 ;
        RECT 628.655 53.795 628.825 53.965 ;
        RECT 629.115 53.795 629.285 53.965 ;
        RECT 629.575 53.795 629.745 53.965 ;
        RECT 630.035 53.795 630.205 53.965 ;
        RECT 630.495 53.795 630.665 53.965 ;
        RECT 630.955 53.795 631.125 53.965 ;
        RECT 83.100 52.945 83.270 53.115 ;
        RECT 77.575 52.265 77.745 52.435 ;
        RECT 78.035 51.585 78.205 51.755 ;
        RECT 82.635 52.605 82.805 52.775 ;
        RECT 84.015 52.265 84.185 52.435 ;
        RECT 83.560 51.925 83.730 52.095 ;
        RECT 85.420 52.945 85.590 53.115 ;
        RECT 84.960 51.925 85.130 52.095 ;
        RECT 86.800 52.945 86.970 53.115 ;
        RECT 86.800 51.925 86.970 52.095 ;
        RECT 99.660 52.945 99.830 53.115 ;
        RECT 99.195 52.265 99.365 52.435 ;
        RECT 89.535 51.585 89.705 51.755 ;
        RECT 100.575 52.605 100.745 52.775 ;
        RECT 100.120 51.925 100.290 52.095 ;
        RECT 101.980 52.945 102.150 53.115 ;
        RECT 101.520 51.925 101.690 52.095 ;
        RECT 103.360 52.945 103.530 53.115 ;
        RECT 103.360 51.925 103.530 52.095 ;
        RECT 112.080 52.945 112.250 53.115 ;
        RECT 111.615 52.265 111.785 52.435 ;
        RECT 106.095 51.585 106.265 51.755 ;
        RECT 112.995 52.605 113.165 52.775 ;
        RECT 112.540 51.925 112.710 52.095 ;
        RECT 114.400 52.945 114.570 53.115 ;
        RECT 113.940 51.925 114.110 52.095 ;
        RECT 115.780 52.945 115.950 53.115 ;
        RECT 115.780 51.925 115.950 52.095 ;
        RECT 127.720 52.945 127.890 53.115 ;
        RECT 127.255 52.265 127.425 52.435 ;
        RECT 118.515 51.585 118.685 51.755 ;
        RECT 128.635 52.265 128.805 52.435 ;
        RECT 128.180 51.925 128.350 52.095 ;
        RECT 130.040 52.945 130.210 53.115 ;
        RECT 129.580 51.925 129.750 52.095 ;
        RECT 131.420 52.945 131.590 53.115 ;
        RECT 131.420 51.925 131.590 52.095 ;
        RECT 140.140 52.945 140.310 53.115 ;
        RECT 139.675 52.265 139.845 52.435 ;
        RECT 141.055 52.265 141.225 52.435 ;
        RECT 140.600 51.925 140.770 52.095 ;
        RECT 142.460 52.945 142.630 53.115 ;
        RECT 142.000 51.925 142.170 52.095 ;
        RECT 143.840 52.945 144.010 53.115 ;
        RECT 143.840 51.925 144.010 52.095 ;
        RECT 155.780 52.945 155.950 53.115 ;
        RECT 155.315 52.605 155.485 52.775 ;
        RECT 156.695 52.605 156.865 52.775 ;
        RECT 156.240 51.925 156.410 52.095 ;
        RECT 158.100 52.945 158.270 53.115 ;
        RECT 157.640 51.925 157.810 52.095 ;
        RECT 159.480 52.945 159.650 53.115 ;
        RECT 159.480 51.925 159.650 52.095 ;
        RECT 162.215 53.285 162.385 53.455 ;
        RECT 170.960 52.945 171.130 53.115 ;
        RECT 170.495 52.265 170.665 52.435 ;
        RECT 171.875 52.605 172.045 52.775 ;
        RECT 171.420 51.925 171.590 52.095 ;
        RECT 173.280 52.945 173.450 53.115 ;
        RECT 172.820 51.925 172.990 52.095 ;
        RECT 174.660 52.945 174.830 53.115 ;
        RECT 174.660 51.925 174.830 52.095 ;
        RECT 185.680 52.945 185.850 53.115 ;
        RECT 185.215 52.265 185.385 52.435 ;
        RECT 186.595 52.605 186.765 52.775 ;
        RECT 186.140 51.925 186.310 52.095 ;
        RECT 188.000 52.945 188.170 53.115 ;
        RECT 187.540 51.925 187.710 52.095 ;
        RECT 189.380 52.945 189.550 53.115 ;
        RECT 189.380 51.925 189.550 52.095 ;
        RECT 198.560 52.945 198.730 53.115 ;
        RECT 198.095 52.265 198.265 52.435 ;
        RECT 192.115 51.585 192.285 51.755 ;
        RECT 199.475 52.265 199.645 52.435 ;
        RECT 199.020 51.925 199.190 52.095 ;
        RECT 200.880 52.945 201.050 53.115 ;
        RECT 200.420 51.925 200.590 52.095 ;
        RECT 202.260 52.945 202.430 53.115 ;
        RECT 202.260 51.925 202.430 52.095 ;
        RECT 210.515 52.605 210.685 52.775 ;
        RECT 212.355 52.605 212.525 52.775 ;
        RECT 213.275 52.265 213.445 52.435 ;
        RECT 214.660 52.605 214.830 52.775 ;
        RECT 204.995 51.585 205.165 51.755 ;
        RECT 215.575 52.265 215.745 52.435 ;
        RECT 216.035 52.265 216.205 52.435 ;
        RECT 217.440 52.605 217.610 52.775 ;
        RECT 226.155 52.605 226.325 52.775 ;
        RECT 223.395 52.265 223.565 52.435 ;
        RECT 225.695 52.265 225.865 52.435 ;
        RECT 218.335 51.585 218.505 51.755 ;
        RECT 234.895 52.605 235.065 52.775 ;
        RECT 231.215 52.265 231.385 52.435 ;
        RECT 232.135 52.265 232.305 52.435 ;
        RECT 232.595 52.265 232.765 52.435 ;
        RECT 239.495 52.265 239.665 52.435 ;
        RECT 240.415 51.585 240.585 51.755 ;
        RECT 245.015 52.265 245.185 52.435 ;
        RECT 245.935 52.265 246.105 52.435 ;
        RECT 247.320 52.605 247.490 52.775 ;
        RECT 248.695 52.265 248.865 52.435 ;
        RECT 249.615 52.265 249.785 52.435 ;
        RECT 250.100 52.605 250.270 52.775 ;
        RECT 256.515 52.605 256.685 52.775 ;
        RECT 256.975 52.265 257.145 52.435 ;
        RECT 258.360 52.605 258.530 52.775 ;
        RECT 259.275 52.265 259.445 52.435 ;
        RECT 259.735 52.265 259.905 52.435 ;
        RECT 261.140 52.605 261.310 52.775 ;
        RECT 262.035 52.605 262.205 52.775 ;
        RECT 250.995 51.585 251.165 51.755 ;
        RECT 273.540 52.605 273.710 52.775 ;
        RECT 272.155 52.265 272.325 52.435 ;
        RECT 272.615 52.265 272.785 52.435 ;
        RECT 274.455 52.265 274.625 52.435 ;
        RECT 274.915 52.265 275.085 52.435 ;
        RECT 276.320 52.605 276.490 52.775 ;
        RECT 277.215 52.605 277.385 52.775 ;
        RECT 284.580 52.605 284.750 52.775 ;
        RECT 283.195 52.265 283.365 52.435 ;
        RECT 283.655 52.265 283.825 52.435 ;
        RECT 285.495 52.265 285.665 52.435 ;
        RECT 285.955 52.265 286.125 52.435 ;
        RECT 287.360 52.605 287.530 52.775 ;
        RECT 288.255 52.605 288.425 52.775 ;
        RECT 296.995 52.265 297.165 52.435 ;
        RECT 298.375 52.265 298.545 52.435 ;
        RECT 308.500 52.605 308.670 52.775 ;
        RECT 307.115 52.265 307.285 52.435 ;
        RECT 307.575 52.265 307.745 52.435 ;
        RECT 309.875 52.265 310.045 52.435 ;
        RECT 310.795 52.265 310.965 52.435 ;
        RECT 311.280 52.605 311.450 52.775 ;
        RECT 296.075 51.585 296.245 51.755 ;
        RECT 317.235 52.265 317.405 52.435 ;
        RECT 312.175 51.585 312.345 51.755 ;
        RECT 318.155 51.585 318.325 51.755 ;
        RECT 323.675 52.265 323.845 52.435 ;
        RECT 324.595 51.585 324.765 51.755 ;
        RECT 329.195 52.265 329.365 52.435 ;
        RECT 330.115 52.265 330.285 52.435 ;
        RECT 331.500 52.605 331.670 52.775 ;
        RECT 332.415 52.265 332.585 52.435 ;
        RECT 332.875 52.265 333.045 52.435 ;
        RECT 334.280 52.605 334.450 52.775 ;
        RECT 335.175 52.605 335.345 52.775 ;
        RECT 340.695 52.605 340.865 52.775 ;
        RECT 341.080 52.265 341.250 52.435 ;
        RECT 342.540 52.605 342.710 52.775 ;
        RECT 343.455 52.265 343.625 52.435 ;
        RECT 343.915 52.265 344.085 52.435 ;
        RECT 345.320 52.605 345.490 52.775 ;
        RECT 346.215 52.605 346.385 52.775 ;
        RECT 352.195 52.605 352.365 52.775 ;
        RECT 352.655 52.265 352.825 52.435 ;
        RECT 354.040 52.605 354.210 52.775 ;
        RECT 354.955 52.265 355.125 52.435 ;
        RECT 355.415 52.265 355.585 52.435 ;
        RECT 356.820 52.605 356.990 52.775 ;
        RECT 357.715 52.605 357.885 52.775 ;
        RECT 365.535 52.605 365.705 52.775 ;
        RECT 364.155 52.265 364.325 52.435 ;
        RECT 365.075 52.265 365.245 52.435 ;
        RECT 371.975 52.265 372.145 52.435 ;
        RECT 372.895 52.265 373.065 52.435 ;
        RECT 371.055 51.585 371.225 51.755 ;
        RECT 380.715 52.605 380.885 52.775 ;
        RECT 385.775 52.945 385.945 53.115 ;
        RECT 390.835 52.265 391.005 52.435 ;
        RECT 624.975 52.265 625.145 52.435 ;
        RECT 42.615 51.075 42.785 51.245 ;
        RECT 43.075 51.075 43.245 51.245 ;
        RECT 43.535 51.075 43.705 51.245 ;
        RECT 43.995 51.075 44.165 51.245 ;
        RECT 44.455 51.075 44.625 51.245 ;
        RECT 44.915 51.075 45.085 51.245 ;
        RECT 45.375 51.075 45.545 51.245 ;
        RECT 45.835 51.075 46.005 51.245 ;
        RECT 46.295 51.075 46.465 51.245 ;
        RECT 46.755 51.075 46.925 51.245 ;
        RECT 47.215 51.075 47.385 51.245 ;
        RECT 47.675 51.075 47.845 51.245 ;
        RECT 48.135 51.075 48.305 51.245 ;
        RECT 48.595 51.075 48.765 51.245 ;
        RECT 49.055 51.075 49.225 51.245 ;
        RECT 49.515 51.075 49.685 51.245 ;
        RECT 49.975 51.075 50.145 51.245 ;
        RECT 50.435 51.075 50.605 51.245 ;
        RECT 50.895 51.075 51.065 51.245 ;
        RECT 51.355 51.075 51.525 51.245 ;
        RECT 51.815 51.075 51.985 51.245 ;
        RECT 52.275 51.075 52.445 51.245 ;
        RECT 52.735 51.075 52.905 51.245 ;
        RECT 53.195 51.075 53.365 51.245 ;
        RECT 53.655 51.075 53.825 51.245 ;
        RECT 54.115 51.075 54.285 51.245 ;
        RECT 54.575 51.075 54.745 51.245 ;
        RECT 55.035 51.075 55.205 51.245 ;
        RECT 55.495 51.075 55.665 51.245 ;
        RECT 55.955 51.075 56.125 51.245 ;
        RECT 56.415 51.075 56.585 51.245 ;
        RECT 56.875 51.075 57.045 51.245 ;
        RECT 57.335 51.075 57.505 51.245 ;
        RECT 57.795 51.075 57.965 51.245 ;
        RECT 58.255 51.075 58.425 51.245 ;
        RECT 58.715 51.075 58.885 51.245 ;
        RECT 59.175 51.075 59.345 51.245 ;
        RECT 59.635 51.075 59.805 51.245 ;
        RECT 60.095 51.075 60.265 51.245 ;
        RECT 60.555 51.075 60.725 51.245 ;
        RECT 61.015 51.075 61.185 51.245 ;
        RECT 61.475 51.075 61.645 51.245 ;
        RECT 61.935 51.075 62.105 51.245 ;
        RECT 62.395 51.075 62.565 51.245 ;
        RECT 62.855 51.075 63.025 51.245 ;
        RECT 63.315 51.075 63.485 51.245 ;
        RECT 63.775 51.075 63.945 51.245 ;
        RECT 64.235 51.075 64.405 51.245 ;
        RECT 64.695 51.075 64.865 51.245 ;
        RECT 65.155 51.075 65.325 51.245 ;
        RECT 65.615 51.075 65.785 51.245 ;
        RECT 66.075 51.075 66.245 51.245 ;
        RECT 66.535 51.075 66.705 51.245 ;
        RECT 66.995 51.075 67.165 51.245 ;
        RECT 67.455 51.075 67.625 51.245 ;
        RECT 67.915 51.075 68.085 51.245 ;
        RECT 68.375 51.075 68.545 51.245 ;
        RECT 68.835 51.075 69.005 51.245 ;
        RECT 69.295 51.075 69.465 51.245 ;
        RECT 69.755 51.075 69.925 51.245 ;
        RECT 70.215 51.075 70.385 51.245 ;
        RECT 70.675 51.075 70.845 51.245 ;
        RECT 71.135 51.075 71.305 51.245 ;
        RECT 71.595 51.075 71.765 51.245 ;
        RECT 72.055 51.075 72.225 51.245 ;
        RECT 72.515 51.075 72.685 51.245 ;
        RECT 72.975 51.075 73.145 51.245 ;
        RECT 73.435 51.075 73.605 51.245 ;
        RECT 73.895 51.075 74.065 51.245 ;
        RECT 74.355 51.075 74.525 51.245 ;
        RECT 74.815 51.075 74.985 51.245 ;
        RECT 75.275 51.075 75.445 51.245 ;
        RECT 75.735 51.075 75.905 51.245 ;
        RECT 76.195 51.075 76.365 51.245 ;
        RECT 76.655 51.075 76.825 51.245 ;
        RECT 77.115 51.075 77.285 51.245 ;
        RECT 77.575 51.075 77.745 51.245 ;
        RECT 78.035 51.075 78.205 51.245 ;
        RECT 78.495 51.075 78.665 51.245 ;
        RECT 78.955 51.075 79.125 51.245 ;
        RECT 79.415 51.075 79.585 51.245 ;
        RECT 79.875 51.075 80.045 51.245 ;
        RECT 80.335 51.075 80.505 51.245 ;
        RECT 80.795 51.075 80.965 51.245 ;
        RECT 81.255 51.075 81.425 51.245 ;
        RECT 81.715 51.075 81.885 51.245 ;
        RECT 82.175 51.075 82.345 51.245 ;
        RECT 82.635 51.075 82.805 51.245 ;
        RECT 83.095 51.075 83.265 51.245 ;
        RECT 83.555 51.075 83.725 51.245 ;
        RECT 84.015 51.075 84.185 51.245 ;
        RECT 84.475 51.075 84.645 51.245 ;
        RECT 84.935 51.075 85.105 51.245 ;
        RECT 85.395 51.075 85.565 51.245 ;
        RECT 85.855 51.075 86.025 51.245 ;
        RECT 86.315 51.075 86.485 51.245 ;
        RECT 86.775 51.075 86.945 51.245 ;
        RECT 87.235 51.075 87.405 51.245 ;
        RECT 87.695 51.075 87.865 51.245 ;
        RECT 88.155 51.075 88.325 51.245 ;
        RECT 88.615 51.075 88.785 51.245 ;
        RECT 89.075 51.075 89.245 51.245 ;
        RECT 89.535 51.075 89.705 51.245 ;
        RECT 89.995 51.075 90.165 51.245 ;
        RECT 90.455 51.075 90.625 51.245 ;
        RECT 90.915 51.075 91.085 51.245 ;
        RECT 91.375 51.075 91.545 51.245 ;
        RECT 91.835 51.075 92.005 51.245 ;
        RECT 92.295 51.075 92.465 51.245 ;
        RECT 92.755 51.075 92.925 51.245 ;
        RECT 93.215 51.075 93.385 51.245 ;
        RECT 93.675 51.075 93.845 51.245 ;
        RECT 94.135 51.075 94.305 51.245 ;
        RECT 94.595 51.075 94.765 51.245 ;
        RECT 95.055 51.075 95.225 51.245 ;
        RECT 95.515 51.075 95.685 51.245 ;
        RECT 95.975 51.075 96.145 51.245 ;
        RECT 96.435 51.075 96.605 51.245 ;
        RECT 96.895 51.075 97.065 51.245 ;
        RECT 97.355 51.075 97.525 51.245 ;
        RECT 97.815 51.075 97.985 51.245 ;
        RECT 98.275 51.075 98.445 51.245 ;
        RECT 98.735 51.075 98.905 51.245 ;
        RECT 99.195 51.075 99.365 51.245 ;
        RECT 99.655 51.075 99.825 51.245 ;
        RECT 100.115 51.075 100.285 51.245 ;
        RECT 100.575 51.075 100.745 51.245 ;
        RECT 101.035 51.075 101.205 51.245 ;
        RECT 101.495 51.075 101.665 51.245 ;
        RECT 101.955 51.075 102.125 51.245 ;
        RECT 102.415 51.075 102.585 51.245 ;
        RECT 102.875 51.075 103.045 51.245 ;
        RECT 103.335 51.075 103.505 51.245 ;
        RECT 103.795 51.075 103.965 51.245 ;
        RECT 104.255 51.075 104.425 51.245 ;
        RECT 104.715 51.075 104.885 51.245 ;
        RECT 105.175 51.075 105.345 51.245 ;
        RECT 105.635 51.075 105.805 51.245 ;
        RECT 106.095 51.075 106.265 51.245 ;
        RECT 106.555 51.075 106.725 51.245 ;
        RECT 107.015 51.075 107.185 51.245 ;
        RECT 107.475 51.075 107.645 51.245 ;
        RECT 107.935 51.075 108.105 51.245 ;
        RECT 108.395 51.075 108.565 51.245 ;
        RECT 108.855 51.075 109.025 51.245 ;
        RECT 109.315 51.075 109.485 51.245 ;
        RECT 109.775 51.075 109.945 51.245 ;
        RECT 110.235 51.075 110.405 51.245 ;
        RECT 110.695 51.075 110.865 51.245 ;
        RECT 111.155 51.075 111.325 51.245 ;
        RECT 111.615 51.075 111.785 51.245 ;
        RECT 112.075 51.075 112.245 51.245 ;
        RECT 112.535 51.075 112.705 51.245 ;
        RECT 112.995 51.075 113.165 51.245 ;
        RECT 113.455 51.075 113.625 51.245 ;
        RECT 113.915 51.075 114.085 51.245 ;
        RECT 114.375 51.075 114.545 51.245 ;
        RECT 114.835 51.075 115.005 51.245 ;
        RECT 115.295 51.075 115.465 51.245 ;
        RECT 115.755 51.075 115.925 51.245 ;
        RECT 116.215 51.075 116.385 51.245 ;
        RECT 116.675 51.075 116.845 51.245 ;
        RECT 117.135 51.075 117.305 51.245 ;
        RECT 117.595 51.075 117.765 51.245 ;
        RECT 118.055 51.075 118.225 51.245 ;
        RECT 118.515 51.075 118.685 51.245 ;
        RECT 118.975 51.075 119.145 51.245 ;
        RECT 119.435 51.075 119.605 51.245 ;
        RECT 119.895 51.075 120.065 51.245 ;
        RECT 120.355 51.075 120.525 51.245 ;
        RECT 120.815 51.075 120.985 51.245 ;
        RECT 121.275 51.075 121.445 51.245 ;
        RECT 121.735 51.075 121.905 51.245 ;
        RECT 122.195 51.075 122.365 51.245 ;
        RECT 122.655 51.075 122.825 51.245 ;
        RECT 123.115 51.075 123.285 51.245 ;
        RECT 123.575 51.075 123.745 51.245 ;
        RECT 124.035 51.075 124.205 51.245 ;
        RECT 124.495 51.075 124.665 51.245 ;
        RECT 124.955 51.075 125.125 51.245 ;
        RECT 125.415 51.075 125.585 51.245 ;
        RECT 125.875 51.075 126.045 51.245 ;
        RECT 126.335 51.075 126.505 51.245 ;
        RECT 126.795 51.075 126.965 51.245 ;
        RECT 127.255 51.075 127.425 51.245 ;
        RECT 127.715 51.075 127.885 51.245 ;
        RECT 128.175 51.075 128.345 51.245 ;
        RECT 128.635 51.075 128.805 51.245 ;
        RECT 129.095 51.075 129.265 51.245 ;
        RECT 129.555 51.075 129.725 51.245 ;
        RECT 130.015 51.075 130.185 51.245 ;
        RECT 130.475 51.075 130.645 51.245 ;
        RECT 130.935 51.075 131.105 51.245 ;
        RECT 131.395 51.075 131.565 51.245 ;
        RECT 131.855 51.075 132.025 51.245 ;
        RECT 132.315 51.075 132.485 51.245 ;
        RECT 132.775 51.075 132.945 51.245 ;
        RECT 133.235 51.075 133.405 51.245 ;
        RECT 133.695 51.075 133.865 51.245 ;
        RECT 134.155 51.075 134.325 51.245 ;
        RECT 134.615 51.075 134.785 51.245 ;
        RECT 135.075 51.075 135.245 51.245 ;
        RECT 135.535 51.075 135.705 51.245 ;
        RECT 135.995 51.075 136.165 51.245 ;
        RECT 136.455 51.075 136.625 51.245 ;
        RECT 136.915 51.075 137.085 51.245 ;
        RECT 137.375 51.075 137.545 51.245 ;
        RECT 137.835 51.075 138.005 51.245 ;
        RECT 138.295 51.075 138.465 51.245 ;
        RECT 138.755 51.075 138.925 51.245 ;
        RECT 139.215 51.075 139.385 51.245 ;
        RECT 139.675 51.075 139.845 51.245 ;
        RECT 140.135 51.075 140.305 51.245 ;
        RECT 140.595 51.075 140.765 51.245 ;
        RECT 141.055 51.075 141.225 51.245 ;
        RECT 141.515 51.075 141.685 51.245 ;
        RECT 141.975 51.075 142.145 51.245 ;
        RECT 142.435 51.075 142.605 51.245 ;
        RECT 142.895 51.075 143.065 51.245 ;
        RECT 143.355 51.075 143.525 51.245 ;
        RECT 143.815 51.075 143.985 51.245 ;
        RECT 144.275 51.075 144.445 51.245 ;
        RECT 144.735 51.075 144.905 51.245 ;
        RECT 145.195 51.075 145.365 51.245 ;
        RECT 145.655 51.075 145.825 51.245 ;
        RECT 146.115 51.075 146.285 51.245 ;
        RECT 146.575 51.075 146.745 51.245 ;
        RECT 147.035 51.075 147.205 51.245 ;
        RECT 147.495 51.075 147.665 51.245 ;
        RECT 147.955 51.075 148.125 51.245 ;
        RECT 148.415 51.075 148.585 51.245 ;
        RECT 148.875 51.075 149.045 51.245 ;
        RECT 149.335 51.075 149.505 51.245 ;
        RECT 149.795 51.075 149.965 51.245 ;
        RECT 150.255 51.075 150.425 51.245 ;
        RECT 150.715 51.075 150.885 51.245 ;
        RECT 151.175 51.075 151.345 51.245 ;
        RECT 151.635 51.075 151.805 51.245 ;
        RECT 152.095 51.075 152.265 51.245 ;
        RECT 152.555 51.075 152.725 51.245 ;
        RECT 153.015 51.075 153.185 51.245 ;
        RECT 153.475 51.075 153.645 51.245 ;
        RECT 153.935 51.075 154.105 51.245 ;
        RECT 154.395 51.075 154.565 51.245 ;
        RECT 154.855 51.075 155.025 51.245 ;
        RECT 155.315 51.075 155.485 51.245 ;
        RECT 155.775 51.075 155.945 51.245 ;
        RECT 156.235 51.075 156.405 51.245 ;
        RECT 156.695 51.075 156.865 51.245 ;
        RECT 157.155 51.075 157.325 51.245 ;
        RECT 157.615 51.075 157.785 51.245 ;
        RECT 158.075 51.075 158.245 51.245 ;
        RECT 158.535 51.075 158.705 51.245 ;
        RECT 158.995 51.075 159.165 51.245 ;
        RECT 159.455 51.075 159.625 51.245 ;
        RECT 159.915 51.075 160.085 51.245 ;
        RECT 160.375 51.075 160.545 51.245 ;
        RECT 160.835 51.075 161.005 51.245 ;
        RECT 161.295 51.075 161.465 51.245 ;
        RECT 161.755 51.075 161.925 51.245 ;
        RECT 162.215 51.075 162.385 51.245 ;
        RECT 162.675 51.075 162.845 51.245 ;
        RECT 163.135 51.075 163.305 51.245 ;
        RECT 163.595 51.075 163.765 51.245 ;
        RECT 164.055 51.075 164.225 51.245 ;
        RECT 164.515 51.075 164.685 51.245 ;
        RECT 164.975 51.075 165.145 51.245 ;
        RECT 165.435 51.075 165.605 51.245 ;
        RECT 165.895 51.075 166.065 51.245 ;
        RECT 166.355 51.075 166.525 51.245 ;
        RECT 166.815 51.075 166.985 51.245 ;
        RECT 167.275 51.075 167.445 51.245 ;
        RECT 167.735 51.075 167.905 51.245 ;
        RECT 168.195 51.075 168.365 51.245 ;
        RECT 168.655 51.075 168.825 51.245 ;
        RECT 169.115 51.075 169.285 51.245 ;
        RECT 169.575 51.075 169.745 51.245 ;
        RECT 170.035 51.075 170.205 51.245 ;
        RECT 170.495 51.075 170.665 51.245 ;
        RECT 170.955 51.075 171.125 51.245 ;
        RECT 171.415 51.075 171.585 51.245 ;
        RECT 171.875 51.075 172.045 51.245 ;
        RECT 172.335 51.075 172.505 51.245 ;
        RECT 172.795 51.075 172.965 51.245 ;
        RECT 173.255 51.075 173.425 51.245 ;
        RECT 173.715 51.075 173.885 51.245 ;
        RECT 174.175 51.075 174.345 51.245 ;
        RECT 174.635 51.075 174.805 51.245 ;
        RECT 175.095 51.075 175.265 51.245 ;
        RECT 175.555 51.075 175.725 51.245 ;
        RECT 176.015 51.075 176.185 51.245 ;
        RECT 176.475 51.075 176.645 51.245 ;
        RECT 176.935 51.075 177.105 51.245 ;
        RECT 177.395 51.075 177.565 51.245 ;
        RECT 177.855 51.075 178.025 51.245 ;
        RECT 178.315 51.075 178.485 51.245 ;
        RECT 178.775 51.075 178.945 51.245 ;
        RECT 179.235 51.075 179.405 51.245 ;
        RECT 179.695 51.075 179.865 51.245 ;
        RECT 180.155 51.075 180.325 51.245 ;
        RECT 180.615 51.075 180.785 51.245 ;
        RECT 181.075 51.075 181.245 51.245 ;
        RECT 181.535 51.075 181.705 51.245 ;
        RECT 181.995 51.075 182.165 51.245 ;
        RECT 182.455 51.075 182.625 51.245 ;
        RECT 182.915 51.075 183.085 51.245 ;
        RECT 183.375 51.075 183.545 51.245 ;
        RECT 183.835 51.075 184.005 51.245 ;
        RECT 184.295 51.075 184.465 51.245 ;
        RECT 184.755 51.075 184.925 51.245 ;
        RECT 185.215 51.075 185.385 51.245 ;
        RECT 185.675 51.075 185.845 51.245 ;
        RECT 186.135 51.075 186.305 51.245 ;
        RECT 186.595 51.075 186.765 51.245 ;
        RECT 187.055 51.075 187.225 51.245 ;
        RECT 187.515 51.075 187.685 51.245 ;
        RECT 187.975 51.075 188.145 51.245 ;
        RECT 188.435 51.075 188.605 51.245 ;
        RECT 188.895 51.075 189.065 51.245 ;
        RECT 189.355 51.075 189.525 51.245 ;
        RECT 189.815 51.075 189.985 51.245 ;
        RECT 190.275 51.075 190.445 51.245 ;
        RECT 190.735 51.075 190.905 51.245 ;
        RECT 191.195 51.075 191.365 51.245 ;
        RECT 191.655 51.075 191.825 51.245 ;
        RECT 192.115 51.075 192.285 51.245 ;
        RECT 192.575 51.075 192.745 51.245 ;
        RECT 193.035 51.075 193.205 51.245 ;
        RECT 193.495 51.075 193.665 51.245 ;
        RECT 193.955 51.075 194.125 51.245 ;
        RECT 194.415 51.075 194.585 51.245 ;
        RECT 194.875 51.075 195.045 51.245 ;
        RECT 195.335 51.075 195.505 51.245 ;
        RECT 195.795 51.075 195.965 51.245 ;
        RECT 196.255 51.075 196.425 51.245 ;
        RECT 196.715 51.075 196.885 51.245 ;
        RECT 197.175 51.075 197.345 51.245 ;
        RECT 197.635 51.075 197.805 51.245 ;
        RECT 198.095 51.075 198.265 51.245 ;
        RECT 198.555 51.075 198.725 51.245 ;
        RECT 199.015 51.075 199.185 51.245 ;
        RECT 199.475 51.075 199.645 51.245 ;
        RECT 199.935 51.075 200.105 51.245 ;
        RECT 200.395 51.075 200.565 51.245 ;
        RECT 200.855 51.075 201.025 51.245 ;
        RECT 201.315 51.075 201.485 51.245 ;
        RECT 201.775 51.075 201.945 51.245 ;
        RECT 202.235 51.075 202.405 51.245 ;
        RECT 202.695 51.075 202.865 51.245 ;
        RECT 203.155 51.075 203.325 51.245 ;
        RECT 203.615 51.075 203.785 51.245 ;
        RECT 204.075 51.075 204.245 51.245 ;
        RECT 204.535 51.075 204.705 51.245 ;
        RECT 204.995 51.075 205.165 51.245 ;
        RECT 205.455 51.075 205.625 51.245 ;
        RECT 205.915 51.075 206.085 51.245 ;
        RECT 206.375 51.075 206.545 51.245 ;
        RECT 206.835 51.075 207.005 51.245 ;
        RECT 207.295 51.075 207.465 51.245 ;
        RECT 207.755 51.075 207.925 51.245 ;
        RECT 208.215 51.075 208.385 51.245 ;
        RECT 208.675 51.075 208.845 51.245 ;
        RECT 209.135 51.075 209.305 51.245 ;
        RECT 209.595 51.075 209.765 51.245 ;
        RECT 210.055 51.075 210.225 51.245 ;
        RECT 210.515 51.075 210.685 51.245 ;
        RECT 210.975 51.075 211.145 51.245 ;
        RECT 211.435 51.075 211.605 51.245 ;
        RECT 211.895 51.075 212.065 51.245 ;
        RECT 212.355 51.075 212.525 51.245 ;
        RECT 212.815 51.075 212.985 51.245 ;
        RECT 213.275 51.075 213.445 51.245 ;
        RECT 213.735 51.075 213.905 51.245 ;
        RECT 214.195 51.075 214.365 51.245 ;
        RECT 214.655 51.075 214.825 51.245 ;
        RECT 215.115 51.075 215.285 51.245 ;
        RECT 215.575 51.075 215.745 51.245 ;
        RECT 216.035 51.075 216.205 51.245 ;
        RECT 216.495 51.075 216.665 51.245 ;
        RECT 216.955 51.075 217.125 51.245 ;
        RECT 217.415 51.075 217.585 51.245 ;
        RECT 217.875 51.075 218.045 51.245 ;
        RECT 218.335 51.075 218.505 51.245 ;
        RECT 218.795 51.075 218.965 51.245 ;
        RECT 219.255 51.075 219.425 51.245 ;
        RECT 219.715 51.075 219.885 51.245 ;
        RECT 220.175 51.075 220.345 51.245 ;
        RECT 220.635 51.075 220.805 51.245 ;
        RECT 221.095 51.075 221.265 51.245 ;
        RECT 221.555 51.075 221.725 51.245 ;
        RECT 222.015 51.075 222.185 51.245 ;
        RECT 222.475 51.075 222.645 51.245 ;
        RECT 222.935 51.075 223.105 51.245 ;
        RECT 223.395 51.075 223.565 51.245 ;
        RECT 223.855 51.075 224.025 51.245 ;
        RECT 224.315 51.075 224.485 51.245 ;
        RECT 224.775 51.075 224.945 51.245 ;
        RECT 225.235 51.075 225.405 51.245 ;
        RECT 225.695 51.075 225.865 51.245 ;
        RECT 226.155 51.075 226.325 51.245 ;
        RECT 226.615 51.075 226.785 51.245 ;
        RECT 227.075 51.075 227.245 51.245 ;
        RECT 227.535 51.075 227.705 51.245 ;
        RECT 227.995 51.075 228.165 51.245 ;
        RECT 228.455 51.075 228.625 51.245 ;
        RECT 228.915 51.075 229.085 51.245 ;
        RECT 229.375 51.075 229.545 51.245 ;
        RECT 229.835 51.075 230.005 51.245 ;
        RECT 230.295 51.075 230.465 51.245 ;
        RECT 230.755 51.075 230.925 51.245 ;
        RECT 231.215 51.075 231.385 51.245 ;
        RECT 231.675 51.075 231.845 51.245 ;
        RECT 232.135 51.075 232.305 51.245 ;
        RECT 232.595 51.075 232.765 51.245 ;
        RECT 233.055 51.075 233.225 51.245 ;
        RECT 233.515 51.075 233.685 51.245 ;
        RECT 233.975 51.075 234.145 51.245 ;
        RECT 234.435 51.075 234.605 51.245 ;
        RECT 234.895 51.075 235.065 51.245 ;
        RECT 235.355 51.075 235.525 51.245 ;
        RECT 235.815 51.075 235.985 51.245 ;
        RECT 236.275 51.075 236.445 51.245 ;
        RECT 236.735 51.075 236.905 51.245 ;
        RECT 237.195 51.075 237.365 51.245 ;
        RECT 237.655 51.075 237.825 51.245 ;
        RECT 238.115 51.075 238.285 51.245 ;
        RECT 238.575 51.075 238.745 51.245 ;
        RECT 239.035 51.075 239.205 51.245 ;
        RECT 239.495 51.075 239.665 51.245 ;
        RECT 239.955 51.075 240.125 51.245 ;
        RECT 240.415 51.075 240.585 51.245 ;
        RECT 240.875 51.075 241.045 51.245 ;
        RECT 241.335 51.075 241.505 51.245 ;
        RECT 241.795 51.075 241.965 51.245 ;
        RECT 242.255 51.075 242.425 51.245 ;
        RECT 242.715 51.075 242.885 51.245 ;
        RECT 243.175 51.075 243.345 51.245 ;
        RECT 243.635 51.075 243.805 51.245 ;
        RECT 244.095 51.075 244.265 51.245 ;
        RECT 244.555 51.075 244.725 51.245 ;
        RECT 245.015 51.075 245.185 51.245 ;
        RECT 245.475 51.075 245.645 51.245 ;
        RECT 245.935 51.075 246.105 51.245 ;
        RECT 246.395 51.075 246.565 51.245 ;
        RECT 246.855 51.075 247.025 51.245 ;
        RECT 247.315 51.075 247.485 51.245 ;
        RECT 247.775 51.075 247.945 51.245 ;
        RECT 248.235 51.075 248.405 51.245 ;
        RECT 248.695 51.075 248.865 51.245 ;
        RECT 249.155 51.075 249.325 51.245 ;
        RECT 249.615 51.075 249.785 51.245 ;
        RECT 250.075 51.075 250.245 51.245 ;
        RECT 250.535 51.075 250.705 51.245 ;
        RECT 250.995 51.075 251.165 51.245 ;
        RECT 251.455 51.075 251.625 51.245 ;
        RECT 251.915 51.075 252.085 51.245 ;
        RECT 252.375 51.075 252.545 51.245 ;
        RECT 252.835 51.075 253.005 51.245 ;
        RECT 253.295 51.075 253.465 51.245 ;
        RECT 253.755 51.075 253.925 51.245 ;
        RECT 254.215 51.075 254.385 51.245 ;
        RECT 254.675 51.075 254.845 51.245 ;
        RECT 255.135 51.075 255.305 51.245 ;
        RECT 255.595 51.075 255.765 51.245 ;
        RECT 256.055 51.075 256.225 51.245 ;
        RECT 256.515 51.075 256.685 51.245 ;
        RECT 256.975 51.075 257.145 51.245 ;
        RECT 257.435 51.075 257.605 51.245 ;
        RECT 257.895 51.075 258.065 51.245 ;
        RECT 258.355 51.075 258.525 51.245 ;
        RECT 258.815 51.075 258.985 51.245 ;
        RECT 259.275 51.075 259.445 51.245 ;
        RECT 259.735 51.075 259.905 51.245 ;
        RECT 260.195 51.075 260.365 51.245 ;
        RECT 260.655 51.075 260.825 51.245 ;
        RECT 261.115 51.075 261.285 51.245 ;
        RECT 261.575 51.075 261.745 51.245 ;
        RECT 262.035 51.075 262.205 51.245 ;
        RECT 262.495 51.075 262.665 51.245 ;
        RECT 262.955 51.075 263.125 51.245 ;
        RECT 263.415 51.075 263.585 51.245 ;
        RECT 263.875 51.075 264.045 51.245 ;
        RECT 264.335 51.075 264.505 51.245 ;
        RECT 264.795 51.075 264.965 51.245 ;
        RECT 265.255 51.075 265.425 51.245 ;
        RECT 265.715 51.075 265.885 51.245 ;
        RECT 266.175 51.075 266.345 51.245 ;
        RECT 266.635 51.075 266.805 51.245 ;
        RECT 267.095 51.075 267.265 51.245 ;
        RECT 267.555 51.075 267.725 51.245 ;
        RECT 268.015 51.075 268.185 51.245 ;
        RECT 268.475 51.075 268.645 51.245 ;
        RECT 268.935 51.075 269.105 51.245 ;
        RECT 269.395 51.075 269.565 51.245 ;
        RECT 269.855 51.075 270.025 51.245 ;
        RECT 270.315 51.075 270.485 51.245 ;
        RECT 270.775 51.075 270.945 51.245 ;
        RECT 271.235 51.075 271.405 51.245 ;
        RECT 271.695 51.075 271.865 51.245 ;
        RECT 272.155 51.075 272.325 51.245 ;
        RECT 272.615 51.075 272.785 51.245 ;
        RECT 273.075 51.075 273.245 51.245 ;
        RECT 273.535 51.075 273.705 51.245 ;
        RECT 273.995 51.075 274.165 51.245 ;
        RECT 274.455 51.075 274.625 51.245 ;
        RECT 274.915 51.075 275.085 51.245 ;
        RECT 275.375 51.075 275.545 51.245 ;
        RECT 275.835 51.075 276.005 51.245 ;
        RECT 276.295 51.075 276.465 51.245 ;
        RECT 276.755 51.075 276.925 51.245 ;
        RECT 277.215 51.075 277.385 51.245 ;
        RECT 277.675 51.075 277.845 51.245 ;
        RECT 278.135 51.075 278.305 51.245 ;
        RECT 278.595 51.075 278.765 51.245 ;
        RECT 279.055 51.075 279.225 51.245 ;
        RECT 279.515 51.075 279.685 51.245 ;
        RECT 279.975 51.075 280.145 51.245 ;
        RECT 280.435 51.075 280.605 51.245 ;
        RECT 280.895 51.075 281.065 51.245 ;
        RECT 281.355 51.075 281.525 51.245 ;
        RECT 281.815 51.075 281.985 51.245 ;
        RECT 282.275 51.075 282.445 51.245 ;
        RECT 282.735 51.075 282.905 51.245 ;
        RECT 283.195 51.075 283.365 51.245 ;
        RECT 283.655 51.075 283.825 51.245 ;
        RECT 284.115 51.075 284.285 51.245 ;
        RECT 284.575 51.075 284.745 51.245 ;
        RECT 285.035 51.075 285.205 51.245 ;
        RECT 285.495 51.075 285.665 51.245 ;
        RECT 285.955 51.075 286.125 51.245 ;
        RECT 286.415 51.075 286.585 51.245 ;
        RECT 286.875 51.075 287.045 51.245 ;
        RECT 287.335 51.075 287.505 51.245 ;
        RECT 287.795 51.075 287.965 51.245 ;
        RECT 288.255 51.075 288.425 51.245 ;
        RECT 288.715 51.075 288.885 51.245 ;
        RECT 289.175 51.075 289.345 51.245 ;
        RECT 289.635 51.075 289.805 51.245 ;
        RECT 290.095 51.075 290.265 51.245 ;
        RECT 290.555 51.075 290.725 51.245 ;
        RECT 291.015 51.075 291.185 51.245 ;
        RECT 291.475 51.075 291.645 51.245 ;
        RECT 291.935 51.075 292.105 51.245 ;
        RECT 292.395 51.075 292.565 51.245 ;
        RECT 292.855 51.075 293.025 51.245 ;
        RECT 293.315 51.075 293.485 51.245 ;
        RECT 293.775 51.075 293.945 51.245 ;
        RECT 294.235 51.075 294.405 51.245 ;
        RECT 294.695 51.075 294.865 51.245 ;
        RECT 295.155 51.075 295.325 51.245 ;
        RECT 295.615 51.075 295.785 51.245 ;
        RECT 296.075 51.075 296.245 51.245 ;
        RECT 296.535 51.075 296.705 51.245 ;
        RECT 296.995 51.075 297.165 51.245 ;
        RECT 297.455 51.075 297.625 51.245 ;
        RECT 297.915 51.075 298.085 51.245 ;
        RECT 298.375 51.075 298.545 51.245 ;
        RECT 298.835 51.075 299.005 51.245 ;
        RECT 299.295 51.075 299.465 51.245 ;
        RECT 299.755 51.075 299.925 51.245 ;
        RECT 300.215 51.075 300.385 51.245 ;
        RECT 300.675 51.075 300.845 51.245 ;
        RECT 301.135 51.075 301.305 51.245 ;
        RECT 301.595 51.075 301.765 51.245 ;
        RECT 302.055 51.075 302.225 51.245 ;
        RECT 302.515 51.075 302.685 51.245 ;
        RECT 302.975 51.075 303.145 51.245 ;
        RECT 303.435 51.075 303.605 51.245 ;
        RECT 303.895 51.075 304.065 51.245 ;
        RECT 304.355 51.075 304.525 51.245 ;
        RECT 304.815 51.075 304.985 51.245 ;
        RECT 305.275 51.075 305.445 51.245 ;
        RECT 305.735 51.075 305.905 51.245 ;
        RECT 306.195 51.075 306.365 51.245 ;
        RECT 306.655 51.075 306.825 51.245 ;
        RECT 307.115 51.075 307.285 51.245 ;
        RECT 307.575 51.075 307.745 51.245 ;
        RECT 308.035 51.075 308.205 51.245 ;
        RECT 308.495 51.075 308.665 51.245 ;
        RECT 308.955 51.075 309.125 51.245 ;
        RECT 309.415 51.075 309.585 51.245 ;
        RECT 309.875 51.075 310.045 51.245 ;
        RECT 310.335 51.075 310.505 51.245 ;
        RECT 310.795 51.075 310.965 51.245 ;
        RECT 311.255 51.075 311.425 51.245 ;
        RECT 311.715 51.075 311.885 51.245 ;
        RECT 312.175 51.075 312.345 51.245 ;
        RECT 312.635 51.075 312.805 51.245 ;
        RECT 313.095 51.075 313.265 51.245 ;
        RECT 313.555 51.075 313.725 51.245 ;
        RECT 314.015 51.075 314.185 51.245 ;
        RECT 314.475 51.075 314.645 51.245 ;
        RECT 314.935 51.075 315.105 51.245 ;
        RECT 315.395 51.075 315.565 51.245 ;
        RECT 315.855 51.075 316.025 51.245 ;
        RECT 316.315 51.075 316.485 51.245 ;
        RECT 316.775 51.075 316.945 51.245 ;
        RECT 317.235 51.075 317.405 51.245 ;
        RECT 317.695 51.075 317.865 51.245 ;
        RECT 318.155 51.075 318.325 51.245 ;
        RECT 318.615 51.075 318.785 51.245 ;
        RECT 319.075 51.075 319.245 51.245 ;
        RECT 319.535 51.075 319.705 51.245 ;
        RECT 319.995 51.075 320.165 51.245 ;
        RECT 320.455 51.075 320.625 51.245 ;
        RECT 320.915 51.075 321.085 51.245 ;
        RECT 321.375 51.075 321.545 51.245 ;
        RECT 321.835 51.075 322.005 51.245 ;
        RECT 322.295 51.075 322.465 51.245 ;
        RECT 322.755 51.075 322.925 51.245 ;
        RECT 323.215 51.075 323.385 51.245 ;
        RECT 323.675 51.075 323.845 51.245 ;
        RECT 324.135 51.075 324.305 51.245 ;
        RECT 324.595 51.075 324.765 51.245 ;
        RECT 325.055 51.075 325.225 51.245 ;
        RECT 325.515 51.075 325.685 51.245 ;
        RECT 325.975 51.075 326.145 51.245 ;
        RECT 326.435 51.075 326.605 51.245 ;
        RECT 326.895 51.075 327.065 51.245 ;
        RECT 327.355 51.075 327.525 51.245 ;
        RECT 327.815 51.075 327.985 51.245 ;
        RECT 328.275 51.075 328.445 51.245 ;
        RECT 328.735 51.075 328.905 51.245 ;
        RECT 329.195 51.075 329.365 51.245 ;
        RECT 329.655 51.075 329.825 51.245 ;
        RECT 330.115 51.075 330.285 51.245 ;
        RECT 330.575 51.075 330.745 51.245 ;
        RECT 331.035 51.075 331.205 51.245 ;
        RECT 331.495 51.075 331.665 51.245 ;
        RECT 331.955 51.075 332.125 51.245 ;
        RECT 332.415 51.075 332.585 51.245 ;
        RECT 332.875 51.075 333.045 51.245 ;
        RECT 333.335 51.075 333.505 51.245 ;
        RECT 333.795 51.075 333.965 51.245 ;
        RECT 334.255 51.075 334.425 51.245 ;
        RECT 334.715 51.075 334.885 51.245 ;
        RECT 335.175 51.075 335.345 51.245 ;
        RECT 335.635 51.075 335.805 51.245 ;
        RECT 336.095 51.075 336.265 51.245 ;
        RECT 336.555 51.075 336.725 51.245 ;
        RECT 337.015 51.075 337.185 51.245 ;
        RECT 337.475 51.075 337.645 51.245 ;
        RECT 337.935 51.075 338.105 51.245 ;
        RECT 338.395 51.075 338.565 51.245 ;
        RECT 338.855 51.075 339.025 51.245 ;
        RECT 339.315 51.075 339.485 51.245 ;
        RECT 339.775 51.075 339.945 51.245 ;
        RECT 340.235 51.075 340.405 51.245 ;
        RECT 340.695 51.075 340.865 51.245 ;
        RECT 341.155 51.075 341.325 51.245 ;
        RECT 341.615 51.075 341.785 51.245 ;
        RECT 342.075 51.075 342.245 51.245 ;
        RECT 342.535 51.075 342.705 51.245 ;
        RECT 342.995 51.075 343.165 51.245 ;
        RECT 343.455 51.075 343.625 51.245 ;
        RECT 343.915 51.075 344.085 51.245 ;
        RECT 344.375 51.075 344.545 51.245 ;
        RECT 344.835 51.075 345.005 51.245 ;
        RECT 345.295 51.075 345.465 51.245 ;
        RECT 345.755 51.075 345.925 51.245 ;
        RECT 346.215 51.075 346.385 51.245 ;
        RECT 346.675 51.075 346.845 51.245 ;
        RECT 347.135 51.075 347.305 51.245 ;
        RECT 347.595 51.075 347.765 51.245 ;
        RECT 348.055 51.075 348.225 51.245 ;
        RECT 348.515 51.075 348.685 51.245 ;
        RECT 348.975 51.075 349.145 51.245 ;
        RECT 349.435 51.075 349.605 51.245 ;
        RECT 349.895 51.075 350.065 51.245 ;
        RECT 350.355 51.075 350.525 51.245 ;
        RECT 350.815 51.075 350.985 51.245 ;
        RECT 351.275 51.075 351.445 51.245 ;
        RECT 351.735 51.075 351.905 51.245 ;
        RECT 352.195 51.075 352.365 51.245 ;
        RECT 352.655 51.075 352.825 51.245 ;
        RECT 353.115 51.075 353.285 51.245 ;
        RECT 353.575 51.075 353.745 51.245 ;
        RECT 354.035 51.075 354.205 51.245 ;
        RECT 354.495 51.075 354.665 51.245 ;
        RECT 354.955 51.075 355.125 51.245 ;
        RECT 355.415 51.075 355.585 51.245 ;
        RECT 355.875 51.075 356.045 51.245 ;
        RECT 356.335 51.075 356.505 51.245 ;
        RECT 356.795 51.075 356.965 51.245 ;
        RECT 357.255 51.075 357.425 51.245 ;
        RECT 357.715 51.075 357.885 51.245 ;
        RECT 358.175 51.075 358.345 51.245 ;
        RECT 358.635 51.075 358.805 51.245 ;
        RECT 359.095 51.075 359.265 51.245 ;
        RECT 359.555 51.075 359.725 51.245 ;
        RECT 360.015 51.075 360.185 51.245 ;
        RECT 360.475 51.075 360.645 51.245 ;
        RECT 360.935 51.075 361.105 51.245 ;
        RECT 361.395 51.075 361.565 51.245 ;
        RECT 361.855 51.075 362.025 51.245 ;
        RECT 362.315 51.075 362.485 51.245 ;
        RECT 362.775 51.075 362.945 51.245 ;
        RECT 363.235 51.075 363.405 51.245 ;
        RECT 363.695 51.075 363.865 51.245 ;
        RECT 364.155 51.075 364.325 51.245 ;
        RECT 364.615 51.075 364.785 51.245 ;
        RECT 365.075 51.075 365.245 51.245 ;
        RECT 365.535 51.075 365.705 51.245 ;
        RECT 365.995 51.075 366.165 51.245 ;
        RECT 366.455 51.075 366.625 51.245 ;
        RECT 366.915 51.075 367.085 51.245 ;
        RECT 367.375 51.075 367.545 51.245 ;
        RECT 367.835 51.075 368.005 51.245 ;
        RECT 368.295 51.075 368.465 51.245 ;
        RECT 368.755 51.075 368.925 51.245 ;
        RECT 369.215 51.075 369.385 51.245 ;
        RECT 369.675 51.075 369.845 51.245 ;
        RECT 370.135 51.075 370.305 51.245 ;
        RECT 370.595 51.075 370.765 51.245 ;
        RECT 371.055 51.075 371.225 51.245 ;
        RECT 371.515 51.075 371.685 51.245 ;
        RECT 371.975 51.075 372.145 51.245 ;
        RECT 372.435 51.075 372.605 51.245 ;
        RECT 372.895 51.075 373.065 51.245 ;
        RECT 373.355 51.075 373.525 51.245 ;
        RECT 373.815 51.075 373.985 51.245 ;
        RECT 374.275 51.075 374.445 51.245 ;
        RECT 374.735 51.075 374.905 51.245 ;
        RECT 375.195 51.075 375.365 51.245 ;
        RECT 375.655 51.075 375.825 51.245 ;
        RECT 376.115 51.075 376.285 51.245 ;
        RECT 376.575 51.075 376.745 51.245 ;
        RECT 377.035 51.075 377.205 51.245 ;
        RECT 377.495 51.075 377.665 51.245 ;
        RECT 377.955 51.075 378.125 51.245 ;
        RECT 378.415 51.075 378.585 51.245 ;
        RECT 378.875 51.075 379.045 51.245 ;
        RECT 379.335 51.075 379.505 51.245 ;
        RECT 379.795 51.075 379.965 51.245 ;
        RECT 380.255 51.075 380.425 51.245 ;
        RECT 380.715 51.075 380.885 51.245 ;
        RECT 381.175 51.075 381.345 51.245 ;
        RECT 381.635 51.075 381.805 51.245 ;
        RECT 382.095 51.075 382.265 51.245 ;
        RECT 382.555 51.075 382.725 51.245 ;
        RECT 383.015 51.075 383.185 51.245 ;
        RECT 383.475 51.075 383.645 51.245 ;
        RECT 383.935 51.075 384.105 51.245 ;
        RECT 384.395 51.075 384.565 51.245 ;
        RECT 384.855 51.075 385.025 51.245 ;
        RECT 385.315 51.075 385.485 51.245 ;
        RECT 385.775 51.075 385.945 51.245 ;
        RECT 386.235 51.075 386.405 51.245 ;
        RECT 386.695 51.075 386.865 51.245 ;
        RECT 387.155 51.075 387.325 51.245 ;
        RECT 387.615 51.075 387.785 51.245 ;
        RECT 388.075 51.075 388.245 51.245 ;
        RECT 388.535 51.075 388.705 51.245 ;
        RECT 388.995 51.075 389.165 51.245 ;
        RECT 389.455 51.075 389.625 51.245 ;
        RECT 389.915 51.075 390.085 51.245 ;
        RECT 390.375 51.075 390.545 51.245 ;
        RECT 390.835 51.075 391.005 51.245 ;
        RECT 391.295 51.075 391.465 51.245 ;
        RECT 391.755 51.075 391.925 51.245 ;
        RECT 392.215 51.075 392.385 51.245 ;
        RECT 392.675 51.075 392.845 51.245 ;
        RECT 393.135 51.075 393.305 51.245 ;
        RECT 393.595 51.075 393.765 51.245 ;
        RECT 394.055 51.075 394.225 51.245 ;
        RECT 394.515 51.075 394.685 51.245 ;
        RECT 394.975 51.075 395.145 51.245 ;
        RECT 395.435 51.075 395.605 51.245 ;
        RECT 395.895 51.075 396.065 51.245 ;
        RECT 396.355 51.075 396.525 51.245 ;
        RECT 396.815 51.075 396.985 51.245 ;
        RECT 397.275 51.075 397.445 51.245 ;
        RECT 397.735 51.075 397.905 51.245 ;
        RECT 398.195 51.075 398.365 51.245 ;
        RECT 398.655 51.075 398.825 51.245 ;
        RECT 399.115 51.075 399.285 51.245 ;
        RECT 399.575 51.075 399.745 51.245 ;
        RECT 400.035 51.075 400.205 51.245 ;
        RECT 400.495 51.075 400.665 51.245 ;
        RECT 400.955 51.075 401.125 51.245 ;
        RECT 401.415 51.075 401.585 51.245 ;
        RECT 401.875 51.075 402.045 51.245 ;
        RECT 402.335 51.075 402.505 51.245 ;
        RECT 402.795 51.075 402.965 51.245 ;
        RECT 403.255 51.075 403.425 51.245 ;
        RECT 403.715 51.075 403.885 51.245 ;
        RECT 404.175 51.075 404.345 51.245 ;
        RECT 404.635 51.075 404.805 51.245 ;
        RECT 405.095 51.075 405.265 51.245 ;
        RECT 405.555 51.075 405.725 51.245 ;
        RECT 406.015 51.075 406.185 51.245 ;
        RECT 406.475 51.075 406.645 51.245 ;
        RECT 406.935 51.075 407.105 51.245 ;
        RECT 407.395 51.075 407.565 51.245 ;
        RECT 407.855 51.075 408.025 51.245 ;
        RECT 408.315 51.075 408.485 51.245 ;
        RECT 408.775 51.075 408.945 51.245 ;
        RECT 409.235 51.075 409.405 51.245 ;
        RECT 409.695 51.075 409.865 51.245 ;
        RECT 410.155 51.075 410.325 51.245 ;
        RECT 410.615 51.075 410.785 51.245 ;
        RECT 411.075 51.075 411.245 51.245 ;
        RECT 411.535 51.075 411.705 51.245 ;
        RECT 411.995 51.075 412.165 51.245 ;
        RECT 412.455 51.075 412.625 51.245 ;
        RECT 412.915 51.075 413.085 51.245 ;
        RECT 413.375 51.075 413.545 51.245 ;
        RECT 413.835 51.075 414.005 51.245 ;
        RECT 414.295 51.075 414.465 51.245 ;
        RECT 414.755 51.075 414.925 51.245 ;
        RECT 415.215 51.075 415.385 51.245 ;
        RECT 415.675 51.075 415.845 51.245 ;
        RECT 416.135 51.075 416.305 51.245 ;
        RECT 416.595 51.075 416.765 51.245 ;
        RECT 417.055 51.075 417.225 51.245 ;
        RECT 417.515 51.075 417.685 51.245 ;
        RECT 417.975 51.075 418.145 51.245 ;
        RECT 418.435 51.075 418.605 51.245 ;
        RECT 418.895 51.075 419.065 51.245 ;
        RECT 419.355 51.075 419.525 51.245 ;
        RECT 419.815 51.075 419.985 51.245 ;
        RECT 420.275 51.075 420.445 51.245 ;
        RECT 420.735 51.075 420.905 51.245 ;
        RECT 421.195 51.075 421.365 51.245 ;
        RECT 421.655 51.075 421.825 51.245 ;
        RECT 422.115 51.075 422.285 51.245 ;
        RECT 422.575 51.075 422.745 51.245 ;
        RECT 423.035 51.075 423.205 51.245 ;
        RECT 423.495 51.075 423.665 51.245 ;
        RECT 423.955 51.075 424.125 51.245 ;
        RECT 424.415 51.075 424.585 51.245 ;
        RECT 424.875 51.075 425.045 51.245 ;
        RECT 425.335 51.075 425.505 51.245 ;
        RECT 425.795 51.075 425.965 51.245 ;
        RECT 426.255 51.075 426.425 51.245 ;
        RECT 426.715 51.075 426.885 51.245 ;
        RECT 427.175 51.075 427.345 51.245 ;
        RECT 427.635 51.075 427.805 51.245 ;
        RECT 428.095 51.075 428.265 51.245 ;
        RECT 428.555 51.075 428.725 51.245 ;
        RECT 429.015 51.075 429.185 51.245 ;
        RECT 429.475 51.075 429.645 51.245 ;
        RECT 429.935 51.075 430.105 51.245 ;
        RECT 430.395 51.075 430.565 51.245 ;
        RECT 430.855 51.075 431.025 51.245 ;
        RECT 431.315 51.075 431.485 51.245 ;
        RECT 431.775 51.075 431.945 51.245 ;
        RECT 432.235 51.075 432.405 51.245 ;
        RECT 432.695 51.075 432.865 51.245 ;
        RECT 433.155 51.075 433.325 51.245 ;
        RECT 433.615 51.075 433.785 51.245 ;
        RECT 434.075 51.075 434.245 51.245 ;
        RECT 434.535 51.075 434.705 51.245 ;
        RECT 434.995 51.075 435.165 51.245 ;
        RECT 435.455 51.075 435.625 51.245 ;
        RECT 435.915 51.075 436.085 51.245 ;
        RECT 436.375 51.075 436.545 51.245 ;
        RECT 436.835 51.075 437.005 51.245 ;
        RECT 437.295 51.075 437.465 51.245 ;
        RECT 437.755 51.075 437.925 51.245 ;
        RECT 438.215 51.075 438.385 51.245 ;
        RECT 438.675 51.075 438.845 51.245 ;
        RECT 439.135 51.075 439.305 51.245 ;
        RECT 439.595 51.075 439.765 51.245 ;
        RECT 440.055 51.075 440.225 51.245 ;
        RECT 440.515 51.075 440.685 51.245 ;
        RECT 440.975 51.075 441.145 51.245 ;
        RECT 441.435 51.075 441.605 51.245 ;
        RECT 441.895 51.075 442.065 51.245 ;
        RECT 442.355 51.075 442.525 51.245 ;
        RECT 442.815 51.075 442.985 51.245 ;
        RECT 443.275 51.075 443.445 51.245 ;
        RECT 443.735 51.075 443.905 51.245 ;
        RECT 444.195 51.075 444.365 51.245 ;
        RECT 444.655 51.075 444.825 51.245 ;
        RECT 445.115 51.075 445.285 51.245 ;
        RECT 445.575 51.075 445.745 51.245 ;
        RECT 446.035 51.075 446.205 51.245 ;
        RECT 446.495 51.075 446.665 51.245 ;
        RECT 446.955 51.075 447.125 51.245 ;
        RECT 447.415 51.075 447.585 51.245 ;
        RECT 447.875 51.075 448.045 51.245 ;
        RECT 448.335 51.075 448.505 51.245 ;
        RECT 448.795 51.075 448.965 51.245 ;
        RECT 449.255 51.075 449.425 51.245 ;
        RECT 449.715 51.075 449.885 51.245 ;
        RECT 450.175 51.075 450.345 51.245 ;
        RECT 450.635 51.075 450.805 51.245 ;
        RECT 451.095 51.075 451.265 51.245 ;
        RECT 451.555 51.075 451.725 51.245 ;
        RECT 452.015 51.075 452.185 51.245 ;
        RECT 452.475 51.075 452.645 51.245 ;
        RECT 452.935 51.075 453.105 51.245 ;
        RECT 453.395 51.075 453.565 51.245 ;
        RECT 453.855 51.075 454.025 51.245 ;
        RECT 454.315 51.075 454.485 51.245 ;
        RECT 454.775 51.075 454.945 51.245 ;
        RECT 455.235 51.075 455.405 51.245 ;
        RECT 455.695 51.075 455.865 51.245 ;
        RECT 456.155 51.075 456.325 51.245 ;
        RECT 456.615 51.075 456.785 51.245 ;
        RECT 457.075 51.075 457.245 51.245 ;
        RECT 457.535 51.075 457.705 51.245 ;
        RECT 457.995 51.075 458.165 51.245 ;
        RECT 458.455 51.075 458.625 51.245 ;
        RECT 458.915 51.075 459.085 51.245 ;
        RECT 459.375 51.075 459.545 51.245 ;
        RECT 459.835 51.075 460.005 51.245 ;
        RECT 460.295 51.075 460.465 51.245 ;
        RECT 460.755 51.075 460.925 51.245 ;
        RECT 461.215 51.075 461.385 51.245 ;
        RECT 461.675 51.075 461.845 51.245 ;
        RECT 462.135 51.075 462.305 51.245 ;
        RECT 462.595 51.075 462.765 51.245 ;
        RECT 463.055 51.075 463.225 51.245 ;
        RECT 463.515 51.075 463.685 51.245 ;
        RECT 463.975 51.075 464.145 51.245 ;
        RECT 464.435 51.075 464.605 51.245 ;
        RECT 464.895 51.075 465.065 51.245 ;
        RECT 465.355 51.075 465.525 51.245 ;
        RECT 465.815 51.075 465.985 51.245 ;
        RECT 466.275 51.075 466.445 51.245 ;
        RECT 466.735 51.075 466.905 51.245 ;
        RECT 467.195 51.075 467.365 51.245 ;
        RECT 467.655 51.075 467.825 51.245 ;
        RECT 468.115 51.075 468.285 51.245 ;
        RECT 468.575 51.075 468.745 51.245 ;
        RECT 469.035 51.075 469.205 51.245 ;
        RECT 469.495 51.075 469.665 51.245 ;
        RECT 469.955 51.075 470.125 51.245 ;
        RECT 470.415 51.075 470.585 51.245 ;
        RECT 470.875 51.075 471.045 51.245 ;
        RECT 471.335 51.075 471.505 51.245 ;
        RECT 471.795 51.075 471.965 51.245 ;
        RECT 472.255 51.075 472.425 51.245 ;
        RECT 472.715 51.075 472.885 51.245 ;
        RECT 473.175 51.075 473.345 51.245 ;
        RECT 473.635 51.075 473.805 51.245 ;
        RECT 474.095 51.075 474.265 51.245 ;
        RECT 474.555 51.075 474.725 51.245 ;
        RECT 475.015 51.075 475.185 51.245 ;
        RECT 475.475 51.075 475.645 51.245 ;
        RECT 475.935 51.075 476.105 51.245 ;
        RECT 476.395 51.075 476.565 51.245 ;
        RECT 476.855 51.075 477.025 51.245 ;
        RECT 477.315 51.075 477.485 51.245 ;
        RECT 477.775 51.075 477.945 51.245 ;
        RECT 478.235 51.075 478.405 51.245 ;
        RECT 478.695 51.075 478.865 51.245 ;
        RECT 479.155 51.075 479.325 51.245 ;
        RECT 479.615 51.075 479.785 51.245 ;
        RECT 480.075 51.075 480.245 51.245 ;
        RECT 480.535 51.075 480.705 51.245 ;
        RECT 480.995 51.075 481.165 51.245 ;
        RECT 481.455 51.075 481.625 51.245 ;
        RECT 481.915 51.075 482.085 51.245 ;
        RECT 482.375 51.075 482.545 51.245 ;
        RECT 482.835 51.075 483.005 51.245 ;
        RECT 483.295 51.075 483.465 51.245 ;
        RECT 483.755 51.075 483.925 51.245 ;
        RECT 484.215 51.075 484.385 51.245 ;
        RECT 484.675 51.075 484.845 51.245 ;
        RECT 485.135 51.075 485.305 51.245 ;
        RECT 485.595 51.075 485.765 51.245 ;
        RECT 486.055 51.075 486.225 51.245 ;
        RECT 486.515 51.075 486.685 51.245 ;
        RECT 486.975 51.075 487.145 51.245 ;
        RECT 487.435 51.075 487.605 51.245 ;
        RECT 487.895 51.075 488.065 51.245 ;
        RECT 488.355 51.075 488.525 51.245 ;
        RECT 488.815 51.075 488.985 51.245 ;
        RECT 489.275 51.075 489.445 51.245 ;
        RECT 489.735 51.075 489.905 51.245 ;
        RECT 490.195 51.075 490.365 51.245 ;
        RECT 490.655 51.075 490.825 51.245 ;
        RECT 491.115 51.075 491.285 51.245 ;
        RECT 491.575 51.075 491.745 51.245 ;
        RECT 492.035 51.075 492.205 51.245 ;
        RECT 492.495 51.075 492.665 51.245 ;
        RECT 492.955 51.075 493.125 51.245 ;
        RECT 493.415 51.075 493.585 51.245 ;
        RECT 493.875 51.075 494.045 51.245 ;
        RECT 494.335 51.075 494.505 51.245 ;
        RECT 494.795 51.075 494.965 51.245 ;
        RECT 495.255 51.075 495.425 51.245 ;
        RECT 495.715 51.075 495.885 51.245 ;
        RECT 496.175 51.075 496.345 51.245 ;
        RECT 496.635 51.075 496.805 51.245 ;
        RECT 497.095 51.075 497.265 51.245 ;
        RECT 497.555 51.075 497.725 51.245 ;
        RECT 498.015 51.075 498.185 51.245 ;
        RECT 498.475 51.075 498.645 51.245 ;
        RECT 498.935 51.075 499.105 51.245 ;
        RECT 499.395 51.075 499.565 51.245 ;
        RECT 499.855 51.075 500.025 51.245 ;
        RECT 500.315 51.075 500.485 51.245 ;
        RECT 500.775 51.075 500.945 51.245 ;
        RECT 501.235 51.075 501.405 51.245 ;
        RECT 501.695 51.075 501.865 51.245 ;
        RECT 502.155 51.075 502.325 51.245 ;
        RECT 502.615 51.075 502.785 51.245 ;
        RECT 503.075 51.075 503.245 51.245 ;
        RECT 503.535 51.075 503.705 51.245 ;
        RECT 503.995 51.075 504.165 51.245 ;
        RECT 504.455 51.075 504.625 51.245 ;
        RECT 504.915 51.075 505.085 51.245 ;
        RECT 505.375 51.075 505.545 51.245 ;
        RECT 505.835 51.075 506.005 51.245 ;
        RECT 506.295 51.075 506.465 51.245 ;
        RECT 506.755 51.075 506.925 51.245 ;
        RECT 507.215 51.075 507.385 51.245 ;
        RECT 507.675 51.075 507.845 51.245 ;
        RECT 508.135 51.075 508.305 51.245 ;
        RECT 508.595 51.075 508.765 51.245 ;
        RECT 509.055 51.075 509.225 51.245 ;
        RECT 509.515 51.075 509.685 51.245 ;
        RECT 509.975 51.075 510.145 51.245 ;
        RECT 510.435 51.075 510.605 51.245 ;
        RECT 510.895 51.075 511.065 51.245 ;
        RECT 511.355 51.075 511.525 51.245 ;
        RECT 511.815 51.075 511.985 51.245 ;
        RECT 512.275 51.075 512.445 51.245 ;
        RECT 512.735 51.075 512.905 51.245 ;
        RECT 513.195 51.075 513.365 51.245 ;
        RECT 513.655 51.075 513.825 51.245 ;
        RECT 514.115 51.075 514.285 51.245 ;
        RECT 514.575 51.075 514.745 51.245 ;
        RECT 515.035 51.075 515.205 51.245 ;
        RECT 515.495 51.075 515.665 51.245 ;
        RECT 515.955 51.075 516.125 51.245 ;
        RECT 516.415 51.075 516.585 51.245 ;
        RECT 516.875 51.075 517.045 51.245 ;
        RECT 517.335 51.075 517.505 51.245 ;
        RECT 517.795 51.075 517.965 51.245 ;
        RECT 518.255 51.075 518.425 51.245 ;
        RECT 518.715 51.075 518.885 51.245 ;
        RECT 519.175 51.075 519.345 51.245 ;
        RECT 519.635 51.075 519.805 51.245 ;
        RECT 520.095 51.075 520.265 51.245 ;
        RECT 520.555 51.075 520.725 51.245 ;
        RECT 521.015 51.075 521.185 51.245 ;
        RECT 521.475 51.075 521.645 51.245 ;
        RECT 521.935 51.075 522.105 51.245 ;
        RECT 522.395 51.075 522.565 51.245 ;
        RECT 522.855 51.075 523.025 51.245 ;
        RECT 523.315 51.075 523.485 51.245 ;
        RECT 523.775 51.075 523.945 51.245 ;
        RECT 524.235 51.075 524.405 51.245 ;
        RECT 524.695 51.075 524.865 51.245 ;
        RECT 525.155 51.075 525.325 51.245 ;
        RECT 525.615 51.075 525.785 51.245 ;
        RECT 526.075 51.075 526.245 51.245 ;
        RECT 526.535 51.075 526.705 51.245 ;
        RECT 526.995 51.075 527.165 51.245 ;
        RECT 527.455 51.075 527.625 51.245 ;
        RECT 527.915 51.075 528.085 51.245 ;
        RECT 528.375 51.075 528.545 51.245 ;
        RECT 528.835 51.075 529.005 51.245 ;
        RECT 529.295 51.075 529.465 51.245 ;
        RECT 529.755 51.075 529.925 51.245 ;
        RECT 530.215 51.075 530.385 51.245 ;
        RECT 530.675 51.075 530.845 51.245 ;
        RECT 531.135 51.075 531.305 51.245 ;
        RECT 531.595 51.075 531.765 51.245 ;
        RECT 532.055 51.075 532.225 51.245 ;
        RECT 532.515 51.075 532.685 51.245 ;
        RECT 532.975 51.075 533.145 51.245 ;
        RECT 533.435 51.075 533.605 51.245 ;
        RECT 533.895 51.075 534.065 51.245 ;
        RECT 534.355 51.075 534.525 51.245 ;
        RECT 534.815 51.075 534.985 51.245 ;
        RECT 535.275 51.075 535.445 51.245 ;
        RECT 535.735 51.075 535.905 51.245 ;
        RECT 536.195 51.075 536.365 51.245 ;
        RECT 536.655 51.075 536.825 51.245 ;
        RECT 537.115 51.075 537.285 51.245 ;
        RECT 537.575 51.075 537.745 51.245 ;
        RECT 538.035 51.075 538.205 51.245 ;
        RECT 538.495 51.075 538.665 51.245 ;
        RECT 538.955 51.075 539.125 51.245 ;
        RECT 539.415 51.075 539.585 51.245 ;
        RECT 539.875 51.075 540.045 51.245 ;
        RECT 540.335 51.075 540.505 51.245 ;
        RECT 540.795 51.075 540.965 51.245 ;
        RECT 541.255 51.075 541.425 51.245 ;
        RECT 541.715 51.075 541.885 51.245 ;
        RECT 542.175 51.075 542.345 51.245 ;
        RECT 542.635 51.075 542.805 51.245 ;
        RECT 543.095 51.075 543.265 51.245 ;
        RECT 543.555 51.075 543.725 51.245 ;
        RECT 544.015 51.075 544.185 51.245 ;
        RECT 544.475 51.075 544.645 51.245 ;
        RECT 544.935 51.075 545.105 51.245 ;
        RECT 545.395 51.075 545.565 51.245 ;
        RECT 545.855 51.075 546.025 51.245 ;
        RECT 546.315 51.075 546.485 51.245 ;
        RECT 546.775 51.075 546.945 51.245 ;
        RECT 547.235 51.075 547.405 51.245 ;
        RECT 547.695 51.075 547.865 51.245 ;
        RECT 548.155 51.075 548.325 51.245 ;
        RECT 548.615 51.075 548.785 51.245 ;
        RECT 549.075 51.075 549.245 51.245 ;
        RECT 549.535 51.075 549.705 51.245 ;
        RECT 549.995 51.075 550.165 51.245 ;
        RECT 550.455 51.075 550.625 51.245 ;
        RECT 550.915 51.075 551.085 51.245 ;
        RECT 551.375 51.075 551.545 51.245 ;
        RECT 551.835 51.075 552.005 51.245 ;
        RECT 552.295 51.075 552.465 51.245 ;
        RECT 552.755 51.075 552.925 51.245 ;
        RECT 553.215 51.075 553.385 51.245 ;
        RECT 553.675 51.075 553.845 51.245 ;
        RECT 554.135 51.075 554.305 51.245 ;
        RECT 554.595 51.075 554.765 51.245 ;
        RECT 555.055 51.075 555.225 51.245 ;
        RECT 555.515 51.075 555.685 51.245 ;
        RECT 555.975 51.075 556.145 51.245 ;
        RECT 556.435 51.075 556.605 51.245 ;
        RECT 556.895 51.075 557.065 51.245 ;
        RECT 557.355 51.075 557.525 51.245 ;
        RECT 557.815 51.075 557.985 51.245 ;
        RECT 558.275 51.075 558.445 51.245 ;
        RECT 558.735 51.075 558.905 51.245 ;
        RECT 559.195 51.075 559.365 51.245 ;
        RECT 559.655 51.075 559.825 51.245 ;
        RECT 560.115 51.075 560.285 51.245 ;
        RECT 560.575 51.075 560.745 51.245 ;
        RECT 561.035 51.075 561.205 51.245 ;
        RECT 561.495 51.075 561.665 51.245 ;
        RECT 561.955 51.075 562.125 51.245 ;
        RECT 562.415 51.075 562.585 51.245 ;
        RECT 562.875 51.075 563.045 51.245 ;
        RECT 563.335 51.075 563.505 51.245 ;
        RECT 563.795 51.075 563.965 51.245 ;
        RECT 564.255 51.075 564.425 51.245 ;
        RECT 564.715 51.075 564.885 51.245 ;
        RECT 565.175 51.075 565.345 51.245 ;
        RECT 565.635 51.075 565.805 51.245 ;
        RECT 566.095 51.075 566.265 51.245 ;
        RECT 566.555 51.075 566.725 51.245 ;
        RECT 567.015 51.075 567.185 51.245 ;
        RECT 567.475 51.075 567.645 51.245 ;
        RECT 567.935 51.075 568.105 51.245 ;
        RECT 568.395 51.075 568.565 51.245 ;
        RECT 568.855 51.075 569.025 51.245 ;
        RECT 569.315 51.075 569.485 51.245 ;
        RECT 569.775 51.075 569.945 51.245 ;
        RECT 570.235 51.075 570.405 51.245 ;
        RECT 570.695 51.075 570.865 51.245 ;
        RECT 571.155 51.075 571.325 51.245 ;
        RECT 571.615 51.075 571.785 51.245 ;
        RECT 572.075 51.075 572.245 51.245 ;
        RECT 572.535 51.075 572.705 51.245 ;
        RECT 572.995 51.075 573.165 51.245 ;
        RECT 573.455 51.075 573.625 51.245 ;
        RECT 573.915 51.075 574.085 51.245 ;
        RECT 574.375 51.075 574.545 51.245 ;
        RECT 574.835 51.075 575.005 51.245 ;
        RECT 575.295 51.075 575.465 51.245 ;
        RECT 575.755 51.075 575.925 51.245 ;
        RECT 576.215 51.075 576.385 51.245 ;
        RECT 576.675 51.075 576.845 51.245 ;
        RECT 577.135 51.075 577.305 51.245 ;
        RECT 577.595 51.075 577.765 51.245 ;
        RECT 578.055 51.075 578.225 51.245 ;
        RECT 578.515 51.075 578.685 51.245 ;
        RECT 578.975 51.075 579.145 51.245 ;
        RECT 579.435 51.075 579.605 51.245 ;
        RECT 579.895 51.075 580.065 51.245 ;
        RECT 580.355 51.075 580.525 51.245 ;
        RECT 580.815 51.075 580.985 51.245 ;
        RECT 581.275 51.075 581.445 51.245 ;
        RECT 581.735 51.075 581.905 51.245 ;
        RECT 582.195 51.075 582.365 51.245 ;
        RECT 582.655 51.075 582.825 51.245 ;
        RECT 583.115 51.075 583.285 51.245 ;
        RECT 583.575 51.075 583.745 51.245 ;
        RECT 584.035 51.075 584.205 51.245 ;
        RECT 584.495 51.075 584.665 51.245 ;
        RECT 584.955 51.075 585.125 51.245 ;
        RECT 585.415 51.075 585.585 51.245 ;
        RECT 585.875 51.075 586.045 51.245 ;
        RECT 586.335 51.075 586.505 51.245 ;
        RECT 586.795 51.075 586.965 51.245 ;
        RECT 587.255 51.075 587.425 51.245 ;
        RECT 587.715 51.075 587.885 51.245 ;
        RECT 588.175 51.075 588.345 51.245 ;
        RECT 588.635 51.075 588.805 51.245 ;
        RECT 589.095 51.075 589.265 51.245 ;
        RECT 589.555 51.075 589.725 51.245 ;
        RECT 590.015 51.075 590.185 51.245 ;
        RECT 590.475 51.075 590.645 51.245 ;
        RECT 590.935 51.075 591.105 51.245 ;
        RECT 591.395 51.075 591.565 51.245 ;
        RECT 591.855 51.075 592.025 51.245 ;
        RECT 592.315 51.075 592.485 51.245 ;
        RECT 592.775 51.075 592.945 51.245 ;
        RECT 593.235 51.075 593.405 51.245 ;
        RECT 593.695 51.075 593.865 51.245 ;
        RECT 594.155 51.075 594.325 51.245 ;
        RECT 594.615 51.075 594.785 51.245 ;
        RECT 595.075 51.075 595.245 51.245 ;
        RECT 595.535 51.075 595.705 51.245 ;
        RECT 595.995 51.075 596.165 51.245 ;
        RECT 596.455 51.075 596.625 51.245 ;
        RECT 596.915 51.075 597.085 51.245 ;
        RECT 597.375 51.075 597.545 51.245 ;
        RECT 597.835 51.075 598.005 51.245 ;
        RECT 598.295 51.075 598.465 51.245 ;
        RECT 598.755 51.075 598.925 51.245 ;
        RECT 599.215 51.075 599.385 51.245 ;
        RECT 599.675 51.075 599.845 51.245 ;
        RECT 600.135 51.075 600.305 51.245 ;
        RECT 600.595 51.075 600.765 51.245 ;
        RECT 601.055 51.075 601.225 51.245 ;
        RECT 601.515 51.075 601.685 51.245 ;
        RECT 601.975 51.075 602.145 51.245 ;
        RECT 602.435 51.075 602.605 51.245 ;
        RECT 602.895 51.075 603.065 51.245 ;
        RECT 603.355 51.075 603.525 51.245 ;
        RECT 603.815 51.075 603.985 51.245 ;
        RECT 604.275 51.075 604.445 51.245 ;
        RECT 604.735 51.075 604.905 51.245 ;
        RECT 605.195 51.075 605.365 51.245 ;
        RECT 605.655 51.075 605.825 51.245 ;
        RECT 606.115 51.075 606.285 51.245 ;
        RECT 606.575 51.075 606.745 51.245 ;
        RECT 607.035 51.075 607.205 51.245 ;
        RECT 607.495 51.075 607.665 51.245 ;
        RECT 607.955 51.075 608.125 51.245 ;
        RECT 608.415 51.075 608.585 51.245 ;
        RECT 608.875 51.075 609.045 51.245 ;
        RECT 609.335 51.075 609.505 51.245 ;
        RECT 609.795 51.075 609.965 51.245 ;
        RECT 610.255 51.075 610.425 51.245 ;
        RECT 610.715 51.075 610.885 51.245 ;
        RECT 611.175 51.075 611.345 51.245 ;
        RECT 611.635 51.075 611.805 51.245 ;
        RECT 612.095 51.075 612.265 51.245 ;
        RECT 612.555 51.075 612.725 51.245 ;
        RECT 613.015 51.075 613.185 51.245 ;
        RECT 613.475 51.075 613.645 51.245 ;
        RECT 613.935 51.075 614.105 51.245 ;
        RECT 614.395 51.075 614.565 51.245 ;
        RECT 614.855 51.075 615.025 51.245 ;
        RECT 615.315 51.075 615.485 51.245 ;
        RECT 615.775 51.075 615.945 51.245 ;
        RECT 616.235 51.075 616.405 51.245 ;
        RECT 616.695 51.075 616.865 51.245 ;
        RECT 617.155 51.075 617.325 51.245 ;
        RECT 617.615 51.075 617.785 51.245 ;
        RECT 618.075 51.075 618.245 51.245 ;
        RECT 618.535 51.075 618.705 51.245 ;
        RECT 618.995 51.075 619.165 51.245 ;
        RECT 619.455 51.075 619.625 51.245 ;
        RECT 619.915 51.075 620.085 51.245 ;
        RECT 620.375 51.075 620.545 51.245 ;
        RECT 620.835 51.075 621.005 51.245 ;
        RECT 621.295 51.075 621.465 51.245 ;
        RECT 621.755 51.075 621.925 51.245 ;
        RECT 622.215 51.075 622.385 51.245 ;
        RECT 622.675 51.075 622.845 51.245 ;
        RECT 623.135 51.075 623.305 51.245 ;
        RECT 623.595 51.075 623.765 51.245 ;
        RECT 624.055 51.075 624.225 51.245 ;
        RECT 624.515 51.075 624.685 51.245 ;
        RECT 624.975 51.075 625.145 51.245 ;
        RECT 625.435 51.075 625.605 51.245 ;
        RECT 625.895 51.075 626.065 51.245 ;
        RECT 626.355 51.075 626.525 51.245 ;
        RECT 626.815 51.075 626.985 51.245 ;
        RECT 627.275 51.075 627.445 51.245 ;
        RECT 627.735 51.075 627.905 51.245 ;
        RECT 628.195 51.075 628.365 51.245 ;
        RECT 628.655 51.075 628.825 51.245 ;
        RECT 629.115 51.075 629.285 51.245 ;
        RECT 629.575 51.075 629.745 51.245 ;
        RECT 630.035 51.075 630.205 51.245 ;
        RECT 630.495 51.075 630.665 51.245 ;
        RECT 630.955 51.075 631.125 51.245 ;
        RECT 73.435 50.565 73.605 50.735 ;
        RECT 72.975 49.885 73.145 50.055 ;
        RECT 78.035 49.885 78.205 50.055 ;
        RECT 78.955 49.885 79.125 50.055 ;
        RECT 80.795 49.885 80.965 50.055 ;
        RECT 85.855 49.885 86.025 50.055 ;
        RECT 86.775 48.865 86.945 49.035 ;
        RECT 91.375 49.545 91.545 49.715 ;
        RECT 91.840 49.205 92.010 49.375 ;
        RECT 92.300 50.225 92.470 50.395 ;
        RECT 92.755 49.885 92.925 50.055 ;
        RECT 93.700 50.225 93.870 50.395 ;
        RECT 95.540 50.225 95.710 50.395 ;
        RECT 94.160 49.205 94.330 49.375 ;
        RECT 95.540 49.205 95.710 49.375 ;
        RECT 105.175 49.885 105.345 50.055 ;
        RECT 107.935 49.885 108.105 50.055 ;
        RECT 108.855 49.885 109.025 50.055 ;
        RECT 99.195 48.865 99.365 49.035 ;
        RECT 113.455 49.885 113.625 50.055 ;
        RECT 113.920 49.205 114.090 49.375 ;
        RECT 114.380 50.225 114.550 50.395 ;
        RECT 114.835 49.885 115.005 50.055 ;
        RECT 115.780 50.225 115.950 50.395 ;
        RECT 117.620 50.225 117.790 50.395 ;
        RECT 116.240 49.205 116.410 49.375 ;
        RECT 117.620 49.205 117.790 49.375 ;
        RECT 120.355 48.865 120.525 49.035 ;
        RECT 125.875 49.545 126.045 49.715 ;
        RECT 126.340 49.205 126.510 49.375 ;
        RECT 126.800 50.225 126.970 50.395 ;
        RECT 127.255 49.885 127.425 50.055 ;
        RECT 128.200 50.225 128.370 50.395 ;
        RECT 130.040 50.225 130.210 50.395 ;
        RECT 128.660 49.205 128.830 49.375 ;
        RECT 130.040 49.205 130.210 49.375 ;
        RECT 133.695 50.565 133.865 50.735 ;
        RECT 141.515 49.885 141.685 50.055 ;
        RECT 141.980 49.205 142.150 49.375 ;
        RECT 142.440 50.225 142.610 50.395 ;
        RECT 142.895 49.885 143.065 50.055 ;
        RECT 143.840 50.225 144.010 50.395 ;
        RECT 145.680 50.225 145.850 50.395 ;
        RECT 144.300 49.205 144.470 49.375 ;
        RECT 145.680 49.205 145.850 49.375 ;
        RECT 153.935 49.545 154.105 49.715 ;
        RECT 154.400 49.205 154.570 49.375 ;
        RECT 154.860 50.225 155.030 50.395 ;
        RECT 155.315 49.885 155.485 50.055 ;
        RECT 156.260 50.225 156.430 50.395 ;
        RECT 158.100 50.225 158.270 50.395 ;
        RECT 156.720 49.205 156.890 49.375 ;
        RECT 158.100 49.205 158.270 49.375 ;
        RECT 169.575 49.885 169.745 50.055 ;
        RECT 160.835 48.865 161.005 49.035 ;
        RECT 170.040 49.205 170.210 49.375 ;
        RECT 170.500 50.225 170.670 50.395 ;
        RECT 170.955 49.885 171.125 50.055 ;
        RECT 171.900 50.225 172.070 50.395 ;
        RECT 173.740 50.225 173.910 50.395 ;
        RECT 172.360 49.205 172.530 49.375 ;
        RECT 173.740 49.205 173.910 49.375 ;
        RECT 176.475 48.865 176.645 49.035 ;
        RECT 181.995 49.885 182.165 50.055 ;
        RECT 182.460 49.205 182.630 49.375 ;
        RECT 182.920 50.225 183.090 50.395 ;
        RECT 183.375 49.885 183.545 50.055 ;
        RECT 184.320 50.225 184.490 50.395 ;
        RECT 186.160 50.225 186.330 50.395 ;
        RECT 184.780 49.205 184.950 49.375 ;
        RECT 186.160 49.205 186.330 49.375 ;
        RECT 188.895 48.865 189.065 49.035 ;
        RECT 195.335 49.885 195.505 50.055 ;
        RECT 194.415 49.205 194.585 49.375 ;
        RECT 197.635 49.545 197.805 49.715 ;
        RECT 198.100 49.205 198.270 49.375 ;
        RECT 198.560 50.225 198.730 50.395 ;
        RECT 199.015 49.885 199.185 50.055 ;
        RECT 199.960 50.225 200.130 50.395 ;
        RECT 201.800 50.225 201.970 50.395 ;
        RECT 200.420 49.205 200.590 49.375 ;
        RECT 201.800 49.205 201.970 49.375 ;
        RECT 204.535 48.865 204.705 49.035 ;
        RECT 210.975 49.885 211.145 50.055 ;
        RECT 210.515 49.545 210.685 49.715 ;
        RECT 212.360 49.545 212.530 49.715 ;
        RECT 213.735 49.885 213.905 50.055 ;
        RECT 214.655 49.885 214.825 50.055 ;
        RECT 215.140 49.545 215.310 49.715 ;
        RECT 230.755 50.225 230.925 50.395 ;
        RECT 216.035 48.865 216.205 49.035 ;
        RECT 230.295 49.885 230.465 50.055 ;
        RECT 231.215 49.885 231.385 50.055 ;
        RECT 232.135 48.865 232.305 49.035 ;
        RECT 238.575 49.885 238.745 50.055 ;
        RECT 238.115 49.545 238.285 49.715 ;
        RECT 239.960 49.545 240.130 49.715 ;
        RECT 241.335 49.885 241.505 50.055 ;
        RECT 242.255 49.885 242.425 50.055 ;
        RECT 242.740 49.545 242.910 49.715 ;
        RECT 259.735 50.565 259.905 50.735 ;
        RECT 253.755 49.885 253.925 50.055 ;
        RECT 254.675 49.885 254.845 50.055 ;
        RECT 243.635 48.865 243.805 49.035 ;
        RECT 256.060 49.545 256.230 49.715 ;
        RECT 256.975 49.885 257.145 50.055 ;
        RECT 257.435 49.885 257.605 50.055 ;
        RECT 258.840 49.545 259.010 49.715 ;
        RECT 264.795 49.885 264.965 50.055 ;
        RECT 265.715 49.205 265.885 49.375 ;
        RECT 271.235 49.885 271.405 50.055 ;
        RECT 270.315 49.545 270.485 49.715 ;
        RECT 272.620 49.545 272.790 49.715 ;
        RECT 273.535 49.885 273.705 50.055 ;
        RECT 273.995 49.885 274.165 50.055 ;
        RECT 275.400 49.545 275.570 49.715 ;
        RECT 283.195 49.885 283.365 50.055 ;
        RECT 284.115 49.885 284.285 50.055 ;
        RECT 276.295 48.865 276.465 49.035 ;
        RECT 284.575 49.545 284.745 49.715 ;
        RECT 290.555 49.885 290.725 50.055 ;
        RECT 290.095 49.545 290.265 49.715 ;
        RECT 291.940 49.545 292.110 49.715 ;
        RECT 293.315 49.885 293.485 50.055 ;
        RECT 294.235 49.885 294.405 50.055 ;
        RECT 294.720 49.545 294.890 49.715 ;
        RECT 300.675 49.885 300.845 50.055 ;
        RECT 303.435 49.885 303.605 50.055 ;
        RECT 302.975 49.545 303.145 49.715 ;
        RECT 314.935 50.565 315.105 50.735 ;
        RECT 315.855 49.885 316.025 50.055 ;
        RECT 317.235 49.885 317.405 50.055 ;
        RECT 324.135 49.885 324.305 50.055 ;
        RECT 323.675 49.545 323.845 49.715 ;
        RECT 325.520 49.545 325.690 49.715 ;
        RECT 326.895 49.885 327.065 50.055 ;
        RECT 327.815 49.885 327.985 50.055 ;
        RECT 328.300 49.545 328.470 49.715 ;
        RECT 337.935 49.885 338.105 50.055 ;
        RECT 349.435 50.565 349.605 50.735 ;
        RECT 344.375 49.885 344.545 50.055 ;
        RECT 343.455 49.545 343.625 49.715 ;
        RECT 345.760 49.545 345.930 49.715 ;
        RECT 346.705 49.885 346.875 50.055 ;
        RECT 347.135 49.885 347.305 50.055 ;
        RECT 354.955 50.565 355.125 50.735 ;
        RECT 348.540 49.545 348.710 49.715 ;
        RECT 355.875 49.885 356.045 50.055 ;
        RECT 356.795 49.885 356.965 50.055 ;
        RECT 367.375 49.885 367.545 50.055 ;
        RECT 368.985 49.885 369.155 50.055 ;
        RECT 375.195 50.565 375.365 50.735 ;
        RECT 368.295 49.545 368.465 49.715 ;
        RECT 374.735 49.885 374.905 50.055 ;
        RECT 376.115 49.885 376.285 50.055 ;
        RECT 382.555 48.865 382.725 49.035 ;
        RECT 387.615 49.205 387.785 49.375 ;
        RECT 394.975 48.865 395.145 49.035 ;
        RECT 400.035 48.865 400.205 49.035 ;
        RECT 405.095 48.865 405.265 49.035 ;
        RECT 414.295 48.865 414.465 49.035 ;
        RECT 429.015 48.865 429.185 49.035 ;
        RECT 436.375 48.865 436.545 49.035 ;
        RECT 451.095 48.865 451.265 49.035 ;
        RECT 458.455 48.865 458.625 49.035 ;
        RECT 469.495 48.865 469.665 49.035 ;
        RECT 480.535 48.865 480.705 49.035 ;
        RECT 487.895 48.865 488.065 49.035 ;
        RECT 513.655 48.865 513.825 49.035 ;
        RECT 521.015 48.865 521.185 49.035 ;
        RECT 535.735 48.865 535.905 49.035 ;
        RECT 543.095 48.865 543.265 49.035 ;
        RECT 554.135 48.865 554.305 49.035 ;
        RECT 564.715 48.865 564.885 49.035 ;
        RECT 572.075 48.865 572.245 49.035 ;
        RECT 597.835 48.865 598.005 49.035 ;
        RECT 619.915 48.865 620.085 49.035 ;
        RECT 624.975 48.865 625.145 49.035 ;
        RECT 42.615 48.355 42.785 48.525 ;
        RECT 43.075 48.355 43.245 48.525 ;
        RECT 43.535 48.355 43.705 48.525 ;
        RECT 43.995 48.355 44.165 48.525 ;
        RECT 44.455 48.355 44.625 48.525 ;
        RECT 44.915 48.355 45.085 48.525 ;
        RECT 45.375 48.355 45.545 48.525 ;
        RECT 45.835 48.355 46.005 48.525 ;
        RECT 46.295 48.355 46.465 48.525 ;
        RECT 46.755 48.355 46.925 48.525 ;
        RECT 47.215 48.355 47.385 48.525 ;
        RECT 47.675 48.355 47.845 48.525 ;
        RECT 48.135 48.355 48.305 48.525 ;
        RECT 48.595 48.355 48.765 48.525 ;
        RECT 49.055 48.355 49.225 48.525 ;
        RECT 49.515 48.355 49.685 48.525 ;
        RECT 49.975 48.355 50.145 48.525 ;
        RECT 50.435 48.355 50.605 48.525 ;
        RECT 50.895 48.355 51.065 48.525 ;
        RECT 51.355 48.355 51.525 48.525 ;
        RECT 51.815 48.355 51.985 48.525 ;
        RECT 52.275 48.355 52.445 48.525 ;
        RECT 52.735 48.355 52.905 48.525 ;
        RECT 53.195 48.355 53.365 48.525 ;
        RECT 53.655 48.355 53.825 48.525 ;
        RECT 54.115 48.355 54.285 48.525 ;
        RECT 54.575 48.355 54.745 48.525 ;
        RECT 55.035 48.355 55.205 48.525 ;
        RECT 55.495 48.355 55.665 48.525 ;
        RECT 55.955 48.355 56.125 48.525 ;
        RECT 56.415 48.355 56.585 48.525 ;
        RECT 56.875 48.355 57.045 48.525 ;
        RECT 57.335 48.355 57.505 48.525 ;
        RECT 57.795 48.355 57.965 48.525 ;
        RECT 58.255 48.355 58.425 48.525 ;
        RECT 58.715 48.355 58.885 48.525 ;
        RECT 59.175 48.355 59.345 48.525 ;
        RECT 59.635 48.355 59.805 48.525 ;
        RECT 60.095 48.355 60.265 48.525 ;
        RECT 60.555 48.355 60.725 48.525 ;
        RECT 61.015 48.355 61.185 48.525 ;
        RECT 61.475 48.355 61.645 48.525 ;
        RECT 61.935 48.355 62.105 48.525 ;
        RECT 62.395 48.355 62.565 48.525 ;
        RECT 62.855 48.355 63.025 48.525 ;
        RECT 63.315 48.355 63.485 48.525 ;
        RECT 63.775 48.355 63.945 48.525 ;
        RECT 64.235 48.355 64.405 48.525 ;
        RECT 64.695 48.355 64.865 48.525 ;
        RECT 65.155 48.355 65.325 48.525 ;
        RECT 65.615 48.355 65.785 48.525 ;
        RECT 66.075 48.355 66.245 48.525 ;
        RECT 66.535 48.355 66.705 48.525 ;
        RECT 66.995 48.355 67.165 48.525 ;
        RECT 67.455 48.355 67.625 48.525 ;
        RECT 67.915 48.355 68.085 48.525 ;
        RECT 68.375 48.355 68.545 48.525 ;
        RECT 68.835 48.355 69.005 48.525 ;
        RECT 69.295 48.355 69.465 48.525 ;
        RECT 69.755 48.355 69.925 48.525 ;
        RECT 70.215 48.355 70.385 48.525 ;
        RECT 70.675 48.355 70.845 48.525 ;
        RECT 71.135 48.355 71.305 48.525 ;
        RECT 71.595 48.355 71.765 48.525 ;
        RECT 72.055 48.355 72.225 48.525 ;
        RECT 72.515 48.355 72.685 48.525 ;
        RECT 72.975 48.355 73.145 48.525 ;
        RECT 73.435 48.355 73.605 48.525 ;
        RECT 73.895 48.355 74.065 48.525 ;
        RECT 74.355 48.355 74.525 48.525 ;
        RECT 74.815 48.355 74.985 48.525 ;
        RECT 75.275 48.355 75.445 48.525 ;
        RECT 75.735 48.355 75.905 48.525 ;
        RECT 76.195 48.355 76.365 48.525 ;
        RECT 76.655 48.355 76.825 48.525 ;
        RECT 77.115 48.355 77.285 48.525 ;
        RECT 77.575 48.355 77.745 48.525 ;
        RECT 78.035 48.355 78.205 48.525 ;
        RECT 78.495 48.355 78.665 48.525 ;
        RECT 78.955 48.355 79.125 48.525 ;
        RECT 79.415 48.355 79.585 48.525 ;
        RECT 79.875 48.355 80.045 48.525 ;
        RECT 80.335 48.355 80.505 48.525 ;
        RECT 80.795 48.355 80.965 48.525 ;
        RECT 81.255 48.355 81.425 48.525 ;
        RECT 81.715 48.355 81.885 48.525 ;
        RECT 82.175 48.355 82.345 48.525 ;
        RECT 82.635 48.355 82.805 48.525 ;
        RECT 83.095 48.355 83.265 48.525 ;
        RECT 83.555 48.355 83.725 48.525 ;
        RECT 84.015 48.355 84.185 48.525 ;
        RECT 84.475 48.355 84.645 48.525 ;
        RECT 84.935 48.355 85.105 48.525 ;
        RECT 85.395 48.355 85.565 48.525 ;
        RECT 85.855 48.355 86.025 48.525 ;
        RECT 86.315 48.355 86.485 48.525 ;
        RECT 86.775 48.355 86.945 48.525 ;
        RECT 87.235 48.355 87.405 48.525 ;
        RECT 87.695 48.355 87.865 48.525 ;
        RECT 88.155 48.355 88.325 48.525 ;
        RECT 88.615 48.355 88.785 48.525 ;
        RECT 89.075 48.355 89.245 48.525 ;
        RECT 89.535 48.355 89.705 48.525 ;
        RECT 89.995 48.355 90.165 48.525 ;
        RECT 90.455 48.355 90.625 48.525 ;
        RECT 90.915 48.355 91.085 48.525 ;
        RECT 91.375 48.355 91.545 48.525 ;
        RECT 91.835 48.355 92.005 48.525 ;
        RECT 92.295 48.355 92.465 48.525 ;
        RECT 92.755 48.355 92.925 48.525 ;
        RECT 93.215 48.355 93.385 48.525 ;
        RECT 93.675 48.355 93.845 48.525 ;
        RECT 94.135 48.355 94.305 48.525 ;
        RECT 94.595 48.355 94.765 48.525 ;
        RECT 95.055 48.355 95.225 48.525 ;
        RECT 95.515 48.355 95.685 48.525 ;
        RECT 95.975 48.355 96.145 48.525 ;
        RECT 96.435 48.355 96.605 48.525 ;
        RECT 96.895 48.355 97.065 48.525 ;
        RECT 97.355 48.355 97.525 48.525 ;
        RECT 97.815 48.355 97.985 48.525 ;
        RECT 98.275 48.355 98.445 48.525 ;
        RECT 98.735 48.355 98.905 48.525 ;
        RECT 99.195 48.355 99.365 48.525 ;
        RECT 99.655 48.355 99.825 48.525 ;
        RECT 100.115 48.355 100.285 48.525 ;
        RECT 100.575 48.355 100.745 48.525 ;
        RECT 101.035 48.355 101.205 48.525 ;
        RECT 101.495 48.355 101.665 48.525 ;
        RECT 101.955 48.355 102.125 48.525 ;
        RECT 102.415 48.355 102.585 48.525 ;
        RECT 102.875 48.355 103.045 48.525 ;
        RECT 103.335 48.355 103.505 48.525 ;
        RECT 103.795 48.355 103.965 48.525 ;
        RECT 104.255 48.355 104.425 48.525 ;
        RECT 104.715 48.355 104.885 48.525 ;
        RECT 105.175 48.355 105.345 48.525 ;
        RECT 105.635 48.355 105.805 48.525 ;
        RECT 106.095 48.355 106.265 48.525 ;
        RECT 106.555 48.355 106.725 48.525 ;
        RECT 107.015 48.355 107.185 48.525 ;
        RECT 107.475 48.355 107.645 48.525 ;
        RECT 107.935 48.355 108.105 48.525 ;
        RECT 108.395 48.355 108.565 48.525 ;
        RECT 108.855 48.355 109.025 48.525 ;
        RECT 109.315 48.355 109.485 48.525 ;
        RECT 109.775 48.355 109.945 48.525 ;
        RECT 110.235 48.355 110.405 48.525 ;
        RECT 110.695 48.355 110.865 48.525 ;
        RECT 111.155 48.355 111.325 48.525 ;
        RECT 111.615 48.355 111.785 48.525 ;
        RECT 112.075 48.355 112.245 48.525 ;
        RECT 112.535 48.355 112.705 48.525 ;
        RECT 112.995 48.355 113.165 48.525 ;
        RECT 113.455 48.355 113.625 48.525 ;
        RECT 113.915 48.355 114.085 48.525 ;
        RECT 114.375 48.355 114.545 48.525 ;
        RECT 114.835 48.355 115.005 48.525 ;
        RECT 115.295 48.355 115.465 48.525 ;
        RECT 115.755 48.355 115.925 48.525 ;
        RECT 116.215 48.355 116.385 48.525 ;
        RECT 116.675 48.355 116.845 48.525 ;
        RECT 117.135 48.355 117.305 48.525 ;
        RECT 117.595 48.355 117.765 48.525 ;
        RECT 118.055 48.355 118.225 48.525 ;
        RECT 118.515 48.355 118.685 48.525 ;
        RECT 118.975 48.355 119.145 48.525 ;
        RECT 119.435 48.355 119.605 48.525 ;
        RECT 119.895 48.355 120.065 48.525 ;
        RECT 120.355 48.355 120.525 48.525 ;
        RECT 120.815 48.355 120.985 48.525 ;
        RECT 121.275 48.355 121.445 48.525 ;
        RECT 121.735 48.355 121.905 48.525 ;
        RECT 122.195 48.355 122.365 48.525 ;
        RECT 122.655 48.355 122.825 48.525 ;
        RECT 123.115 48.355 123.285 48.525 ;
        RECT 123.575 48.355 123.745 48.525 ;
        RECT 124.035 48.355 124.205 48.525 ;
        RECT 124.495 48.355 124.665 48.525 ;
        RECT 124.955 48.355 125.125 48.525 ;
        RECT 125.415 48.355 125.585 48.525 ;
        RECT 125.875 48.355 126.045 48.525 ;
        RECT 126.335 48.355 126.505 48.525 ;
        RECT 126.795 48.355 126.965 48.525 ;
        RECT 127.255 48.355 127.425 48.525 ;
        RECT 127.715 48.355 127.885 48.525 ;
        RECT 128.175 48.355 128.345 48.525 ;
        RECT 128.635 48.355 128.805 48.525 ;
        RECT 129.095 48.355 129.265 48.525 ;
        RECT 129.555 48.355 129.725 48.525 ;
        RECT 130.015 48.355 130.185 48.525 ;
        RECT 130.475 48.355 130.645 48.525 ;
        RECT 130.935 48.355 131.105 48.525 ;
        RECT 131.395 48.355 131.565 48.525 ;
        RECT 131.855 48.355 132.025 48.525 ;
        RECT 132.315 48.355 132.485 48.525 ;
        RECT 132.775 48.355 132.945 48.525 ;
        RECT 133.235 48.355 133.405 48.525 ;
        RECT 133.695 48.355 133.865 48.525 ;
        RECT 134.155 48.355 134.325 48.525 ;
        RECT 134.615 48.355 134.785 48.525 ;
        RECT 135.075 48.355 135.245 48.525 ;
        RECT 135.535 48.355 135.705 48.525 ;
        RECT 135.995 48.355 136.165 48.525 ;
        RECT 136.455 48.355 136.625 48.525 ;
        RECT 136.915 48.355 137.085 48.525 ;
        RECT 137.375 48.355 137.545 48.525 ;
        RECT 137.835 48.355 138.005 48.525 ;
        RECT 138.295 48.355 138.465 48.525 ;
        RECT 138.755 48.355 138.925 48.525 ;
        RECT 139.215 48.355 139.385 48.525 ;
        RECT 139.675 48.355 139.845 48.525 ;
        RECT 140.135 48.355 140.305 48.525 ;
        RECT 140.595 48.355 140.765 48.525 ;
        RECT 141.055 48.355 141.225 48.525 ;
        RECT 141.515 48.355 141.685 48.525 ;
        RECT 141.975 48.355 142.145 48.525 ;
        RECT 142.435 48.355 142.605 48.525 ;
        RECT 142.895 48.355 143.065 48.525 ;
        RECT 143.355 48.355 143.525 48.525 ;
        RECT 143.815 48.355 143.985 48.525 ;
        RECT 144.275 48.355 144.445 48.525 ;
        RECT 144.735 48.355 144.905 48.525 ;
        RECT 145.195 48.355 145.365 48.525 ;
        RECT 145.655 48.355 145.825 48.525 ;
        RECT 146.115 48.355 146.285 48.525 ;
        RECT 146.575 48.355 146.745 48.525 ;
        RECT 147.035 48.355 147.205 48.525 ;
        RECT 147.495 48.355 147.665 48.525 ;
        RECT 147.955 48.355 148.125 48.525 ;
        RECT 148.415 48.355 148.585 48.525 ;
        RECT 148.875 48.355 149.045 48.525 ;
        RECT 149.335 48.355 149.505 48.525 ;
        RECT 149.795 48.355 149.965 48.525 ;
        RECT 150.255 48.355 150.425 48.525 ;
        RECT 150.715 48.355 150.885 48.525 ;
        RECT 151.175 48.355 151.345 48.525 ;
        RECT 151.635 48.355 151.805 48.525 ;
        RECT 152.095 48.355 152.265 48.525 ;
        RECT 152.555 48.355 152.725 48.525 ;
        RECT 153.015 48.355 153.185 48.525 ;
        RECT 153.475 48.355 153.645 48.525 ;
        RECT 153.935 48.355 154.105 48.525 ;
        RECT 154.395 48.355 154.565 48.525 ;
        RECT 154.855 48.355 155.025 48.525 ;
        RECT 155.315 48.355 155.485 48.525 ;
        RECT 155.775 48.355 155.945 48.525 ;
        RECT 156.235 48.355 156.405 48.525 ;
        RECT 156.695 48.355 156.865 48.525 ;
        RECT 157.155 48.355 157.325 48.525 ;
        RECT 157.615 48.355 157.785 48.525 ;
        RECT 158.075 48.355 158.245 48.525 ;
        RECT 158.535 48.355 158.705 48.525 ;
        RECT 158.995 48.355 159.165 48.525 ;
        RECT 159.455 48.355 159.625 48.525 ;
        RECT 159.915 48.355 160.085 48.525 ;
        RECT 160.375 48.355 160.545 48.525 ;
        RECT 160.835 48.355 161.005 48.525 ;
        RECT 161.295 48.355 161.465 48.525 ;
        RECT 161.755 48.355 161.925 48.525 ;
        RECT 162.215 48.355 162.385 48.525 ;
        RECT 162.675 48.355 162.845 48.525 ;
        RECT 163.135 48.355 163.305 48.525 ;
        RECT 163.595 48.355 163.765 48.525 ;
        RECT 164.055 48.355 164.225 48.525 ;
        RECT 164.515 48.355 164.685 48.525 ;
        RECT 164.975 48.355 165.145 48.525 ;
        RECT 165.435 48.355 165.605 48.525 ;
        RECT 165.895 48.355 166.065 48.525 ;
        RECT 166.355 48.355 166.525 48.525 ;
        RECT 166.815 48.355 166.985 48.525 ;
        RECT 167.275 48.355 167.445 48.525 ;
        RECT 167.735 48.355 167.905 48.525 ;
        RECT 168.195 48.355 168.365 48.525 ;
        RECT 168.655 48.355 168.825 48.525 ;
        RECT 169.115 48.355 169.285 48.525 ;
        RECT 169.575 48.355 169.745 48.525 ;
        RECT 170.035 48.355 170.205 48.525 ;
        RECT 170.495 48.355 170.665 48.525 ;
        RECT 170.955 48.355 171.125 48.525 ;
        RECT 171.415 48.355 171.585 48.525 ;
        RECT 171.875 48.355 172.045 48.525 ;
        RECT 172.335 48.355 172.505 48.525 ;
        RECT 172.795 48.355 172.965 48.525 ;
        RECT 173.255 48.355 173.425 48.525 ;
        RECT 173.715 48.355 173.885 48.525 ;
        RECT 174.175 48.355 174.345 48.525 ;
        RECT 174.635 48.355 174.805 48.525 ;
        RECT 175.095 48.355 175.265 48.525 ;
        RECT 175.555 48.355 175.725 48.525 ;
        RECT 176.015 48.355 176.185 48.525 ;
        RECT 176.475 48.355 176.645 48.525 ;
        RECT 176.935 48.355 177.105 48.525 ;
        RECT 177.395 48.355 177.565 48.525 ;
        RECT 177.855 48.355 178.025 48.525 ;
        RECT 178.315 48.355 178.485 48.525 ;
        RECT 178.775 48.355 178.945 48.525 ;
        RECT 179.235 48.355 179.405 48.525 ;
        RECT 179.695 48.355 179.865 48.525 ;
        RECT 180.155 48.355 180.325 48.525 ;
        RECT 180.615 48.355 180.785 48.525 ;
        RECT 181.075 48.355 181.245 48.525 ;
        RECT 181.535 48.355 181.705 48.525 ;
        RECT 181.995 48.355 182.165 48.525 ;
        RECT 182.455 48.355 182.625 48.525 ;
        RECT 182.915 48.355 183.085 48.525 ;
        RECT 183.375 48.355 183.545 48.525 ;
        RECT 183.835 48.355 184.005 48.525 ;
        RECT 184.295 48.355 184.465 48.525 ;
        RECT 184.755 48.355 184.925 48.525 ;
        RECT 185.215 48.355 185.385 48.525 ;
        RECT 185.675 48.355 185.845 48.525 ;
        RECT 186.135 48.355 186.305 48.525 ;
        RECT 186.595 48.355 186.765 48.525 ;
        RECT 187.055 48.355 187.225 48.525 ;
        RECT 187.515 48.355 187.685 48.525 ;
        RECT 187.975 48.355 188.145 48.525 ;
        RECT 188.435 48.355 188.605 48.525 ;
        RECT 188.895 48.355 189.065 48.525 ;
        RECT 189.355 48.355 189.525 48.525 ;
        RECT 189.815 48.355 189.985 48.525 ;
        RECT 190.275 48.355 190.445 48.525 ;
        RECT 190.735 48.355 190.905 48.525 ;
        RECT 191.195 48.355 191.365 48.525 ;
        RECT 191.655 48.355 191.825 48.525 ;
        RECT 192.115 48.355 192.285 48.525 ;
        RECT 192.575 48.355 192.745 48.525 ;
        RECT 193.035 48.355 193.205 48.525 ;
        RECT 193.495 48.355 193.665 48.525 ;
        RECT 193.955 48.355 194.125 48.525 ;
        RECT 194.415 48.355 194.585 48.525 ;
        RECT 194.875 48.355 195.045 48.525 ;
        RECT 195.335 48.355 195.505 48.525 ;
        RECT 195.795 48.355 195.965 48.525 ;
        RECT 196.255 48.355 196.425 48.525 ;
        RECT 196.715 48.355 196.885 48.525 ;
        RECT 197.175 48.355 197.345 48.525 ;
        RECT 197.635 48.355 197.805 48.525 ;
        RECT 198.095 48.355 198.265 48.525 ;
        RECT 198.555 48.355 198.725 48.525 ;
        RECT 199.015 48.355 199.185 48.525 ;
        RECT 199.475 48.355 199.645 48.525 ;
        RECT 199.935 48.355 200.105 48.525 ;
        RECT 200.395 48.355 200.565 48.525 ;
        RECT 200.855 48.355 201.025 48.525 ;
        RECT 201.315 48.355 201.485 48.525 ;
        RECT 201.775 48.355 201.945 48.525 ;
        RECT 202.235 48.355 202.405 48.525 ;
        RECT 202.695 48.355 202.865 48.525 ;
        RECT 203.155 48.355 203.325 48.525 ;
        RECT 203.615 48.355 203.785 48.525 ;
        RECT 204.075 48.355 204.245 48.525 ;
        RECT 204.535 48.355 204.705 48.525 ;
        RECT 204.995 48.355 205.165 48.525 ;
        RECT 205.455 48.355 205.625 48.525 ;
        RECT 205.915 48.355 206.085 48.525 ;
        RECT 206.375 48.355 206.545 48.525 ;
        RECT 206.835 48.355 207.005 48.525 ;
        RECT 207.295 48.355 207.465 48.525 ;
        RECT 207.755 48.355 207.925 48.525 ;
        RECT 208.215 48.355 208.385 48.525 ;
        RECT 208.675 48.355 208.845 48.525 ;
        RECT 209.135 48.355 209.305 48.525 ;
        RECT 209.595 48.355 209.765 48.525 ;
        RECT 210.055 48.355 210.225 48.525 ;
        RECT 210.515 48.355 210.685 48.525 ;
        RECT 210.975 48.355 211.145 48.525 ;
        RECT 211.435 48.355 211.605 48.525 ;
        RECT 211.895 48.355 212.065 48.525 ;
        RECT 212.355 48.355 212.525 48.525 ;
        RECT 212.815 48.355 212.985 48.525 ;
        RECT 213.275 48.355 213.445 48.525 ;
        RECT 213.735 48.355 213.905 48.525 ;
        RECT 214.195 48.355 214.365 48.525 ;
        RECT 214.655 48.355 214.825 48.525 ;
        RECT 215.115 48.355 215.285 48.525 ;
        RECT 215.575 48.355 215.745 48.525 ;
        RECT 216.035 48.355 216.205 48.525 ;
        RECT 216.495 48.355 216.665 48.525 ;
        RECT 216.955 48.355 217.125 48.525 ;
        RECT 217.415 48.355 217.585 48.525 ;
        RECT 217.875 48.355 218.045 48.525 ;
        RECT 218.335 48.355 218.505 48.525 ;
        RECT 218.795 48.355 218.965 48.525 ;
        RECT 219.255 48.355 219.425 48.525 ;
        RECT 219.715 48.355 219.885 48.525 ;
        RECT 220.175 48.355 220.345 48.525 ;
        RECT 220.635 48.355 220.805 48.525 ;
        RECT 221.095 48.355 221.265 48.525 ;
        RECT 221.555 48.355 221.725 48.525 ;
        RECT 222.015 48.355 222.185 48.525 ;
        RECT 222.475 48.355 222.645 48.525 ;
        RECT 222.935 48.355 223.105 48.525 ;
        RECT 223.395 48.355 223.565 48.525 ;
        RECT 223.855 48.355 224.025 48.525 ;
        RECT 224.315 48.355 224.485 48.525 ;
        RECT 224.775 48.355 224.945 48.525 ;
        RECT 225.235 48.355 225.405 48.525 ;
        RECT 225.695 48.355 225.865 48.525 ;
        RECT 226.155 48.355 226.325 48.525 ;
        RECT 226.615 48.355 226.785 48.525 ;
        RECT 227.075 48.355 227.245 48.525 ;
        RECT 227.535 48.355 227.705 48.525 ;
        RECT 227.995 48.355 228.165 48.525 ;
        RECT 228.455 48.355 228.625 48.525 ;
        RECT 228.915 48.355 229.085 48.525 ;
        RECT 229.375 48.355 229.545 48.525 ;
        RECT 229.835 48.355 230.005 48.525 ;
        RECT 230.295 48.355 230.465 48.525 ;
        RECT 230.755 48.355 230.925 48.525 ;
        RECT 231.215 48.355 231.385 48.525 ;
        RECT 231.675 48.355 231.845 48.525 ;
        RECT 232.135 48.355 232.305 48.525 ;
        RECT 232.595 48.355 232.765 48.525 ;
        RECT 233.055 48.355 233.225 48.525 ;
        RECT 233.515 48.355 233.685 48.525 ;
        RECT 233.975 48.355 234.145 48.525 ;
        RECT 234.435 48.355 234.605 48.525 ;
        RECT 234.895 48.355 235.065 48.525 ;
        RECT 235.355 48.355 235.525 48.525 ;
        RECT 235.815 48.355 235.985 48.525 ;
        RECT 236.275 48.355 236.445 48.525 ;
        RECT 236.735 48.355 236.905 48.525 ;
        RECT 237.195 48.355 237.365 48.525 ;
        RECT 237.655 48.355 237.825 48.525 ;
        RECT 238.115 48.355 238.285 48.525 ;
        RECT 238.575 48.355 238.745 48.525 ;
        RECT 239.035 48.355 239.205 48.525 ;
        RECT 239.495 48.355 239.665 48.525 ;
        RECT 239.955 48.355 240.125 48.525 ;
        RECT 240.415 48.355 240.585 48.525 ;
        RECT 240.875 48.355 241.045 48.525 ;
        RECT 241.335 48.355 241.505 48.525 ;
        RECT 241.795 48.355 241.965 48.525 ;
        RECT 242.255 48.355 242.425 48.525 ;
        RECT 242.715 48.355 242.885 48.525 ;
        RECT 243.175 48.355 243.345 48.525 ;
        RECT 243.635 48.355 243.805 48.525 ;
        RECT 244.095 48.355 244.265 48.525 ;
        RECT 244.555 48.355 244.725 48.525 ;
        RECT 245.015 48.355 245.185 48.525 ;
        RECT 245.475 48.355 245.645 48.525 ;
        RECT 245.935 48.355 246.105 48.525 ;
        RECT 246.395 48.355 246.565 48.525 ;
        RECT 246.855 48.355 247.025 48.525 ;
        RECT 247.315 48.355 247.485 48.525 ;
        RECT 247.775 48.355 247.945 48.525 ;
        RECT 248.235 48.355 248.405 48.525 ;
        RECT 248.695 48.355 248.865 48.525 ;
        RECT 249.155 48.355 249.325 48.525 ;
        RECT 249.615 48.355 249.785 48.525 ;
        RECT 250.075 48.355 250.245 48.525 ;
        RECT 250.535 48.355 250.705 48.525 ;
        RECT 250.995 48.355 251.165 48.525 ;
        RECT 251.455 48.355 251.625 48.525 ;
        RECT 251.915 48.355 252.085 48.525 ;
        RECT 252.375 48.355 252.545 48.525 ;
        RECT 252.835 48.355 253.005 48.525 ;
        RECT 253.295 48.355 253.465 48.525 ;
        RECT 253.755 48.355 253.925 48.525 ;
        RECT 254.215 48.355 254.385 48.525 ;
        RECT 254.675 48.355 254.845 48.525 ;
        RECT 255.135 48.355 255.305 48.525 ;
        RECT 255.595 48.355 255.765 48.525 ;
        RECT 256.055 48.355 256.225 48.525 ;
        RECT 256.515 48.355 256.685 48.525 ;
        RECT 256.975 48.355 257.145 48.525 ;
        RECT 257.435 48.355 257.605 48.525 ;
        RECT 257.895 48.355 258.065 48.525 ;
        RECT 258.355 48.355 258.525 48.525 ;
        RECT 258.815 48.355 258.985 48.525 ;
        RECT 259.275 48.355 259.445 48.525 ;
        RECT 259.735 48.355 259.905 48.525 ;
        RECT 260.195 48.355 260.365 48.525 ;
        RECT 260.655 48.355 260.825 48.525 ;
        RECT 261.115 48.355 261.285 48.525 ;
        RECT 261.575 48.355 261.745 48.525 ;
        RECT 262.035 48.355 262.205 48.525 ;
        RECT 262.495 48.355 262.665 48.525 ;
        RECT 262.955 48.355 263.125 48.525 ;
        RECT 263.415 48.355 263.585 48.525 ;
        RECT 263.875 48.355 264.045 48.525 ;
        RECT 264.335 48.355 264.505 48.525 ;
        RECT 264.795 48.355 264.965 48.525 ;
        RECT 265.255 48.355 265.425 48.525 ;
        RECT 265.715 48.355 265.885 48.525 ;
        RECT 266.175 48.355 266.345 48.525 ;
        RECT 266.635 48.355 266.805 48.525 ;
        RECT 267.095 48.355 267.265 48.525 ;
        RECT 267.555 48.355 267.725 48.525 ;
        RECT 268.015 48.355 268.185 48.525 ;
        RECT 268.475 48.355 268.645 48.525 ;
        RECT 268.935 48.355 269.105 48.525 ;
        RECT 269.395 48.355 269.565 48.525 ;
        RECT 269.855 48.355 270.025 48.525 ;
        RECT 270.315 48.355 270.485 48.525 ;
        RECT 270.775 48.355 270.945 48.525 ;
        RECT 271.235 48.355 271.405 48.525 ;
        RECT 271.695 48.355 271.865 48.525 ;
        RECT 272.155 48.355 272.325 48.525 ;
        RECT 272.615 48.355 272.785 48.525 ;
        RECT 273.075 48.355 273.245 48.525 ;
        RECT 273.535 48.355 273.705 48.525 ;
        RECT 273.995 48.355 274.165 48.525 ;
        RECT 274.455 48.355 274.625 48.525 ;
        RECT 274.915 48.355 275.085 48.525 ;
        RECT 275.375 48.355 275.545 48.525 ;
        RECT 275.835 48.355 276.005 48.525 ;
        RECT 276.295 48.355 276.465 48.525 ;
        RECT 276.755 48.355 276.925 48.525 ;
        RECT 277.215 48.355 277.385 48.525 ;
        RECT 277.675 48.355 277.845 48.525 ;
        RECT 278.135 48.355 278.305 48.525 ;
        RECT 278.595 48.355 278.765 48.525 ;
        RECT 279.055 48.355 279.225 48.525 ;
        RECT 279.515 48.355 279.685 48.525 ;
        RECT 279.975 48.355 280.145 48.525 ;
        RECT 280.435 48.355 280.605 48.525 ;
        RECT 280.895 48.355 281.065 48.525 ;
        RECT 281.355 48.355 281.525 48.525 ;
        RECT 281.815 48.355 281.985 48.525 ;
        RECT 282.275 48.355 282.445 48.525 ;
        RECT 282.735 48.355 282.905 48.525 ;
        RECT 283.195 48.355 283.365 48.525 ;
        RECT 283.655 48.355 283.825 48.525 ;
        RECT 284.115 48.355 284.285 48.525 ;
        RECT 284.575 48.355 284.745 48.525 ;
        RECT 285.035 48.355 285.205 48.525 ;
        RECT 285.495 48.355 285.665 48.525 ;
        RECT 285.955 48.355 286.125 48.525 ;
        RECT 286.415 48.355 286.585 48.525 ;
        RECT 286.875 48.355 287.045 48.525 ;
        RECT 287.335 48.355 287.505 48.525 ;
        RECT 287.795 48.355 287.965 48.525 ;
        RECT 288.255 48.355 288.425 48.525 ;
        RECT 288.715 48.355 288.885 48.525 ;
        RECT 289.175 48.355 289.345 48.525 ;
        RECT 289.635 48.355 289.805 48.525 ;
        RECT 290.095 48.355 290.265 48.525 ;
        RECT 290.555 48.355 290.725 48.525 ;
        RECT 291.015 48.355 291.185 48.525 ;
        RECT 291.475 48.355 291.645 48.525 ;
        RECT 291.935 48.355 292.105 48.525 ;
        RECT 292.395 48.355 292.565 48.525 ;
        RECT 292.855 48.355 293.025 48.525 ;
        RECT 293.315 48.355 293.485 48.525 ;
        RECT 293.775 48.355 293.945 48.525 ;
        RECT 294.235 48.355 294.405 48.525 ;
        RECT 294.695 48.355 294.865 48.525 ;
        RECT 295.155 48.355 295.325 48.525 ;
        RECT 295.615 48.355 295.785 48.525 ;
        RECT 296.075 48.355 296.245 48.525 ;
        RECT 296.535 48.355 296.705 48.525 ;
        RECT 296.995 48.355 297.165 48.525 ;
        RECT 297.455 48.355 297.625 48.525 ;
        RECT 297.915 48.355 298.085 48.525 ;
        RECT 298.375 48.355 298.545 48.525 ;
        RECT 298.835 48.355 299.005 48.525 ;
        RECT 299.295 48.355 299.465 48.525 ;
        RECT 299.755 48.355 299.925 48.525 ;
        RECT 300.215 48.355 300.385 48.525 ;
        RECT 300.675 48.355 300.845 48.525 ;
        RECT 301.135 48.355 301.305 48.525 ;
        RECT 301.595 48.355 301.765 48.525 ;
        RECT 302.055 48.355 302.225 48.525 ;
        RECT 302.515 48.355 302.685 48.525 ;
        RECT 302.975 48.355 303.145 48.525 ;
        RECT 303.435 48.355 303.605 48.525 ;
        RECT 303.895 48.355 304.065 48.525 ;
        RECT 304.355 48.355 304.525 48.525 ;
        RECT 304.815 48.355 304.985 48.525 ;
        RECT 305.275 48.355 305.445 48.525 ;
        RECT 305.735 48.355 305.905 48.525 ;
        RECT 306.195 48.355 306.365 48.525 ;
        RECT 306.655 48.355 306.825 48.525 ;
        RECT 307.115 48.355 307.285 48.525 ;
        RECT 307.575 48.355 307.745 48.525 ;
        RECT 308.035 48.355 308.205 48.525 ;
        RECT 308.495 48.355 308.665 48.525 ;
        RECT 308.955 48.355 309.125 48.525 ;
        RECT 309.415 48.355 309.585 48.525 ;
        RECT 309.875 48.355 310.045 48.525 ;
        RECT 310.335 48.355 310.505 48.525 ;
        RECT 310.795 48.355 310.965 48.525 ;
        RECT 311.255 48.355 311.425 48.525 ;
        RECT 311.715 48.355 311.885 48.525 ;
        RECT 312.175 48.355 312.345 48.525 ;
        RECT 312.635 48.355 312.805 48.525 ;
        RECT 313.095 48.355 313.265 48.525 ;
        RECT 313.555 48.355 313.725 48.525 ;
        RECT 314.015 48.355 314.185 48.525 ;
        RECT 314.475 48.355 314.645 48.525 ;
        RECT 314.935 48.355 315.105 48.525 ;
        RECT 315.395 48.355 315.565 48.525 ;
        RECT 315.855 48.355 316.025 48.525 ;
        RECT 316.315 48.355 316.485 48.525 ;
        RECT 316.775 48.355 316.945 48.525 ;
        RECT 317.235 48.355 317.405 48.525 ;
        RECT 317.695 48.355 317.865 48.525 ;
        RECT 318.155 48.355 318.325 48.525 ;
        RECT 318.615 48.355 318.785 48.525 ;
        RECT 319.075 48.355 319.245 48.525 ;
        RECT 319.535 48.355 319.705 48.525 ;
        RECT 319.995 48.355 320.165 48.525 ;
        RECT 320.455 48.355 320.625 48.525 ;
        RECT 320.915 48.355 321.085 48.525 ;
        RECT 321.375 48.355 321.545 48.525 ;
        RECT 321.835 48.355 322.005 48.525 ;
        RECT 322.295 48.355 322.465 48.525 ;
        RECT 322.755 48.355 322.925 48.525 ;
        RECT 323.215 48.355 323.385 48.525 ;
        RECT 323.675 48.355 323.845 48.525 ;
        RECT 324.135 48.355 324.305 48.525 ;
        RECT 324.595 48.355 324.765 48.525 ;
        RECT 325.055 48.355 325.225 48.525 ;
        RECT 325.515 48.355 325.685 48.525 ;
        RECT 325.975 48.355 326.145 48.525 ;
        RECT 326.435 48.355 326.605 48.525 ;
        RECT 326.895 48.355 327.065 48.525 ;
        RECT 327.355 48.355 327.525 48.525 ;
        RECT 327.815 48.355 327.985 48.525 ;
        RECT 328.275 48.355 328.445 48.525 ;
        RECT 328.735 48.355 328.905 48.525 ;
        RECT 329.195 48.355 329.365 48.525 ;
        RECT 329.655 48.355 329.825 48.525 ;
        RECT 330.115 48.355 330.285 48.525 ;
        RECT 330.575 48.355 330.745 48.525 ;
        RECT 331.035 48.355 331.205 48.525 ;
        RECT 331.495 48.355 331.665 48.525 ;
        RECT 331.955 48.355 332.125 48.525 ;
        RECT 332.415 48.355 332.585 48.525 ;
        RECT 332.875 48.355 333.045 48.525 ;
        RECT 333.335 48.355 333.505 48.525 ;
        RECT 333.795 48.355 333.965 48.525 ;
        RECT 334.255 48.355 334.425 48.525 ;
        RECT 334.715 48.355 334.885 48.525 ;
        RECT 335.175 48.355 335.345 48.525 ;
        RECT 335.635 48.355 335.805 48.525 ;
        RECT 336.095 48.355 336.265 48.525 ;
        RECT 336.555 48.355 336.725 48.525 ;
        RECT 337.015 48.355 337.185 48.525 ;
        RECT 337.475 48.355 337.645 48.525 ;
        RECT 337.935 48.355 338.105 48.525 ;
        RECT 338.395 48.355 338.565 48.525 ;
        RECT 338.855 48.355 339.025 48.525 ;
        RECT 339.315 48.355 339.485 48.525 ;
        RECT 339.775 48.355 339.945 48.525 ;
        RECT 340.235 48.355 340.405 48.525 ;
        RECT 340.695 48.355 340.865 48.525 ;
        RECT 341.155 48.355 341.325 48.525 ;
        RECT 341.615 48.355 341.785 48.525 ;
        RECT 342.075 48.355 342.245 48.525 ;
        RECT 342.535 48.355 342.705 48.525 ;
        RECT 342.995 48.355 343.165 48.525 ;
        RECT 343.455 48.355 343.625 48.525 ;
        RECT 343.915 48.355 344.085 48.525 ;
        RECT 344.375 48.355 344.545 48.525 ;
        RECT 344.835 48.355 345.005 48.525 ;
        RECT 345.295 48.355 345.465 48.525 ;
        RECT 345.755 48.355 345.925 48.525 ;
        RECT 346.215 48.355 346.385 48.525 ;
        RECT 346.675 48.355 346.845 48.525 ;
        RECT 347.135 48.355 347.305 48.525 ;
        RECT 347.595 48.355 347.765 48.525 ;
        RECT 348.055 48.355 348.225 48.525 ;
        RECT 348.515 48.355 348.685 48.525 ;
        RECT 348.975 48.355 349.145 48.525 ;
        RECT 349.435 48.355 349.605 48.525 ;
        RECT 349.895 48.355 350.065 48.525 ;
        RECT 350.355 48.355 350.525 48.525 ;
        RECT 350.815 48.355 350.985 48.525 ;
        RECT 351.275 48.355 351.445 48.525 ;
        RECT 351.735 48.355 351.905 48.525 ;
        RECT 352.195 48.355 352.365 48.525 ;
        RECT 352.655 48.355 352.825 48.525 ;
        RECT 353.115 48.355 353.285 48.525 ;
        RECT 353.575 48.355 353.745 48.525 ;
        RECT 354.035 48.355 354.205 48.525 ;
        RECT 354.495 48.355 354.665 48.525 ;
        RECT 354.955 48.355 355.125 48.525 ;
        RECT 355.415 48.355 355.585 48.525 ;
        RECT 355.875 48.355 356.045 48.525 ;
        RECT 356.335 48.355 356.505 48.525 ;
        RECT 356.795 48.355 356.965 48.525 ;
        RECT 357.255 48.355 357.425 48.525 ;
        RECT 357.715 48.355 357.885 48.525 ;
        RECT 358.175 48.355 358.345 48.525 ;
        RECT 358.635 48.355 358.805 48.525 ;
        RECT 359.095 48.355 359.265 48.525 ;
        RECT 359.555 48.355 359.725 48.525 ;
        RECT 360.015 48.355 360.185 48.525 ;
        RECT 360.475 48.355 360.645 48.525 ;
        RECT 360.935 48.355 361.105 48.525 ;
        RECT 361.395 48.355 361.565 48.525 ;
        RECT 361.855 48.355 362.025 48.525 ;
        RECT 362.315 48.355 362.485 48.525 ;
        RECT 362.775 48.355 362.945 48.525 ;
        RECT 363.235 48.355 363.405 48.525 ;
        RECT 363.695 48.355 363.865 48.525 ;
        RECT 364.155 48.355 364.325 48.525 ;
        RECT 364.615 48.355 364.785 48.525 ;
        RECT 365.075 48.355 365.245 48.525 ;
        RECT 365.535 48.355 365.705 48.525 ;
        RECT 365.995 48.355 366.165 48.525 ;
        RECT 366.455 48.355 366.625 48.525 ;
        RECT 366.915 48.355 367.085 48.525 ;
        RECT 367.375 48.355 367.545 48.525 ;
        RECT 367.835 48.355 368.005 48.525 ;
        RECT 368.295 48.355 368.465 48.525 ;
        RECT 368.755 48.355 368.925 48.525 ;
        RECT 369.215 48.355 369.385 48.525 ;
        RECT 369.675 48.355 369.845 48.525 ;
        RECT 370.135 48.355 370.305 48.525 ;
        RECT 370.595 48.355 370.765 48.525 ;
        RECT 371.055 48.355 371.225 48.525 ;
        RECT 371.515 48.355 371.685 48.525 ;
        RECT 371.975 48.355 372.145 48.525 ;
        RECT 372.435 48.355 372.605 48.525 ;
        RECT 372.895 48.355 373.065 48.525 ;
        RECT 373.355 48.355 373.525 48.525 ;
        RECT 373.815 48.355 373.985 48.525 ;
        RECT 374.275 48.355 374.445 48.525 ;
        RECT 374.735 48.355 374.905 48.525 ;
        RECT 375.195 48.355 375.365 48.525 ;
        RECT 375.655 48.355 375.825 48.525 ;
        RECT 376.115 48.355 376.285 48.525 ;
        RECT 376.575 48.355 376.745 48.525 ;
        RECT 377.035 48.355 377.205 48.525 ;
        RECT 377.495 48.355 377.665 48.525 ;
        RECT 377.955 48.355 378.125 48.525 ;
        RECT 378.415 48.355 378.585 48.525 ;
        RECT 378.875 48.355 379.045 48.525 ;
        RECT 379.335 48.355 379.505 48.525 ;
        RECT 379.795 48.355 379.965 48.525 ;
        RECT 380.255 48.355 380.425 48.525 ;
        RECT 380.715 48.355 380.885 48.525 ;
        RECT 381.175 48.355 381.345 48.525 ;
        RECT 381.635 48.355 381.805 48.525 ;
        RECT 382.095 48.355 382.265 48.525 ;
        RECT 382.555 48.355 382.725 48.525 ;
        RECT 383.015 48.355 383.185 48.525 ;
        RECT 383.475 48.355 383.645 48.525 ;
        RECT 383.935 48.355 384.105 48.525 ;
        RECT 384.395 48.355 384.565 48.525 ;
        RECT 384.855 48.355 385.025 48.525 ;
        RECT 385.315 48.355 385.485 48.525 ;
        RECT 385.775 48.355 385.945 48.525 ;
        RECT 386.235 48.355 386.405 48.525 ;
        RECT 386.695 48.355 386.865 48.525 ;
        RECT 387.155 48.355 387.325 48.525 ;
        RECT 387.615 48.355 387.785 48.525 ;
        RECT 388.075 48.355 388.245 48.525 ;
        RECT 388.535 48.355 388.705 48.525 ;
        RECT 388.995 48.355 389.165 48.525 ;
        RECT 389.455 48.355 389.625 48.525 ;
        RECT 389.915 48.355 390.085 48.525 ;
        RECT 390.375 48.355 390.545 48.525 ;
        RECT 390.835 48.355 391.005 48.525 ;
        RECT 391.295 48.355 391.465 48.525 ;
        RECT 391.755 48.355 391.925 48.525 ;
        RECT 392.215 48.355 392.385 48.525 ;
        RECT 392.675 48.355 392.845 48.525 ;
        RECT 393.135 48.355 393.305 48.525 ;
        RECT 393.595 48.355 393.765 48.525 ;
        RECT 394.055 48.355 394.225 48.525 ;
        RECT 394.515 48.355 394.685 48.525 ;
        RECT 394.975 48.355 395.145 48.525 ;
        RECT 395.435 48.355 395.605 48.525 ;
        RECT 395.895 48.355 396.065 48.525 ;
        RECT 396.355 48.355 396.525 48.525 ;
        RECT 396.815 48.355 396.985 48.525 ;
        RECT 397.275 48.355 397.445 48.525 ;
        RECT 397.735 48.355 397.905 48.525 ;
        RECT 398.195 48.355 398.365 48.525 ;
        RECT 398.655 48.355 398.825 48.525 ;
        RECT 399.115 48.355 399.285 48.525 ;
        RECT 399.575 48.355 399.745 48.525 ;
        RECT 400.035 48.355 400.205 48.525 ;
        RECT 400.495 48.355 400.665 48.525 ;
        RECT 400.955 48.355 401.125 48.525 ;
        RECT 401.415 48.355 401.585 48.525 ;
        RECT 401.875 48.355 402.045 48.525 ;
        RECT 402.335 48.355 402.505 48.525 ;
        RECT 402.795 48.355 402.965 48.525 ;
        RECT 403.255 48.355 403.425 48.525 ;
        RECT 403.715 48.355 403.885 48.525 ;
        RECT 404.175 48.355 404.345 48.525 ;
        RECT 404.635 48.355 404.805 48.525 ;
        RECT 405.095 48.355 405.265 48.525 ;
        RECT 405.555 48.355 405.725 48.525 ;
        RECT 406.015 48.355 406.185 48.525 ;
        RECT 406.475 48.355 406.645 48.525 ;
        RECT 406.935 48.355 407.105 48.525 ;
        RECT 407.395 48.355 407.565 48.525 ;
        RECT 407.855 48.355 408.025 48.525 ;
        RECT 408.315 48.355 408.485 48.525 ;
        RECT 408.775 48.355 408.945 48.525 ;
        RECT 409.235 48.355 409.405 48.525 ;
        RECT 409.695 48.355 409.865 48.525 ;
        RECT 410.155 48.355 410.325 48.525 ;
        RECT 410.615 48.355 410.785 48.525 ;
        RECT 411.075 48.355 411.245 48.525 ;
        RECT 411.535 48.355 411.705 48.525 ;
        RECT 411.995 48.355 412.165 48.525 ;
        RECT 412.455 48.355 412.625 48.525 ;
        RECT 412.915 48.355 413.085 48.525 ;
        RECT 413.375 48.355 413.545 48.525 ;
        RECT 413.835 48.355 414.005 48.525 ;
        RECT 414.295 48.355 414.465 48.525 ;
        RECT 414.755 48.355 414.925 48.525 ;
        RECT 415.215 48.355 415.385 48.525 ;
        RECT 415.675 48.355 415.845 48.525 ;
        RECT 416.135 48.355 416.305 48.525 ;
        RECT 416.595 48.355 416.765 48.525 ;
        RECT 417.055 48.355 417.225 48.525 ;
        RECT 417.515 48.355 417.685 48.525 ;
        RECT 417.975 48.355 418.145 48.525 ;
        RECT 418.435 48.355 418.605 48.525 ;
        RECT 418.895 48.355 419.065 48.525 ;
        RECT 419.355 48.355 419.525 48.525 ;
        RECT 419.815 48.355 419.985 48.525 ;
        RECT 420.275 48.355 420.445 48.525 ;
        RECT 420.735 48.355 420.905 48.525 ;
        RECT 421.195 48.355 421.365 48.525 ;
        RECT 421.655 48.355 421.825 48.525 ;
        RECT 422.115 48.355 422.285 48.525 ;
        RECT 422.575 48.355 422.745 48.525 ;
        RECT 423.035 48.355 423.205 48.525 ;
        RECT 423.495 48.355 423.665 48.525 ;
        RECT 423.955 48.355 424.125 48.525 ;
        RECT 424.415 48.355 424.585 48.525 ;
        RECT 424.875 48.355 425.045 48.525 ;
        RECT 425.335 48.355 425.505 48.525 ;
        RECT 425.795 48.355 425.965 48.525 ;
        RECT 426.255 48.355 426.425 48.525 ;
        RECT 426.715 48.355 426.885 48.525 ;
        RECT 427.175 48.355 427.345 48.525 ;
        RECT 427.635 48.355 427.805 48.525 ;
        RECT 428.095 48.355 428.265 48.525 ;
        RECT 428.555 48.355 428.725 48.525 ;
        RECT 429.015 48.355 429.185 48.525 ;
        RECT 429.475 48.355 429.645 48.525 ;
        RECT 429.935 48.355 430.105 48.525 ;
        RECT 430.395 48.355 430.565 48.525 ;
        RECT 430.855 48.355 431.025 48.525 ;
        RECT 431.315 48.355 431.485 48.525 ;
        RECT 431.775 48.355 431.945 48.525 ;
        RECT 432.235 48.355 432.405 48.525 ;
        RECT 432.695 48.355 432.865 48.525 ;
        RECT 433.155 48.355 433.325 48.525 ;
        RECT 433.615 48.355 433.785 48.525 ;
        RECT 434.075 48.355 434.245 48.525 ;
        RECT 434.535 48.355 434.705 48.525 ;
        RECT 434.995 48.355 435.165 48.525 ;
        RECT 435.455 48.355 435.625 48.525 ;
        RECT 435.915 48.355 436.085 48.525 ;
        RECT 436.375 48.355 436.545 48.525 ;
        RECT 436.835 48.355 437.005 48.525 ;
        RECT 437.295 48.355 437.465 48.525 ;
        RECT 437.755 48.355 437.925 48.525 ;
        RECT 438.215 48.355 438.385 48.525 ;
        RECT 438.675 48.355 438.845 48.525 ;
        RECT 439.135 48.355 439.305 48.525 ;
        RECT 439.595 48.355 439.765 48.525 ;
        RECT 440.055 48.355 440.225 48.525 ;
        RECT 440.515 48.355 440.685 48.525 ;
        RECT 440.975 48.355 441.145 48.525 ;
        RECT 441.435 48.355 441.605 48.525 ;
        RECT 441.895 48.355 442.065 48.525 ;
        RECT 442.355 48.355 442.525 48.525 ;
        RECT 442.815 48.355 442.985 48.525 ;
        RECT 443.275 48.355 443.445 48.525 ;
        RECT 443.735 48.355 443.905 48.525 ;
        RECT 444.195 48.355 444.365 48.525 ;
        RECT 444.655 48.355 444.825 48.525 ;
        RECT 445.115 48.355 445.285 48.525 ;
        RECT 445.575 48.355 445.745 48.525 ;
        RECT 446.035 48.355 446.205 48.525 ;
        RECT 446.495 48.355 446.665 48.525 ;
        RECT 446.955 48.355 447.125 48.525 ;
        RECT 447.415 48.355 447.585 48.525 ;
        RECT 447.875 48.355 448.045 48.525 ;
        RECT 448.335 48.355 448.505 48.525 ;
        RECT 448.795 48.355 448.965 48.525 ;
        RECT 449.255 48.355 449.425 48.525 ;
        RECT 449.715 48.355 449.885 48.525 ;
        RECT 450.175 48.355 450.345 48.525 ;
        RECT 450.635 48.355 450.805 48.525 ;
        RECT 451.095 48.355 451.265 48.525 ;
        RECT 451.555 48.355 451.725 48.525 ;
        RECT 452.015 48.355 452.185 48.525 ;
        RECT 452.475 48.355 452.645 48.525 ;
        RECT 452.935 48.355 453.105 48.525 ;
        RECT 453.395 48.355 453.565 48.525 ;
        RECT 453.855 48.355 454.025 48.525 ;
        RECT 454.315 48.355 454.485 48.525 ;
        RECT 454.775 48.355 454.945 48.525 ;
        RECT 455.235 48.355 455.405 48.525 ;
        RECT 455.695 48.355 455.865 48.525 ;
        RECT 456.155 48.355 456.325 48.525 ;
        RECT 456.615 48.355 456.785 48.525 ;
        RECT 457.075 48.355 457.245 48.525 ;
        RECT 457.535 48.355 457.705 48.525 ;
        RECT 457.995 48.355 458.165 48.525 ;
        RECT 458.455 48.355 458.625 48.525 ;
        RECT 458.915 48.355 459.085 48.525 ;
        RECT 459.375 48.355 459.545 48.525 ;
        RECT 459.835 48.355 460.005 48.525 ;
        RECT 460.295 48.355 460.465 48.525 ;
        RECT 460.755 48.355 460.925 48.525 ;
        RECT 461.215 48.355 461.385 48.525 ;
        RECT 461.675 48.355 461.845 48.525 ;
        RECT 462.135 48.355 462.305 48.525 ;
        RECT 462.595 48.355 462.765 48.525 ;
        RECT 463.055 48.355 463.225 48.525 ;
        RECT 463.515 48.355 463.685 48.525 ;
        RECT 463.975 48.355 464.145 48.525 ;
        RECT 464.435 48.355 464.605 48.525 ;
        RECT 464.895 48.355 465.065 48.525 ;
        RECT 465.355 48.355 465.525 48.525 ;
        RECT 465.815 48.355 465.985 48.525 ;
        RECT 466.275 48.355 466.445 48.525 ;
        RECT 466.735 48.355 466.905 48.525 ;
        RECT 467.195 48.355 467.365 48.525 ;
        RECT 467.655 48.355 467.825 48.525 ;
        RECT 468.115 48.355 468.285 48.525 ;
        RECT 468.575 48.355 468.745 48.525 ;
        RECT 469.035 48.355 469.205 48.525 ;
        RECT 469.495 48.355 469.665 48.525 ;
        RECT 469.955 48.355 470.125 48.525 ;
        RECT 470.415 48.355 470.585 48.525 ;
        RECT 470.875 48.355 471.045 48.525 ;
        RECT 471.335 48.355 471.505 48.525 ;
        RECT 471.795 48.355 471.965 48.525 ;
        RECT 472.255 48.355 472.425 48.525 ;
        RECT 472.715 48.355 472.885 48.525 ;
        RECT 473.175 48.355 473.345 48.525 ;
        RECT 473.635 48.355 473.805 48.525 ;
        RECT 474.095 48.355 474.265 48.525 ;
        RECT 474.555 48.355 474.725 48.525 ;
        RECT 475.015 48.355 475.185 48.525 ;
        RECT 475.475 48.355 475.645 48.525 ;
        RECT 475.935 48.355 476.105 48.525 ;
        RECT 476.395 48.355 476.565 48.525 ;
        RECT 476.855 48.355 477.025 48.525 ;
        RECT 477.315 48.355 477.485 48.525 ;
        RECT 477.775 48.355 477.945 48.525 ;
        RECT 478.235 48.355 478.405 48.525 ;
        RECT 478.695 48.355 478.865 48.525 ;
        RECT 479.155 48.355 479.325 48.525 ;
        RECT 479.615 48.355 479.785 48.525 ;
        RECT 480.075 48.355 480.245 48.525 ;
        RECT 480.535 48.355 480.705 48.525 ;
        RECT 480.995 48.355 481.165 48.525 ;
        RECT 481.455 48.355 481.625 48.525 ;
        RECT 481.915 48.355 482.085 48.525 ;
        RECT 482.375 48.355 482.545 48.525 ;
        RECT 482.835 48.355 483.005 48.525 ;
        RECT 483.295 48.355 483.465 48.525 ;
        RECT 483.755 48.355 483.925 48.525 ;
        RECT 484.215 48.355 484.385 48.525 ;
        RECT 484.675 48.355 484.845 48.525 ;
        RECT 485.135 48.355 485.305 48.525 ;
        RECT 485.595 48.355 485.765 48.525 ;
        RECT 486.055 48.355 486.225 48.525 ;
        RECT 486.515 48.355 486.685 48.525 ;
        RECT 486.975 48.355 487.145 48.525 ;
        RECT 487.435 48.355 487.605 48.525 ;
        RECT 487.895 48.355 488.065 48.525 ;
        RECT 488.355 48.355 488.525 48.525 ;
        RECT 488.815 48.355 488.985 48.525 ;
        RECT 489.275 48.355 489.445 48.525 ;
        RECT 489.735 48.355 489.905 48.525 ;
        RECT 490.195 48.355 490.365 48.525 ;
        RECT 490.655 48.355 490.825 48.525 ;
        RECT 491.115 48.355 491.285 48.525 ;
        RECT 491.575 48.355 491.745 48.525 ;
        RECT 492.035 48.355 492.205 48.525 ;
        RECT 492.495 48.355 492.665 48.525 ;
        RECT 492.955 48.355 493.125 48.525 ;
        RECT 493.415 48.355 493.585 48.525 ;
        RECT 493.875 48.355 494.045 48.525 ;
        RECT 494.335 48.355 494.505 48.525 ;
        RECT 494.795 48.355 494.965 48.525 ;
        RECT 495.255 48.355 495.425 48.525 ;
        RECT 495.715 48.355 495.885 48.525 ;
        RECT 496.175 48.355 496.345 48.525 ;
        RECT 496.635 48.355 496.805 48.525 ;
        RECT 497.095 48.355 497.265 48.525 ;
        RECT 497.555 48.355 497.725 48.525 ;
        RECT 498.015 48.355 498.185 48.525 ;
        RECT 498.475 48.355 498.645 48.525 ;
        RECT 498.935 48.355 499.105 48.525 ;
        RECT 499.395 48.355 499.565 48.525 ;
        RECT 499.855 48.355 500.025 48.525 ;
        RECT 500.315 48.355 500.485 48.525 ;
        RECT 500.775 48.355 500.945 48.525 ;
        RECT 501.235 48.355 501.405 48.525 ;
        RECT 501.695 48.355 501.865 48.525 ;
        RECT 502.155 48.355 502.325 48.525 ;
        RECT 502.615 48.355 502.785 48.525 ;
        RECT 503.075 48.355 503.245 48.525 ;
        RECT 503.535 48.355 503.705 48.525 ;
        RECT 503.995 48.355 504.165 48.525 ;
        RECT 504.455 48.355 504.625 48.525 ;
        RECT 504.915 48.355 505.085 48.525 ;
        RECT 505.375 48.355 505.545 48.525 ;
        RECT 505.835 48.355 506.005 48.525 ;
        RECT 506.295 48.355 506.465 48.525 ;
        RECT 506.755 48.355 506.925 48.525 ;
        RECT 507.215 48.355 507.385 48.525 ;
        RECT 507.675 48.355 507.845 48.525 ;
        RECT 508.135 48.355 508.305 48.525 ;
        RECT 508.595 48.355 508.765 48.525 ;
        RECT 509.055 48.355 509.225 48.525 ;
        RECT 509.515 48.355 509.685 48.525 ;
        RECT 509.975 48.355 510.145 48.525 ;
        RECT 510.435 48.355 510.605 48.525 ;
        RECT 510.895 48.355 511.065 48.525 ;
        RECT 511.355 48.355 511.525 48.525 ;
        RECT 511.815 48.355 511.985 48.525 ;
        RECT 512.275 48.355 512.445 48.525 ;
        RECT 512.735 48.355 512.905 48.525 ;
        RECT 513.195 48.355 513.365 48.525 ;
        RECT 513.655 48.355 513.825 48.525 ;
        RECT 514.115 48.355 514.285 48.525 ;
        RECT 514.575 48.355 514.745 48.525 ;
        RECT 515.035 48.355 515.205 48.525 ;
        RECT 515.495 48.355 515.665 48.525 ;
        RECT 515.955 48.355 516.125 48.525 ;
        RECT 516.415 48.355 516.585 48.525 ;
        RECT 516.875 48.355 517.045 48.525 ;
        RECT 517.335 48.355 517.505 48.525 ;
        RECT 517.795 48.355 517.965 48.525 ;
        RECT 518.255 48.355 518.425 48.525 ;
        RECT 518.715 48.355 518.885 48.525 ;
        RECT 519.175 48.355 519.345 48.525 ;
        RECT 519.635 48.355 519.805 48.525 ;
        RECT 520.095 48.355 520.265 48.525 ;
        RECT 520.555 48.355 520.725 48.525 ;
        RECT 521.015 48.355 521.185 48.525 ;
        RECT 521.475 48.355 521.645 48.525 ;
        RECT 521.935 48.355 522.105 48.525 ;
        RECT 522.395 48.355 522.565 48.525 ;
        RECT 522.855 48.355 523.025 48.525 ;
        RECT 523.315 48.355 523.485 48.525 ;
        RECT 523.775 48.355 523.945 48.525 ;
        RECT 524.235 48.355 524.405 48.525 ;
        RECT 524.695 48.355 524.865 48.525 ;
        RECT 525.155 48.355 525.325 48.525 ;
        RECT 525.615 48.355 525.785 48.525 ;
        RECT 526.075 48.355 526.245 48.525 ;
        RECT 526.535 48.355 526.705 48.525 ;
        RECT 526.995 48.355 527.165 48.525 ;
        RECT 527.455 48.355 527.625 48.525 ;
        RECT 527.915 48.355 528.085 48.525 ;
        RECT 528.375 48.355 528.545 48.525 ;
        RECT 528.835 48.355 529.005 48.525 ;
        RECT 529.295 48.355 529.465 48.525 ;
        RECT 529.755 48.355 529.925 48.525 ;
        RECT 530.215 48.355 530.385 48.525 ;
        RECT 530.675 48.355 530.845 48.525 ;
        RECT 531.135 48.355 531.305 48.525 ;
        RECT 531.595 48.355 531.765 48.525 ;
        RECT 532.055 48.355 532.225 48.525 ;
        RECT 532.515 48.355 532.685 48.525 ;
        RECT 532.975 48.355 533.145 48.525 ;
        RECT 533.435 48.355 533.605 48.525 ;
        RECT 533.895 48.355 534.065 48.525 ;
        RECT 534.355 48.355 534.525 48.525 ;
        RECT 534.815 48.355 534.985 48.525 ;
        RECT 535.275 48.355 535.445 48.525 ;
        RECT 535.735 48.355 535.905 48.525 ;
        RECT 536.195 48.355 536.365 48.525 ;
        RECT 536.655 48.355 536.825 48.525 ;
        RECT 537.115 48.355 537.285 48.525 ;
        RECT 537.575 48.355 537.745 48.525 ;
        RECT 538.035 48.355 538.205 48.525 ;
        RECT 538.495 48.355 538.665 48.525 ;
        RECT 538.955 48.355 539.125 48.525 ;
        RECT 539.415 48.355 539.585 48.525 ;
        RECT 539.875 48.355 540.045 48.525 ;
        RECT 540.335 48.355 540.505 48.525 ;
        RECT 540.795 48.355 540.965 48.525 ;
        RECT 541.255 48.355 541.425 48.525 ;
        RECT 541.715 48.355 541.885 48.525 ;
        RECT 542.175 48.355 542.345 48.525 ;
        RECT 542.635 48.355 542.805 48.525 ;
        RECT 543.095 48.355 543.265 48.525 ;
        RECT 543.555 48.355 543.725 48.525 ;
        RECT 544.015 48.355 544.185 48.525 ;
        RECT 544.475 48.355 544.645 48.525 ;
        RECT 544.935 48.355 545.105 48.525 ;
        RECT 545.395 48.355 545.565 48.525 ;
        RECT 545.855 48.355 546.025 48.525 ;
        RECT 546.315 48.355 546.485 48.525 ;
        RECT 546.775 48.355 546.945 48.525 ;
        RECT 547.235 48.355 547.405 48.525 ;
        RECT 547.695 48.355 547.865 48.525 ;
        RECT 548.155 48.355 548.325 48.525 ;
        RECT 548.615 48.355 548.785 48.525 ;
        RECT 549.075 48.355 549.245 48.525 ;
        RECT 549.535 48.355 549.705 48.525 ;
        RECT 549.995 48.355 550.165 48.525 ;
        RECT 550.455 48.355 550.625 48.525 ;
        RECT 550.915 48.355 551.085 48.525 ;
        RECT 551.375 48.355 551.545 48.525 ;
        RECT 551.835 48.355 552.005 48.525 ;
        RECT 552.295 48.355 552.465 48.525 ;
        RECT 552.755 48.355 552.925 48.525 ;
        RECT 553.215 48.355 553.385 48.525 ;
        RECT 553.675 48.355 553.845 48.525 ;
        RECT 554.135 48.355 554.305 48.525 ;
        RECT 554.595 48.355 554.765 48.525 ;
        RECT 555.055 48.355 555.225 48.525 ;
        RECT 555.515 48.355 555.685 48.525 ;
        RECT 555.975 48.355 556.145 48.525 ;
        RECT 556.435 48.355 556.605 48.525 ;
        RECT 556.895 48.355 557.065 48.525 ;
        RECT 557.355 48.355 557.525 48.525 ;
        RECT 557.815 48.355 557.985 48.525 ;
        RECT 558.275 48.355 558.445 48.525 ;
        RECT 558.735 48.355 558.905 48.525 ;
        RECT 559.195 48.355 559.365 48.525 ;
        RECT 559.655 48.355 559.825 48.525 ;
        RECT 560.115 48.355 560.285 48.525 ;
        RECT 560.575 48.355 560.745 48.525 ;
        RECT 561.035 48.355 561.205 48.525 ;
        RECT 561.495 48.355 561.665 48.525 ;
        RECT 561.955 48.355 562.125 48.525 ;
        RECT 562.415 48.355 562.585 48.525 ;
        RECT 562.875 48.355 563.045 48.525 ;
        RECT 563.335 48.355 563.505 48.525 ;
        RECT 563.795 48.355 563.965 48.525 ;
        RECT 564.255 48.355 564.425 48.525 ;
        RECT 564.715 48.355 564.885 48.525 ;
        RECT 565.175 48.355 565.345 48.525 ;
        RECT 565.635 48.355 565.805 48.525 ;
        RECT 566.095 48.355 566.265 48.525 ;
        RECT 566.555 48.355 566.725 48.525 ;
        RECT 567.015 48.355 567.185 48.525 ;
        RECT 567.475 48.355 567.645 48.525 ;
        RECT 567.935 48.355 568.105 48.525 ;
        RECT 568.395 48.355 568.565 48.525 ;
        RECT 568.855 48.355 569.025 48.525 ;
        RECT 569.315 48.355 569.485 48.525 ;
        RECT 569.775 48.355 569.945 48.525 ;
        RECT 570.235 48.355 570.405 48.525 ;
        RECT 570.695 48.355 570.865 48.525 ;
        RECT 571.155 48.355 571.325 48.525 ;
        RECT 571.615 48.355 571.785 48.525 ;
        RECT 572.075 48.355 572.245 48.525 ;
        RECT 572.535 48.355 572.705 48.525 ;
        RECT 572.995 48.355 573.165 48.525 ;
        RECT 573.455 48.355 573.625 48.525 ;
        RECT 573.915 48.355 574.085 48.525 ;
        RECT 574.375 48.355 574.545 48.525 ;
        RECT 574.835 48.355 575.005 48.525 ;
        RECT 575.295 48.355 575.465 48.525 ;
        RECT 575.755 48.355 575.925 48.525 ;
        RECT 576.215 48.355 576.385 48.525 ;
        RECT 576.675 48.355 576.845 48.525 ;
        RECT 577.135 48.355 577.305 48.525 ;
        RECT 577.595 48.355 577.765 48.525 ;
        RECT 578.055 48.355 578.225 48.525 ;
        RECT 578.515 48.355 578.685 48.525 ;
        RECT 578.975 48.355 579.145 48.525 ;
        RECT 579.435 48.355 579.605 48.525 ;
        RECT 579.895 48.355 580.065 48.525 ;
        RECT 580.355 48.355 580.525 48.525 ;
        RECT 580.815 48.355 580.985 48.525 ;
        RECT 581.275 48.355 581.445 48.525 ;
        RECT 581.735 48.355 581.905 48.525 ;
        RECT 582.195 48.355 582.365 48.525 ;
        RECT 582.655 48.355 582.825 48.525 ;
        RECT 583.115 48.355 583.285 48.525 ;
        RECT 583.575 48.355 583.745 48.525 ;
        RECT 584.035 48.355 584.205 48.525 ;
        RECT 584.495 48.355 584.665 48.525 ;
        RECT 584.955 48.355 585.125 48.525 ;
        RECT 585.415 48.355 585.585 48.525 ;
        RECT 585.875 48.355 586.045 48.525 ;
        RECT 586.335 48.355 586.505 48.525 ;
        RECT 586.795 48.355 586.965 48.525 ;
        RECT 587.255 48.355 587.425 48.525 ;
        RECT 587.715 48.355 587.885 48.525 ;
        RECT 588.175 48.355 588.345 48.525 ;
        RECT 588.635 48.355 588.805 48.525 ;
        RECT 589.095 48.355 589.265 48.525 ;
        RECT 589.555 48.355 589.725 48.525 ;
        RECT 590.015 48.355 590.185 48.525 ;
        RECT 590.475 48.355 590.645 48.525 ;
        RECT 590.935 48.355 591.105 48.525 ;
        RECT 591.395 48.355 591.565 48.525 ;
        RECT 591.855 48.355 592.025 48.525 ;
        RECT 592.315 48.355 592.485 48.525 ;
        RECT 592.775 48.355 592.945 48.525 ;
        RECT 593.235 48.355 593.405 48.525 ;
        RECT 593.695 48.355 593.865 48.525 ;
        RECT 594.155 48.355 594.325 48.525 ;
        RECT 594.615 48.355 594.785 48.525 ;
        RECT 595.075 48.355 595.245 48.525 ;
        RECT 595.535 48.355 595.705 48.525 ;
        RECT 595.995 48.355 596.165 48.525 ;
        RECT 596.455 48.355 596.625 48.525 ;
        RECT 596.915 48.355 597.085 48.525 ;
        RECT 597.375 48.355 597.545 48.525 ;
        RECT 597.835 48.355 598.005 48.525 ;
        RECT 598.295 48.355 598.465 48.525 ;
        RECT 598.755 48.355 598.925 48.525 ;
        RECT 599.215 48.355 599.385 48.525 ;
        RECT 599.675 48.355 599.845 48.525 ;
        RECT 600.135 48.355 600.305 48.525 ;
        RECT 600.595 48.355 600.765 48.525 ;
        RECT 601.055 48.355 601.225 48.525 ;
        RECT 601.515 48.355 601.685 48.525 ;
        RECT 601.975 48.355 602.145 48.525 ;
        RECT 602.435 48.355 602.605 48.525 ;
        RECT 602.895 48.355 603.065 48.525 ;
        RECT 603.355 48.355 603.525 48.525 ;
        RECT 603.815 48.355 603.985 48.525 ;
        RECT 604.275 48.355 604.445 48.525 ;
        RECT 604.735 48.355 604.905 48.525 ;
        RECT 605.195 48.355 605.365 48.525 ;
        RECT 605.655 48.355 605.825 48.525 ;
        RECT 606.115 48.355 606.285 48.525 ;
        RECT 606.575 48.355 606.745 48.525 ;
        RECT 607.035 48.355 607.205 48.525 ;
        RECT 607.495 48.355 607.665 48.525 ;
        RECT 607.955 48.355 608.125 48.525 ;
        RECT 608.415 48.355 608.585 48.525 ;
        RECT 608.875 48.355 609.045 48.525 ;
        RECT 609.335 48.355 609.505 48.525 ;
        RECT 609.795 48.355 609.965 48.525 ;
        RECT 610.255 48.355 610.425 48.525 ;
        RECT 610.715 48.355 610.885 48.525 ;
        RECT 611.175 48.355 611.345 48.525 ;
        RECT 611.635 48.355 611.805 48.525 ;
        RECT 612.095 48.355 612.265 48.525 ;
        RECT 612.555 48.355 612.725 48.525 ;
        RECT 613.015 48.355 613.185 48.525 ;
        RECT 613.475 48.355 613.645 48.525 ;
        RECT 613.935 48.355 614.105 48.525 ;
        RECT 614.395 48.355 614.565 48.525 ;
        RECT 614.855 48.355 615.025 48.525 ;
        RECT 615.315 48.355 615.485 48.525 ;
        RECT 615.775 48.355 615.945 48.525 ;
        RECT 616.235 48.355 616.405 48.525 ;
        RECT 616.695 48.355 616.865 48.525 ;
        RECT 617.155 48.355 617.325 48.525 ;
        RECT 617.615 48.355 617.785 48.525 ;
        RECT 618.075 48.355 618.245 48.525 ;
        RECT 618.535 48.355 618.705 48.525 ;
        RECT 618.995 48.355 619.165 48.525 ;
        RECT 619.455 48.355 619.625 48.525 ;
        RECT 619.915 48.355 620.085 48.525 ;
        RECT 620.375 48.355 620.545 48.525 ;
        RECT 620.835 48.355 621.005 48.525 ;
        RECT 621.295 48.355 621.465 48.525 ;
        RECT 621.755 48.355 621.925 48.525 ;
        RECT 622.215 48.355 622.385 48.525 ;
        RECT 622.675 48.355 622.845 48.525 ;
        RECT 623.135 48.355 623.305 48.525 ;
        RECT 623.595 48.355 623.765 48.525 ;
        RECT 624.055 48.355 624.225 48.525 ;
        RECT 624.515 48.355 624.685 48.525 ;
        RECT 624.975 48.355 625.145 48.525 ;
        RECT 625.435 48.355 625.605 48.525 ;
        RECT 625.895 48.355 626.065 48.525 ;
        RECT 626.355 48.355 626.525 48.525 ;
        RECT 626.815 48.355 626.985 48.525 ;
        RECT 627.275 48.355 627.445 48.525 ;
        RECT 627.735 48.355 627.905 48.525 ;
        RECT 628.195 48.355 628.365 48.525 ;
        RECT 628.655 48.355 628.825 48.525 ;
        RECT 629.115 48.355 629.285 48.525 ;
        RECT 629.575 48.355 629.745 48.525 ;
        RECT 630.035 48.355 630.205 48.525 ;
        RECT 630.495 48.355 630.665 48.525 ;
        RECT 630.955 48.355 631.125 48.525 ;
        RECT 72.515 46.825 72.685 46.995 ;
        RECT 72.975 46.145 73.145 46.315 ;
        RECT 77.575 47.165 77.745 47.335 ;
        RECT 78.035 46.825 78.205 46.995 ;
        RECT 80.335 46.485 80.505 46.655 ;
        RECT 85.395 46.825 85.565 46.995 ;
        RECT 86.315 46.145 86.485 46.315 ;
        RECT 94.595 47.165 94.765 47.335 ;
        RECT 90.915 46.825 91.085 46.995 ;
        RECT 93.215 46.825 93.385 46.995 ;
        RECT 103.335 46.825 103.505 46.995 ;
        RECT 106.095 46.825 106.265 46.995 ;
        RECT 114.835 47.165 115.005 47.335 ;
        RECT 111.615 46.825 111.785 46.995 ;
        RECT 113.915 46.825 114.085 46.995 ;
        RECT 104.715 46.145 104.885 46.315 ;
        RECT 118.975 46.485 119.145 46.655 ;
        RECT 120.355 47.505 120.525 47.675 ;
        RECT 119.710 46.825 119.880 46.995 ;
        RECT 120.815 47.165 120.985 47.335 ;
        RECT 122.655 46.825 122.825 46.995 ;
        RECT 128.180 47.505 128.350 47.675 ;
        RECT 127.750 47.165 127.920 47.335 ;
        RECT 129.095 47.165 129.265 47.335 ;
        RECT 128.640 46.485 128.810 46.655 ;
        RECT 130.500 47.505 130.670 47.675 ;
        RECT 130.040 46.485 130.210 46.655 ;
        RECT 131.880 47.505 132.050 47.675 ;
        RECT 131.880 46.485 132.050 46.655 ;
        RECT 134.615 47.505 134.785 47.675 ;
        RECT 149.795 47.845 149.965 48.015 ;
        RECT 146.120 47.165 146.290 47.335 ;
        RECT 144.735 46.825 144.905 46.995 ;
        RECT 145.195 46.825 145.365 46.995 ;
        RECT 147.035 46.825 147.205 46.995 ;
        RECT 147.495 46.825 147.665 46.995 ;
        RECT 148.900 47.165 149.070 47.335 ;
        RECT 155.780 47.505 155.950 47.675 ;
        RECT 155.315 47.165 155.485 47.335 ;
        RECT 156.695 46.825 156.865 46.995 ;
        RECT 156.240 46.485 156.410 46.655 ;
        RECT 158.100 47.505 158.270 47.675 ;
        RECT 157.640 46.485 157.810 46.655 ;
        RECT 159.480 47.505 159.650 47.675 ;
        RECT 159.480 46.485 159.650 46.655 ;
        RECT 169.580 47.505 169.750 47.675 ;
        RECT 162.215 46.145 162.385 46.315 ;
        RECT 169.115 46.825 169.285 46.995 ;
        RECT 170.465 47.165 170.635 47.335 ;
        RECT 170.040 46.485 170.210 46.655 ;
        RECT 171.900 47.505 172.070 47.675 ;
        RECT 171.440 46.485 171.610 46.655 ;
        RECT 173.280 47.505 173.450 47.675 ;
        RECT 173.280 46.485 173.450 46.655 ;
        RECT 185.220 47.505 185.390 47.675 ;
        RECT 184.755 46.825 184.925 46.995 ;
        RECT 186.135 47.165 186.305 47.335 ;
        RECT 185.680 46.485 185.850 46.655 ;
        RECT 187.540 47.505 187.710 47.675 ;
        RECT 187.080 46.485 187.250 46.655 ;
        RECT 188.920 47.505 189.090 47.675 ;
        RECT 188.920 46.485 189.090 46.655 ;
        RECT 191.655 47.505 191.825 47.675 ;
        RECT 197.640 47.505 197.810 47.675 ;
        RECT 197.175 46.825 197.345 46.995 ;
        RECT 198.555 46.825 198.725 46.995 ;
        RECT 198.100 46.485 198.270 46.655 ;
        RECT 199.960 47.505 200.130 47.675 ;
        RECT 199.500 46.485 199.670 46.655 ;
        RECT 201.340 47.505 201.510 47.675 ;
        RECT 201.340 46.485 201.510 46.655 ;
        RECT 205.455 46.485 205.625 46.655 ;
        RECT 211.435 46.485 211.605 46.655 ;
        RECT 212.815 47.845 212.985 48.015 ;
        RECT 214.655 47.505 214.825 47.675 ;
        RECT 212.170 46.825 212.340 46.995 ;
        RECT 213.130 46.825 213.300 46.995 ;
        RECT 219.255 47.505 219.425 47.675 ;
        RECT 222.935 47.165 223.105 47.335 ;
        RECT 220.175 46.825 220.345 46.995 ;
        RECT 220.635 46.825 220.805 46.995 ;
        RECT 230.755 46.485 230.925 46.655 ;
        RECT 232.135 47.845 232.305 48.015 ;
        RECT 231.490 47.165 231.660 47.335 ;
        RECT 232.595 47.165 232.765 47.335 ;
        RECT 234.435 47.165 234.605 47.335 ;
        RECT 239.495 47.165 239.665 47.335 ;
        RECT 240.415 46.825 240.585 46.995 ;
        RECT 241.800 47.165 241.970 47.335 ;
        RECT 242.745 46.825 242.915 46.995 ;
        RECT 243.175 46.825 243.345 46.995 ;
        RECT 244.580 47.165 244.750 47.335 ;
        RECT 245.475 47.165 245.645 47.335 ;
        RECT 250.535 46.825 250.705 46.995 ;
        RECT 251.915 47.505 252.085 47.675 ;
        RECT 252.375 47.165 252.545 47.335 ;
        RECT 258.355 46.485 258.525 46.655 ;
        RECT 259.275 46.825 259.445 46.995 ;
        RECT 261.115 46.825 261.285 46.995 ;
        RECT 268.475 47.845 268.645 48.015 ;
        RECT 267.555 46.825 267.725 46.995 ;
        RECT 274.455 46.825 274.625 46.995 ;
        RECT 275.835 46.825 276.005 46.995 ;
        RECT 273.535 46.145 273.705 46.315 ;
        RECT 284.115 46.825 284.285 46.995 ;
        RECT 287.335 46.825 287.505 46.995 ;
        RECT 288.255 46.825 288.425 46.995 ;
        RECT 290.095 46.825 290.265 46.995 ;
        RECT 291.015 46.825 291.185 46.995 ;
        RECT 285.495 46.145 285.665 46.315 ;
        RECT 297.915 47.165 298.085 47.335 ;
        RECT 298.375 46.825 298.545 46.995 ;
        RECT 304.815 46.825 304.985 46.995 ;
        RECT 306.195 46.825 306.365 46.995 ;
        RECT 311.255 46.825 311.425 46.995 ;
        RECT 314.015 46.825 314.185 46.995 ;
        RECT 303.895 46.145 304.065 46.315 ;
        RECT 325.055 46.825 325.225 46.995 ;
        RECT 326.435 46.825 326.605 46.995 ;
        RECT 312.635 46.145 312.805 46.315 ;
        RECT 332.875 46.825 333.045 46.995 ;
        RECT 333.795 46.825 333.965 46.995 ;
        RECT 324.135 46.145 324.305 46.315 ;
        RECT 335.175 46.485 335.345 46.655 ;
        RECT 340.695 46.825 340.865 46.995 ;
        RECT 342.075 46.825 342.245 46.995 ;
        RECT 353.115 46.825 353.285 46.995 ;
        RECT 354.035 46.825 354.205 46.995 ;
        RECT 339.775 46.145 339.945 46.315 ;
        RECT 360.935 46.825 361.105 46.995 ;
        RECT 361.855 46.825 362.025 46.995 ;
        RECT 352.195 46.145 352.365 46.315 ;
        RECT 370.595 47.165 370.765 47.335 ;
        RECT 368.755 46.825 368.925 46.995 ;
        RECT 369.675 46.825 369.845 46.995 ;
        RECT 360.015 46.145 360.185 46.315 ;
        RECT 390.835 47.505 391.005 47.675 ;
        RECT 385.775 46.825 385.945 46.995 ;
        RECT 400.955 46.825 401.125 46.995 ;
        RECT 408.775 46.825 408.945 46.995 ;
        RECT 413.835 46.825 414.005 46.995 ;
        RECT 418.895 46.825 419.065 46.995 ;
        RECT 423.955 46.825 424.125 46.995 ;
        RECT 429.015 46.825 429.185 46.995 ;
        RECT 441.895 46.825 442.065 46.995 ;
        RECT 446.955 46.825 447.125 46.995 ;
        RECT 452.015 46.825 452.185 46.995 ;
        RECT 457.075 46.825 457.245 46.995 ;
        RECT 469.955 46.825 470.125 46.995 ;
        RECT 475.015 46.825 475.185 46.995 ;
        RECT 480.075 46.825 480.245 46.995 ;
        RECT 485.135 46.825 485.305 46.995 ;
        RECT 492.955 46.825 493.125 46.995 ;
        RECT 498.015 46.825 498.185 46.995 ;
        RECT 503.075 46.825 503.245 46.995 ;
        RECT 508.135 46.825 508.305 46.995 ;
        RECT 521.015 46.825 521.185 46.995 ;
        RECT 526.075 46.825 526.245 46.995 ;
        RECT 531.135 46.825 531.305 46.995 ;
        RECT 536.195 46.825 536.365 46.995 ;
        RECT 541.255 46.825 541.425 46.995 ;
        RECT 549.075 46.825 549.245 46.995 ;
        RECT 554.135 46.825 554.305 46.995 ;
        RECT 559.195 46.825 559.365 46.995 ;
        RECT 564.255 46.825 564.425 46.995 ;
        RECT 569.315 46.825 569.485 46.995 ;
        RECT 577.135 46.825 577.305 46.995 ;
        RECT 582.195 46.825 582.365 46.995 ;
        RECT 587.255 46.825 587.425 46.995 ;
        RECT 592.315 46.825 592.485 46.995 ;
        RECT 597.375 46.825 597.545 46.995 ;
        RECT 605.195 46.825 605.365 46.995 ;
        RECT 610.255 46.825 610.425 46.995 ;
        RECT 615.315 46.825 615.485 46.995 ;
        RECT 620.375 46.825 620.545 46.995 ;
        RECT 625.435 46.825 625.605 46.995 ;
        RECT 42.615 45.635 42.785 45.805 ;
        RECT 43.075 45.635 43.245 45.805 ;
        RECT 43.535 45.635 43.705 45.805 ;
        RECT 43.995 45.635 44.165 45.805 ;
        RECT 44.455 45.635 44.625 45.805 ;
        RECT 44.915 45.635 45.085 45.805 ;
        RECT 45.375 45.635 45.545 45.805 ;
        RECT 45.835 45.635 46.005 45.805 ;
        RECT 46.295 45.635 46.465 45.805 ;
        RECT 46.755 45.635 46.925 45.805 ;
        RECT 47.215 45.635 47.385 45.805 ;
        RECT 47.675 45.635 47.845 45.805 ;
        RECT 48.135 45.635 48.305 45.805 ;
        RECT 48.595 45.635 48.765 45.805 ;
        RECT 49.055 45.635 49.225 45.805 ;
        RECT 49.515 45.635 49.685 45.805 ;
        RECT 49.975 45.635 50.145 45.805 ;
        RECT 50.435 45.635 50.605 45.805 ;
        RECT 50.895 45.635 51.065 45.805 ;
        RECT 51.355 45.635 51.525 45.805 ;
        RECT 51.815 45.635 51.985 45.805 ;
        RECT 52.275 45.635 52.445 45.805 ;
        RECT 52.735 45.635 52.905 45.805 ;
        RECT 53.195 45.635 53.365 45.805 ;
        RECT 53.655 45.635 53.825 45.805 ;
        RECT 54.115 45.635 54.285 45.805 ;
        RECT 54.575 45.635 54.745 45.805 ;
        RECT 55.035 45.635 55.205 45.805 ;
        RECT 55.495 45.635 55.665 45.805 ;
        RECT 55.955 45.635 56.125 45.805 ;
        RECT 56.415 45.635 56.585 45.805 ;
        RECT 56.875 45.635 57.045 45.805 ;
        RECT 57.335 45.635 57.505 45.805 ;
        RECT 57.795 45.635 57.965 45.805 ;
        RECT 58.255 45.635 58.425 45.805 ;
        RECT 58.715 45.635 58.885 45.805 ;
        RECT 59.175 45.635 59.345 45.805 ;
        RECT 59.635 45.635 59.805 45.805 ;
        RECT 60.095 45.635 60.265 45.805 ;
        RECT 60.555 45.635 60.725 45.805 ;
        RECT 61.015 45.635 61.185 45.805 ;
        RECT 61.475 45.635 61.645 45.805 ;
        RECT 61.935 45.635 62.105 45.805 ;
        RECT 62.395 45.635 62.565 45.805 ;
        RECT 62.855 45.635 63.025 45.805 ;
        RECT 63.315 45.635 63.485 45.805 ;
        RECT 63.775 45.635 63.945 45.805 ;
        RECT 64.235 45.635 64.405 45.805 ;
        RECT 64.695 45.635 64.865 45.805 ;
        RECT 65.155 45.635 65.325 45.805 ;
        RECT 65.615 45.635 65.785 45.805 ;
        RECT 66.075 45.635 66.245 45.805 ;
        RECT 66.535 45.635 66.705 45.805 ;
        RECT 66.995 45.635 67.165 45.805 ;
        RECT 67.455 45.635 67.625 45.805 ;
        RECT 67.915 45.635 68.085 45.805 ;
        RECT 68.375 45.635 68.545 45.805 ;
        RECT 68.835 45.635 69.005 45.805 ;
        RECT 69.295 45.635 69.465 45.805 ;
        RECT 69.755 45.635 69.925 45.805 ;
        RECT 70.215 45.635 70.385 45.805 ;
        RECT 70.675 45.635 70.845 45.805 ;
        RECT 71.135 45.635 71.305 45.805 ;
        RECT 71.595 45.635 71.765 45.805 ;
        RECT 72.055 45.635 72.225 45.805 ;
        RECT 72.515 45.635 72.685 45.805 ;
        RECT 72.975 45.635 73.145 45.805 ;
        RECT 73.435 45.635 73.605 45.805 ;
        RECT 73.895 45.635 74.065 45.805 ;
        RECT 74.355 45.635 74.525 45.805 ;
        RECT 74.815 45.635 74.985 45.805 ;
        RECT 75.275 45.635 75.445 45.805 ;
        RECT 75.735 45.635 75.905 45.805 ;
        RECT 76.195 45.635 76.365 45.805 ;
        RECT 76.655 45.635 76.825 45.805 ;
        RECT 77.115 45.635 77.285 45.805 ;
        RECT 77.575 45.635 77.745 45.805 ;
        RECT 78.035 45.635 78.205 45.805 ;
        RECT 78.495 45.635 78.665 45.805 ;
        RECT 78.955 45.635 79.125 45.805 ;
        RECT 79.415 45.635 79.585 45.805 ;
        RECT 79.875 45.635 80.045 45.805 ;
        RECT 80.335 45.635 80.505 45.805 ;
        RECT 80.795 45.635 80.965 45.805 ;
        RECT 81.255 45.635 81.425 45.805 ;
        RECT 81.715 45.635 81.885 45.805 ;
        RECT 82.175 45.635 82.345 45.805 ;
        RECT 82.635 45.635 82.805 45.805 ;
        RECT 83.095 45.635 83.265 45.805 ;
        RECT 83.555 45.635 83.725 45.805 ;
        RECT 84.015 45.635 84.185 45.805 ;
        RECT 84.475 45.635 84.645 45.805 ;
        RECT 84.935 45.635 85.105 45.805 ;
        RECT 85.395 45.635 85.565 45.805 ;
        RECT 85.855 45.635 86.025 45.805 ;
        RECT 86.315 45.635 86.485 45.805 ;
        RECT 86.775 45.635 86.945 45.805 ;
        RECT 87.235 45.635 87.405 45.805 ;
        RECT 87.695 45.635 87.865 45.805 ;
        RECT 88.155 45.635 88.325 45.805 ;
        RECT 88.615 45.635 88.785 45.805 ;
        RECT 89.075 45.635 89.245 45.805 ;
        RECT 89.535 45.635 89.705 45.805 ;
        RECT 89.995 45.635 90.165 45.805 ;
        RECT 90.455 45.635 90.625 45.805 ;
        RECT 90.915 45.635 91.085 45.805 ;
        RECT 91.375 45.635 91.545 45.805 ;
        RECT 91.835 45.635 92.005 45.805 ;
        RECT 92.295 45.635 92.465 45.805 ;
        RECT 92.755 45.635 92.925 45.805 ;
        RECT 93.215 45.635 93.385 45.805 ;
        RECT 93.675 45.635 93.845 45.805 ;
        RECT 94.135 45.635 94.305 45.805 ;
        RECT 94.595 45.635 94.765 45.805 ;
        RECT 95.055 45.635 95.225 45.805 ;
        RECT 95.515 45.635 95.685 45.805 ;
        RECT 95.975 45.635 96.145 45.805 ;
        RECT 96.435 45.635 96.605 45.805 ;
        RECT 96.895 45.635 97.065 45.805 ;
        RECT 97.355 45.635 97.525 45.805 ;
        RECT 97.815 45.635 97.985 45.805 ;
        RECT 98.275 45.635 98.445 45.805 ;
        RECT 98.735 45.635 98.905 45.805 ;
        RECT 99.195 45.635 99.365 45.805 ;
        RECT 99.655 45.635 99.825 45.805 ;
        RECT 100.115 45.635 100.285 45.805 ;
        RECT 100.575 45.635 100.745 45.805 ;
        RECT 101.035 45.635 101.205 45.805 ;
        RECT 101.495 45.635 101.665 45.805 ;
        RECT 101.955 45.635 102.125 45.805 ;
        RECT 102.415 45.635 102.585 45.805 ;
        RECT 102.875 45.635 103.045 45.805 ;
        RECT 103.335 45.635 103.505 45.805 ;
        RECT 103.795 45.635 103.965 45.805 ;
        RECT 104.255 45.635 104.425 45.805 ;
        RECT 104.715 45.635 104.885 45.805 ;
        RECT 105.175 45.635 105.345 45.805 ;
        RECT 105.635 45.635 105.805 45.805 ;
        RECT 106.095 45.635 106.265 45.805 ;
        RECT 106.555 45.635 106.725 45.805 ;
        RECT 107.015 45.635 107.185 45.805 ;
        RECT 107.475 45.635 107.645 45.805 ;
        RECT 107.935 45.635 108.105 45.805 ;
        RECT 108.395 45.635 108.565 45.805 ;
        RECT 108.855 45.635 109.025 45.805 ;
        RECT 109.315 45.635 109.485 45.805 ;
        RECT 109.775 45.635 109.945 45.805 ;
        RECT 110.235 45.635 110.405 45.805 ;
        RECT 110.695 45.635 110.865 45.805 ;
        RECT 111.155 45.635 111.325 45.805 ;
        RECT 111.615 45.635 111.785 45.805 ;
        RECT 112.075 45.635 112.245 45.805 ;
        RECT 112.535 45.635 112.705 45.805 ;
        RECT 112.995 45.635 113.165 45.805 ;
        RECT 113.455 45.635 113.625 45.805 ;
        RECT 113.915 45.635 114.085 45.805 ;
        RECT 114.375 45.635 114.545 45.805 ;
        RECT 114.835 45.635 115.005 45.805 ;
        RECT 115.295 45.635 115.465 45.805 ;
        RECT 115.755 45.635 115.925 45.805 ;
        RECT 116.215 45.635 116.385 45.805 ;
        RECT 116.675 45.635 116.845 45.805 ;
        RECT 117.135 45.635 117.305 45.805 ;
        RECT 117.595 45.635 117.765 45.805 ;
        RECT 118.055 45.635 118.225 45.805 ;
        RECT 118.515 45.635 118.685 45.805 ;
        RECT 118.975 45.635 119.145 45.805 ;
        RECT 119.435 45.635 119.605 45.805 ;
        RECT 119.895 45.635 120.065 45.805 ;
        RECT 120.355 45.635 120.525 45.805 ;
        RECT 120.815 45.635 120.985 45.805 ;
        RECT 121.275 45.635 121.445 45.805 ;
        RECT 121.735 45.635 121.905 45.805 ;
        RECT 122.195 45.635 122.365 45.805 ;
        RECT 122.655 45.635 122.825 45.805 ;
        RECT 123.115 45.635 123.285 45.805 ;
        RECT 123.575 45.635 123.745 45.805 ;
        RECT 124.035 45.635 124.205 45.805 ;
        RECT 124.495 45.635 124.665 45.805 ;
        RECT 124.955 45.635 125.125 45.805 ;
        RECT 125.415 45.635 125.585 45.805 ;
        RECT 125.875 45.635 126.045 45.805 ;
        RECT 126.335 45.635 126.505 45.805 ;
        RECT 126.795 45.635 126.965 45.805 ;
        RECT 127.255 45.635 127.425 45.805 ;
        RECT 127.715 45.635 127.885 45.805 ;
        RECT 128.175 45.635 128.345 45.805 ;
        RECT 128.635 45.635 128.805 45.805 ;
        RECT 129.095 45.635 129.265 45.805 ;
        RECT 129.555 45.635 129.725 45.805 ;
        RECT 130.015 45.635 130.185 45.805 ;
        RECT 130.475 45.635 130.645 45.805 ;
        RECT 130.935 45.635 131.105 45.805 ;
        RECT 131.395 45.635 131.565 45.805 ;
        RECT 131.855 45.635 132.025 45.805 ;
        RECT 132.315 45.635 132.485 45.805 ;
        RECT 132.775 45.635 132.945 45.805 ;
        RECT 133.235 45.635 133.405 45.805 ;
        RECT 133.695 45.635 133.865 45.805 ;
        RECT 134.155 45.635 134.325 45.805 ;
        RECT 134.615 45.635 134.785 45.805 ;
        RECT 135.075 45.635 135.245 45.805 ;
        RECT 135.535 45.635 135.705 45.805 ;
        RECT 135.995 45.635 136.165 45.805 ;
        RECT 136.455 45.635 136.625 45.805 ;
        RECT 136.915 45.635 137.085 45.805 ;
        RECT 137.375 45.635 137.545 45.805 ;
        RECT 137.835 45.635 138.005 45.805 ;
        RECT 138.295 45.635 138.465 45.805 ;
        RECT 138.755 45.635 138.925 45.805 ;
        RECT 139.215 45.635 139.385 45.805 ;
        RECT 139.675 45.635 139.845 45.805 ;
        RECT 140.135 45.635 140.305 45.805 ;
        RECT 140.595 45.635 140.765 45.805 ;
        RECT 141.055 45.635 141.225 45.805 ;
        RECT 141.515 45.635 141.685 45.805 ;
        RECT 141.975 45.635 142.145 45.805 ;
        RECT 142.435 45.635 142.605 45.805 ;
        RECT 142.895 45.635 143.065 45.805 ;
        RECT 143.355 45.635 143.525 45.805 ;
        RECT 143.815 45.635 143.985 45.805 ;
        RECT 144.275 45.635 144.445 45.805 ;
        RECT 144.735 45.635 144.905 45.805 ;
        RECT 145.195 45.635 145.365 45.805 ;
        RECT 145.655 45.635 145.825 45.805 ;
        RECT 146.115 45.635 146.285 45.805 ;
        RECT 146.575 45.635 146.745 45.805 ;
        RECT 147.035 45.635 147.205 45.805 ;
        RECT 147.495 45.635 147.665 45.805 ;
        RECT 147.955 45.635 148.125 45.805 ;
        RECT 148.415 45.635 148.585 45.805 ;
        RECT 148.875 45.635 149.045 45.805 ;
        RECT 149.335 45.635 149.505 45.805 ;
        RECT 149.795 45.635 149.965 45.805 ;
        RECT 150.255 45.635 150.425 45.805 ;
        RECT 150.715 45.635 150.885 45.805 ;
        RECT 151.175 45.635 151.345 45.805 ;
        RECT 151.635 45.635 151.805 45.805 ;
        RECT 152.095 45.635 152.265 45.805 ;
        RECT 152.555 45.635 152.725 45.805 ;
        RECT 153.015 45.635 153.185 45.805 ;
        RECT 153.475 45.635 153.645 45.805 ;
        RECT 153.935 45.635 154.105 45.805 ;
        RECT 154.395 45.635 154.565 45.805 ;
        RECT 154.855 45.635 155.025 45.805 ;
        RECT 155.315 45.635 155.485 45.805 ;
        RECT 155.775 45.635 155.945 45.805 ;
        RECT 156.235 45.635 156.405 45.805 ;
        RECT 156.695 45.635 156.865 45.805 ;
        RECT 157.155 45.635 157.325 45.805 ;
        RECT 157.615 45.635 157.785 45.805 ;
        RECT 158.075 45.635 158.245 45.805 ;
        RECT 158.535 45.635 158.705 45.805 ;
        RECT 158.995 45.635 159.165 45.805 ;
        RECT 159.455 45.635 159.625 45.805 ;
        RECT 159.915 45.635 160.085 45.805 ;
        RECT 160.375 45.635 160.545 45.805 ;
        RECT 160.835 45.635 161.005 45.805 ;
        RECT 161.295 45.635 161.465 45.805 ;
        RECT 161.755 45.635 161.925 45.805 ;
        RECT 162.215 45.635 162.385 45.805 ;
        RECT 162.675 45.635 162.845 45.805 ;
        RECT 163.135 45.635 163.305 45.805 ;
        RECT 163.595 45.635 163.765 45.805 ;
        RECT 164.055 45.635 164.225 45.805 ;
        RECT 164.515 45.635 164.685 45.805 ;
        RECT 164.975 45.635 165.145 45.805 ;
        RECT 165.435 45.635 165.605 45.805 ;
        RECT 165.895 45.635 166.065 45.805 ;
        RECT 166.355 45.635 166.525 45.805 ;
        RECT 166.815 45.635 166.985 45.805 ;
        RECT 167.275 45.635 167.445 45.805 ;
        RECT 167.735 45.635 167.905 45.805 ;
        RECT 168.195 45.635 168.365 45.805 ;
        RECT 168.655 45.635 168.825 45.805 ;
        RECT 169.115 45.635 169.285 45.805 ;
        RECT 169.575 45.635 169.745 45.805 ;
        RECT 170.035 45.635 170.205 45.805 ;
        RECT 170.495 45.635 170.665 45.805 ;
        RECT 170.955 45.635 171.125 45.805 ;
        RECT 171.415 45.635 171.585 45.805 ;
        RECT 171.875 45.635 172.045 45.805 ;
        RECT 172.335 45.635 172.505 45.805 ;
        RECT 172.795 45.635 172.965 45.805 ;
        RECT 173.255 45.635 173.425 45.805 ;
        RECT 173.715 45.635 173.885 45.805 ;
        RECT 174.175 45.635 174.345 45.805 ;
        RECT 174.635 45.635 174.805 45.805 ;
        RECT 175.095 45.635 175.265 45.805 ;
        RECT 175.555 45.635 175.725 45.805 ;
        RECT 176.015 45.635 176.185 45.805 ;
        RECT 176.475 45.635 176.645 45.805 ;
        RECT 176.935 45.635 177.105 45.805 ;
        RECT 177.395 45.635 177.565 45.805 ;
        RECT 177.855 45.635 178.025 45.805 ;
        RECT 178.315 45.635 178.485 45.805 ;
        RECT 178.775 45.635 178.945 45.805 ;
        RECT 179.235 45.635 179.405 45.805 ;
        RECT 179.695 45.635 179.865 45.805 ;
        RECT 180.155 45.635 180.325 45.805 ;
        RECT 180.615 45.635 180.785 45.805 ;
        RECT 181.075 45.635 181.245 45.805 ;
        RECT 181.535 45.635 181.705 45.805 ;
        RECT 181.995 45.635 182.165 45.805 ;
        RECT 182.455 45.635 182.625 45.805 ;
        RECT 182.915 45.635 183.085 45.805 ;
        RECT 183.375 45.635 183.545 45.805 ;
        RECT 183.835 45.635 184.005 45.805 ;
        RECT 184.295 45.635 184.465 45.805 ;
        RECT 184.755 45.635 184.925 45.805 ;
        RECT 185.215 45.635 185.385 45.805 ;
        RECT 185.675 45.635 185.845 45.805 ;
        RECT 186.135 45.635 186.305 45.805 ;
        RECT 186.595 45.635 186.765 45.805 ;
        RECT 187.055 45.635 187.225 45.805 ;
        RECT 187.515 45.635 187.685 45.805 ;
        RECT 187.975 45.635 188.145 45.805 ;
        RECT 188.435 45.635 188.605 45.805 ;
        RECT 188.895 45.635 189.065 45.805 ;
        RECT 189.355 45.635 189.525 45.805 ;
        RECT 189.815 45.635 189.985 45.805 ;
        RECT 190.275 45.635 190.445 45.805 ;
        RECT 190.735 45.635 190.905 45.805 ;
        RECT 191.195 45.635 191.365 45.805 ;
        RECT 191.655 45.635 191.825 45.805 ;
        RECT 192.115 45.635 192.285 45.805 ;
        RECT 192.575 45.635 192.745 45.805 ;
        RECT 193.035 45.635 193.205 45.805 ;
        RECT 193.495 45.635 193.665 45.805 ;
        RECT 193.955 45.635 194.125 45.805 ;
        RECT 194.415 45.635 194.585 45.805 ;
        RECT 194.875 45.635 195.045 45.805 ;
        RECT 195.335 45.635 195.505 45.805 ;
        RECT 195.795 45.635 195.965 45.805 ;
        RECT 196.255 45.635 196.425 45.805 ;
        RECT 196.715 45.635 196.885 45.805 ;
        RECT 197.175 45.635 197.345 45.805 ;
        RECT 197.635 45.635 197.805 45.805 ;
        RECT 198.095 45.635 198.265 45.805 ;
        RECT 198.555 45.635 198.725 45.805 ;
        RECT 199.015 45.635 199.185 45.805 ;
        RECT 199.475 45.635 199.645 45.805 ;
        RECT 199.935 45.635 200.105 45.805 ;
        RECT 200.395 45.635 200.565 45.805 ;
        RECT 200.855 45.635 201.025 45.805 ;
        RECT 201.315 45.635 201.485 45.805 ;
        RECT 201.775 45.635 201.945 45.805 ;
        RECT 202.235 45.635 202.405 45.805 ;
        RECT 202.695 45.635 202.865 45.805 ;
        RECT 203.155 45.635 203.325 45.805 ;
        RECT 203.615 45.635 203.785 45.805 ;
        RECT 204.075 45.635 204.245 45.805 ;
        RECT 204.535 45.635 204.705 45.805 ;
        RECT 204.995 45.635 205.165 45.805 ;
        RECT 205.455 45.635 205.625 45.805 ;
        RECT 205.915 45.635 206.085 45.805 ;
        RECT 206.375 45.635 206.545 45.805 ;
        RECT 206.835 45.635 207.005 45.805 ;
        RECT 207.295 45.635 207.465 45.805 ;
        RECT 207.755 45.635 207.925 45.805 ;
        RECT 208.215 45.635 208.385 45.805 ;
        RECT 208.675 45.635 208.845 45.805 ;
        RECT 209.135 45.635 209.305 45.805 ;
        RECT 209.595 45.635 209.765 45.805 ;
        RECT 210.055 45.635 210.225 45.805 ;
        RECT 210.515 45.635 210.685 45.805 ;
        RECT 210.975 45.635 211.145 45.805 ;
        RECT 211.435 45.635 211.605 45.805 ;
        RECT 211.895 45.635 212.065 45.805 ;
        RECT 212.355 45.635 212.525 45.805 ;
        RECT 212.815 45.635 212.985 45.805 ;
        RECT 213.275 45.635 213.445 45.805 ;
        RECT 213.735 45.635 213.905 45.805 ;
        RECT 214.195 45.635 214.365 45.805 ;
        RECT 214.655 45.635 214.825 45.805 ;
        RECT 215.115 45.635 215.285 45.805 ;
        RECT 215.575 45.635 215.745 45.805 ;
        RECT 216.035 45.635 216.205 45.805 ;
        RECT 216.495 45.635 216.665 45.805 ;
        RECT 216.955 45.635 217.125 45.805 ;
        RECT 217.415 45.635 217.585 45.805 ;
        RECT 217.875 45.635 218.045 45.805 ;
        RECT 218.335 45.635 218.505 45.805 ;
        RECT 218.795 45.635 218.965 45.805 ;
        RECT 219.255 45.635 219.425 45.805 ;
        RECT 219.715 45.635 219.885 45.805 ;
        RECT 220.175 45.635 220.345 45.805 ;
        RECT 220.635 45.635 220.805 45.805 ;
        RECT 221.095 45.635 221.265 45.805 ;
        RECT 221.555 45.635 221.725 45.805 ;
        RECT 222.015 45.635 222.185 45.805 ;
        RECT 222.475 45.635 222.645 45.805 ;
        RECT 222.935 45.635 223.105 45.805 ;
        RECT 223.395 45.635 223.565 45.805 ;
        RECT 223.855 45.635 224.025 45.805 ;
        RECT 224.315 45.635 224.485 45.805 ;
        RECT 224.775 45.635 224.945 45.805 ;
        RECT 225.235 45.635 225.405 45.805 ;
        RECT 225.695 45.635 225.865 45.805 ;
        RECT 226.155 45.635 226.325 45.805 ;
        RECT 226.615 45.635 226.785 45.805 ;
        RECT 227.075 45.635 227.245 45.805 ;
        RECT 227.535 45.635 227.705 45.805 ;
        RECT 227.995 45.635 228.165 45.805 ;
        RECT 228.455 45.635 228.625 45.805 ;
        RECT 228.915 45.635 229.085 45.805 ;
        RECT 229.375 45.635 229.545 45.805 ;
        RECT 229.835 45.635 230.005 45.805 ;
        RECT 230.295 45.635 230.465 45.805 ;
        RECT 230.755 45.635 230.925 45.805 ;
        RECT 231.215 45.635 231.385 45.805 ;
        RECT 231.675 45.635 231.845 45.805 ;
        RECT 232.135 45.635 232.305 45.805 ;
        RECT 232.595 45.635 232.765 45.805 ;
        RECT 233.055 45.635 233.225 45.805 ;
        RECT 233.515 45.635 233.685 45.805 ;
        RECT 233.975 45.635 234.145 45.805 ;
        RECT 234.435 45.635 234.605 45.805 ;
        RECT 234.895 45.635 235.065 45.805 ;
        RECT 235.355 45.635 235.525 45.805 ;
        RECT 235.815 45.635 235.985 45.805 ;
        RECT 236.275 45.635 236.445 45.805 ;
        RECT 236.735 45.635 236.905 45.805 ;
        RECT 237.195 45.635 237.365 45.805 ;
        RECT 237.655 45.635 237.825 45.805 ;
        RECT 238.115 45.635 238.285 45.805 ;
        RECT 238.575 45.635 238.745 45.805 ;
        RECT 239.035 45.635 239.205 45.805 ;
        RECT 239.495 45.635 239.665 45.805 ;
        RECT 239.955 45.635 240.125 45.805 ;
        RECT 240.415 45.635 240.585 45.805 ;
        RECT 240.875 45.635 241.045 45.805 ;
        RECT 241.335 45.635 241.505 45.805 ;
        RECT 241.795 45.635 241.965 45.805 ;
        RECT 242.255 45.635 242.425 45.805 ;
        RECT 242.715 45.635 242.885 45.805 ;
        RECT 243.175 45.635 243.345 45.805 ;
        RECT 243.635 45.635 243.805 45.805 ;
        RECT 244.095 45.635 244.265 45.805 ;
        RECT 244.555 45.635 244.725 45.805 ;
        RECT 245.015 45.635 245.185 45.805 ;
        RECT 245.475 45.635 245.645 45.805 ;
        RECT 245.935 45.635 246.105 45.805 ;
        RECT 246.395 45.635 246.565 45.805 ;
        RECT 246.855 45.635 247.025 45.805 ;
        RECT 247.315 45.635 247.485 45.805 ;
        RECT 247.775 45.635 247.945 45.805 ;
        RECT 248.235 45.635 248.405 45.805 ;
        RECT 248.695 45.635 248.865 45.805 ;
        RECT 249.155 45.635 249.325 45.805 ;
        RECT 249.615 45.635 249.785 45.805 ;
        RECT 250.075 45.635 250.245 45.805 ;
        RECT 250.535 45.635 250.705 45.805 ;
        RECT 250.995 45.635 251.165 45.805 ;
        RECT 251.455 45.635 251.625 45.805 ;
        RECT 251.915 45.635 252.085 45.805 ;
        RECT 252.375 45.635 252.545 45.805 ;
        RECT 252.835 45.635 253.005 45.805 ;
        RECT 253.295 45.635 253.465 45.805 ;
        RECT 253.755 45.635 253.925 45.805 ;
        RECT 254.215 45.635 254.385 45.805 ;
        RECT 254.675 45.635 254.845 45.805 ;
        RECT 255.135 45.635 255.305 45.805 ;
        RECT 255.595 45.635 255.765 45.805 ;
        RECT 256.055 45.635 256.225 45.805 ;
        RECT 256.515 45.635 256.685 45.805 ;
        RECT 256.975 45.635 257.145 45.805 ;
        RECT 257.435 45.635 257.605 45.805 ;
        RECT 257.895 45.635 258.065 45.805 ;
        RECT 258.355 45.635 258.525 45.805 ;
        RECT 258.815 45.635 258.985 45.805 ;
        RECT 259.275 45.635 259.445 45.805 ;
        RECT 259.735 45.635 259.905 45.805 ;
        RECT 260.195 45.635 260.365 45.805 ;
        RECT 260.655 45.635 260.825 45.805 ;
        RECT 261.115 45.635 261.285 45.805 ;
        RECT 261.575 45.635 261.745 45.805 ;
        RECT 262.035 45.635 262.205 45.805 ;
        RECT 262.495 45.635 262.665 45.805 ;
        RECT 262.955 45.635 263.125 45.805 ;
        RECT 263.415 45.635 263.585 45.805 ;
        RECT 263.875 45.635 264.045 45.805 ;
        RECT 264.335 45.635 264.505 45.805 ;
        RECT 264.795 45.635 264.965 45.805 ;
        RECT 265.255 45.635 265.425 45.805 ;
        RECT 265.715 45.635 265.885 45.805 ;
        RECT 266.175 45.635 266.345 45.805 ;
        RECT 266.635 45.635 266.805 45.805 ;
        RECT 267.095 45.635 267.265 45.805 ;
        RECT 267.555 45.635 267.725 45.805 ;
        RECT 268.015 45.635 268.185 45.805 ;
        RECT 268.475 45.635 268.645 45.805 ;
        RECT 268.935 45.635 269.105 45.805 ;
        RECT 269.395 45.635 269.565 45.805 ;
        RECT 269.855 45.635 270.025 45.805 ;
        RECT 270.315 45.635 270.485 45.805 ;
        RECT 270.775 45.635 270.945 45.805 ;
        RECT 271.235 45.635 271.405 45.805 ;
        RECT 271.695 45.635 271.865 45.805 ;
        RECT 272.155 45.635 272.325 45.805 ;
        RECT 272.615 45.635 272.785 45.805 ;
        RECT 273.075 45.635 273.245 45.805 ;
        RECT 273.535 45.635 273.705 45.805 ;
        RECT 273.995 45.635 274.165 45.805 ;
        RECT 274.455 45.635 274.625 45.805 ;
        RECT 274.915 45.635 275.085 45.805 ;
        RECT 275.375 45.635 275.545 45.805 ;
        RECT 275.835 45.635 276.005 45.805 ;
        RECT 276.295 45.635 276.465 45.805 ;
        RECT 276.755 45.635 276.925 45.805 ;
        RECT 277.215 45.635 277.385 45.805 ;
        RECT 277.675 45.635 277.845 45.805 ;
        RECT 278.135 45.635 278.305 45.805 ;
        RECT 278.595 45.635 278.765 45.805 ;
        RECT 279.055 45.635 279.225 45.805 ;
        RECT 279.515 45.635 279.685 45.805 ;
        RECT 279.975 45.635 280.145 45.805 ;
        RECT 280.435 45.635 280.605 45.805 ;
        RECT 280.895 45.635 281.065 45.805 ;
        RECT 281.355 45.635 281.525 45.805 ;
        RECT 281.815 45.635 281.985 45.805 ;
        RECT 282.275 45.635 282.445 45.805 ;
        RECT 282.735 45.635 282.905 45.805 ;
        RECT 283.195 45.635 283.365 45.805 ;
        RECT 283.655 45.635 283.825 45.805 ;
        RECT 284.115 45.635 284.285 45.805 ;
        RECT 284.575 45.635 284.745 45.805 ;
        RECT 285.035 45.635 285.205 45.805 ;
        RECT 285.495 45.635 285.665 45.805 ;
        RECT 285.955 45.635 286.125 45.805 ;
        RECT 286.415 45.635 286.585 45.805 ;
        RECT 286.875 45.635 287.045 45.805 ;
        RECT 287.335 45.635 287.505 45.805 ;
        RECT 287.795 45.635 287.965 45.805 ;
        RECT 288.255 45.635 288.425 45.805 ;
        RECT 288.715 45.635 288.885 45.805 ;
        RECT 289.175 45.635 289.345 45.805 ;
        RECT 289.635 45.635 289.805 45.805 ;
        RECT 290.095 45.635 290.265 45.805 ;
        RECT 290.555 45.635 290.725 45.805 ;
        RECT 291.015 45.635 291.185 45.805 ;
        RECT 291.475 45.635 291.645 45.805 ;
        RECT 291.935 45.635 292.105 45.805 ;
        RECT 292.395 45.635 292.565 45.805 ;
        RECT 292.855 45.635 293.025 45.805 ;
        RECT 293.315 45.635 293.485 45.805 ;
        RECT 293.775 45.635 293.945 45.805 ;
        RECT 294.235 45.635 294.405 45.805 ;
        RECT 294.695 45.635 294.865 45.805 ;
        RECT 295.155 45.635 295.325 45.805 ;
        RECT 295.615 45.635 295.785 45.805 ;
        RECT 296.075 45.635 296.245 45.805 ;
        RECT 296.535 45.635 296.705 45.805 ;
        RECT 296.995 45.635 297.165 45.805 ;
        RECT 297.455 45.635 297.625 45.805 ;
        RECT 297.915 45.635 298.085 45.805 ;
        RECT 298.375 45.635 298.545 45.805 ;
        RECT 298.835 45.635 299.005 45.805 ;
        RECT 299.295 45.635 299.465 45.805 ;
        RECT 299.755 45.635 299.925 45.805 ;
        RECT 300.215 45.635 300.385 45.805 ;
        RECT 300.675 45.635 300.845 45.805 ;
        RECT 301.135 45.635 301.305 45.805 ;
        RECT 301.595 45.635 301.765 45.805 ;
        RECT 302.055 45.635 302.225 45.805 ;
        RECT 302.515 45.635 302.685 45.805 ;
        RECT 302.975 45.635 303.145 45.805 ;
        RECT 303.435 45.635 303.605 45.805 ;
        RECT 303.895 45.635 304.065 45.805 ;
        RECT 304.355 45.635 304.525 45.805 ;
        RECT 304.815 45.635 304.985 45.805 ;
        RECT 305.275 45.635 305.445 45.805 ;
        RECT 305.735 45.635 305.905 45.805 ;
        RECT 306.195 45.635 306.365 45.805 ;
        RECT 306.655 45.635 306.825 45.805 ;
        RECT 307.115 45.635 307.285 45.805 ;
        RECT 307.575 45.635 307.745 45.805 ;
        RECT 308.035 45.635 308.205 45.805 ;
        RECT 308.495 45.635 308.665 45.805 ;
        RECT 308.955 45.635 309.125 45.805 ;
        RECT 309.415 45.635 309.585 45.805 ;
        RECT 309.875 45.635 310.045 45.805 ;
        RECT 310.335 45.635 310.505 45.805 ;
        RECT 310.795 45.635 310.965 45.805 ;
        RECT 311.255 45.635 311.425 45.805 ;
        RECT 311.715 45.635 311.885 45.805 ;
        RECT 312.175 45.635 312.345 45.805 ;
        RECT 312.635 45.635 312.805 45.805 ;
        RECT 313.095 45.635 313.265 45.805 ;
        RECT 313.555 45.635 313.725 45.805 ;
        RECT 314.015 45.635 314.185 45.805 ;
        RECT 314.475 45.635 314.645 45.805 ;
        RECT 314.935 45.635 315.105 45.805 ;
        RECT 315.395 45.635 315.565 45.805 ;
        RECT 315.855 45.635 316.025 45.805 ;
        RECT 316.315 45.635 316.485 45.805 ;
        RECT 316.775 45.635 316.945 45.805 ;
        RECT 317.235 45.635 317.405 45.805 ;
        RECT 317.695 45.635 317.865 45.805 ;
        RECT 318.155 45.635 318.325 45.805 ;
        RECT 318.615 45.635 318.785 45.805 ;
        RECT 319.075 45.635 319.245 45.805 ;
        RECT 319.535 45.635 319.705 45.805 ;
        RECT 319.995 45.635 320.165 45.805 ;
        RECT 320.455 45.635 320.625 45.805 ;
        RECT 320.915 45.635 321.085 45.805 ;
        RECT 321.375 45.635 321.545 45.805 ;
        RECT 321.835 45.635 322.005 45.805 ;
        RECT 322.295 45.635 322.465 45.805 ;
        RECT 322.755 45.635 322.925 45.805 ;
        RECT 323.215 45.635 323.385 45.805 ;
        RECT 323.675 45.635 323.845 45.805 ;
        RECT 324.135 45.635 324.305 45.805 ;
        RECT 324.595 45.635 324.765 45.805 ;
        RECT 325.055 45.635 325.225 45.805 ;
        RECT 325.515 45.635 325.685 45.805 ;
        RECT 325.975 45.635 326.145 45.805 ;
        RECT 326.435 45.635 326.605 45.805 ;
        RECT 326.895 45.635 327.065 45.805 ;
        RECT 327.355 45.635 327.525 45.805 ;
        RECT 327.815 45.635 327.985 45.805 ;
        RECT 328.275 45.635 328.445 45.805 ;
        RECT 328.735 45.635 328.905 45.805 ;
        RECT 329.195 45.635 329.365 45.805 ;
        RECT 329.655 45.635 329.825 45.805 ;
        RECT 330.115 45.635 330.285 45.805 ;
        RECT 330.575 45.635 330.745 45.805 ;
        RECT 331.035 45.635 331.205 45.805 ;
        RECT 331.495 45.635 331.665 45.805 ;
        RECT 331.955 45.635 332.125 45.805 ;
        RECT 332.415 45.635 332.585 45.805 ;
        RECT 332.875 45.635 333.045 45.805 ;
        RECT 333.335 45.635 333.505 45.805 ;
        RECT 333.795 45.635 333.965 45.805 ;
        RECT 334.255 45.635 334.425 45.805 ;
        RECT 334.715 45.635 334.885 45.805 ;
        RECT 335.175 45.635 335.345 45.805 ;
        RECT 335.635 45.635 335.805 45.805 ;
        RECT 336.095 45.635 336.265 45.805 ;
        RECT 336.555 45.635 336.725 45.805 ;
        RECT 337.015 45.635 337.185 45.805 ;
        RECT 337.475 45.635 337.645 45.805 ;
        RECT 337.935 45.635 338.105 45.805 ;
        RECT 338.395 45.635 338.565 45.805 ;
        RECT 338.855 45.635 339.025 45.805 ;
        RECT 339.315 45.635 339.485 45.805 ;
        RECT 339.775 45.635 339.945 45.805 ;
        RECT 340.235 45.635 340.405 45.805 ;
        RECT 340.695 45.635 340.865 45.805 ;
        RECT 341.155 45.635 341.325 45.805 ;
        RECT 341.615 45.635 341.785 45.805 ;
        RECT 342.075 45.635 342.245 45.805 ;
        RECT 342.535 45.635 342.705 45.805 ;
        RECT 342.995 45.635 343.165 45.805 ;
        RECT 343.455 45.635 343.625 45.805 ;
        RECT 343.915 45.635 344.085 45.805 ;
        RECT 344.375 45.635 344.545 45.805 ;
        RECT 344.835 45.635 345.005 45.805 ;
        RECT 345.295 45.635 345.465 45.805 ;
        RECT 345.755 45.635 345.925 45.805 ;
        RECT 346.215 45.635 346.385 45.805 ;
        RECT 346.675 45.635 346.845 45.805 ;
        RECT 347.135 45.635 347.305 45.805 ;
        RECT 347.595 45.635 347.765 45.805 ;
        RECT 348.055 45.635 348.225 45.805 ;
        RECT 348.515 45.635 348.685 45.805 ;
        RECT 348.975 45.635 349.145 45.805 ;
        RECT 349.435 45.635 349.605 45.805 ;
        RECT 349.895 45.635 350.065 45.805 ;
        RECT 350.355 45.635 350.525 45.805 ;
        RECT 350.815 45.635 350.985 45.805 ;
        RECT 351.275 45.635 351.445 45.805 ;
        RECT 351.735 45.635 351.905 45.805 ;
        RECT 352.195 45.635 352.365 45.805 ;
        RECT 352.655 45.635 352.825 45.805 ;
        RECT 353.115 45.635 353.285 45.805 ;
        RECT 353.575 45.635 353.745 45.805 ;
        RECT 354.035 45.635 354.205 45.805 ;
        RECT 354.495 45.635 354.665 45.805 ;
        RECT 354.955 45.635 355.125 45.805 ;
        RECT 355.415 45.635 355.585 45.805 ;
        RECT 355.875 45.635 356.045 45.805 ;
        RECT 356.335 45.635 356.505 45.805 ;
        RECT 356.795 45.635 356.965 45.805 ;
        RECT 357.255 45.635 357.425 45.805 ;
        RECT 357.715 45.635 357.885 45.805 ;
        RECT 358.175 45.635 358.345 45.805 ;
        RECT 358.635 45.635 358.805 45.805 ;
        RECT 359.095 45.635 359.265 45.805 ;
        RECT 359.555 45.635 359.725 45.805 ;
        RECT 360.015 45.635 360.185 45.805 ;
        RECT 360.475 45.635 360.645 45.805 ;
        RECT 360.935 45.635 361.105 45.805 ;
        RECT 361.395 45.635 361.565 45.805 ;
        RECT 361.855 45.635 362.025 45.805 ;
        RECT 362.315 45.635 362.485 45.805 ;
        RECT 362.775 45.635 362.945 45.805 ;
        RECT 363.235 45.635 363.405 45.805 ;
        RECT 363.695 45.635 363.865 45.805 ;
        RECT 364.155 45.635 364.325 45.805 ;
        RECT 364.615 45.635 364.785 45.805 ;
        RECT 365.075 45.635 365.245 45.805 ;
        RECT 365.535 45.635 365.705 45.805 ;
        RECT 365.995 45.635 366.165 45.805 ;
        RECT 366.455 45.635 366.625 45.805 ;
        RECT 366.915 45.635 367.085 45.805 ;
        RECT 367.375 45.635 367.545 45.805 ;
        RECT 367.835 45.635 368.005 45.805 ;
        RECT 368.295 45.635 368.465 45.805 ;
        RECT 368.755 45.635 368.925 45.805 ;
        RECT 369.215 45.635 369.385 45.805 ;
        RECT 369.675 45.635 369.845 45.805 ;
        RECT 370.135 45.635 370.305 45.805 ;
        RECT 370.595 45.635 370.765 45.805 ;
        RECT 371.055 45.635 371.225 45.805 ;
        RECT 371.515 45.635 371.685 45.805 ;
        RECT 371.975 45.635 372.145 45.805 ;
        RECT 372.435 45.635 372.605 45.805 ;
        RECT 372.895 45.635 373.065 45.805 ;
        RECT 373.355 45.635 373.525 45.805 ;
        RECT 373.815 45.635 373.985 45.805 ;
        RECT 374.275 45.635 374.445 45.805 ;
        RECT 374.735 45.635 374.905 45.805 ;
        RECT 375.195 45.635 375.365 45.805 ;
        RECT 375.655 45.635 375.825 45.805 ;
        RECT 376.115 45.635 376.285 45.805 ;
        RECT 376.575 45.635 376.745 45.805 ;
        RECT 377.035 45.635 377.205 45.805 ;
        RECT 377.495 45.635 377.665 45.805 ;
        RECT 377.955 45.635 378.125 45.805 ;
        RECT 378.415 45.635 378.585 45.805 ;
        RECT 378.875 45.635 379.045 45.805 ;
        RECT 379.335 45.635 379.505 45.805 ;
        RECT 379.795 45.635 379.965 45.805 ;
        RECT 380.255 45.635 380.425 45.805 ;
        RECT 380.715 45.635 380.885 45.805 ;
        RECT 381.175 45.635 381.345 45.805 ;
        RECT 381.635 45.635 381.805 45.805 ;
        RECT 382.095 45.635 382.265 45.805 ;
        RECT 382.555 45.635 382.725 45.805 ;
        RECT 383.015 45.635 383.185 45.805 ;
        RECT 383.475 45.635 383.645 45.805 ;
        RECT 383.935 45.635 384.105 45.805 ;
        RECT 384.395 45.635 384.565 45.805 ;
        RECT 384.855 45.635 385.025 45.805 ;
        RECT 385.315 45.635 385.485 45.805 ;
        RECT 385.775 45.635 385.945 45.805 ;
        RECT 386.235 45.635 386.405 45.805 ;
        RECT 386.695 45.635 386.865 45.805 ;
        RECT 387.155 45.635 387.325 45.805 ;
        RECT 387.615 45.635 387.785 45.805 ;
        RECT 388.075 45.635 388.245 45.805 ;
        RECT 388.535 45.635 388.705 45.805 ;
        RECT 388.995 45.635 389.165 45.805 ;
        RECT 389.455 45.635 389.625 45.805 ;
        RECT 389.915 45.635 390.085 45.805 ;
        RECT 390.375 45.635 390.545 45.805 ;
        RECT 390.835 45.635 391.005 45.805 ;
        RECT 391.295 45.635 391.465 45.805 ;
        RECT 391.755 45.635 391.925 45.805 ;
        RECT 392.215 45.635 392.385 45.805 ;
        RECT 392.675 45.635 392.845 45.805 ;
        RECT 393.135 45.635 393.305 45.805 ;
        RECT 393.595 45.635 393.765 45.805 ;
        RECT 394.055 45.635 394.225 45.805 ;
        RECT 394.515 45.635 394.685 45.805 ;
        RECT 394.975 45.635 395.145 45.805 ;
        RECT 395.435 45.635 395.605 45.805 ;
        RECT 395.895 45.635 396.065 45.805 ;
        RECT 396.355 45.635 396.525 45.805 ;
        RECT 396.815 45.635 396.985 45.805 ;
        RECT 397.275 45.635 397.445 45.805 ;
        RECT 397.735 45.635 397.905 45.805 ;
        RECT 398.195 45.635 398.365 45.805 ;
        RECT 398.655 45.635 398.825 45.805 ;
        RECT 399.115 45.635 399.285 45.805 ;
        RECT 399.575 45.635 399.745 45.805 ;
        RECT 400.035 45.635 400.205 45.805 ;
        RECT 400.495 45.635 400.665 45.805 ;
        RECT 400.955 45.635 401.125 45.805 ;
        RECT 401.415 45.635 401.585 45.805 ;
        RECT 401.875 45.635 402.045 45.805 ;
        RECT 402.335 45.635 402.505 45.805 ;
        RECT 402.795 45.635 402.965 45.805 ;
        RECT 403.255 45.635 403.425 45.805 ;
        RECT 403.715 45.635 403.885 45.805 ;
        RECT 404.175 45.635 404.345 45.805 ;
        RECT 404.635 45.635 404.805 45.805 ;
        RECT 405.095 45.635 405.265 45.805 ;
        RECT 405.555 45.635 405.725 45.805 ;
        RECT 406.015 45.635 406.185 45.805 ;
        RECT 406.475 45.635 406.645 45.805 ;
        RECT 406.935 45.635 407.105 45.805 ;
        RECT 407.395 45.635 407.565 45.805 ;
        RECT 407.855 45.635 408.025 45.805 ;
        RECT 408.315 45.635 408.485 45.805 ;
        RECT 408.775 45.635 408.945 45.805 ;
        RECT 409.235 45.635 409.405 45.805 ;
        RECT 409.695 45.635 409.865 45.805 ;
        RECT 410.155 45.635 410.325 45.805 ;
        RECT 410.615 45.635 410.785 45.805 ;
        RECT 411.075 45.635 411.245 45.805 ;
        RECT 411.535 45.635 411.705 45.805 ;
        RECT 411.995 45.635 412.165 45.805 ;
        RECT 412.455 45.635 412.625 45.805 ;
        RECT 412.915 45.635 413.085 45.805 ;
        RECT 413.375 45.635 413.545 45.805 ;
        RECT 413.835 45.635 414.005 45.805 ;
        RECT 414.295 45.635 414.465 45.805 ;
        RECT 414.755 45.635 414.925 45.805 ;
        RECT 415.215 45.635 415.385 45.805 ;
        RECT 415.675 45.635 415.845 45.805 ;
        RECT 416.135 45.635 416.305 45.805 ;
        RECT 416.595 45.635 416.765 45.805 ;
        RECT 417.055 45.635 417.225 45.805 ;
        RECT 417.515 45.635 417.685 45.805 ;
        RECT 417.975 45.635 418.145 45.805 ;
        RECT 418.435 45.635 418.605 45.805 ;
        RECT 418.895 45.635 419.065 45.805 ;
        RECT 419.355 45.635 419.525 45.805 ;
        RECT 419.815 45.635 419.985 45.805 ;
        RECT 420.275 45.635 420.445 45.805 ;
        RECT 420.735 45.635 420.905 45.805 ;
        RECT 421.195 45.635 421.365 45.805 ;
        RECT 421.655 45.635 421.825 45.805 ;
        RECT 422.115 45.635 422.285 45.805 ;
        RECT 422.575 45.635 422.745 45.805 ;
        RECT 423.035 45.635 423.205 45.805 ;
        RECT 423.495 45.635 423.665 45.805 ;
        RECT 423.955 45.635 424.125 45.805 ;
        RECT 424.415 45.635 424.585 45.805 ;
        RECT 424.875 45.635 425.045 45.805 ;
        RECT 425.335 45.635 425.505 45.805 ;
        RECT 425.795 45.635 425.965 45.805 ;
        RECT 426.255 45.635 426.425 45.805 ;
        RECT 426.715 45.635 426.885 45.805 ;
        RECT 427.175 45.635 427.345 45.805 ;
        RECT 427.635 45.635 427.805 45.805 ;
        RECT 428.095 45.635 428.265 45.805 ;
        RECT 428.555 45.635 428.725 45.805 ;
        RECT 429.015 45.635 429.185 45.805 ;
        RECT 429.475 45.635 429.645 45.805 ;
        RECT 429.935 45.635 430.105 45.805 ;
        RECT 430.395 45.635 430.565 45.805 ;
        RECT 430.855 45.635 431.025 45.805 ;
        RECT 431.315 45.635 431.485 45.805 ;
        RECT 431.775 45.635 431.945 45.805 ;
        RECT 432.235 45.635 432.405 45.805 ;
        RECT 432.695 45.635 432.865 45.805 ;
        RECT 433.155 45.635 433.325 45.805 ;
        RECT 433.615 45.635 433.785 45.805 ;
        RECT 434.075 45.635 434.245 45.805 ;
        RECT 434.535 45.635 434.705 45.805 ;
        RECT 434.995 45.635 435.165 45.805 ;
        RECT 435.455 45.635 435.625 45.805 ;
        RECT 435.915 45.635 436.085 45.805 ;
        RECT 436.375 45.635 436.545 45.805 ;
        RECT 436.835 45.635 437.005 45.805 ;
        RECT 437.295 45.635 437.465 45.805 ;
        RECT 437.755 45.635 437.925 45.805 ;
        RECT 438.215 45.635 438.385 45.805 ;
        RECT 438.675 45.635 438.845 45.805 ;
        RECT 439.135 45.635 439.305 45.805 ;
        RECT 439.595 45.635 439.765 45.805 ;
        RECT 440.055 45.635 440.225 45.805 ;
        RECT 440.515 45.635 440.685 45.805 ;
        RECT 440.975 45.635 441.145 45.805 ;
        RECT 441.435 45.635 441.605 45.805 ;
        RECT 441.895 45.635 442.065 45.805 ;
        RECT 442.355 45.635 442.525 45.805 ;
        RECT 442.815 45.635 442.985 45.805 ;
        RECT 443.275 45.635 443.445 45.805 ;
        RECT 443.735 45.635 443.905 45.805 ;
        RECT 444.195 45.635 444.365 45.805 ;
        RECT 444.655 45.635 444.825 45.805 ;
        RECT 445.115 45.635 445.285 45.805 ;
        RECT 445.575 45.635 445.745 45.805 ;
        RECT 446.035 45.635 446.205 45.805 ;
        RECT 446.495 45.635 446.665 45.805 ;
        RECT 446.955 45.635 447.125 45.805 ;
        RECT 447.415 45.635 447.585 45.805 ;
        RECT 447.875 45.635 448.045 45.805 ;
        RECT 448.335 45.635 448.505 45.805 ;
        RECT 448.795 45.635 448.965 45.805 ;
        RECT 449.255 45.635 449.425 45.805 ;
        RECT 449.715 45.635 449.885 45.805 ;
        RECT 450.175 45.635 450.345 45.805 ;
        RECT 450.635 45.635 450.805 45.805 ;
        RECT 451.095 45.635 451.265 45.805 ;
        RECT 451.555 45.635 451.725 45.805 ;
        RECT 452.015 45.635 452.185 45.805 ;
        RECT 452.475 45.635 452.645 45.805 ;
        RECT 452.935 45.635 453.105 45.805 ;
        RECT 453.395 45.635 453.565 45.805 ;
        RECT 453.855 45.635 454.025 45.805 ;
        RECT 454.315 45.635 454.485 45.805 ;
        RECT 454.775 45.635 454.945 45.805 ;
        RECT 455.235 45.635 455.405 45.805 ;
        RECT 455.695 45.635 455.865 45.805 ;
        RECT 456.155 45.635 456.325 45.805 ;
        RECT 456.615 45.635 456.785 45.805 ;
        RECT 457.075 45.635 457.245 45.805 ;
        RECT 457.535 45.635 457.705 45.805 ;
        RECT 457.995 45.635 458.165 45.805 ;
        RECT 458.455 45.635 458.625 45.805 ;
        RECT 458.915 45.635 459.085 45.805 ;
        RECT 459.375 45.635 459.545 45.805 ;
        RECT 459.835 45.635 460.005 45.805 ;
        RECT 460.295 45.635 460.465 45.805 ;
        RECT 460.755 45.635 460.925 45.805 ;
        RECT 461.215 45.635 461.385 45.805 ;
        RECT 461.675 45.635 461.845 45.805 ;
        RECT 462.135 45.635 462.305 45.805 ;
        RECT 462.595 45.635 462.765 45.805 ;
        RECT 463.055 45.635 463.225 45.805 ;
        RECT 463.515 45.635 463.685 45.805 ;
        RECT 463.975 45.635 464.145 45.805 ;
        RECT 464.435 45.635 464.605 45.805 ;
        RECT 464.895 45.635 465.065 45.805 ;
        RECT 465.355 45.635 465.525 45.805 ;
        RECT 465.815 45.635 465.985 45.805 ;
        RECT 466.275 45.635 466.445 45.805 ;
        RECT 466.735 45.635 466.905 45.805 ;
        RECT 467.195 45.635 467.365 45.805 ;
        RECT 467.655 45.635 467.825 45.805 ;
        RECT 468.115 45.635 468.285 45.805 ;
        RECT 468.575 45.635 468.745 45.805 ;
        RECT 469.035 45.635 469.205 45.805 ;
        RECT 469.495 45.635 469.665 45.805 ;
        RECT 469.955 45.635 470.125 45.805 ;
        RECT 470.415 45.635 470.585 45.805 ;
        RECT 470.875 45.635 471.045 45.805 ;
        RECT 471.335 45.635 471.505 45.805 ;
        RECT 471.795 45.635 471.965 45.805 ;
        RECT 472.255 45.635 472.425 45.805 ;
        RECT 472.715 45.635 472.885 45.805 ;
        RECT 473.175 45.635 473.345 45.805 ;
        RECT 473.635 45.635 473.805 45.805 ;
        RECT 474.095 45.635 474.265 45.805 ;
        RECT 474.555 45.635 474.725 45.805 ;
        RECT 475.015 45.635 475.185 45.805 ;
        RECT 475.475 45.635 475.645 45.805 ;
        RECT 475.935 45.635 476.105 45.805 ;
        RECT 476.395 45.635 476.565 45.805 ;
        RECT 476.855 45.635 477.025 45.805 ;
        RECT 477.315 45.635 477.485 45.805 ;
        RECT 477.775 45.635 477.945 45.805 ;
        RECT 478.235 45.635 478.405 45.805 ;
        RECT 478.695 45.635 478.865 45.805 ;
        RECT 479.155 45.635 479.325 45.805 ;
        RECT 479.615 45.635 479.785 45.805 ;
        RECT 480.075 45.635 480.245 45.805 ;
        RECT 480.535 45.635 480.705 45.805 ;
        RECT 480.995 45.635 481.165 45.805 ;
        RECT 481.455 45.635 481.625 45.805 ;
        RECT 481.915 45.635 482.085 45.805 ;
        RECT 482.375 45.635 482.545 45.805 ;
        RECT 482.835 45.635 483.005 45.805 ;
        RECT 483.295 45.635 483.465 45.805 ;
        RECT 483.755 45.635 483.925 45.805 ;
        RECT 484.215 45.635 484.385 45.805 ;
        RECT 484.675 45.635 484.845 45.805 ;
        RECT 485.135 45.635 485.305 45.805 ;
        RECT 485.595 45.635 485.765 45.805 ;
        RECT 486.055 45.635 486.225 45.805 ;
        RECT 486.515 45.635 486.685 45.805 ;
        RECT 486.975 45.635 487.145 45.805 ;
        RECT 487.435 45.635 487.605 45.805 ;
        RECT 487.895 45.635 488.065 45.805 ;
        RECT 488.355 45.635 488.525 45.805 ;
        RECT 488.815 45.635 488.985 45.805 ;
        RECT 489.275 45.635 489.445 45.805 ;
        RECT 489.735 45.635 489.905 45.805 ;
        RECT 490.195 45.635 490.365 45.805 ;
        RECT 490.655 45.635 490.825 45.805 ;
        RECT 491.115 45.635 491.285 45.805 ;
        RECT 491.575 45.635 491.745 45.805 ;
        RECT 492.035 45.635 492.205 45.805 ;
        RECT 492.495 45.635 492.665 45.805 ;
        RECT 492.955 45.635 493.125 45.805 ;
        RECT 493.415 45.635 493.585 45.805 ;
        RECT 493.875 45.635 494.045 45.805 ;
        RECT 494.335 45.635 494.505 45.805 ;
        RECT 494.795 45.635 494.965 45.805 ;
        RECT 495.255 45.635 495.425 45.805 ;
        RECT 495.715 45.635 495.885 45.805 ;
        RECT 496.175 45.635 496.345 45.805 ;
        RECT 496.635 45.635 496.805 45.805 ;
        RECT 497.095 45.635 497.265 45.805 ;
        RECT 497.555 45.635 497.725 45.805 ;
        RECT 498.015 45.635 498.185 45.805 ;
        RECT 498.475 45.635 498.645 45.805 ;
        RECT 498.935 45.635 499.105 45.805 ;
        RECT 499.395 45.635 499.565 45.805 ;
        RECT 499.855 45.635 500.025 45.805 ;
        RECT 500.315 45.635 500.485 45.805 ;
        RECT 500.775 45.635 500.945 45.805 ;
        RECT 501.235 45.635 501.405 45.805 ;
        RECT 501.695 45.635 501.865 45.805 ;
        RECT 502.155 45.635 502.325 45.805 ;
        RECT 502.615 45.635 502.785 45.805 ;
        RECT 503.075 45.635 503.245 45.805 ;
        RECT 503.535 45.635 503.705 45.805 ;
        RECT 503.995 45.635 504.165 45.805 ;
        RECT 504.455 45.635 504.625 45.805 ;
        RECT 504.915 45.635 505.085 45.805 ;
        RECT 505.375 45.635 505.545 45.805 ;
        RECT 505.835 45.635 506.005 45.805 ;
        RECT 506.295 45.635 506.465 45.805 ;
        RECT 506.755 45.635 506.925 45.805 ;
        RECT 507.215 45.635 507.385 45.805 ;
        RECT 507.675 45.635 507.845 45.805 ;
        RECT 508.135 45.635 508.305 45.805 ;
        RECT 508.595 45.635 508.765 45.805 ;
        RECT 509.055 45.635 509.225 45.805 ;
        RECT 509.515 45.635 509.685 45.805 ;
        RECT 509.975 45.635 510.145 45.805 ;
        RECT 510.435 45.635 510.605 45.805 ;
        RECT 510.895 45.635 511.065 45.805 ;
        RECT 511.355 45.635 511.525 45.805 ;
        RECT 511.815 45.635 511.985 45.805 ;
        RECT 512.275 45.635 512.445 45.805 ;
        RECT 512.735 45.635 512.905 45.805 ;
        RECT 513.195 45.635 513.365 45.805 ;
        RECT 513.655 45.635 513.825 45.805 ;
        RECT 514.115 45.635 514.285 45.805 ;
        RECT 514.575 45.635 514.745 45.805 ;
        RECT 515.035 45.635 515.205 45.805 ;
        RECT 515.495 45.635 515.665 45.805 ;
        RECT 515.955 45.635 516.125 45.805 ;
        RECT 516.415 45.635 516.585 45.805 ;
        RECT 516.875 45.635 517.045 45.805 ;
        RECT 517.335 45.635 517.505 45.805 ;
        RECT 517.795 45.635 517.965 45.805 ;
        RECT 518.255 45.635 518.425 45.805 ;
        RECT 518.715 45.635 518.885 45.805 ;
        RECT 519.175 45.635 519.345 45.805 ;
        RECT 519.635 45.635 519.805 45.805 ;
        RECT 520.095 45.635 520.265 45.805 ;
        RECT 520.555 45.635 520.725 45.805 ;
        RECT 521.015 45.635 521.185 45.805 ;
        RECT 521.475 45.635 521.645 45.805 ;
        RECT 521.935 45.635 522.105 45.805 ;
        RECT 522.395 45.635 522.565 45.805 ;
        RECT 522.855 45.635 523.025 45.805 ;
        RECT 523.315 45.635 523.485 45.805 ;
        RECT 523.775 45.635 523.945 45.805 ;
        RECT 524.235 45.635 524.405 45.805 ;
        RECT 524.695 45.635 524.865 45.805 ;
        RECT 525.155 45.635 525.325 45.805 ;
        RECT 525.615 45.635 525.785 45.805 ;
        RECT 526.075 45.635 526.245 45.805 ;
        RECT 526.535 45.635 526.705 45.805 ;
        RECT 526.995 45.635 527.165 45.805 ;
        RECT 527.455 45.635 527.625 45.805 ;
        RECT 527.915 45.635 528.085 45.805 ;
        RECT 528.375 45.635 528.545 45.805 ;
        RECT 528.835 45.635 529.005 45.805 ;
        RECT 529.295 45.635 529.465 45.805 ;
        RECT 529.755 45.635 529.925 45.805 ;
        RECT 530.215 45.635 530.385 45.805 ;
        RECT 530.675 45.635 530.845 45.805 ;
        RECT 531.135 45.635 531.305 45.805 ;
        RECT 531.595 45.635 531.765 45.805 ;
        RECT 532.055 45.635 532.225 45.805 ;
        RECT 532.515 45.635 532.685 45.805 ;
        RECT 532.975 45.635 533.145 45.805 ;
        RECT 533.435 45.635 533.605 45.805 ;
        RECT 533.895 45.635 534.065 45.805 ;
        RECT 534.355 45.635 534.525 45.805 ;
        RECT 534.815 45.635 534.985 45.805 ;
        RECT 535.275 45.635 535.445 45.805 ;
        RECT 535.735 45.635 535.905 45.805 ;
        RECT 536.195 45.635 536.365 45.805 ;
        RECT 536.655 45.635 536.825 45.805 ;
        RECT 537.115 45.635 537.285 45.805 ;
        RECT 537.575 45.635 537.745 45.805 ;
        RECT 538.035 45.635 538.205 45.805 ;
        RECT 538.495 45.635 538.665 45.805 ;
        RECT 538.955 45.635 539.125 45.805 ;
        RECT 539.415 45.635 539.585 45.805 ;
        RECT 539.875 45.635 540.045 45.805 ;
        RECT 540.335 45.635 540.505 45.805 ;
        RECT 540.795 45.635 540.965 45.805 ;
        RECT 541.255 45.635 541.425 45.805 ;
        RECT 541.715 45.635 541.885 45.805 ;
        RECT 542.175 45.635 542.345 45.805 ;
        RECT 542.635 45.635 542.805 45.805 ;
        RECT 543.095 45.635 543.265 45.805 ;
        RECT 543.555 45.635 543.725 45.805 ;
        RECT 544.015 45.635 544.185 45.805 ;
        RECT 544.475 45.635 544.645 45.805 ;
        RECT 544.935 45.635 545.105 45.805 ;
        RECT 545.395 45.635 545.565 45.805 ;
        RECT 545.855 45.635 546.025 45.805 ;
        RECT 546.315 45.635 546.485 45.805 ;
        RECT 546.775 45.635 546.945 45.805 ;
        RECT 547.235 45.635 547.405 45.805 ;
        RECT 547.695 45.635 547.865 45.805 ;
        RECT 548.155 45.635 548.325 45.805 ;
        RECT 548.615 45.635 548.785 45.805 ;
        RECT 549.075 45.635 549.245 45.805 ;
        RECT 549.535 45.635 549.705 45.805 ;
        RECT 549.995 45.635 550.165 45.805 ;
        RECT 550.455 45.635 550.625 45.805 ;
        RECT 550.915 45.635 551.085 45.805 ;
        RECT 551.375 45.635 551.545 45.805 ;
        RECT 551.835 45.635 552.005 45.805 ;
        RECT 552.295 45.635 552.465 45.805 ;
        RECT 552.755 45.635 552.925 45.805 ;
        RECT 553.215 45.635 553.385 45.805 ;
        RECT 553.675 45.635 553.845 45.805 ;
        RECT 554.135 45.635 554.305 45.805 ;
        RECT 554.595 45.635 554.765 45.805 ;
        RECT 555.055 45.635 555.225 45.805 ;
        RECT 555.515 45.635 555.685 45.805 ;
        RECT 555.975 45.635 556.145 45.805 ;
        RECT 556.435 45.635 556.605 45.805 ;
        RECT 556.895 45.635 557.065 45.805 ;
        RECT 557.355 45.635 557.525 45.805 ;
        RECT 557.815 45.635 557.985 45.805 ;
        RECT 558.275 45.635 558.445 45.805 ;
        RECT 558.735 45.635 558.905 45.805 ;
        RECT 559.195 45.635 559.365 45.805 ;
        RECT 559.655 45.635 559.825 45.805 ;
        RECT 560.115 45.635 560.285 45.805 ;
        RECT 560.575 45.635 560.745 45.805 ;
        RECT 561.035 45.635 561.205 45.805 ;
        RECT 561.495 45.635 561.665 45.805 ;
        RECT 561.955 45.635 562.125 45.805 ;
        RECT 562.415 45.635 562.585 45.805 ;
        RECT 562.875 45.635 563.045 45.805 ;
        RECT 563.335 45.635 563.505 45.805 ;
        RECT 563.795 45.635 563.965 45.805 ;
        RECT 564.255 45.635 564.425 45.805 ;
        RECT 564.715 45.635 564.885 45.805 ;
        RECT 565.175 45.635 565.345 45.805 ;
        RECT 565.635 45.635 565.805 45.805 ;
        RECT 566.095 45.635 566.265 45.805 ;
        RECT 566.555 45.635 566.725 45.805 ;
        RECT 567.015 45.635 567.185 45.805 ;
        RECT 567.475 45.635 567.645 45.805 ;
        RECT 567.935 45.635 568.105 45.805 ;
        RECT 568.395 45.635 568.565 45.805 ;
        RECT 568.855 45.635 569.025 45.805 ;
        RECT 569.315 45.635 569.485 45.805 ;
        RECT 569.775 45.635 569.945 45.805 ;
        RECT 570.235 45.635 570.405 45.805 ;
        RECT 570.695 45.635 570.865 45.805 ;
        RECT 571.155 45.635 571.325 45.805 ;
        RECT 571.615 45.635 571.785 45.805 ;
        RECT 572.075 45.635 572.245 45.805 ;
        RECT 572.535 45.635 572.705 45.805 ;
        RECT 572.995 45.635 573.165 45.805 ;
        RECT 573.455 45.635 573.625 45.805 ;
        RECT 573.915 45.635 574.085 45.805 ;
        RECT 574.375 45.635 574.545 45.805 ;
        RECT 574.835 45.635 575.005 45.805 ;
        RECT 575.295 45.635 575.465 45.805 ;
        RECT 575.755 45.635 575.925 45.805 ;
        RECT 576.215 45.635 576.385 45.805 ;
        RECT 576.675 45.635 576.845 45.805 ;
        RECT 577.135 45.635 577.305 45.805 ;
        RECT 577.595 45.635 577.765 45.805 ;
        RECT 578.055 45.635 578.225 45.805 ;
        RECT 578.515 45.635 578.685 45.805 ;
        RECT 578.975 45.635 579.145 45.805 ;
        RECT 579.435 45.635 579.605 45.805 ;
        RECT 579.895 45.635 580.065 45.805 ;
        RECT 580.355 45.635 580.525 45.805 ;
        RECT 580.815 45.635 580.985 45.805 ;
        RECT 581.275 45.635 581.445 45.805 ;
        RECT 581.735 45.635 581.905 45.805 ;
        RECT 582.195 45.635 582.365 45.805 ;
        RECT 582.655 45.635 582.825 45.805 ;
        RECT 583.115 45.635 583.285 45.805 ;
        RECT 583.575 45.635 583.745 45.805 ;
        RECT 584.035 45.635 584.205 45.805 ;
        RECT 584.495 45.635 584.665 45.805 ;
        RECT 584.955 45.635 585.125 45.805 ;
        RECT 585.415 45.635 585.585 45.805 ;
        RECT 585.875 45.635 586.045 45.805 ;
        RECT 586.335 45.635 586.505 45.805 ;
        RECT 586.795 45.635 586.965 45.805 ;
        RECT 587.255 45.635 587.425 45.805 ;
        RECT 587.715 45.635 587.885 45.805 ;
        RECT 588.175 45.635 588.345 45.805 ;
        RECT 588.635 45.635 588.805 45.805 ;
        RECT 589.095 45.635 589.265 45.805 ;
        RECT 589.555 45.635 589.725 45.805 ;
        RECT 590.015 45.635 590.185 45.805 ;
        RECT 590.475 45.635 590.645 45.805 ;
        RECT 590.935 45.635 591.105 45.805 ;
        RECT 591.395 45.635 591.565 45.805 ;
        RECT 591.855 45.635 592.025 45.805 ;
        RECT 592.315 45.635 592.485 45.805 ;
        RECT 592.775 45.635 592.945 45.805 ;
        RECT 593.235 45.635 593.405 45.805 ;
        RECT 593.695 45.635 593.865 45.805 ;
        RECT 594.155 45.635 594.325 45.805 ;
        RECT 594.615 45.635 594.785 45.805 ;
        RECT 595.075 45.635 595.245 45.805 ;
        RECT 595.535 45.635 595.705 45.805 ;
        RECT 595.995 45.635 596.165 45.805 ;
        RECT 596.455 45.635 596.625 45.805 ;
        RECT 596.915 45.635 597.085 45.805 ;
        RECT 597.375 45.635 597.545 45.805 ;
        RECT 597.835 45.635 598.005 45.805 ;
        RECT 598.295 45.635 598.465 45.805 ;
        RECT 598.755 45.635 598.925 45.805 ;
        RECT 599.215 45.635 599.385 45.805 ;
        RECT 599.675 45.635 599.845 45.805 ;
        RECT 600.135 45.635 600.305 45.805 ;
        RECT 600.595 45.635 600.765 45.805 ;
        RECT 601.055 45.635 601.225 45.805 ;
        RECT 601.515 45.635 601.685 45.805 ;
        RECT 601.975 45.635 602.145 45.805 ;
        RECT 602.435 45.635 602.605 45.805 ;
        RECT 602.895 45.635 603.065 45.805 ;
        RECT 603.355 45.635 603.525 45.805 ;
        RECT 603.815 45.635 603.985 45.805 ;
        RECT 604.275 45.635 604.445 45.805 ;
        RECT 604.735 45.635 604.905 45.805 ;
        RECT 605.195 45.635 605.365 45.805 ;
        RECT 605.655 45.635 605.825 45.805 ;
        RECT 606.115 45.635 606.285 45.805 ;
        RECT 606.575 45.635 606.745 45.805 ;
        RECT 607.035 45.635 607.205 45.805 ;
        RECT 607.495 45.635 607.665 45.805 ;
        RECT 607.955 45.635 608.125 45.805 ;
        RECT 608.415 45.635 608.585 45.805 ;
        RECT 608.875 45.635 609.045 45.805 ;
        RECT 609.335 45.635 609.505 45.805 ;
        RECT 609.795 45.635 609.965 45.805 ;
        RECT 610.255 45.635 610.425 45.805 ;
        RECT 610.715 45.635 610.885 45.805 ;
        RECT 611.175 45.635 611.345 45.805 ;
        RECT 611.635 45.635 611.805 45.805 ;
        RECT 612.095 45.635 612.265 45.805 ;
        RECT 612.555 45.635 612.725 45.805 ;
        RECT 613.015 45.635 613.185 45.805 ;
        RECT 613.475 45.635 613.645 45.805 ;
        RECT 613.935 45.635 614.105 45.805 ;
        RECT 614.395 45.635 614.565 45.805 ;
        RECT 614.855 45.635 615.025 45.805 ;
        RECT 615.315 45.635 615.485 45.805 ;
        RECT 615.775 45.635 615.945 45.805 ;
        RECT 616.235 45.635 616.405 45.805 ;
        RECT 616.695 45.635 616.865 45.805 ;
        RECT 617.155 45.635 617.325 45.805 ;
        RECT 617.615 45.635 617.785 45.805 ;
        RECT 618.075 45.635 618.245 45.805 ;
        RECT 618.535 45.635 618.705 45.805 ;
        RECT 618.995 45.635 619.165 45.805 ;
        RECT 619.455 45.635 619.625 45.805 ;
        RECT 619.915 45.635 620.085 45.805 ;
        RECT 620.375 45.635 620.545 45.805 ;
        RECT 620.835 45.635 621.005 45.805 ;
        RECT 621.295 45.635 621.465 45.805 ;
        RECT 621.755 45.635 621.925 45.805 ;
        RECT 622.215 45.635 622.385 45.805 ;
        RECT 622.675 45.635 622.845 45.805 ;
        RECT 623.135 45.635 623.305 45.805 ;
        RECT 623.595 45.635 623.765 45.805 ;
        RECT 624.055 45.635 624.225 45.805 ;
        RECT 624.515 45.635 624.685 45.805 ;
        RECT 624.975 45.635 625.145 45.805 ;
        RECT 625.435 45.635 625.605 45.805 ;
        RECT 625.895 45.635 626.065 45.805 ;
        RECT 626.355 45.635 626.525 45.805 ;
        RECT 626.815 45.635 626.985 45.805 ;
        RECT 627.275 45.635 627.445 45.805 ;
        RECT 627.735 45.635 627.905 45.805 ;
        RECT 628.195 45.635 628.365 45.805 ;
        RECT 628.655 45.635 628.825 45.805 ;
        RECT 629.115 45.635 629.285 45.805 ;
        RECT 629.575 45.635 629.745 45.805 ;
        RECT 630.035 45.635 630.205 45.805 ;
        RECT 630.495 45.635 630.665 45.805 ;
        RECT 630.955 45.635 631.125 45.805 ;
        RECT 78.495 44.785 78.665 44.955 ;
        RECT 81.255 44.785 81.425 44.955 ;
        RECT 79.415 44.445 79.585 44.615 ;
        RECT 86.735 44.445 86.905 44.615 ;
        RECT 87.235 44.445 87.405 44.615 ;
        RECT 95.515 44.785 95.685 44.955 ;
        RECT 94.135 44.445 94.305 44.615 ;
        RECT 101.495 45.125 101.665 45.295 ;
        RECT 100.575 44.445 100.745 44.615 ;
        RECT 106.095 44.785 106.265 44.955 ;
        RECT 109.775 44.785 109.945 44.955 ;
        RECT 107.935 44.105 108.105 44.275 ;
        RECT 115.295 44.445 115.465 44.615 ;
        RECT 107.475 43.425 107.645 43.595 ;
        RECT 118.515 45.125 118.685 45.295 ;
        RECT 117.135 44.105 117.305 44.275 ;
        RECT 123.115 44.445 123.285 44.615 ;
        RECT 128.635 44.785 128.805 44.955 ;
        RECT 116.675 43.425 116.845 43.595 ;
        RECT 123.575 43.425 123.745 43.595 ;
        RECT 129.370 44.105 129.540 44.275 ;
        RECT 130.475 44.105 130.645 44.275 ;
        RECT 136.915 44.445 137.085 44.615 ;
        RECT 130.015 43.765 130.185 43.935 ;
        RECT 131.855 43.425 132.025 43.595 ;
        RECT 137.835 43.765 138.005 43.935 ;
        RECT 143.355 44.445 143.525 44.615 ;
        RECT 150.255 45.125 150.425 45.295 ;
        RECT 144.275 43.425 144.445 43.595 ;
        RECT 148.875 44.445 149.045 44.615 ;
        RECT 151.175 44.445 151.345 44.615 ;
        RECT 157.155 44.445 157.325 44.615 ;
        RECT 157.620 43.765 157.790 43.935 ;
        RECT 158.080 44.785 158.250 44.955 ;
        RECT 158.535 44.105 158.705 44.275 ;
        RECT 159.480 44.785 159.650 44.955 ;
        RECT 161.320 44.785 161.490 44.955 ;
        RECT 159.940 43.765 160.110 43.935 ;
        RECT 161.320 43.765 161.490 43.935 ;
        RECT 164.055 43.425 164.225 43.595 ;
        RECT 174.635 44.445 174.805 44.615 ;
        RECT 174.175 44.105 174.345 44.275 ;
        RECT 176.020 44.105 176.190 44.275 ;
        RECT 177.395 44.445 177.565 44.615 ;
        RECT 178.315 44.445 178.485 44.615 ;
        RECT 178.800 44.105 178.970 44.275 ;
        RECT 186.135 44.445 186.305 44.615 ;
        RECT 179.235 43.765 179.405 43.935 ;
        RECT 186.600 43.765 186.770 43.935 ;
        RECT 187.060 44.785 187.230 44.955 ;
        RECT 187.515 44.445 187.685 44.615 ;
        RECT 188.460 44.785 188.630 44.955 ;
        RECT 190.300 44.785 190.470 44.955 ;
        RECT 188.920 43.765 189.090 43.935 ;
        RECT 190.300 43.765 190.470 43.935 ;
        RECT 193.035 45.125 193.205 45.295 ;
        RECT 206.375 44.445 206.545 44.615 ;
        RECT 204.075 44.105 204.245 44.275 ;
        RECT 208.215 44.445 208.385 44.615 ;
        RECT 208.675 44.105 208.845 44.275 ;
        RECT 214.655 44.445 214.825 44.615 ;
        RECT 215.115 44.445 215.285 44.615 ;
        RECT 215.780 44.445 215.950 44.615 ;
        RECT 217.875 44.445 218.045 44.615 ;
        RECT 222.935 45.125 223.105 45.295 ;
        RECT 222.045 44.445 222.215 44.615 ;
        RECT 228.455 44.445 228.625 44.615 ;
        RECT 229.835 44.445 230.005 44.615 ;
        RECT 228.915 43.765 229.085 43.935 ;
        RECT 230.755 44.105 230.925 44.275 ;
        RECT 237.195 45.125 237.365 45.295 ;
        RECT 236.275 44.445 236.445 44.615 ;
        RECT 242.715 44.445 242.885 44.615 ;
        RECT 243.635 44.445 243.805 44.615 ;
        RECT 249.615 44.785 249.785 44.955 ;
        RECT 245.475 44.105 245.645 44.275 ;
        RECT 250.535 44.445 250.705 44.615 ;
        RECT 256.975 44.785 257.145 44.955 ;
        RECT 258.355 45.125 258.525 45.295 ;
        RECT 250.995 43.425 251.165 43.595 ;
        RECT 257.895 44.445 258.065 44.615 ;
        RECT 263.875 44.445 264.045 44.615 ;
        RECT 264.795 43.425 264.965 43.595 ;
        RECT 271.235 44.445 271.405 44.615 ;
        RECT 277.215 45.125 277.385 45.295 ;
        RECT 272.155 43.765 272.325 43.935 ;
        RECT 278.135 44.445 278.305 44.615 ;
        RECT 279.055 44.445 279.225 44.615 ;
        RECT 286.875 44.445 287.045 44.615 ;
        RECT 288.485 44.445 288.655 44.615 ;
        RECT 294.235 45.125 294.405 45.295 ;
        RECT 287.795 44.105 287.965 44.275 ;
        RECT 293.315 44.445 293.485 44.615 ;
        RECT 301.135 44.445 301.305 44.615 ;
        RECT 302.515 44.445 302.685 44.615 ;
        RECT 302.055 44.105 302.225 44.275 ;
        RECT 307.575 44.445 307.745 44.615 ;
        RECT 308.495 43.425 308.665 43.595 ;
        RECT 315.395 44.445 315.565 44.615 ;
        RECT 316.775 44.445 316.945 44.615 ;
        RECT 316.315 44.105 316.485 44.275 ;
        RECT 321.835 44.445 322.005 44.615 ;
        RECT 328.735 45.125 328.905 45.295 ;
        RECT 322.755 43.425 322.925 43.595 ;
        RECT 329.655 44.445 329.825 44.615 ;
        RECT 330.575 44.445 330.745 44.615 ;
        RECT 336.095 44.445 336.265 44.615 ;
        RECT 337.015 43.425 337.185 43.595 ;
        RECT 345.295 44.445 345.465 44.615 ;
        RECT 345.755 44.105 345.925 44.275 ;
        RECT 348.055 44.445 348.225 44.615 ;
        RECT 348.975 44.445 349.145 44.615 ;
        RECT 350.815 44.445 350.985 44.615 ;
        RECT 351.735 44.445 351.905 44.615 ;
        RECT 357.255 45.125 357.425 45.295 ;
        RECT 358.175 44.445 358.345 44.615 ;
        RECT 359.095 44.445 359.265 44.615 ;
        RECT 364.615 44.445 364.785 44.615 ;
        RECT 371.515 45.125 371.685 45.295 ;
        RECT 365.075 43.765 365.245 43.935 ;
        RECT 372.435 44.445 372.605 44.615 ;
        RECT 373.355 44.445 373.525 44.615 ;
        RECT 379.795 43.425 379.965 43.595 ;
        RECT 386.235 44.445 386.405 44.615 ;
        RECT 391.295 43.765 391.465 43.935 ;
        RECT 502.615 43.425 502.785 43.595 ;
        RECT 586.795 43.425 586.965 43.595 ;
        RECT 42.615 42.915 42.785 43.085 ;
        RECT 43.075 42.915 43.245 43.085 ;
        RECT 43.535 42.915 43.705 43.085 ;
        RECT 43.995 42.915 44.165 43.085 ;
        RECT 44.455 42.915 44.625 43.085 ;
        RECT 44.915 42.915 45.085 43.085 ;
        RECT 45.375 42.915 45.545 43.085 ;
        RECT 45.835 42.915 46.005 43.085 ;
        RECT 46.295 42.915 46.465 43.085 ;
        RECT 46.755 42.915 46.925 43.085 ;
        RECT 47.215 42.915 47.385 43.085 ;
        RECT 47.675 42.915 47.845 43.085 ;
        RECT 48.135 42.915 48.305 43.085 ;
        RECT 48.595 42.915 48.765 43.085 ;
        RECT 49.055 42.915 49.225 43.085 ;
        RECT 49.515 42.915 49.685 43.085 ;
        RECT 49.975 42.915 50.145 43.085 ;
        RECT 50.435 42.915 50.605 43.085 ;
        RECT 50.895 42.915 51.065 43.085 ;
        RECT 51.355 42.915 51.525 43.085 ;
        RECT 51.815 42.915 51.985 43.085 ;
        RECT 52.275 42.915 52.445 43.085 ;
        RECT 52.735 42.915 52.905 43.085 ;
        RECT 53.195 42.915 53.365 43.085 ;
        RECT 53.655 42.915 53.825 43.085 ;
        RECT 54.115 42.915 54.285 43.085 ;
        RECT 54.575 42.915 54.745 43.085 ;
        RECT 55.035 42.915 55.205 43.085 ;
        RECT 55.495 42.915 55.665 43.085 ;
        RECT 55.955 42.915 56.125 43.085 ;
        RECT 56.415 42.915 56.585 43.085 ;
        RECT 56.875 42.915 57.045 43.085 ;
        RECT 57.335 42.915 57.505 43.085 ;
        RECT 57.795 42.915 57.965 43.085 ;
        RECT 58.255 42.915 58.425 43.085 ;
        RECT 58.715 42.915 58.885 43.085 ;
        RECT 59.175 42.915 59.345 43.085 ;
        RECT 59.635 42.915 59.805 43.085 ;
        RECT 60.095 42.915 60.265 43.085 ;
        RECT 60.555 42.915 60.725 43.085 ;
        RECT 61.015 42.915 61.185 43.085 ;
        RECT 61.475 42.915 61.645 43.085 ;
        RECT 61.935 42.915 62.105 43.085 ;
        RECT 62.395 42.915 62.565 43.085 ;
        RECT 62.855 42.915 63.025 43.085 ;
        RECT 63.315 42.915 63.485 43.085 ;
        RECT 63.775 42.915 63.945 43.085 ;
        RECT 64.235 42.915 64.405 43.085 ;
        RECT 64.695 42.915 64.865 43.085 ;
        RECT 65.155 42.915 65.325 43.085 ;
        RECT 65.615 42.915 65.785 43.085 ;
        RECT 66.075 42.915 66.245 43.085 ;
        RECT 66.535 42.915 66.705 43.085 ;
        RECT 66.995 42.915 67.165 43.085 ;
        RECT 67.455 42.915 67.625 43.085 ;
        RECT 67.915 42.915 68.085 43.085 ;
        RECT 68.375 42.915 68.545 43.085 ;
        RECT 68.835 42.915 69.005 43.085 ;
        RECT 69.295 42.915 69.465 43.085 ;
        RECT 69.755 42.915 69.925 43.085 ;
        RECT 70.215 42.915 70.385 43.085 ;
        RECT 70.675 42.915 70.845 43.085 ;
        RECT 71.135 42.915 71.305 43.085 ;
        RECT 71.595 42.915 71.765 43.085 ;
        RECT 72.055 42.915 72.225 43.085 ;
        RECT 72.515 42.915 72.685 43.085 ;
        RECT 72.975 42.915 73.145 43.085 ;
        RECT 73.435 42.915 73.605 43.085 ;
        RECT 73.895 42.915 74.065 43.085 ;
        RECT 74.355 42.915 74.525 43.085 ;
        RECT 74.815 42.915 74.985 43.085 ;
        RECT 75.275 42.915 75.445 43.085 ;
        RECT 75.735 42.915 75.905 43.085 ;
        RECT 76.195 42.915 76.365 43.085 ;
        RECT 76.655 42.915 76.825 43.085 ;
        RECT 77.115 42.915 77.285 43.085 ;
        RECT 77.575 42.915 77.745 43.085 ;
        RECT 78.035 42.915 78.205 43.085 ;
        RECT 78.495 42.915 78.665 43.085 ;
        RECT 78.955 42.915 79.125 43.085 ;
        RECT 79.415 42.915 79.585 43.085 ;
        RECT 79.875 42.915 80.045 43.085 ;
        RECT 80.335 42.915 80.505 43.085 ;
        RECT 80.795 42.915 80.965 43.085 ;
        RECT 81.255 42.915 81.425 43.085 ;
        RECT 81.715 42.915 81.885 43.085 ;
        RECT 82.175 42.915 82.345 43.085 ;
        RECT 82.635 42.915 82.805 43.085 ;
        RECT 83.095 42.915 83.265 43.085 ;
        RECT 83.555 42.915 83.725 43.085 ;
        RECT 84.015 42.915 84.185 43.085 ;
        RECT 84.475 42.915 84.645 43.085 ;
        RECT 84.935 42.915 85.105 43.085 ;
        RECT 85.395 42.915 85.565 43.085 ;
        RECT 85.855 42.915 86.025 43.085 ;
        RECT 86.315 42.915 86.485 43.085 ;
        RECT 86.775 42.915 86.945 43.085 ;
        RECT 87.235 42.915 87.405 43.085 ;
        RECT 87.695 42.915 87.865 43.085 ;
        RECT 88.155 42.915 88.325 43.085 ;
        RECT 88.615 42.915 88.785 43.085 ;
        RECT 89.075 42.915 89.245 43.085 ;
        RECT 89.535 42.915 89.705 43.085 ;
        RECT 89.995 42.915 90.165 43.085 ;
        RECT 90.455 42.915 90.625 43.085 ;
        RECT 90.915 42.915 91.085 43.085 ;
        RECT 91.375 42.915 91.545 43.085 ;
        RECT 91.835 42.915 92.005 43.085 ;
        RECT 92.295 42.915 92.465 43.085 ;
        RECT 92.755 42.915 92.925 43.085 ;
        RECT 93.215 42.915 93.385 43.085 ;
        RECT 93.675 42.915 93.845 43.085 ;
        RECT 94.135 42.915 94.305 43.085 ;
        RECT 94.595 42.915 94.765 43.085 ;
        RECT 95.055 42.915 95.225 43.085 ;
        RECT 95.515 42.915 95.685 43.085 ;
        RECT 95.975 42.915 96.145 43.085 ;
        RECT 96.435 42.915 96.605 43.085 ;
        RECT 96.895 42.915 97.065 43.085 ;
        RECT 97.355 42.915 97.525 43.085 ;
        RECT 97.815 42.915 97.985 43.085 ;
        RECT 98.275 42.915 98.445 43.085 ;
        RECT 98.735 42.915 98.905 43.085 ;
        RECT 99.195 42.915 99.365 43.085 ;
        RECT 99.655 42.915 99.825 43.085 ;
        RECT 100.115 42.915 100.285 43.085 ;
        RECT 100.575 42.915 100.745 43.085 ;
        RECT 101.035 42.915 101.205 43.085 ;
        RECT 101.495 42.915 101.665 43.085 ;
        RECT 101.955 42.915 102.125 43.085 ;
        RECT 102.415 42.915 102.585 43.085 ;
        RECT 102.875 42.915 103.045 43.085 ;
        RECT 103.335 42.915 103.505 43.085 ;
        RECT 103.795 42.915 103.965 43.085 ;
        RECT 104.255 42.915 104.425 43.085 ;
        RECT 104.715 42.915 104.885 43.085 ;
        RECT 105.175 42.915 105.345 43.085 ;
        RECT 105.635 42.915 105.805 43.085 ;
        RECT 106.095 42.915 106.265 43.085 ;
        RECT 106.555 42.915 106.725 43.085 ;
        RECT 107.015 42.915 107.185 43.085 ;
        RECT 107.475 42.915 107.645 43.085 ;
        RECT 107.935 42.915 108.105 43.085 ;
        RECT 108.395 42.915 108.565 43.085 ;
        RECT 108.855 42.915 109.025 43.085 ;
        RECT 109.315 42.915 109.485 43.085 ;
        RECT 109.775 42.915 109.945 43.085 ;
        RECT 110.235 42.915 110.405 43.085 ;
        RECT 110.695 42.915 110.865 43.085 ;
        RECT 111.155 42.915 111.325 43.085 ;
        RECT 111.615 42.915 111.785 43.085 ;
        RECT 112.075 42.915 112.245 43.085 ;
        RECT 112.535 42.915 112.705 43.085 ;
        RECT 112.995 42.915 113.165 43.085 ;
        RECT 113.455 42.915 113.625 43.085 ;
        RECT 113.915 42.915 114.085 43.085 ;
        RECT 114.375 42.915 114.545 43.085 ;
        RECT 114.835 42.915 115.005 43.085 ;
        RECT 115.295 42.915 115.465 43.085 ;
        RECT 115.755 42.915 115.925 43.085 ;
        RECT 116.215 42.915 116.385 43.085 ;
        RECT 116.675 42.915 116.845 43.085 ;
        RECT 117.135 42.915 117.305 43.085 ;
        RECT 117.595 42.915 117.765 43.085 ;
        RECT 118.055 42.915 118.225 43.085 ;
        RECT 118.515 42.915 118.685 43.085 ;
        RECT 118.975 42.915 119.145 43.085 ;
        RECT 119.435 42.915 119.605 43.085 ;
        RECT 119.895 42.915 120.065 43.085 ;
        RECT 120.355 42.915 120.525 43.085 ;
        RECT 120.815 42.915 120.985 43.085 ;
        RECT 121.275 42.915 121.445 43.085 ;
        RECT 121.735 42.915 121.905 43.085 ;
        RECT 122.195 42.915 122.365 43.085 ;
        RECT 122.655 42.915 122.825 43.085 ;
        RECT 123.115 42.915 123.285 43.085 ;
        RECT 123.575 42.915 123.745 43.085 ;
        RECT 124.035 42.915 124.205 43.085 ;
        RECT 124.495 42.915 124.665 43.085 ;
        RECT 124.955 42.915 125.125 43.085 ;
        RECT 125.415 42.915 125.585 43.085 ;
        RECT 125.875 42.915 126.045 43.085 ;
        RECT 126.335 42.915 126.505 43.085 ;
        RECT 126.795 42.915 126.965 43.085 ;
        RECT 127.255 42.915 127.425 43.085 ;
        RECT 127.715 42.915 127.885 43.085 ;
        RECT 128.175 42.915 128.345 43.085 ;
        RECT 128.635 42.915 128.805 43.085 ;
        RECT 129.095 42.915 129.265 43.085 ;
        RECT 129.555 42.915 129.725 43.085 ;
        RECT 130.015 42.915 130.185 43.085 ;
        RECT 130.475 42.915 130.645 43.085 ;
        RECT 130.935 42.915 131.105 43.085 ;
        RECT 131.395 42.915 131.565 43.085 ;
        RECT 131.855 42.915 132.025 43.085 ;
        RECT 132.315 42.915 132.485 43.085 ;
        RECT 132.775 42.915 132.945 43.085 ;
        RECT 133.235 42.915 133.405 43.085 ;
        RECT 133.695 42.915 133.865 43.085 ;
        RECT 134.155 42.915 134.325 43.085 ;
        RECT 134.615 42.915 134.785 43.085 ;
        RECT 135.075 42.915 135.245 43.085 ;
        RECT 135.535 42.915 135.705 43.085 ;
        RECT 135.995 42.915 136.165 43.085 ;
        RECT 136.455 42.915 136.625 43.085 ;
        RECT 136.915 42.915 137.085 43.085 ;
        RECT 137.375 42.915 137.545 43.085 ;
        RECT 137.835 42.915 138.005 43.085 ;
        RECT 138.295 42.915 138.465 43.085 ;
        RECT 138.755 42.915 138.925 43.085 ;
        RECT 139.215 42.915 139.385 43.085 ;
        RECT 139.675 42.915 139.845 43.085 ;
        RECT 140.135 42.915 140.305 43.085 ;
        RECT 140.595 42.915 140.765 43.085 ;
        RECT 141.055 42.915 141.225 43.085 ;
        RECT 141.515 42.915 141.685 43.085 ;
        RECT 141.975 42.915 142.145 43.085 ;
        RECT 142.435 42.915 142.605 43.085 ;
        RECT 142.895 42.915 143.065 43.085 ;
        RECT 143.355 42.915 143.525 43.085 ;
        RECT 143.815 42.915 143.985 43.085 ;
        RECT 144.275 42.915 144.445 43.085 ;
        RECT 144.735 42.915 144.905 43.085 ;
        RECT 145.195 42.915 145.365 43.085 ;
        RECT 145.655 42.915 145.825 43.085 ;
        RECT 146.115 42.915 146.285 43.085 ;
        RECT 146.575 42.915 146.745 43.085 ;
        RECT 147.035 42.915 147.205 43.085 ;
        RECT 147.495 42.915 147.665 43.085 ;
        RECT 147.955 42.915 148.125 43.085 ;
        RECT 148.415 42.915 148.585 43.085 ;
        RECT 148.875 42.915 149.045 43.085 ;
        RECT 149.335 42.915 149.505 43.085 ;
        RECT 149.795 42.915 149.965 43.085 ;
        RECT 150.255 42.915 150.425 43.085 ;
        RECT 150.715 42.915 150.885 43.085 ;
        RECT 151.175 42.915 151.345 43.085 ;
        RECT 151.635 42.915 151.805 43.085 ;
        RECT 152.095 42.915 152.265 43.085 ;
        RECT 152.555 42.915 152.725 43.085 ;
        RECT 153.015 42.915 153.185 43.085 ;
        RECT 153.475 42.915 153.645 43.085 ;
        RECT 153.935 42.915 154.105 43.085 ;
        RECT 154.395 42.915 154.565 43.085 ;
        RECT 154.855 42.915 155.025 43.085 ;
        RECT 155.315 42.915 155.485 43.085 ;
        RECT 155.775 42.915 155.945 43.085 ;
        RECT 156.235 42.915 156.405 43.085 ;
        RECT 156.695 42.915 156.865 43.085 ;
        RECT 157.155 42.915 157.325 43.085 ;
        RECT 157.615 42.915 157.785 43.085 ;
        RECT 158.075 42.915 158.245 43.085 ;
        RECT 158.535 42.915 158.705 43.085 ;
        RECT 158.995 42.915 159.165 43.085 ;
        RECT 159.455 42.915 159.625 43.085 ;
        RECT 159.915 42.915 160.085 43.085 ;
        RECT 160.375 42.915 160.545 43.085 ;
        RECT 160.835 42.915 161.005 43.085 ;
        RECT 161.295 42.915 161.465 43.085 ;
        RECT 161.755 42.915 161.925 43.085 ;
        RECT 162.215 42.915 162.385 43.085 ;
        RECT 162.675 42.915 162.845 43.085 ;
        RECT 163.135 42.915 163.305 43.085 ;
        RECT 163.595 42.915 163.765 43.085 ;
        RECT 164.055 42.915 164.225 43.085 ;
        RECT 164.515 42.915 164.685 43.085 ;
        RECT 164.975 42.915 165.145 43.085 ;
        RECT 165.435 42.915 165.605 43.085 ;
        RECT 165.895 42.915 166.065 43.085 ;
        RECT 166.355 42.915 166.525 43.085 ;
        RECT 166.815 42.915 166.985 43.085 ;
        RECT 167.275 42.915 167.445 43.085 ;
        RECT 167.735 42.915 167.905 43.085 ;
        RECT 168.195 42.915 168.365 43.085 ;
        RECT 168.655 42.915 168.825 43.085 ;
        RECT 169.115 42.915 169.285 43.085 ;
        RECT 169.575 42.915 169.745 43.085 ;
        RECT 170.035 42.915 170.205 43.085 ;
        RECT 170.495 42.915 170.665 43.085 ;
        RECT 170.955 42.915 171.125 43.085 ;
        RECT 171.415 42.915 171.585 43.085 ;
        RECT 171.875 42.915 172.045 43.085 ;
        RECT 172.335 42.915 172.505 43.085 ;
        RECT 172.795 42.915 172.965 43.085 ;
        RECT 173.255 42.915 173.425 43.085 ;
        RECT 173.715 42.915 173.885 43.085 ;
        RECT 174.175 42.915 174.345 43.085 ;
        RECT 174.635 42.915 174.805 43.085 ;
        RECT 175.095 42.915 175.265 43.085 ;
        RECT 175.555 42.915 175.725 43.085 ;
        RECT 176.015 42.915 176.185 43.085 ;
        RECT 176.475 42.915 176.645 43.085 ;
        RECT 176.935 42.915 177.105 43.085 ;
        RECT 177.395 42.915 177.565 43.085 ;
        RECT 177.855 42.915 178.025 43.085 ;
        RECT 178.315 42.915 178.485 43.085 ;
        RECT 178.775 42.915 178.945 43.085 ;
        RECT 179.235 42.915 179.405 43.085 ;
        RECT 179.695 42.915 179.865 43.085 ;
        RECT 180.155 42.915 180.325 43.085 ;
        RECT 180.615 42.915 180.785 43.085 ;
        RECT 181.075 42.915 181.245 43.085 ;
        RECT 181.535 42.915 181.705 43.085 ;
        RECT 181.995 42.915 182.165 43.085 ;
        RECT 182.455 42.915 182.625 43.085 ;
        RECT 182.915 42.915 183.085 43.085 ;
        RECT 183.375 42.915 183.545 43.085 ;
        RECT 183.835 42.915 184.005 43.085 ;
        RECT 184.295 42.915 184.465 43.085 ;
        RECT 184.755 42.915 184.925 43.085 ;
        RECT 185.215 42.915 185.385 43.085 ;
        RECT 185.675 42.915 185.845 43.085 ;
        RECT 186.135 42.915 186.305 43.085 ;
        RECT 186.595 42.915 186.765 43.085 ;
        RECT 187.055 42.915 187.225 43.085 ;
        RECT 187.515 42.915 187.685 43.085 ;
        RECT 187.975 42.915 188.145 43.085 ;
        RECT 188.435 42.915 188.605 43.085 ;
        RECT 188.895 42.915 189.065 43.085 ;
        RECT 189.355 42.915 189.525 43.085 ;
        RECT 189.815 42.915 189.985 43.085 ;
        RECT 190.275 42.915 190.445 43.085 ;
        RECT 190.735 42.915 190.905 43.085 ;
        RECT 191.195 42.915 191.365 43.085 ;
        RECT 191.655 42.915 191.825 43.085 ;
        RECT 192.115 42.915 192.285 43.085 ;
        RECT 192.575 42.915 192.745 43.085 ;
        RECT 193.035 42.915 193.205 43.085 ;
        RECT 193.495 42.915 193.665 43.085 ;
        RECT 193.955 42.915 194.125 43.085 ;
        RECT 194.415 42.915 194.585 43.085 ;
        RECT 194.875 42.915 195.045 43.085 ;
        RECT 195.335 42.915 195.505 43.085 ;
        RECT 195.795 42.915 195.965 43.085 ;
        RECT 196.255 42.915 196.425 43.085 ;
        RECT 196.715 42.915 196.885 43.085 ;
        RECT 197.175 42.915 197.345 43.085 ;
        RECT 197.635 42.915 197.805 43.085 ;
        RECT 198.095 42.915 198.265 43.085 ;
        RECT 198.555 42.915 198.725 43.085 ;
        RECT 199.015 42.915 199.185 43.085 ;
        RECT 199.475 42.915 199.645 43.085 ;
        RECT 199.935 42.915 200.105 43.085 ;
        RECT 200.395 42.915 200.565 43.085 ;
        RECT 200.855 42.915 201.025 43.085 ;
        RECT 201.315 42.915 201.485 43.085 ;
        RECT 201.775 42.915 201.945 43.085 ;
        RECT 202.235 42.915 202.405 43.085 ;
        RECT 202.695 42.915 202.865 43.085 ;
        RECT 203.155 42.915 203.325 43.085 ;
        RECT 203.615 42.915 203.785 43.085 ;
        RECT 204.075 42.915 204.245 43.085 ;
        RECT 204.535 42.915 204.705 43.085 ;
        RECT 204.995 42.915 205.165 43.085 ;
        RECT 205.455 42.915 205.625 43.085 ;
        RECT 205.915 42.915 206.085 43.085 ;
        RECT 206.375 42.915 206.545 43.085 ;
        RECT 206.835 42.915 207.005 43.085 ;
        RECT 207.295 42.915 207.465 43.085 ;
        RECT 207.755 42.915 207.925 43.085 ;
        RECT 208.215 42.915 208.385 43.085 ;
        RECT 208.675 42.915 208.845 43.085 ;
        RECT 209.135 42.915 209.305 43.085 ;
        RECT 209.595 42.915 209.765 43.085 ;
        RECT 210.055 42.915 210.225 43.085 ;
        RECT 210.515 42.915 210.685 43.085 ;
        RECT 210.975 42.915 211.145 43.085 ;
        RECT 211.435 42.915 211.605 43.085 ;
        RECT 211.895 42.915 212.065 43.085 ;
        RECT 212.355 42.915 212.525 43.085 ;
        RECT 212.815 42.915 212.985 43.085 ;
        RECT 213.275 42.915 213.445 43.085 ;
        RECT 213.735 42.915 213.905 43.085 ;
        RECT 214.195 42.915 214.365 43.085 ;
        RECT 214.655 42.915 214.825 43.085 ;
        RECT 215.115 42.915 215.285 43.085 ;
        RECT 215.575 42.915 215.745 43.085 ;
        RECT 216.035 42.915 216.205 43.085 ;
        RECT 216.495 42.915 216.665 43.085 ;
        RECT 216.955 42.915 217.125 43.085 ;
        RECT 217.415 42.915 217.585 43.085 ;
        RECT 217.875 42.915 218.045 43.085 ;
        RECT 218.335 42.915 218.505 43.085 ;
        RECT 218.795 42.915 218.965 43.085 ;
        RECT 219.255 42.915 219.425 43.085 ;
        RECT 219.715 42.915 219.885 43.085 ;
        RECT 220.175 42.915 220.345 43.085 ;
        RECT 220.635 42.915 220.805 43.085 ;
        RECT 221.095 42.915 221.265 43.085 ;
        RECT 221.555 42.915 221.725 43.085 ;
        RECT 222.015 42.915 222.185 43.085 ;
        RECT 222.475 42.915 222.645 43.085 ;
        RECT 222.935 42.915 223.105 43.085 ;
        RECT 223.395 42.915 223.565 43.085 ;
        RECT 223.855 42.915 224.025 43.085 ;
        RECT 224.315 42.915 224.485 43.085 ;
        RECT 224.775 42.915 224.945 43.085 ;
        RECT 225.235 42.915 225.405 43.085 ;
        RECT 225.695 42.915 225.865 43.085 ;
        RECT 226.155 42.915 226.325 43.085 ;
        RECT 226.615 42.915 226.785 43.085 ;
        RECT 227.075 42.915 227.245 43.085 ;
        RECT 227.535 42.915 227.705 43.085 ;
        RECT 227.995 42.915 228.165 43.085 ;
        RECT 228.455 42.915 228.625 43.085 ;
        RECT 228.915 42.915 229.085 43.085 ;
        RECT 229.375 42.915 229.545 43.085 ;
        RECT 229.835 42.915 230.005 43.085 ;
        RECT 230.295 42.915 230.465 43.085 ;
        RECT 230.755 42.915 230.925 43.085 ;
        RECT 231.215 42.915 231.385 43.085 ;
        RECT 231.675 42.915 231.845 43.085 ;
        RECT 232.135 42.915 232.305 43.085 ;
        RECT 232.595 42.915 232.765 43.085 ;
        RECT 233.055 42.915 233.225 43.085 ;
        RECT 233.515 42.915 233.685 43.085 ;
        RECT 233.975 42.915 234.145 43.085 ;
        RECT 234.435 42.915 234.605 43.085 ;
        RECT 234.895 42.915 235.065 43.085 ;
        RECT 235.355 42.915 235.525 43.085 ;
        RECT 235.815 42.915 235.985 43.085 ;
        RECT 236.275 42.915 236.445 43.085 ;
        RECT 236.735 42.915 236.905 43.085 ;
        RECT 237.195 42.915 237.365 43.085 ;
        RECT 237.655 42.915 237.825 43.085 ;
        RECT 238.115 42.915 238.285 43.085 ;
        RECT 238.575 42.915 238.745 43.085 ;
        RECT 239.035 42.915 239.205 43.085 ;
        RECT 239.495 42.915 239.665 43.085 ;
        RECT 239.955 42.915 240.125 43.085 ;
        RECT 240.415 42.915 240.585 43.085 ;
        RECT 240.875 42.915 241.045 43.085 ;
        RECT 241.335 42.915 241.505 43.085 ;
        RECT 241.795 42.915 241.965 43.085 ;
        RECT 242.255 42.915 242.425 43.085 ;
        RECT 242.715 42.915 242.885 43.085 ;
        RECT 243.175 42.915 243.345 43.085 ;
        RECT 243.635 42.915 243.805 43.085 ;
        RECT 244.095 42.915 244.265 43.085 ;
        RECT 244.555 42.915 244.725 43.085 ;
        RECT 245.015 42.915 245.185 43.085 ;
        RECT 245.475 42.915 245.645 43.085 ;
        RECT 245.935 42.915 246.105 43.085 ;
        RECT 246.395 42.915 246.565 43.085 ;
        RECT 246.855 42.915 247.025 43.085 ;
        RECT 247.315 42.915 247.485 43.085 ;
        RECT 247.775 42.915 247.945 43.085 ;
        RECT 248.235 42.915 248.405 43.085 ;
        RECT 248.695 42.915 248.865 43.085 ;
        RECT 249.155 42.915 249.325 43.085 ;
        RECT 249.615 42.915 249.785 43.085 ;
        RECT 250.075 42.915 250.245 43.085 ;
        RECT 250.535 42.915 250.705 43.085 ;
        RECT 250.995 42.915 251.165 43.085 ;
        RECT 251.455 42.915 251.625 43.085 ;
        RECT 251.915 42.915 252.085 43.085 ;
        RECT 252.375 42.915 252.545 43.085 ;
        RECT 252.835 42.915 253.005 43.085 ;
        RECT 253.295 42.915 253.465 43.085 ;
        RECT 253.755 42.915 253.925 43.085 ;
        RECT 254.215 42.915 254.385 43.085 ;
        RECT 254.675 42.915 254.845 43.085 ;
        RECT 255.135 42.915 255.305 43.085 ;
        RECT 255.595 42.915 255.765 43.085 ;
        RECT 256.055 42.915 256.225 43.085 ;
        RECT 256.515 42.915 256.685 43.085 ;
        RECT 256.975 42.915 257.145 43.085 ;
        RECT 257.435 42.915 257.605 43.085 ;
        RECT 257.895 42.915 258.065 43.085 ;
        RECT 258.355 42.915 258.525 43.085 ;
        RECT 258.815 42.915 258.985 43.085 ;
        RECT 259.275 42.915 259.445 43.085 ;
        RECT 259.735 42.915 259.905 43.085 ;
        RECT 260.195 42.915 260.365 43.085 ;
        RECT 260.655 42.915 260.825 43.085 ;
        RECT 261.115 42.915 261.285 43.085 ;
        RECT 261.575 42.915 261.745 43.085 ;
        RECT 262.035 42.915 262.205 43.085 ;
        RECT 262.495 42.915 262.665 43.085 ;
        RECT 262.955 42.915 263.125 43.085 ;
        RECT 263.415 42.915 263.585 43.085 ;
        RECT 263.875 42.915 264.045 43.085 ;
        RECT 264.335 42.915 264.505 43.085 ;
        RECT 264.795 42.915 264.965 43.085 ;
        RECT 265.255 42.915 265.425 43.085 ;
        RECT 265.715 42.915 265.885 43.085 ;
        RECT 266.175 42.915 266.345 43.085 ;
        RECT 266.635 42.915 266.805 43.085 ;
        RECT 267.095 42.915 267.265 43.085 ;
        RECT 267.555 42.915 267.725 43.085 ;
        RECT 268.015 42.915 268.185 43.085 ;
        RECT 268.475 42.915 268.645 43.085 ;
        RECT 268.935 42.915 269.105 43.085 ;
        RECT 269.395 42.915 269.565 43.085 ;
        RECT 269.855 42.915 270.025 43.085 ;
        RECT 270.315 42.915 270.485 43.085 ;
        RECT 270.775 42.915 270.945 43.085 ;
        RECT 271.235 42.915 271.405 43.085 ;
        RECT 271.695 42.915 271.865 43.085 ;
        RECT 272.155 42.915 272.325 43.085 ;
        RECT 272.615 42.915 272.785 43.085 ;
        RECT 273.075 42.915 273.245 43.085 ;
        RECT 273.535 42.915 273.705 43.085 ;
        RECT 273.995 42.915 274.165 43.085 ;
        RECT 274.455 42.915 274.625 43.085 ;
        RECT 274.915 42.915 275.085 43.085 ;
        RECT 275.375 42.915 275.545 43.085 ;
        RECT 275.835 42.915 276.005 43.085 ;
        RECT 276.295 42.915 276.465 43.085 ;
        RECT 276.755 42.915 276.925 43.085 ;
        RECT 277.215 42.915 277.385 43.085 ;
        RECT 277.675 42.915 277.845 43.085 ;
        RECT 278.135 42.915 278.305 43.085 ;
        RECT 278.595 42.915 278.765 43.085 ;
        RECT 279.055 42.915 279.225 43.085 ;
        RECT 279.515 42.915 279.685 43.085 ;
        RECT 279.975 42.915 280.145 43.085 ;
        RECT 280.435 42.915 280.605 43.085 ;
        RECT 280.895 42.915 281.065 43.085 ;
        RECT 281.355 42.915 281.525 43.085 ;
        RECT 281.815 42.915 281.985 43.085 ;
        RECT 282.275 42.915 282.445 43.085 ;
        RECT 282.735 42.915 282.905 43.085 ;
        RECT 283.195 42.915 283.365 43.085 ;
        RECT 283.655 42.915 283.825 43.085 ;
        RECT 284.115 42.915 284.285 43.085 ;
        RECT 284.575 42.915 284.745 43.085 ;
        RECT 285.035 42.915 285.205 43.085 ;
        RECT 285.495 42.915 285.665 43.085 ;
        RECT 285.955 42.915 286.125 43.085 ;
        RECT 286.415 42.915 286.585 43.085 ;
        RECT 286.875 42.915 287.045 43.085 ;
        RECT 287.335 42.915 287.505 43.085 ;
        RECT 287.795 42.915 287.965 43.085 ;
        RECT 288.255 42.915 288.425 43.085 ;
        RECT 288.715 42.915 288.885 43.085 ;
        RECT 289.175 42.915 289.345 43.085 ;
        RECT 289.635 42.915 289.805 43.085 ;
        RECT 290.095 42.915 290.265 43.085 ;
        RECT 290.555 42.915 290.725 43.085 ;
        RECT 291.015 42.915 291.185 43.085 ;
        RECT 291.475 42.915 291.645 43.085 ;
        RECT 291.935 42.915 292.105 43.085 ;
        RECT 292.395 42.915 292.565 43.085 ;
        RECT 292.855 42.915 293.025 43.085 ;
        RECT 293.315 42.915 293.485 43.085 ;
        RECT 293.775 42.915 293.945 43.085 ;
        RECT 294.235 42.915 294.405 43.085 ;
        RECT 294.695 42.915 294.865 43.085 ;
        RECT 295.155 42.915 295.325 43.085 ;
        RECT 295.615 42.915 295.785 43.085 ;
        RECT 296.075 42.915 296.245 43.085 ;
        RECT 296.535 42.915 296.705 43.085 ;
        RECT 296.995 42.915 297.165 43.085 ;
        RECT 297.455 42.915 297.625 43.085 ;
        RECT 297.915 42.915 298.085 43.085 ;
        RECT 298.375 42.915 298.545 43.085 ;
        RECT 298.835 42.915 299.005 43.085 ;
        RECT 299.295 42.915 299.465 43.085 ;
        RECT 299.755 42.915 299.925 43.085 ;
        RECT 300.215 42.915 300.385 43.085 ;
        RECT 300.675 42.915 300.845 43.085 ;
        RECT 301.135 42.915 301.305 43.085 ;
        RECT 301.595 42.915 301.765 43.085 ;
        RECT 302.055 42.915 302.225 43.085 ;
        RECT 302.515 42.915 302.685 43.085 ;
        RECT 302.975 42.915 303.145 43.085 ;
        RECT 303.435 42.915 303.605 43.085 ;
        RECT 303.895 42.915 304.065 43.085 ;
        RECT 304.355 42.915 304.525 43.085 ;
        RECT 304.815 42.915 304.985 43.085 ;
        RECT 305.275 42.915 305.445 43.085 ;
        RECT 305.735 42.915 305.905 43.085 ;
        RECT 306.195 42.915 306.365 43.085 ;
        RECT 306.655 42.915 306.825 43.085 ;
        RECT 307.115 42.915 307.285 43.085 ;
        RECT 307.575 42.915 307.745 43.085 ;
        RECT 308.035 42.915 308.205 43.085 ;
        RECT 308.495 42.915 308.665 43.085 ;
        RECT 308.955 42.915 309.125 43.085 ;
        RECT 309.415 42.915 309.585 43.085 ;
        RECT 309.875 42.915 310.045 43.085 ;
        RECT 310.335 42.915 310.505 43.085 ;
        RECT 310.795 42.915 310.965 43.085 ;
        RECT 311.255 42.915 311.425 43.085 ;
        RECT 311.715 42.915 311.885 43.085 ;
        RECT 312.175 42.915 312.345 43.085 ;
        RECT 312.635 42.915 312.805 43.085 ;
        RECT 313.095 42.915 313.265 43.085 ;
        RECT 313.555 42.915 313.725 43.085 ;
        RECT 314.015 42.915 314.185 43.085 ;
        RECT 314.475 42.915 314.645 43.085 ;
        RECT 314.935 42.915 315.105 43.085 ;
        RECT 315.395 42.915 315.565 43.085 ;
        RECT 315.855 42.915 316.025 43.085 ;
        RECT 316.315 42.915 316.485 43.085 ;
        RECT 316.775 42.915 316.945 43.085 ;
        RECT 317.235 42.915 317.405 43.085 ;
        RECT 317.695 42.915 317.865 43.085 ;
        RECT 318.155 42.915 318.325 43.085 ;
        RECT 318.615 42.915 318.785 43.085 ;
        RECT 319.075 42.915 319.245 43.085 ;
        RECT 319.535 42.915 319.705 43.085 ;
        RECT 319.995 42.915 320.165 43.085 ;
        RECT 320.455 42.915 320.625 43.085 ;
        RECT 320.915 42.915 321.085 43.085 ;
        RECT 321.375 42.915 321.545 43.085 ;
        RECT 321.835 42.915 322.005 43.085 ;
        RECT 322.295 42.915 322.465 43.085 ;
        RECT 322.755 42.915 322.925 43.085 ;
        RECT 323.215 42.915 323.385 43.085 ;
        RECT 323.675 42.915 323.845 43.085 ;
        RECT 324.135 42.915 324.305 43.085 ;
        RECT 324.595 42.915 324.765 43.085 ;
        RECT 325.055 42.915 325.225 43.085 ;
        RECT 325.515 42.915 325.685 43.085 ;
        RECT 325.975 42.915 326.145 43.085 ;
        RECT 326.435 42.915 326.605 43.085 ;
        RECT 326.895 42.915 327.065 43.085 ;
        RECT 327.355 42.915 327.525 43.085 ;
        RECT 327.815 42.915 327.985 43.085 ;
        RECT 328.275 42.915 328.445 43.085 ;
        RECT 328.735 42.915 328.905 43.085 ;
        RECT 329.195 42.915 329.365 43.085 ;
        RECT 329.655 42.915 329.825 43.085 ;
        RECT 330.115 42.915 330.285 43.085 ;
        RECT 330.575 42.915 330.745 43.085 ;
        RECT 331.035 42.915 331.205 43.085 ;
        RECT 331.495 42.915 331.665 43.085 ;
        RECT 331.955 42.915 332.125 43.085 ;
        RECT 332.415 42.915 332.585 43.085 ;
        RECT 332.875 42.915 333.045 43.085 ;
        RECT 333.335 42.915 333.505 43.085 ;
        RECT 333.795 42.915 333.965 43.085 ;
        RECT 334.255 42.915 334.425 43.085 ;
        RECT 334.715 42.915 334.885 43.085 ;
        RECT 335.175 42.915 335.345 43.085 ;
        RECT 335.635 42.915 335.805 43.085 ;
        RECT 336.095 42.915 336.265 43.085 ;
        RECT 336.555 42.915 336.725 43.085 ;
        RECT 337.015 42.915 337.185 43.085 ;
        RECT 337.475 42.915 337.645 43.085 ;
        RECT 337.935 42.915 338.105 43.085 ;
        RECT 338.395 42.915 338.565 43.085 ;
        RECT 338.855 42.915 339.025 43.085 ;
        RECT 339.315 42.915 339.485 43.085 ;
        RECT 339.775 42.915 339.945 43.085 ;
        RECT 340.235 42.915 340.405 43.085 ;
        RECT 340.695 42.915 340.865 43.085 ;
        RECT 341.155 42.915 341.325 43.085 ;
        RECT 341.615 42.915 341.785 43.085 ;
        RECT 342.075 42.915 342.245 43.085 ;
        RECT 342.535 42.915 342.705 43.085 ;
        RECT 342.995 42.915 343.165 43.085 ;
        RECT 343.455 42.915 343.625 43.085 ;
        RECT 343.915 42.915 344.085 43.085 ;
        RECT 344.375 42.915 344.545 43.085 ;
        RECT 344.835 42.915 345.005 43.085 ;
        RECT 345.295 42.915 345.465 43.085 ;
        RECT 345.755 42.915 345.925 43.085 ;
        RECT 346.215 42.915 346.385 43.085 ;
        RECT 346.675 42.915 346.845 43.085 ;
        RECT 347.135 42.915 347.305 43.085 ;
        RECT 347.595 42.915 347.765 43.085 ;
        RECT 348.055 42.915 348.225 43.085 ;
        RECT 348.515 42.915 348.685 43.085 ;
        RECT 348.975 42.915 349.145 43.085 ;
        RECT 349.435 42.915 349.605 43.085 ;
        RECT 349.895 42.915 350.065 43.085 ;
        RECT 350.355 42.915 350.525 43.085 ;
        RECT 350.815 42.915 350.985 43.085 ;
        RECT 351.275 42.915 351.445 43.085 ;
        RECT 351.735 42.915 351.905 43.085 ;
        RECT 352.195 42.915 352.365 43.085 ;
        RECT 352.655 42.915 352.825 43.085 ;
        RECT 353.115 42.915 353.285 43.085 ;
        RECT 353.575 42.915 353.745 43.085 ;
        RECT 354.035 42.915 354.205 43.085 ;
        RECT 354.495 42.915 354.665 43.085 ;
        RECT 354.955 42.915 355.125 43.085 ;
        RECT 355.415 42.915 355.585 43.085 ;
        RECT 355.875 42.915 356.045 43.085 ;
        RECT 356.335 42.915 356.505 43.085 ;
        RECT 356.795 42.915 356.965 43.085 ;
        RECT 357.255 42.915 357.425 43.085 ;
        RECT 357.715 42.915 357.885 43.085 ;
        RECT 358.175 42.915 358.345 43.085 ;
        RECT 358.635 42.915 358.805 43.085 ;
        RECT 359.095 42.915 359.265 43.085 ;
        RECT 359.555 42.915 359.725 43.085 ;
        RECT 360.015 42.915 360.185 43.085 ;
        RECT 360.475 42.915 360.645 43.085 ;
        RECT 360.935 42.915 361.105 43.085 ;
        RECT 361.395 42.915 361.565 43.085 ;
        RECT 361.855 42.915 362.025 43.085 ;
        RECT 362.315 42.915 362.485 43.085 ;
        RECT 362.775 42.915 362.945 43.085 ;
        RECT 363.235 42.915 363.405 43.085 ;
        RECT 363.695 42.915 363.865 43.085 ;
        RECT 364.155 42.915 364.325 43.085 ;
        RECT 364.615 42.915 364.785 43.085 ;
        RECT 365.075 42.915 365.245 43.085 ;
        RECT 365.535 42.915 365.705 43.085 ;
        RECT 365.995 42.915 366.165 43.085 ;
        RECT 366.455 42.915 366.625 43.085 ;
        RECT 366.915 42.915 367.085 43.085 ;
        RECT 367.375 42.915 367.545 43.085 ;
        RECT 367.835 42.915 368.005 43.085 ;
        RECT 368.295 42.915 368.465 43.085 ;
        RECT 368.755 42.915 368.925 43.085 ;
        RECT 369.215 42.915 369.385 43.085 ;
        RECT 369.675 42.915 369.845 43.085 ;
        RECT 370.135 42.915 370.305 43.085 ;
        RECT 370.595 42.915 370.765 43.085 ;
        RECT 371.055 42.915 371.225 43.085 ;
        RECT 371.515 42.915 371.685 43.085 ;
        RECT 371.975 42.915 372.145 43.085 ;
        RECT 372.435 42.915 372.605 43.085 ;
        RECT 372.895 42.915 373.065 43.085 ;
        RECT 373.355 42.915 373.525 43.085 ;
        RECT 373.815 42.915 373.985 43.085 ;
        RECT 374.275 42.915 374.445 43.085 ;
        RECT 374.735 42.915 374.905 43.085 ;
        RECT 375.195 42.915 375.365 43.085 ;
        RECT 375.655 42.915 375.825 43.085 ;
        RECT 376.115 42.915 376.285 43.085 ;
        RECT 376.575 42.915 376.745 43.085 ;
        RECT 377.035 42.915 377.205 43.085 ;
        RECT 377.495 42.915 377.665 43.085 ;
        RECT 377.955 42.915 378.125 43.085 ;
        RECT 378.415 42.915 378.585 43.085 ;
        RECT 378.875 42.915 379.045 43.085 ;
        RECT 379.335 42.915 379.505 43.085 ;
        RECT 379.795 42.915 379.965 43.085 ;
        RECT 380.255 42.915 380.425 43.085 ;
        RECT 380.715 42.915 380.885 43.085 ;
        RECT 381.175 42.915 381.345 43.085 ;
        RECT 381.635 42.915 381.805 43.085 ;
        RECT 382.095 42.915 382.265 43.085 ;
        RECT 382.555 42.915 382.725 43.085 ;
        RECT 383.015 42.915 383.185 43.085 ;
        RECT 383.475 42.915 383.645 43.085 ;
        RECT 383.935 42.915 384.105 43.085 ;
        RECT 384.395 42.915 384.565 43.085 ;
        RECT 384.855 42.915 385.025 43.085 ;
        RECT 385.315 42.915 385.485 43.085 ;
        RECT 385.775 42.915 385.945 43.085 ;
        RECT 386.235 42.915 386.405 43.085 ;
        RECT 386.695 42.915 386.865 43.085 ;
        RECT 387.155 42.915 387.325 43.085 ;
        RECT 387.615 42.915 387.785 43.085 ;
        RECT 388.075 42.915 388.245 43.085 ;
        RECT 388.535 42.915 388.705 43.085 ;
        RECT 388.995 42.915 389.165 43.085 ;
        RECT 389.455 42.915 389.625 43.085 ;
        RECT 389.915 42.915 390.085 43.085 ;
        RECT 390.375 42.915 390.545 43.085 ;
        RECT 390.835 42.915 391.005 43.085 ;
        RECT 391.295 42.915 391.465 43.085 ;
        RECT 391.755 42.915 391.925 43.085 ;
        RECT 392.215 42.915 392.385 43.085 ;
        RECT 392.675 42.915 392.845 43.085 ;
        RECT 393.135 42.915 393.305 43.085 ;
        RECT 393.595 42.915 393.765 43.085 ;
        RECT 394.055 42.915 394.225 43.085 ;
        RECT 394.515 42.915 394.685 43.085 ;
        RECT 394.975 42.915 395.145 43.085 ;
        RECT 395.435 42.915 395.605 43.085 ;
        RECT 395.895 42.915 396.065 43.085 ;
        RECT 396.355 42.915 396.525 43.085 ;
        RECT 396.815 42.915 396.985 43.085 ;
        RECT 397.275 42.915 397.445 43.085 ;
        RECT 397.735 42.915 397.905 43.085 ;
        RECT 398.195 42.915 398.365 43.085 ;
        RECT 398.655 42.915 398.825 43.085 ;
        RECT 399.115 42.915 399.285 43.085 ;
        RECT 399.575 42.915 399.745 43.085 ;
        RECT 400.035 42.915 400.205 43.085 ;
        RECT 400.495 42.915 400.665 43.085 ;
        RECT 400.955 42.915 401.125 43.085 ;
        RECT 401.415 42.915 401.585 43.085 ;
        RECT 401.875 42.915 402.045 43.085 ;
        RECT 402.335 42.915 402.505 43.085 ;
        RECT 402.795 42.915 402.965 43.085 ;
        RECT 403.255 42.915 403.425 43.085 ;
        RECT 403.715 42.915 403.885 43.085 ;
        RECT 404.175 42.915 404.345 43.085 ;
        RECT 404.635 42.915 404.805 43.085 ;
        RECT 405.095 42.915 405.265 43.085 ;
        RECT 405.555 42.915 405.725 43.085 ;
        RECT 406.015 42.915 406.185 43.085 ;
        RECT 406.475 42.915 406.645 43.085 ;
        RECT 406.935 42.915 407.105 43.085 ;
        RECT 407.395 42.915 407.565 43.085 ;
        RECT 407.855 42.915 408.025 43.085 ;
        RECT 408.315 42.915 408.485 43.085 ;
        RECT 408.775 42.915 408.945 43.085 ;
        RECT 409.235 42.915 409.405 43.085 ;
        RECT 409.695 42.915 409.865 43.085 ;
        RECT 410.155 42.915 410.325 43.085 ;
        RECT 410.615 42.915 410.785 43.085 ;
        RECT 411.075 42.915 411.245 43.085 ;
        RECT 411.535 42.915 411.705 43.085 ;
        RECT 411.995 42.915 412.165 43.085 ;
        RECT 412.455 42.915 412.625 43.085 ;
        RECT 412.915 42.915 413.085 43.085 ;
        RECT 413.375 42.915 413.545 43.085 ;
        RECT 413.835 42.915 414.005 43.085 ;
        RECT 414.295 42.915 414.465 43.085 ;
        RECT 414.755 42.915 414.925 43.085 ;
        RECT 415.215 42.915 415.385 43.085 ;
        RECT 415.675 42.915 415.845 43.085 ;
        RECT 416.135 42.915 416.305 43.085 ;
        RECT 416.595 42.915 416.765 43.085 ;
        RECT 417.055 42.915 417.225 43.085 ;
        RECT 417.515 42.915 417.685 43.085 ;
        RECT 417.975 42.915 418.145 43.085 ;
        RECT 418.435 42.915 418.605 43.085 ;
        RECT 418.895 42.915 419.065 43.085 ;
        RECT 419.355 42.915 419.525 43.085 ;
        RECT 419.815 42.915 419.985 43.085 ;
        RECT 420.275 42.915 420.445 43.085 ;
        RECT 420.735 42.915 420.905 43.085 ;
        RECT 421.195 42.915 421.365 43.085 ;
        RECT 421.655 42.915 421.825 43.085 ;
        RECT 422.115 42.915 422.285 43.085 ;
        RECT 422.575 42.915 422.745 43.085 ;
        RECT 423.035 42.915 423.205 43.085 ;
        RECT 423.495 42.915 423.665 43.085 ;
        RECT 423.955 42.915 424.125 43.085 ;
        RECT 424.415 42.915 424.585 43.085 ;
        RECT 424.875 42.915 425.045 43.085 ;
        RECT 425.335 42.915 425.505 43.085 ;
        RECT 425.795 42.915 425.965 43.085 ;
        RECT 426.255 42.915 426.425 43.085 ;
        RECT 426.715 42.915 426.885 43.085 ;
        RECT 427.175 42.915 427.345 43.085 ;
        RECT 427.635 42.915 427.805 43.085 ;
        RECT 428.095 42.915 428.265 43.085 ;
        RECT 428.555 42.915 428.725 43.085 ;
        RECT 429.015 42.915 429.185 43.085 ;
        RECT 429.475 42.915 429.645 43.085 ;
        RECT 429.935 42.915 430.105 43.085 ;
        RECT 430.395 42.915 430.565 43.085 ;
        RECT 430.855 42.915 431.025 43.085 ;
        RECT 431.315 42.915 431.485 43.085 ;
        RECT 431.775 42.915 431.945 43.085 ;
        RECT 432.235 42.915 432.405 43.085 ;
        RECT 432.695 42.915 432.865 43.085 ;
        RECT 433.155 42.915 433.325 43.085 ;
        RECT 433.615 42.915 433.785 43.085 ;
        RECT 434.075 42.915 434.245 43.085 ;
        RECT 434.535 42.915 434.705 43.085 ;
        RECT 434.995 42.915 435.165 43.085 ;
        RECT 435.455 42.915 435.625 43.085 ;
        RECT 435.915 42.915 436.085 43.085 ;
        RECT 436.375 42.915 436.545 43.085 ;
        RECT 436.835 42.915 437.005 43.085 ;
        RECT 437.295 42.915 437.465 43.085 ;
        RECT 437.755 42.915 437.925 43.085 ;
        RECT 438.215 42.915 438.385 43.085 ;
        RECT 438.675 42.915 438.845 43.085 ;
        RECT 439.135 42.915 439.305 43.085 ;
        RECT 439.595 42.915 439.765 43.085 ;
        RECT 440.055 42.915 440.225 43.085 ;
        RECT 440.515 42.915 440.685 43.085 ;
        RECT 440.975 42.915 441.145 43.085 ;
        RECT 441.435 42.915 441.605 43.085 ;
        RECT 441.895 42.915 442.065 43.085 ;
        RECT 442.355 42.915 442.525 43.085 ;
        RECT 442.815 42.915 442.985 43.085 ;
        RECT 443.275 42.915 443.445 43.085 ;
        RECT 443.735 42.915 443.905 43.085 ;
        RECT 444.195 42.915 444.365 43.085 ;
        RECT 444.655 42.915 444.825 43.085 ;
        RECT 445.115 42.915 445.285 43.085 ;
        RECT 445.575 42.915 445.745 43.085 ;
        RECT 446.035 42.915 446.205 43.085 ;
        RECT 446.495 42.915 446.665 43.085 ;
        RECT 446.955 42.915 447.125 43.085 ;
        RECT 447.415 42.915 447.585 43.085 ;
        RECT 447.875 42.915 448.045 43.085 ;
        RECT 448.335 42.915 448.505 43.085 ;
        RECT 448.795 42.915 448.965 43.085 ;
        RECT 449.255 42.915 449.425 43.085 ;
        RECT 449.715 42.915 449.885 43.085 ;
        RECT 450.175 42.915 450.345 43.085 ;
        RECT 450.635 42.915 450.805 43.085 ;
        RECT 451.095 42.915 451.265 43.085 ;
        RECT 451.555 42.915 451.725 43.085 ;
        RECT 452.015 42.915 452.185 43.085 ;
        RECT 452.475 42.915 452.645 43.085 ;
        RECT 452.935 42.915 453.105 43.085 ;
        RECT 453.395 42.915 453.565 43.085 ;
        RECT 453.855 42.915 454.025 43.085 ;
        RECT 454.315 42.915 454.485 43.085 ;
        RECT 454.775 42.915 454.945 43.085 ;
        RECT 455.235 42.915 455.405 43.085 ;
        RECT 455.695 42.915 455.865 43.085 ;
        RECT 456.155 42.915 456.325 43.085 ;
        RECT 456.615 42.915 456.785 43.085 ;
        RECT 457.075 42.915 457.245 43.085 ;
        RECT 457.535 42.915 457.705 43.085 ;
        RECT 457.995 42.915 458.165 43.085 ;
        RECT 458.455 42.915 458.625 43.085 ;
        RECT 458.915 42.915 459.085 43.085 ;
        RECT 459.375 42.915 459.545 43.085 ;
        RECT 459.835 42.915 460.005 43.085 ;
        RECT 460.295 42.915 460.465 43.085 ;
        RECT 460.755 42.915 460.925 43.085 ;
        RECT 461.215 42.915 461.385 43.085 ;
        RECT 461.675 42.915 461.845 43.085 ;
        RECT 462.135 42.915 462.305 43.085 ;
        RECT 462.595 42.915 462.765 43.085 ;
        RECT 463.055 42.915 463.225 43.085 ;
        RECT 463.515 42.915 463.685 43.085 ;
        RECT 463.975 42.915 464.145 43.085 ;
        RECT 464.435 42.915 464.605 43.085 ;
        RECT 464.895 42.915 465.065 43.085 ;
        RECT 465.355 42.915 465.525 43.085 ;
        RECT 465.815 42.915 465.985 43.085 ;
        RECT 466.275 42.915 466.445 43.085 ;
        RECT 466.735 42.915 466.905 43.085 ;
        RECT 467.195 42.915 467.365 43.085 ;
        RECT 467.655 42.915 467.825 43.085 ;
        RECT 468.115 42.915 468.285 43.085 ;
        RECT 468.575 42.915 468.745 43.085 ;
        RECT 469.035 42.915 469.205 43.085 ;
        RECT 469.495 42.915 469.665 43.085 ;
        RECT 469.955 42.915 470.125 43.085 ;
        RECT 470.415 42.915 470.585 43.085 ;
        RECT 470.875 42.915 471.045 43.085 ;
        RECT 471.335 42.915 471.505 43.085 ;
        RECT 471.795 42.915 471.965 43.085 ;
        RECT 472.255 42.915 472.425 43.085 ;
        RECT 472.715 42.915 472.885 43.085 ;
        RECT 473.175 42.915 473.345 43.085 ;
        RECT 473.635 42.915 473.805 43.085 ;
        RECT 474.095 42.915 474.265 43.085 ;
        RECT 474.555 42.915 474.725 43.085 ;
        RECT 475.015 42.915 475.185 43.085 ;
        RECT 475.475 42.915 475.645 43.085 ;
        RECT 475.935 42.915 476.105 43.085 ;
        RECT 476.395 42.915 476.565 43.085 ;
        RECT 476.855 42.915 477.025 43.085 ;
        RECT 477.315 42.915 477.485 43.085 ;
        RECT 477.775 42.915 477.945 43.085 ;
        RECT 478.235 42.915 478.405 43.085 ;
        RECT 478.695 42.915 478.865 43.085 ;
        RECT 479.155 42.915 479.325 43.085 ;
        RECT 479.615 42.915 479.785 43.085 ;
        RECT 480.075 42.915 480.245 43.085 ;
        RECT 480.535 42.915 480.705 43.085 ;
        RECT 480.995 42.915 481.165 43.085 ;
        RECT 481.455 42.915 481.625 43.085 ;
        RECT 481.915 42.915 482.085 43.085 ;
        RECT 482.375 42.915 482.545 43.085 ;
        RECT 482.835 42.915 483.005 43.085 ;
        RECT 483.295 42.915 483.465 43.085 ;
        RECT 483.755 42.915 483.925 43.085 ;
        RECT 484.215 42.915 484.385 43.085 ;
        RECT 484.675 42.915 484.845 43.085 ;
        RECT 485.135 42.915 485.305 43.085 ;
        RECT 485.595 42.915 485.765 43.085 ;
        RECT 486.055 42.915 486.225 43.085 ;
        RECT 486.515 42.915 486.685 43.085 ;
        RECT 486.975 42.915 487.145 43.085 ;
        RECT 487.435 42.915 487.605 43.085 ;
        RECT 487.895 42.915 488.065 43.085 ;
        RECT 488.355 42.915 488.525 43.085 ;
        RECT 488.815 42.915 488.985 43.085 ;
        RECT 489.275 42.915 489.445 43.085 ;
        RECT 489.735 42.915 489.905 43.085 ;
        RECT 490.195 42.915 490.365 43.085 ;
        RECT 490.655 42.915 490.825 43.085 ;
        RECT 491.115 42.915 491.285 43.085 ;
        RECT 491.575 42.915 491.745 43.085 ;
        RECT 492.035 42.915 492.205 43.085 ;
        RECT 492.495 42.915 492.665 43.085 ;
        RECT 492.955 42.915 493.125 43.085 ;
        RECT 493.415 42.915 493.585 43.085 ;
        RECT 493.875 42.915 494.045 43.085 ;
        RECT 494.335 42.915 494.505 43.085 ;
        RECT 494.795 42.915 494.965 43.085 ;
        RECT 495.255 42.915 495.425 43.085 ;
        RECT 495.715 42.915 495.885 43.085 ;
        RECT 496.175 42.915 496.345 43.085 ;
        RECT 496.635 42.915 496.805 43.085 ;
        RECT 497.095 42.915 497.265 43.085 ;
        RECT 497.555 42.915 497.725 43.085 ;
        RECT 498.015 42.915 498.185 43.085 ;
        RECT 498.475 42.915 498.645 43.085 ;
        RECT 498.935 42.915 499.105 43.085 ;
        RECT 499.395 42.915 499.565 43.085 ;
        RECT 499.855 42.915 500.025 43.085 ;
        RECT 500.315 42.915 500.485 43.085 ;
        RECT 500.775 42.915 500.945 43.085 ;
        RECT 501.235 42.915 501.405 43.085 ;
        RECT 501.695 42.915 501.865 43.085 ;
        RECT 502.155 42.915 502.325 43.085 ;
        RECT 502.615 42.915 502.785 43.085 ;
        RECT 503.075 42.915 503.245 43.085 ;
        RECT 503.535 42.915 503.705 43.085 ;
        RECT 503.995 42.915 504.165 43.085 ;
        RECT 504.455 42.915 504.625 43.085 ;
        RECT 504.915 42.915 505.085 43.085 ;
        RECT 505.375 42.915 505.545 43.085 ;
        RECT 505.835 42.915 506.005 43.085 ;
        RECT 506.295 42.915 506.465 43.085 ;
        RECT 506.755 42.915 506.925 43.085 ;
        RECT 507.215 42.915 507.385 43.085 ;
        RECT 507.675 42.915 507.845 43.085 ;
        RECT 508.135 42.915 508.305 43.085 ;
        RECT 508.595 42.915 508.765 43.085 ;
        RECT 509.055 42.915 509.225 43.085 ;
        RECT 509.515 42.915 509.685 43.085 ;
        RECT 509.975 42.915 510.145 43.085 ;
        RECT 510.435 42.915 510.605 43.085 ;
        RECT 510.895 42.915 511.065 43.085 ;
        RECT 511.355 42.915 511.525 43.085 ;
        RECT 511.815 42.915 511.985 43.085 ;
        RECT 512.275 42.915 512.445 43.085 ;
        RECT 512.735 42.915 512.905 43.085 ;
        RECT 513.195 42.915 513.365 43.085 ;
        RECT 513.655 42.915 513.825 43.085 ;
        RECT 514.115 42.915 514.285 43.085 ;
        RECT 514.575 42.915 514.745 43.085 ;
        RECT 515.035 42.915 515.205 43.085 ;
        RECT 515.495 42.915 515.665 43.085 ;
        RECT 515.955 42.915 516.125 43.085 ;
        RECT 516.415 42.915 516.585 43.085 ;
        RECT 516.875 42.915 517.045 43.085 ;
        RECT 517.335 42.915 517.505 43.085 ;
        RECT 517.795 42.915 517.965 43.085 ;
        RECT 518.255 42.915 518.425 43.085 ;
        RECT 518.715 42.915 518.885 43.085 ;
        RECT 519.175 42.915 519.345 43.085 ;
        RECT 519.635 42.915 519.805 43.085 ;
        RECT 520.095 42.915 520.265 43.085 ;
        RECT 520.555 42.915 520.725 43.085 ;
        RECT 521.015 42.915 521.185 43.085 ;
        RECT 521.475 42.915 521.645 43.085 ;
        RECT 521.935 42.915 522.105 43.085 ;
        RECT 522.395 42.915 522.565 43.085 ;
        RECT 522.855 42.915 523.025 43.085 ;
        RECT 523.315 42.915 523.485 43.085 ;
        RECT 523.775 42.915 523.945 43.085 ;
        RECT 524.235 42.915 524.405 43.085 ;
        RECT 524.695 42.915 524.865 43.085 ;
        RECT 525.155 42.915 525.325 43.085 ;
        RECT 525.615 42.915 525.785 43.085 ;
        RECT 526.075 42.915 526.245 43.085 ;
        RECT 526.535 42.915 526.705 43.085 ;
        RECT 526.995 42.915 527.165 43.085 ;
        RECT 527.455 42.915 527.625 43.085 ;
        RECT 527.915 42.915 528.085 43.085 ;
        RECT 528.375 42.915 528.545 43.085 ;
        RECT 528.835 42.915 529.005 43.085 ;
        RECT 529.295 42.915 529.465 43.085 ;
        RECT 529.755 42.915 529.925 43.085 ;
        RECT 530.215 42.915 530.385 43.085 ;
        RECT 530.675 42.915 530.845 43.085 ;
        RECT 531.135 42.915 531.305 43.085 ;
        RECT 531.595 42.915 531.765 43.085 ;
        RECT 532.055 42.915 532.225 43.085 ;
        RECT 532.515 42.915 532.685 43.085 ;
        RECT 532.975 42.915 533.145 43.085 ;
        RECT 533.435 42.915 533.605 43.085 ;
        RECT 533.895 42.915 534.065 43.085 ;
        RECT 534.355 42.915 534.525 43.085 ;
        RECT 534.815 42.915 534.985 43.085 ;
        RECT 535.275 42.915 535.445 43.085 ;
        RECT 535.735 42.915 535.905 43.085 ;
        RECT 536.195 42.915 536.365 43.085 ;
        RECT 536.655 42.915 536.825 43.085 ;
        RECT 537.115 42.915 537.285 43.085 ;
        RECT 537.575 42.915 537.745 43.085 ;
        RECT 538.035 42.915 538.205 43.085 ;
        RECT 538.495 42.915 538.665 43.085 ;
        RECT 538.955 42.915 539.125 43.085 ;
        RECT 539.415 42.915 539.585 43.085 ;
        RECT 539.875 42.915 540.045 43.085 ;
        RECT 540.335 42.915 540.505 43.085 ;
        RECT 540.795 42.915 540.965 43.085 ;
        RECT 541.255 42.915 541.425 43.085 ;
        RECT 541.715 42.915 541.885 43.085 ;
        RECT 542.175 42.915 542.345 43.085 ;
        RECT 542.635 42.915 542.805 43.085 ;
        RECT 543.095 42.915 543.265 43.085 ;
        RECT 543.555 42.915 543.725 43.085 ;
        RECT 544.015 42.915 544.185 43.085 ;
        RECT 544.475 42.915 544.645 43.085 ;
        RECT 544.935 42.915 545.105 43.085 ;
        RECT 545.395 42.915 545.565 43.085 ;
        RECT 545.855 42.915 546.025 43.085 ;
        RECT 546.315 42.915 546.485 43.085 ;
        RECT 546.775 42.915 546.945 43.085 ;
        RECT 547.235 42.915 547.405 43.085 ;
        RECT 547.695 42.915 547.865 43.085 ;
        RECT 548.155 42.915 548.325 43.085 ;
        RECT 548.615 42.915 548.785 43.085 ;
        RECT 549.075 42.915 549.245 43.085 ;
        RECT 549.535 42.915 549.705 43.085 ;
        RECT 549.995 42.915 550.165 43.085 ;
        RECT 550.455 42.915 550.625 43.085 ;
        RECT 550.915 42.915 551.085 43.085 ;
        RECT 551.375 42.915 551.545 43.085 ;
        RECT 551.835 42.915 552.005 43.085 ;
        RECT 552.295 42.915 552.465 43.085 ;
        RECT 552.755 42.915 552.925 43.085 ;
        RECT 553.215 42.915 553.385 43.085 ;
        RECT 553.675 42.915 553.845 43.085 ;
        RECT 554.135 42.915 554.305 43.085 ;
        RECT 554.595 42.915 554.765 43.085 ;
        RECT 555.055 42.915 555.225 43.085 ;
        RECT 555.515 42.915 555.685 43.085 ;
        RECT 555.975 42.915 556.145 43.085 ;
        RECT 556.435 42.915 556.605 43.085 ;
        RECT 556.895 42.915 557.065 43.085 ;
        RECT 557.355 42.915 557.525 43.085 ;
        RECT 557.815 42.915 557.985 43.085 ;
        RECT 558.275 42.915 558.445 43.085 ;
        RECT 558.735 42.915 558.905 43.085 ;
        RECT 559.195 42.915 559.365 43.085 ;
        RECT 559.655 42.915 559.825 43.085 ;
        RECT 560.115 42.915 560.285 43.085 ;
        RECT 560.575 42.915 560.745 43.085 ;
        RECT 561.035 42.915 561.205 43.085 ;
        RECT 561.495 42.915 561.665 43.085 ;
        RECT 561.955 42.915 562.125 43.085 ;
        RECT 562.415 42.915 562.585 43.085 ;
        RECT 562.875 42.915 563.045 43.085 ;
        RECT 563.335 42.915 563.505 43.085 ;
        RECT 563.795 42.915 563.965 43.085 ;
        RECT 564.255 42.915 564.425 43.085 ;
        RECT 564.715 42.915 564.885 43.085 ;
        RECT 565.175 42.915 565.345 43.085 ;
        RECT 565.635 42.915 565.805 43.085 ;
        RECT 566.095 42.915 566.265 43.085 ;
        RECT 566.555 42.915 566.725 43.085 ;
        RECT 567.015 42.915 567.185 43.085 ;
        RECT 567.475 42.915 567.645 43.085 ;
        RECT 567.935 42.915 568.105 43.085 ;
        RECT 568.395 42.915 568.565 43.085 ;
        RECT 568.855 42.915 569.025 43.085 ;
        RECT 569.315 42.915 569.485 43.085 ;
        RECT 569.775 42.915 569.945 43.085 ;
        RECT 570.235 42.915 570.405 43.085 ;
        RECT 570.695 42.915 570.865 43.085 ;
        RECT 571.155 42.915 571.325 43.085 ;
        RECT 571.615 42.915 571.785 43.085 ;
        RECT 572.075 42.915 572.245 43.085 ;
        RECT 572.535 42.915 572.705 43.085 ;
        RECT 572.995 42.915 573.165 43.085 ;
        RECT 573.455 42.915 573.625 43.085 ;
        RECT 573.915 42.915 574.085 43.085 ;
        RECT 574.375 42.915 574.545 43.085 ;
        RECT 574.835 42.915 575.005 43.085 ;
        RECT 575.295 42.915 575.465 43.085 ;
        RECT 575.755 42.915 575.925 43.085 ;
        RECT 576.215 42.915 576.385 43.085 ;
        RECT 576.675 42.915 576.845 43.085 ;
        RECT 577.135 42.915 577.305 43.085 ;
        RECT 577.595 42.915 577.765 43.085 ;
        RECT 578.055 42.915 578.225 43.085 ;
        RECT 578.515 42.915 578.685 43.085 ;
        RECT 578.975 42.915 579.145 43.085 ;
        RECT 579.435 42.915 579.605 43.085 ;
        RECT 579.895 42.915 580.065 43.085 ;
        RECT 580.355 42.915 580.525 43.085 ;
        RECT 580.815 42.915 580.985 43.085 ;
        RECT 581.275 42.915 581.445 43.085 ;
        RECT 581.735 42.915 581.905 43.085 ;
        RECT 582.195 42.915 582.365 43.085 ;
        RECT 582.655 42.915 582.825 43.085 ;
        RECT 583.115 42.915 583.285 43.085 ;
        RECT 583.575 42.915 583.745 43.085 ;
        RECT 584.035 42.915 584.205 43.085 ;
        RECT 584.495 42.915 584.665 43.085 ;
        RECT 584.955 42.915 585.125 43.085 ;
        RECT 585.415 42.915 585.585 43.085 ;
        RECT 585.875 42.915 586.045 43.085 ;
        RECT 586.335 42.915 586.505 43.085 ;
        RECT 586.795 42.915 586.965 43.085 ;
        RECT 587.255 42.915 587.425 43.085 ;
        RECT 587.715 42.915 587.885 43.085 ;
        RECT 588.175 42.915 588.345 43.085 ;
        RECT 588.635 42.915 588.805 43.085 ;
        RECT 589.095 42.915 589.265 43.085 ;
        RECT 589.555 42.915 589.725 43.085 ;
        RECT 590.015 42.915 590.185 43.085 ;
        RECT 590.475 42.915 590.645 43.085 ;
        RECT 590.935 42.915 591.105 43.085 ;
        RECT 591.395 42.915 591.565 43.085 ;
        RECT 591.855 42.915 592.025 43.085 ;
        RECT 592.315 42.915 592.485 43.085 ;
        RECT 592.775 42.915 592.945 43.085 ;
        RECT 593.235 42.915 593.405 43.085 ;
        RECT 593.695 42.915 593.865 43.085 ;
        RECT 594.155 42.915 594.325 43.085 ;
        RECT 594.615 42.915 594.785 43.085 ;
        RECT 595.075 42.915 595.245 43.085 ;
        RECT 595.535 42.915 595.705 43.085 ;
        RECT 595.995 42.915 596.165 43.085 ;
        RECT 596.455 42.915 596.625 43.085 ;
        RECT 596.915 42.915 597.085 43.085 ;
        RECT 597.375 42.915 597.545 43.085 ;
        RECT 597.835 42.915 598.005 43.085 ;
        RECT 598.295 42.915 598.465 43.085 ;
        RECT 598.755 42.915 598.925 43.085 ;
        RECT 599.215 42.915 599.385 43.085 ;
        RECT 599.675 42.915 599.845 43.085 ;
        RECT 600.135 42.915 600.305 43.085 ;
        RECT 600.595 42.915 600.765 43.085 ;
        RECT 601.055 42.915 601.225 43.085 ;
        RECT 601.515 42.915 601.685 43.085 ;
        RECT 601.975 42.915 602.145 43.085 ;
        RECT 602.435 42.915 602.605 43.085 ;
        RECT 602.895 42.915 603.065 43.085 ;
        RECT 603.355 42.915 603.525 43.085 ;
        RECT 603.815 42.915 603.985 43.085 ;
        RECT 604.275 42.915 604.445 43.085 ;
        RECT 604.735 42.915 604.905 43.085 ;
        RECT 605.195 42.915 605.365 43.085 ;
        RECT 605.655 42.915 605.825 43.085 ;
        RECT 606.115 42.915 606.285 43.085 ;
        RECT 606.575 42.915 606.745 43.085 ;
        RECT 607.035 42.915 607.205 43.085 ;
        RECT 607.495 42.915 607.665 43.085 ;
        RECT 607.955 42.915 608.125 43.085 ;
        RECT 608.415 42.915 608.585 43.085 ;
        RECT 608.875 42.915 609.045 43.085 ;
        RECT 609.335 42.915 609.505 43.085 ;
        RECT 609.795 42.915 609.965 43.085 ;
        RECT 610.255 42.915 610.425 43.085 ;
        RECT 610.715 42.915 610.885 43.085 ;
        RECT 611.175 42.915 611.345 43.085 ;
        RECT 611.635 42.915 611.805 43.085 ;
        RECT 612.095 42.915 612.265 43.085 ;
        RECT 612.555 42.915 612.725 43.085 ;
        RECT 613.015 42.915 613.185 43.085 ;
        RECT 613.475 42.915 613.645 43.085 ;
        RECT 613.935 42.915 614.105 43.085 ;
        RECT 614.395 42.915 614.565 43.085 ;
        RECT 614.855 42.915 615.025 43.085 ;
        RECT 615.315 42.915 615.485 43.085 ;
        RECT 615.775 42.915 615.945 43.085 ;
        RECT 616.235 42.915 616.405 43.085 ;
        RECT 616.695 42.915 616.865 43.085 ;
        RECT 617.155 42.915 617.325 43.085 ;
        RECT 617.615 42.915 617.785 43.085 ;
        RECT 618.075 42.915 618.245 43.085 ;
        RECT 618.535 42.915 618.705 43.085 ;
        RECT 618.995 42.915 619.165 43.085 ;
        RECT 619.455 42.915 619.625 43.085 ;
        RECT 619.915 42.915 620.085 43.085 ;
        RECT 620.375 42.915 620.545 43.085 ;
        RECT 620.835 42.915 621.005 43.085 ;
        RECT 621.295 42.915 621.465 43.085 ;
        RECT 621.755 42.915 621.925 43.085 ;
        RECT 622.215 42.915 622.385 43.085 ;
        RECT 622.675 42.915 622.845 43.085 ;
        RECT 623.135 42.915 623.305 43.085 ;
        RECT 623.595 42.915 623.765 43.085 ;
        RECT 624.055 42.915 624.225 43.085 ;
        RECT 624.515 42.915 624.685 43.085 ;
        RECT 624.975 42.915 625.145 43.085 ;
        RECT 625.435 42.915 625.605 43.085 ;
        RECT 625.895 42.915 626.065 43.085 ;
        RECT 626.355 42.915 626.525 43.085 ;
        RECT 626.815 42.915 626.985 43.085 ;
        RECT 627.275 42.915 627.445 43.085 ;
        RECT 627.735 42.915 627.905 43.085 ;
        RECT 628.195 42.915 628.365 43.085 ;
        RECT 628.655 42.915 628.825 43.085 ;
        RECT 629.115 42.915 629.285 43.085 ;
        RECT 629.575 42.915 629.745 43.085 ;
        RECT 630.035 42.915 630.205 43.085 ;
        RECT 630.495 42.915 630.665 43.085 ;
        RECT 630.955 42.915 631.125 43.085 ;
        RECT 215.115 42.405 215.285 42.575 ;
        RECT 155.775 42.065 155.945 42.235 ;
        RECT 163.135 41.725 163.305 41.895 ;
        RECT 175.095 41.725 175.265 41.895 ;
        RECT 221.555 42.405 221.725 42.575 ;
        RECT 224.775 42.065 224.945 42.235 ;
        RECT 224.315 41.725 224.485 41.895 ;
        RECT 258.355 40.705 258.525 40.875 ;
        RECT 42.615 619.555 42.785 619.725 ;
        RECT 43.075 619.555 43.245 619.725 ;
        RECT 43.535 619.555 43.705 619.725 ;
        RECT 43.995 619.555 44.165 619.725 ;
        RECT 44.455 619.555 44.625 619.725 ;
        RECT 44.915 619.555 45.085 619.725 ;
        RECT 45.375 619.555 45.545 619.725 ;
        RECT 45.835 619.555 46.005 619.725 ;
        RECT 46.295 619.555 46.465 619.725 ;
        RECT 46.755 619.555 46.925 619.725 ;
        RECT 47.215 619.555 47.385 619.725 ;
        RECT 47.675 619.555 47.845 619.725 ;
        RECT 48.135 619.555 48.305 619.725 ;
        RECT 48.595 619.555 48.765 619.725 ;
        RECT 49.055 619.555 49.225 619.725 ;
        RECT 49.515 619.555 49.685 619.725 ;
        RECT 49.975 619.555 50.145 619.725 ;
        RECT 50.435 619.555 50.605 619.725 ;
        RECT 50.895 619.555 51.065 619.725 ;
        RECT 51.355 619.555 51.525 619.725 ;
        RECT 51.815 619.555 51.985 619.725 ;
        RECT 52.275 619.555 52.445 619.725 ;
        RECT 52.735 619.555 52.905 619.725 ;
        RECT 53.195 619.555 53.365 619.725 ;
        RECT 53.655 619.555 53.825 619.725 ;
        RECT 42.615 616.835 42.785 617.005 ;
        RECT 43.075 616.835 43.245 617.005 ;
        RECT 43.535 616.835 43.705 617.005 ;
        RECT 43.995 616.835 44.165 617.005 ;
        RECT 44.455 616.835 44.625 617.005 ;
        RECT 44.915 616.835 45.085 617.005 ;
        RECT 45.375 616.835 45.545 617.005 ;
        RECT 45.835 616.835 46.005 617.005 ;
        RECT 46.295 616.835 46.465 617.005 ;
        RECT 46.755 616.835 46.925 617.005 ;
        RECT 47.215 616.835 47.385 617.005 ;
        RECT 47.675 616.835 47.845 617.005 ;
        RECT 48.135 616.835 48.305 617.005 ;
        RECT 48.595 616.835 48.765 617.005 ;
        RECT 49.055 616.835 49.225 617.005 ;
        RECT 49.515 616.835 49.685 617.005 ;
        RECT 49.975 616.835 50.145 617.005 ;
        RECT 50.435 616.835 50.605 617.005 ;
        RECT 50.895 616.835 51.065 617.005 ;
        RECT 51.355 616.835 51.525 617.005 ;
        RECT 51.815 616.835 51.985 617.005 ;
        RECT 52.275 616.835 52.445 617.005 ;
        RECT 52.735 616.835 52.905 617.005 ;
        RECT 53.195 616.835 53.365 617.005 ;
        RECT 53.655 616.835 53.825 617.005 ;
        RECT 42.615 614.115 42.785 614.285 ;
        RECT 43.075 614.115 43.245 614.285 ;
        RECT 43.535 614.115 43.705 614.285 ;
        RECT 43.995 614.115 44.165 614.285 ;
        RECT 44.455 614.115 44.625 614.285 ;
        RECT 44.915 614.115 45.085 614.285 ;
        RECT 45.375 614.115 45.545 614.285 ;
        RECT 45.835 614.115 46.005 614.285 ;
        RECT 46.295 614.115 46.465 614.285 ;
        RECT 46.755 614.115 46.925 614.285 ;
        RECT 47.215 614.115 47.385 614.285 ;
        RECT 47.675 614.115 47.845 614.285 ;
        RECT 48.135 614.115 48.305 614.285 ;
        RECT 48.595 614.115 48.765 614.285 ;
        RECT 49.055 614.115 49.225 614.285 ;
        RECT 49.515 614.115 49.685 614.285 ;
        RECT 49.975 614.115 50.145 614.285 ;
        RECT 50.435 614.115 50.605 614.285 ;
        RECT 50.895 614.115 51.065 614.285 ;
        RECT 51.355 614.115 51.525 614.285 ;
        RECT 51.815 614.115 51.985 614.285 ;
        RECT 52.275 614.115 52.445 614.285 ;
        RECT 52.735 614.115 52.905 614.285 ;
        RECT 53.195 614.115 53.365 614.285 ;
        RECT 53.655 614.115 53.825 614.285 ;
        RECT 42.615 611.395 42.785 611.565 ;
        RECT 43.075 611.395 43.245 611.565 ;
        RECT 43.535 611.395 43.705 611.565 ;
        RECT 43.995 611.395 44.165 611.565 ;
        RECT 44.455 611.395 44.625 611.565 ;
        RECT 44.915 611.395 45.085 611.565 ;
        RECT 45.375 611.395 45.545 611.565 ;
        RECT 45.835 611.395 46.005 611.565 ;
        RECT 46.295 611.395 46.465 611.565 ;
        RECT 46.755 611.395 46.925 611.565 ;
        RECT 47.215 611.395 47.385 611.565 ;
        RECT 47.675 611.395 47.845 611.565 ;
        RECT 48.135 611.395 48.305 611.565 ;
        RECT 48.595 611.395 48.765 611.565 ;
        RECT 49.055 611.395 49.225 611.565 ;
        RECT 49.515 611.395 49.685 611.565 ;
        RECT 49.975 611.395 50.145 611.565 ;
        RECT 50.435 611.395 50.605 611.565 ;
        RECT 50.895 611.395 51.065 611.565 ;
        RECT 51.355 611.395 51.525 611.565 ;
        RECT 51.815 611.395 51.985 611.565 ;
        RECT 52.275 611.395 52.445 611.565 ;
        RECT 52.735 611.395 52.905 611.565 ;
        RECT 53.195 611.395 53.365 611.565 ;
        RECT 53.655 611.395 53.825 611.565 ;
        RECT 42.615 608.675 42.785 608.845 ;
        RECT 43.075 608.675 43.245 608.845 ;
        RECT 43.535 608.675 43.705 608.845 ;
        RECT 43.995 608.675 44.165 608.845 ;
        RECT 44.455 608.675 44.625 608.845 ;
        RECT 44.915 608.675 45.085 608.845 ;
        RECT 45.375 608.675 45.545 608.845 ;
        RECT 45.835 608.675 46.005 608.845 ;
        RECT 46.295 608.675 46.465 608.845 ;
        RECT 46.755 608.675 46.925 608.845 ;
        RECT 47.215 608.675 47.385 608.845 ;
        RECT 47.675 608.675 47.845 608.845 ;
        RECT 48.135 608.675 48.305 608.845 ;
        RECT 48.595 608.675 48.765 608.845 ;
        RECT 49.055 608.675 49.225 608.845 ;
        RECT 49.515 608.675 49.685 608.845 ;
        RECT 49.975 608.675 50.145 608.845 ;
        RECT 50.435 608.675 50.605 608.845 ;
        RECT 50.895 608.675 51.065 608.845 ;
        RECT 51.355 608.675 51.525 608.845 ;
        RECT 51.815 608.675 51.985 608.845 ;
        RECT 52.275 608.675 52.445 608.845 ;
        RECT 52.735 608.675 52.905 608.845 ;
        RECT 53.195 608.675 53.365 608.845 ;
        RECT 53.655 608.675 53.825 608.845 ;
        RECT 42.615 605.955 42.785 606.125 ;
        RECT 43.075 605.955 43.245 606.125 ;
        RECT 43.535 605.955 43.705 606.125 ;
        RECT 43.995 605.955 44.165 606.125 ;
        RECT 44.455 605.955 44.625 606.125 ;
        RECT 44.915 605.955 45.085 606.125 ;
        RECT 45.375 605.955 45.545 606.125 ;
        RECT 45.835 605.955 46.005 606.125 ;
        RECT 46.295 605.955 46.465 606.125 ;
        RECT 46.755 605.955 46.925 606.125 ;
        RECT 47.215 605.955 47.385 606.125 ;
        RECT 47.675 605.955 47.845 606.125 ;
        RECT 48.135 605.955 48.305 606.125 ;
        RECT 48.595 605.955 48.765 606.125 ;
        RECT 49.055 605.955 49.225 606.125 ;
        RECT 49.515 605.955 49.685 606.125 ;
        RECT 49.975 605.955 50.145 606.125 ;
        RECT 50.435 605.955 50.605 606.125 ;
        RECT 50.895 605.955 51.065 606.125 ;
        RECT 51.355 605.955 51.525 606.125 ;
        RECT 51.815 605.955 51.985 606.125 ;
        RECT 52.275 605.955 52.445 606.125 ;
        RECT 52.735 605.955 52.905 606.125 ;
        RECT 53.195 605.955 53.365 606.125 ;
        RECT 53.655 605.955 53.825 606.125 ;
        RECT 42.615 603.235 42.785 603.405 ;
        RECT 43.075 603.235 43.245 603.405 ;
        RECT 43.535 603.235 43.705 603.405 ;
        RECT 43.995 603.235 44.165 603.405 ;
        RECT 44.455 603.235 44.625 603.405 ;
        RECT 44.915 603.235 45.085 603.405 ;
        RECT 45.375 603.235 45.545 603.405 ;
        RECT 45.835 603.235 46.005 603.405 ;
        RECT 46.295 603.235 46.465 603.405 ;
        RECT 46.755 603.235 46.925 603.405 ;
        RECT 47.215 603.235 47.385 603.405 ;
        RECT 47.675 603.235 47.845 603.405 ;
        RECT 48.135 603.235 48.305 603.405 ;
        RECT 48.595 603.235 48.765 603.405 ;
        RECT 49.055 603.235 49.225 603.405 ;
        RECT 49.515 603.235 49.685 603.405 ;
        RECT 49.975 603.235 50.145 603.405 ;
        RECT 50.435 603.235 50.605 603.405 ;
        RECT 50.895 603.235 51.065 603.405 ;
        RECT 51.355 603.235 51.525 603.405 ;
        RECT 51.815 603.235 51.985 603.405 ;
        RECT 52.275 603.235 52.445 603.405 ;
        RECT 52.735 603.235 52.905 603.405 ;
        RECT 53.195 603.235 53.365 603.405 ;
        RECT 53.655 603.235 53.825 603.405 ;
        RECT 42.615 600.515 42.785 600.685 ;
        RECT 43.075 600.515 43.245 600.685 ;
        RECT 43.535 600.515 43.705 600.685 ;
        RECT 43.995 600.515 44.165 600.685 ;
        RECT 44.455 600.515 44.625 600.685 ;
        RECT 44.915 600.515 45.085 600.685 ;
        RECT 45.375 600.515 45.545 600.685 ;
        RECT 45.835 600.515 46.005 600.685 ;
        RECT 46.295 600.515 46.465 600.685 ;
        RECT 46.755 600.515 46.925 600.685 ;
        RECT 47.215 600.515 47.385 600.685 ;
        RECT 47.675 600.515 47.845 600.685 ;
        RECT 48.135 600.515 48.305 600.685 ;
        RECT 48.595 600.515 48.765 600.685 ;
        RECT 49.055 600.515 49.225 600.685 ;
        RECT 49.515 600.515 49.685 600.685 ;
        RECT 49.975 600.515 50.145 600.685 ;
        RECT 50.435 600.515 50.605 600.685 ;
        RECT 50.895 600.515 51.065 600.685 ;
        RECT 51.355 600.515 51.525 600.685 ;
        RECT 51.815 600.515 51.985 600.685 ;
        RECT 52.275 600.515 52.445 600.685 ;
        RECT 52.735 600.515 52.905 600.685 ;
        RECT 53.195 600.515 53.365 600.685 ;
        RECT 53.655 600.515 53.825 600.685 ;
        RECT 42.615 597.795 42.785 597.965 ;
        RECT 43.075 597.795 43.245 597.965 ;
        RECT 43.535 597.795 43.705 597.965 ;
        RECT 43.995 597.795 44.165 597.965 ;
        RECT 44.455 597.795 44.625 597.965 ;
        RECT 44.915 597.795 45.085 597.965 ;
        RECT 45.375 597.795 45.545 597.965 ;
        RECT 45.835 597.795 46.005 597.965 ;
        RECT 46.295 597.795 46.465 597.965 ;
        RECT 46.755 597.795 46.925 597.965 ;
        RECT 47.215 597.795 47.385 597.965 ;
        RECT 47.675 597.795 47.845 597.965 ;
        RECT 48.135 597.795 48.305 597.965 ;
        RECT 48.595 597.795 48.765 597.965 ;
        RECT 49.055 597.795 49.225 597.965 ;
        RECT 49.515 597.795 49.685 597.965 ;
        RECT 49.975 597.795 50.145 597.965 ;
        RECT 50.435 597.795 50.605 597.965 ;
        RECT 50.895 597.795 51.065 597.965 ;
        RECT 51.355 597.795 51.525 597.965 ;
        RECT 51.815 597.795 51.985 597.965 ;
        RECT 52.275 597.795 52.445 597.965 ;
        RECT 52.735 597.795 52.905 597.965 ;
        RECT 53.195 597.795 53.365 597.965 ;
        RECT 53.655 597.795 53.825 597.965 ;
        RECT 42.615 595.075 42.785 595.245 ;
        RECT 43.075 595.075 43.245 595.245 ;
        RECT 43.535 595.075 43.705 595.245 ;
        RECT 43.995 595.075 44.165 595.245 ;
        RECT 44.455 595.075 44.625 595.245 ;
        RECT 44.915 595.075 45.085 595.245 ;
        RECT 45.375 595.075 45.545 595.245 ;
        RECT 45.835 595.075 46.005 595.245 ;
        RECT 46.295 595.075 46.465 595.245 ;
        RECT 46.755 595.075 46.925 595.245 ;
        RECT 47.215 595.075 47.385 595.245 ;
        RECT 47.675 595.075 47.845 595.245 ;
        RECT 48.135 595.075 48.305 595.245 ;
        RECT 48.595 595.075 48.765 595.245 ;
        RECT 49.055 595.075 49.225 595.245 ;
        RECT 49.515 595.075 49.685 595.245 ;
        RECT 49.975 595.075 50.145 595.245 ;
        RECT 50.435 595.075 50.605 595.245 ;
        RECT 50.895 595.075 51.065 595.245 ;
        RECT 51.355 595.075 51.525 595.245 ;
        RECT 51.815 595.075 51.985 595.245 ;
        RECT 52.275 595.075 52.445 595.245 ;
        RECT 52.735 595.075 52.905 595.245 ;
        RECT 53.195 595.075 53.365 595.245 ;
        RECT 53.655 595.075 53.825 595.245 ;
        RECT 42.615 592.355 42.785 592.525 ;
        RECT 43.075 592.355 43.245 592.525 ;
        RECT 43.535 592.355 43.705 592.525 ;
        RECT 43.995 592.355 44.165 592.525 ;
        RECT 44.455 592.355 44.625 592.525 ;
        RECT 44.915 592.355 45.085 592.525 ;
        RECT 45.375 592.355 45.545 592.525 ;
        RECT 45.835 592.355 46.005 592.525 ;
        RECT 46.295 592.355 46.465 592.525 ;
        RECT 46.755 592.355 46.925 592.525 ;
        RECT 47.215 592.355 47.385 592.525 ;
        RECT 47.675 592.355 47.845 592.525 ;
        RECT 48.135 592.355 48.305 592.525 ;
        RECT 48.595 592.355 48.765 592.525 ;
        RECT 49.055 592.355 49.225 592.525 ;
        RECT 49.515 592.355 49.685 592.525 ;
        RECT 49.975 592.355 50.145 592.525 ;
        RECT 50.435 592.355 50.605 592.525 ;
        RECT 50.895 592.355 51.065 592.525 ;
        RECT 51.355 592.355 51.525 592.525 ;
        RECT 51.815 592.355 51.985 592.525 ;
        RECT 52.275 592.355 52.445 592.525 ;
        RECT 52.735 592.355 52.905 592.525 ;
        RECT 53.195 592.355 53.365 592.525 ;
        RECT 53.655 592.355 53.825 592.525 ;
        RECT 42.615 589.635 42.785 589.805 ;
        RECT 43.075 589.635 43.245 589.805 ;
        RECT 43.535 589.635 43.705 589.805 ;
        RECT 43.995 589.635 44.165 589.805 ;
        RECT 44.455 589.635 44.625 589.805 ;
        RECT 44.915 589.635 45.085 589.805 ;
        RECT 45.375 589.635 45.545 589.805 ;
        RECT 45.835 589.635 46.005 589.805 ;
        RECT 46.295 589.635 46.465 589.805 ;
        RECT 46.755 589.635 46.925 589.805 ;
        RECT 47.215 589.635 47.385 589.805 ;
        RECT 47.675 589.635 47.845 589.805 ;
        RECT 48.135 589.635 48.305 589.805 ;
        RECT 48.595 589.635 48.765 589.805 ;
        RECT 49.055 589.635 49.225 589.805 ;
        RECT 49.515 589.635 49.685 589.805 ;
        RECT 49.975 589.635 50.145 589.805 ;
        RECT 50.435 589.635 50.605 589.805 ;
        RECT 50.895 589.635 51.065 589.805 ;
        RECT 51.355 589.635 51.525 589.805 ;
        RECT 51.815 589.635 51.985 589.805 ;
        RECT 52.275 589.635 52.445 589.805 ;
        RECT 52.735 589.635 52.905 589.805 ;
        RECT 53.195 589.635 53.365 589.805 ;
        RECT 53.655 589.635 53.825 589.805 ;
        RECT 42.615 586.915 42.785 587.085 ;
        RECT 43.075 586.915 43.245 587.085 ;
        RECT 43.535 586.915 43.705 587.085 ;
        RECT 43.995 586.915 44.165 587.085 ;
        RECT 44.455 586.915 44.625 587.085 ;
        RECT 44.915 586.915 45.085 587.085 ;
        RECT 45.375 586.915 45.545 587.085 ;
        RECT 45.835 586.915 46.005 587.085 ;
        RECT 46.295 586.915 46.465 587.085 ;
        RECT 46.755 586.915 46.925 587.085 ;
        RECT 47.215 586.915 47.385 587.085 ;
        RECT 47.675 586.915 47.845 587.085 ;
        RECT 48.135 586.915 48.305 587.085 ;
        RECT 48.595 586.915 48.765 587.085 ;
        RECT 49.055 586.915 49.225 587.085 ;
        RECT 49.515 586.915 49.685 587.085 ;
        RECT 49.975 586.915 50.145 587.085 ;
        RECT 50.435 586.915 50.605 587.085 ;
        RECT 50.895 586.915 51.065 587.085 ;
        RECT 51.355 586.915 51.525 587.085 ;
        RECT 51.815 586.915 51.985 587.085 ;
        RECT 52.275 586.915 52.445 587.085 ;
        RECT 52.735 586.915 52.905 587.085 ;
        RECT 53.195 586.915 53.365 587.085 ;
        RECT 53.655 586.915 53.825 587.085 ;
        RECT 42.615 584.195 42.785 584.365 ;
        RECT 43.075 584.195 43.245 584.365 ;
        RECT 43.535 584.195 43.705 584.365 ;
        RECT 43.995 584.195 44.165 584.365 ;
        RECT 44.455 584.195 44.625 584.365 ;
        RECT 44.915 584.195 45.085 584.365 ;
        RECT 45.375 584.195 45.545 584.365 ;
        RECT 45.835 584.195 46.005 584.365 ;
        RECT 46.295 584.195 46.465 584.365 ;
        RECT 46.755 584.195 46.925 584.365 ;
        RECT 47.215 584.195 47.385 584.365 ;
        RECT 47.675 584.195 47.845 584.365 ;
        RECT 48.135 584.195 48.305 584.365 ;
        RECT 48.595 584.195 48.765 584.365 ;
        RECT 49.055 584.195 49.225 584.365 ;
        RECT 49.515 584.195 49.685 584.365 ;
        RECT 49.975 584.195 50.145 584.365 ;
        RECT 50.435 584.195 50.605 584.365 ;
        RECT 50.895 584.195 51.065 584.365 ;
        RECT 51.355 584.195 51.525 584.365 ;
        RECT 51.815 584.195 51.985 584.365 ;
        RECT 52.275 584.195 52.445 584.365 ;
        RECT 52.735 584.195 52.905 584.365 ;
        RECT 53.195 584.195 53.365 584.365 ;
        RECT 53.655 584.195 53.825 584.365 ;
        RECT 42.615 581.475 42.785 581.645 ;
        RECT 43.075 581.475 43.245 581.645 ;
        RECT 43.535 581.475 43.705 581.645 ;
        RECT 43.995 581.475 44.165 581.645 ;
        RECT 44.455 581.475 44.625 581.645 ;
        RECT 44.915 581.475 45.085 581.645 ;
        RECT 45.375 581.475 45.545 581.645 ;
        RECT 45.835 581.475 46.005 581.645 ;
        RECT 46.295 581.475 46.465 581.645 ;
        RECT 46.755 581.475 46.925 581.645 ;
        RECT 47.215 581.475 47.385 581.645 ;
        RECT 47.675 581.475 47.845 581.645 ;
        RECT 48.135 581.475 48.305 581.645 ;
        RECT 48.595 581.475 48.765 581.645 ;
        RECT 49.055 581.475 49.225 581.645 ;
        RECT 49.515 581.475 49.685 581.645 ;
        RECT 49.975 581.475 50.145 581.645 ;
        RECT 50.435 581.475 50.605 581.645 ;
        RECT 50.895 581.475 51.065 581.645 ;
        RECT 51.355 581.475 51.525 581.645 ;
        RECT 51.815 581.475 51.985 581.645 ;
        RECT 52.275 581.475 52.445 581.645 ;
        RECT 52.735 581.475 52.905 581.645 ;
        RECT 53.195 581.475 53.365 581.645 ;
        RECT 53.655 581.475 53.825 581.645 ;
        RECT 42.615 578.755 42.785 578.925 ;
        RECT 43.075 578.755 43.245 578.925 ;
        RECT 43.535 578.755 43.705 578.925 ;
        RECT 43.995 578.755 44.165 578.925 ;
        RECT 44.455 578.755 44.625 578.925 ;
        RECT 44.915 578.755 45.085 578.925 ;
        RECT 45.375 578.755 45.545 578.925 ;
        RECT 45.835 578.755 46.005 578.925 ;
        RECT 46.295 578.755 46.465 578.925 ;
        RECT 46.755 578.755 46.925 578.925 ;
        RECT 47.215 578.755 47.385 578.925 ;
        RECT 47.675 578.755 47.845 578.925 ;
        RECT 48.135 578.755 48.305 578.925 ;
        RECT 48.595 578.755 48.765 578.925 ;
        RECT 49.055 578.755 49.225 578.925 ;
        RECT 49.515 578.755 49.685 578.925 ;
        RECT 49.975 578.755 50.145 578.925 ;
        RECT 50.435 578.755 50.605 578.925 ;
        RECT 50.895 578.755 51.065 578.925 ;
        RECT 51.355 578.755 51.525 578.925 ;
        RECT 51.815 578.755 51.985 578.925 ;
        RECT 52.275 578.755 52.445 578.925 ;
        RECT 52.735 578.755 52.905 578.925 ;
        RECT 53.195 578.755 53.365 578.925 ;
        RECT 53.655 578.755 53.825 578.925 ;
        RECT 42.615 576.035 42.785 576.205 ;
        RECT 43.075 576.035 43.245 576.205 ;
        RECT 43.535 576.035 43.705 576.205 ;
        RECT 43.995 576.035 44.165 576.205 ;
        RECT 44.455 576.035 44.625 576.205 ;
        RECT 44.915 576.035 45.085 576.205 ;
        RECT 45.375 576.035 45.545 576.205 ;
        RECT 45.835 576.035 46.005 576.205 ;
        RECT 46.295 576.035 46.465 576.205 ;
        RECT 46.755 576.035 46.925 576.205 ;
        RECT 47.215 576.035 47.385 576.205 ;
        RECT 47.675 576.035 47.845 576.205 ;
        RECT 48.135 576.035 48.305 576.205 ;
        RECT 48.595 576.035 48.765 576.205 ;
        RECT 49.055 576.035 49.225 576.205 ;
        RECT 49.515 576.035 49.685 576.205 ;
        RECT 49.975 576.035 50.145 576.205 ;
        RECT 50.435 576.035 50.605 576.205 ;
        RECT 50.895 576.035 51.065 576.205 ;
        RECT 51.355 576.035 51.525 576.205 ;
        RECT 51.815 576.035 51.985 576.205 ;
        RECT 52.275 576.035 52.445 576.205 ;
        RECT 52.735 576.035 52.905 576.205 ;
        RECT 53.195 576.035 53.365 576.205 ;
        RECT 53.655 576.035 53.825 576.205 ;
        RECT 42.615 573.315 42.785 573.485 ;
        RECT 43.075 573.315 43.245 573.485 ;
        RECT 43.535 573.315 43.705 573.485 ;
        RECT 43.995 573.315 44.165 573.485 ;
        RECT 44.455 573.315 44.625 573.485 ;
        RECT 44.915 573.315 45.085 573.485 ;
        RECT 45.375 573.315 45.545 573.485 ;
        RECT 45.835 573.315 46.005 573.485 ;
        RECT 46.295 573.315 46.465 573.485 ;
        RECT 46.755 573.315 46.925 573.485 ;
        RECT 47.215 573.315 47.385 573.485 ;
        RECT 47.675 573.315 47.845 573.485 ;
        RECT 48.135 573.315 48.305 573.485 ;
        RECT 48.595 573.315 48.765 573.485 ;
        RECT 49.055 573.315 49.225 573.485 ;
        RECT 49.515 573.315 49.685 573.485 ;
        RECT 49.975 573.315 50.145 573.485 ;
        RECT 50.435 573.315 50.605 573.485 ;
        RECT 50.895 573.315 51.065 573.485 ;
        RECT 51.355 573.315 51.525 573.485 ;
        RECT 51.815 573.315 51.985 573.485 ;
        RECT 52.275 573.315 52.445 573.485 ;
        RECT 52.735 573.315 52.905 573.485 ;
        RECT 53.195 573.315 53.365 573.485 ;
        RECT 53.655 573.315 53.825 573.485 ;
        RECT 42.615 570.595 42.785 570.765 ;
        RECT 43.075 570.595 43.245 570.765 ;
        RECT 43.535 570.595 43.705 570.765 ;
        RECT 43.995 570.595 44.165 570.765 ;
        RECT 44.455 570.595 44.625 570.765 ;
        RECT 44.915 570.595 45.085 570.765 ;
        RECT 45.375 570.595 45.545 570.765 ;
        RECT 45.835 570.595 46.005 570.765 ;
        RECT 46.295 570.595 46.465 570.765 ;
        RECT 46.755 570.595 46.925 570.765 ;
        RECT 47.215 570.595 47.385 570.765 ;
        RECT 47.675 570.595 47.845 570.765 ;
        RECT 48.135 570.595 48.305 570.765 ;
        RECT 48.595 570.595 48.765 570.765 ;
        RECT 49.055 570.595 49.225 570.765 ;
        RECT 49.515 570.595 49.685 570.765 ;
        RECT 49.975 570.595 50.145 570.765 ;
        RECT 50.435 570.595 50.605 570.765 ;
        RECT 50.895 570.595 51.065 570.765 ;
        RECT 51.355 570.595 51.525 570.765 ;
        RECT 51.815 570.595 51.985 570.765 ;
        RECT 52.275 570.595 52.445 570.765 ;
        RECT 52.735 570.595 52.905 570.765 ;
        RECT 53.195 570.595 53.365 570.765 ;
        RECT 53.655 570.595 53.825 570.765 ;
        RECT 42.615 567.875 42.785 568.045 ;
        RECT 43.075 567.875 43.245 568.045 ;
        RECT 43.535 567.875 43.705 568.045 ;
        RECT 43.995 567.875 44.165 568.045 ;
        RECT 44.455 567.875 44.625 568.045 ;
        RECT 44.915 567.875 45.085 568.045 ;
        RECT 45.375 567.875 45.545 568.045 ;
        RECT 45.835 567.875 46.005 568.045 ;
        RECT 46.295 567.875 46.465 568.045 ;
        RECT 46.755 567.875 46.925 568.045 ;
        RECT 47.215 567.875 47.385 568.045 ;
        RECT 47.675 567.875 47.845 568.045 ;
        RECT 48.135 567.875 48.305 568.045 ;
        RECT 48.595 567.875 48.765 568.045 ;
        RECT 49.055 567.875 49.225 568.045 ;
        RECT 49.515 567.875 49.685 568.045 ;
        RECT 49.975 567.875 50.145 568.045 ;
        RECT 50.435 567.875 50.605 568.045 ;
        RECT 50.895 567.875 51.065 568.045 ;
        RECT 51.355 567.875 51.525 568.045 ;
        RECT 51.815 567.875 51.985 568.045 ;
        RECT 52.275 567.875 52.445 568.045 ;
        RECT 52.735 567.875 52.905 568.045 ;
        RECT 53.195 567.875 53.365 568.045 ;
        RECT 53.655 567.875 53.825 568.045 ;
        RECT 42.615 565.155 42.785 565.325 ;
        RECT 43.075 565.155 43.245 565.325 ;
        RECT 43.535 565.155 43.705 565.325 ;
        RECT 43.995 565.155 44.165 565.325 ;
        RECT 44.455 565.155 44.625 565.325 ;
        RECT 44.915 565.155 45.085 565.325 ;
        RECT 45.375 565.155 45.545 565.325 ;
        RECT 45.835 565.155 46.005 565.325 ;
        RECT 46.295 565.155 46.465 565.325 ;
        RECT 46.755 565.155 46.925 565.325 ;
        RECT 47.215 565.155 47.385 565.325 ;
        RECT 47.675 565.155 47.845 565.325 ;
        RECT 48.135 565.155 48.305 565.325 ;
        RECT 48.595 565.155 48.765 565.325 ;
        RECT 49.055 565.155 49.225 565.325 ;
        RECT 49.515 565.155 49.685 565.325 ;
        RECT 49.975 565.155 50.145 565.325 ;
        RECT 50.435 565.155 50.605 565.325 ;
        RECT 50.895 565.155 51.065 565.325 ;
        RECT 51.355 565.155 51.525 565.325 ;
        RECT 51.815 565.155 51.985 565.325 ;
        RECT 52.275 565.155 52.445 565.325 ;
        RECT 52.735 565.155 52.905 565.325 ;
        RECT 53.195 565.155 53.365 565.325 ;
        RECT 53.655 565.155 53.825 565.325 ;
        RECT 42.615 562.435 42.785 562.605 ;
        RECT 43.075 562.435 43.245 562.605 ;
        RECT 43.535 562.435 43.705 562.605 ;
        RECT 43.995 562.435 44.165 562.605 ;
        RECT 44.455 562.435 44.625 562.605 ;
        RECT 44.915 562.435 45.085 562.605 ;
        RECT 45.375 562.435 45.545 562.605 ;
        RECT 45.835 562.435 46.005 562.605 ;
        RECT 46.295 562.435 46.465 562.605 ;
        RECT 46.755 562.435 46.925 562.605 ;
        RECT 47.215 562.435 47.385 562.605 ;
        RECT 47.675 562.435 47.845 562.605 ;
        RECT 48.135 562.435 48.305 562.605 ;
        RECT 48.595 562.435 48.765 562.605 ;
        RECT 49.055 562.435 49.225 562.605 ;
        RECT 49.515 562.435 49.685 562.605 ;
        RECT 49.975 562.435 50.145 562.605 ;
        RECT 50.435 562.435 50.605 562.605 ;
        RECT 50.895 562.435 51.065 562.605 ;
        RECT 51.355 562.435 51.525 562.605 ;
        RECT 51.815 562.435 51.985 562.605 ;
        RECT 52.275 562.435 52.445 562.605 ;
        RECT 52.735 562.435 52.905 562.605 ;
        RECT 53.195 562.435 53.365 562.605 ;
        RECT 53.655 562.435 53.825 562.605 ;
        RECT 42.615 559.715 42.785 559.885 ;
        RECT 43.075 559.715 43.245 559.885 ;
        RECT 43.535 559.715 43.705 559.885 ;
        RECT 43.995 559.715 44.165 559.885 ;
        RECT 44.455 559.715 44.625 559.885 ;
        RECT 44.915 559.715 45.085 559.885 ;
        RECT 45.375 559.715 45.545 559.885 ;
        RECT 45.835 559.715 46.005 559.885 ;
        RECT 46.295 559.715 46.465 559.885 ;
        RECT 46.755 559.715 46.925 559.885 ;
        RECT 47.215 559.715 47.385 559.885 ;
        RECT 47.675 559.715 47.845 559.885 ;
        RECT 48.135 559.715 48.305 559.885 ;
        RECT 48.595 559.715 48.765 559.885 ;
        RECT 49.055 559.715 49.225 559.885 ;
        RECT 49.515 559.715 49.685 559.885 ;
        RECT 49.975 559.715 50.145 559.885 ;
        RECT 50.435 559.715 50.605 559.885 ;
        RECT 50.895 559.715 51.065 559.885 ;
        RECT 51.355 559.715 51.525 559.885 ;
        RECT 51.815 559.715 51.985 559.885 ;
        RECT 52.275 559.715 52.445 559.885 ;
        RECT 52.735 559.715 52.905 559.885 ;
        RECT 53.195 559.715 53.365 559.885 ;
        RECT 53.655 559.715 53.825 559.885 ;
        RECT 42.615 556.995 42.785 557.165 ;
        RECT 43.075 556.995 43.245 557.165 ;
        RECT 43.535 556.995 43.705 557.165 ;
        RECT 43.995 556.995 44.165 557.165 ;
        RECT 44.455 556.995 44.625 557.165 ;
        RECT 44.915 556.995 45.085 557.165 ;
        RECT 45.375 556.995 45.545 557.165 ;
        RECT 45.835 556.995 46.005 557.165 ;
        RECT 46.295 556.995 46.465 557.165 ;
        RECT 46.755 556.995 46.925 557.165 ;
        RECT 47.215 556.995 47.385 557.165 ;
        RECT 47.675 556.995 47.845 557.165 ;
        RECT 48.135 556.995 48.305 557.165 ;
        RECT 48.595 556.995 48.765 557.165 ;
        RECT 49.055 556.995 49.225 557.165 ;
        RECT 49.515 556.995 49.685 557.165 ;
        RECT 49.975 556.995 50.145 557.165 ;
        RECT 50.435 556.995 50.605 557.165 ;
        RECT 50.895 556.995 51.065 557.165 ;
        RECT 51.355 556.995 51.525 557.165 ;
        RECT 51.815 556.995 51.985 557.165 ;
        RECT 52.275 556.995 52.445 557.165 ;
        RECT 52.735 556.995 52.905 557.165 ;
        RECT 53.195 556.995 53.365 557.165 ;
        RECT 53.655 556.995 53.825 557.165 ;
        RECT 42.615 554.275 42.785 554.445 ;
        RECT 43.075 554.275 43.245 554.445 ;
        RECT 43.535 554.275 43.705 554.445 ;
        RECT 43.995 554.275 44.165 554.445 ;
        RECT 44.455 554.275 44.625 554.445 ;
        RECT 44.915 554.275 45.085 554.445 ;
        RECT 45.375 554.275 45.545 554.445 ;
        RECT 45.835 554.275 46.005 554.445 ;
        RECT 46.295 554.275 46.465 554.445 ;
        RECT 46.755 554.275 46.925 554.445 ;
        RECT 47.215 554.275 47.385 554.445 ;
        RECT 47.675 554.275 47.845 554.445 ;
        RECT 48.135 554.275 48.305 554.445 ;
        RECT 48.595 554.275 48.765 554.445 ;
        RECT 49.055 554.275 49.225 554.445 ;
        RECT 49.515 554.275 49.685 554.445 ;
        RECT 49.975 554.275 50.145 554.445 ;
        RECT 50.435 554.275 50.605 554.445 ;
        RECT 50.895 554.275 51.065 554.445 ;
        RECT 51.355 554.275 51.525 554.445 ;
        RECT 51.815 554.275 51.985 554.445 ;
        RECT 52.275 554.275 52.445 554.445 ;
        RECT 52.735 554.275 52.905 554.445 ;
        RECT 53.195 554.275 53.365 554.445 ;
        RECT 53.655 554.275 53.825 554.445 ;
        RECT 42.615 551.555 42.785 551.725 ;
        RECT 43.075 551.555 43.245 551.725 ;
        RECT 43.535 551.555 43.705 551.725 ;
        RECT 43.995 551.555 44.165 551.725 ;
        RECT 44.455 551.555 44.625 551.725 ;
        RECT 44.915 551.555 45.085 551.725 ;
        RECT 45.375 551.555 45.545 551.725 ;
        RECT 45.835 551.555 46.005 551.725 ;
        RECT 46.295 551.555 46.465 551.725 ;
        RECT 46.755 551.555 46.925 551.725 ;
        RECT 47.215 551.555 47.385 551.725 ;
        RECT 47.675 551.555 47.845 551.725 ;
        RECT 48.135 551.555 48.305 551.725 ;
        RECT 48.595 551.555 48.765 551.725 ;
        RECT 49.055 551.555 49.225 551.725 ;
        RECT 49.515 551.555 49.685 551.725 ;
        RECT 49.975 551.555 50.145 551.725 ;
        RECT 50.435 551.555 50.605 551.725 ;
        RECT 50.895 551.555 51.065 551.725 ;
        RECT 51.355 551.555 51.525 551.725 ;
        RECT 51.815 551.555 51.985 551.725 ;
        RECT 52.275 551.555 52.445 551.725 ;
        RECT 52.735 551.555 52.905 551.725 ;
        RECT 53.195 551.555 53.365 551.725 ;
        RECT 53.655 551.555 53.825 551.725 ;
        RECT 42.615 548.835 42.785 549.005 ;
        RECT 43.075 548.835 43.245 549.005 ;
        RECT 43.535 548.835 43.705 549.005 ;
        RECT 43.995 548.835 44.165 549.005 ;
        RECT 44.455 548.835 44.625 549.005 ;
        RECT 44.915 548.835 45.085 549.005 ;
        RECT 45.375 548.835 45.545 549.005 ;
        RECT 45.835 548.835 46.005 549.005 ;
        RECT 46.295 548.835 46.465 549.005 ;
        RECT 46.755 548.835 46.925 549.005 ;
        RECT 47.215 548.835 47.385 549.005 ;
        RECT 47.675 548.835 47.845 549.005 ;
        RECT 48.135 548.835 48.305 549.005 ;
        RECT 48.595 548.835 48.765 549.005 ;
        RECT 49.055 548.835 49.225 549.005 ;
        RECT 49.515 548.835 49.685 549.005 ;
        RECT 49.975 548.835 50.145 549.005 ;
        RECT 50.435 548.835 50.605 549.005 ;
        RECT 50.895 548.835 51.065 549.005 ;
        RECT 51.355 548.835 51.525 549.005 ;
        RECT 51.815 548.835 51.985 549.005 ;
        RECT 52.275 548.835 52.445 549.005 ;
        RECT 52.735 548.835 52.905 549.005 ;
        RECT 53.195 548.835 53.365 549.005 ;
        RECT 53.655 548.835 53.825 549.005 ;
        RECT 42.615 546.115 42.785 546.285 ;
        RECT 43.075 546.115 43.245 546.285 ;
        RECT 43.535 546.115 43.705 546.285 ;
        RECT 43.995 546.115 44.165 546.285 ;
        RECT 44.455 546.115 44.625 546.285 ;
        RECT 44.915 546.115 45.085 546.285 ;
        RECT 45.375 546.115 45.545 546.285 ;
        RECT 45.835 546.115 46.005 546.285 ;
        RECT 46.295 546.115 46.465 546.285 ;
        RECT 46.755 546.115 46.925 546.285 ;
        RECT 47.215 546.115 47.385 546.285 ;
        RECT 47.675 546.115 47.845 546.285 ;
        RECT 48.135 546.115 48.305 546.285 ;
        RECT 48.595 546.115 48.765 546.285 ;
        RECT 49.055 546.115 49.225 546.285 ;
        RECT 49.515 546.115 49.685 546.285 ;
        RECT 49.975 546.115 50.145 546.285 ;
        RECT 50.435 546.115 50.605 546.285 ;
        RECT 50.895 546.115 51.065 546.285 ;
        RECT 51.355 546.115 51.525 546.285 ;
        RECT 51.815 546.115 51.985 546.285 ;
        RECT 52.275 546.115 52.445 546.285 ;
        RECT 52.735 546.115 52.905 546.285 ;
        RECT 53.195 546.115 53.365 546.285 ;
        RECT 53.655 546.115 53.825 546.285 ;
        RECT 42.615 543.395 42.785 543.565 ;
        RECT 43.075 543.395 43.245 543.565 ;
        RECT 43.535 543.395 43.705 543.565 ;
        RECT 43.995 543.395 44.165 543.565 ;
        RECT 44.455 543.395 44.625 543.565 ;
        RECT 44.915 543.395 45.085 543.565 ;
        RECT 45.375 543.395 45.545 543.565 ;
        RECT 45.835 543.395 46.005 543.565 ;
        RECT 46.295 543.395 46.465 543.565 ;
        RECT 46.755 543.395 46.925 543.565 ;
        RECT 47.215 543.395 47.385 543.565 ;
        RECT 47.675 543.395 47.845 543.565 ;
        RECT 48.135 543.395 48.305 543.565 ;
        RECT 48.595 543.395 48.765 543.565 ;
        RECT 49.055 543.395 49.225 543.565 ;
        RECT 49.515 543.395 49.685 543.565 ;
        RECT 49.975 543.395 50.145 543.565 ;
        RECT 50.435 543.395 50.605 543.565 ;
        RECT 50.895 543.395 51.065 543.565 ;
        RECT 51.355 543.395 51.525 543.565 ;
        RECT 51.815 543.395 51.985 543.565 ;
        RECT 52.275 543.395 52.445 543.565 ;
        RECT 52.735 543.395 52.905 543.565 ;
        RECT 53.195 543.395 53.365 543.565 ;
        RECT 53.655 543.395 53.825 543.565 ;
        RECT 42.615 540.675 42.785 540.845 ;
        RECT 43.075 540.675 43.245 540.845 ;
        RECT 43.535 540.675 43.705 540.845 ;
        RECT 43.995 540.675 44.165 540.845 ;
        RECT 44.455 540.675 44.625 540.845 ;
        RECT 44.915 540.675 45.085 540.845 ;
        RECT 45.375 540.675 45.545 540.845 ;
        RECT 45.835 540.675 46.005 540.845 ;
        RECT 46.295 540.675 46.465 540.845 ;
        RECT 46.755 540.675 46.925 540.845 ;
        RECT 47.215 540.675 47.385 540.845 ;
        RECT 47.675 540.675 47.845 540.845 ;
        RECT 48.135 540.675 48.305 540.845 ;
        RECT 48.595 540.675 48.765 540.845 ;
        RECT 49.055 540.675 49.225 540.845 ;
        RECT 49.515 540.675 49.685 540.845 ;
        RECT 49.975 540.675 50.145 540.845 ;
        RECT 50.435 540.675 50.605 540.845 ;
        RECT 50.895 540.675 51.065 540.845 ;
        RECT 51.355 540.675 51.525 540.845 ;
        RECT 51.815 540.675 51.985 540.845 ;
        RECT 52.275 540.675 52.445 540.845 ;
        RECT 52.735 540.675 52.905 540.845 ;
        RECT 53.195 540.675 53.365 540.845 ;
        RECT 53.655 540.675 53.825 540.845 ;
        RECT 42.615 537.955 42.785 538.125 ;
        RECT 43.075 537.955 43.245 538.125 ;
        RECT 43.535 537.955 43.705 538.125 ;
        RECT 43.995 537.955 44.165 538.125 ;
        RECT 44.455 537.955 44.625 538.125 ;
        RECT 44.915 537.955 45.085 538.125 ;
        RECT 45.375 537.955 45.545 538.125 ;
        RECT 45.835 537.955 46.005 538.125 ;
        RECT 46.295 537.955 46.465 538.125 ;
        RECT 46.755 537.955 46.925 538.125 ;
        RECT 47.215 537.955 47.385 538.125 ;
        RECT 47.675 537.955 47.845 538.125 ;
        RECT 48.135 537.955 48.305 538.125 ;
        RECT 48.595 537.955 48.765 538.125 ;
        RECT 49.055 537.955 49.225 538.125 ;
        RECT 49.515 537.955 49.685 538.125 ;
        RECT 49.975 537.955 50.145 538.125 ;
        RECT 50.435 537.955 50.605 538.125 ;
        RECT 50.895 537.955 51.065 538.125 ;
        RECT 51.355 537.955 51.525 538.125 ;
        RECT 51.815 537.955 51.985 538.125 ;
        RECT 52.275 537.955 52.445 538.125 ;
        RECT 52.735 537.955 52.905 538.125 ;
        RECT 53.195 537.955 53.365 538.125 ;
        RECT 53.655 537.955 53.825 538.125 ;
        RECT 42.615 535.235 42.785 535.405 ;
        RECT 43.075 535.235 43.245 535.405 ;
        RECT 43.535 535.235 43.705 535.405 ;
        RECT 43.995 535.235 44.165 535.405 ;
        RECT 44.455 535.235 44.625 535.405 ;
        RECT 44.915 535.235 45.085 535.405 ;
        RECT 45.375 535.235 45.545 535.405 ;
        RECT 45.835 535.235 46.005 535.405 ;
        RECT 46.295 535.235 46.465 535.405 ;
        RECT 46.755 535.235 46.925 535.405 ;
        RECT 47.215 535.235 47.385 535.405 ;
        RECT 47.675 535.235 47.845 535.405 ;
        RECT 48.135 535.235 48.305 535.405 ;
        RECT 48.595 535.235 48.765 535.405 ;
        RECT 49.055 535.235 49.225 535.405 ;
        RECT 49.515 535.235 49.685 535.405 ;
        RECT 49.975 535.235 50.145 535.405 ;
        RECT 50.435 535.235 50.605 535.405 ;
        RECT 50.895 535.235 51.065 535.405 ;
        RECT 51.355 535.235 51.525 535.405 ;
        RECT 51.815 535.235 51.985 535.405 ;
        RECT 52.275 535.235 52.445 535.405 ;
        RECT 52.735 535.235 52.905 535.405 ;
        RECT 53.195 535.235 53.365 535.405 ;
        RECT 53.655 535.235 53.825 535.405 ;
        RECT 42.615 532.515 42.785 532.685 ;
        RECT 43.075 532.515 43.245 532.685 ;
        RECT 43.535 532.515 43.705 532.685 ;
        RECT 43.995 532.515 44.165 532.685 ;
        RECT 44.455 532.515 44.625 532.685 ;
        RECT 44.915 532.515 45.085 532.685 ;
        RECT 45.375 532.515 45.545 532.685 ;
        RECT 45.835 532.515 46.005 532.685 ;
        RECT 46.295 532.515 46.465 532.685 ;
        RECT 46.755 532.515 46.925 532.685 ;
        RECT 47.215 532.515 47.385 532.685 ;
        RECT 47.675 532.515 47.845 532.685 ;
        RECT 48.135 532.515 48.305 532.685 ;
        RECT 48.595 532.515 48.765 532.685 ;
        RECT 49.055 532.515 49.225 532.685 ;
        RECT 49.515 532.515 49.685 532.685 ;
        RECT 49.975 532.515 50.145 532.685 ;
        RECT 50.435 532.515 50.605 532.685 ;
        RECT 50.895 532.515 51.065 532.685 ;
        RECT 51.355 532.515 51.525 532.685 ;
        RECT 51.815 532.515 51.985 532.685 ;
        RECT 52.275 532.515 52.445 532.685 ;
        RECT 52.735 532.515 52.905 532.685 ;
        RECT 53.195 532.515 53.365 532.685 ;
        RECT 53.655 532.515 53.825 532.685 ;
        RECT 42.615 529.795 42.785 529.965 ;
        RECT 43.075 529.795 43.245 529.965 ;
        RECT 43.535 529.795 43.705 529.965 ;
        RECT 43.995 529.795 44.165 529.965 ;
        RECT 44.455 529.795 44.625 529.965 ;
        RECT 44.915 529.795 45.085 529.965 ;
        RECT 45.375 529.795 45.545 529.965 ;
        RECT 45.835 529.795 46.005 529.965 ;
        RECT 46.295 529.795 46.465 529.965 ;
        RECT 46.755 529.795 46.925 529.965 ;
        RECT 47.215 529.795 47.385 529.965 ;
        RECT 47.675 529.795 47.845 529.965 ;
        RECT 48.135 529.795 48.305 529.965 ;
        RECT 48.595 529.795 48.765 529.965 ;
        RECT 49.055 529.795 49.225 529.965 ;
        RECT 49.515 529.795 49.685 529.965 ;
        RECT 49.975 529.795 50.145 529.965 ;
        RECT 50.435 529.795 50.605 529.965 ;
        RECT 50.895 529.795 51.065 529.965 ;
        RECT 51.355 529.795 51.525 529.965 ;
        RECT 51.815 529.795 51.985 529.965 ;
        RECT 52.275 529.795 52.445 529.965 ;
        RECT 52.735 529.795 52.905 529.965 ;
        RECT 53.195 529.795 53.365 529.965 ;
        RECT 53.655 529.795 53.825 529.965 ;
        RECT 42.615 527.075 42.785 527.245 ;
        RECT 43.075 527.075 43.245 527.245 ;
        RECT 43.535 527.075 43.705 527.245 ;
        RECT 43.995 527.075 44.165 527.245 ;
        RECT 44.455 527.075 44.625 527.245 ;
        RECT 44.915 527.075 45.085 527.245 ;
        RECT 45.375 527.075 45.545 527.245 ;
        RECT 45.835 527.075 46.005 527.245 ;
        RECT 46.295 527.075 46.465 527.245 ;
        RECT 46.755 527.075 46.925 527.245 ;
        RECT 47.215 527.075 47.385 527.245 ;
        RECT 47.675 527.075 47.845 527.245 ;
        RECT 48.135 527.075 48.305 527.245 ;
        RECT 48.595 527.075 48.765 527.245 ;
        RECT 49.055 527.075 49.225 527.245 ;
        RECT 49.515 527.075 49.685 527.245 ;
        RECT 49.975 527.075 50.145 527.245 ;
        RECT 50.435 527.075 50.605 527.245 ;
        RECT 50.895 527.075 51.065 527.245 ;
        RECT 51.355 527.075 51.525 527.245 ;
        RECT 51.815 527.075 51.985 527.245 ;
        RECT 52.275 527.075 52.445 527.245 ;
        RECT 52.735 527.075 52.905 527.245 ;
        RECT 53.195 527.075 53.365 527.245 ;
        RECT 53.655 527.075 53.825 527.245 ;
        RECT 42.615 524.355 42.785 524.525 ;
        RECT 43.075 524.355 43.245 524.525 ;
        RECT 43.535 524.355 43.705 524.525 ;
        RECT 43.995 524.355 44.165 524.525 ;
        RECT 44.455 524.355 44.625 524.525 ;
        RECT 44.915 524.355 45.085 524.525 ;
        RECT 45.375 524.355 45.545 524.525 ;
        RECT 45.835 524.355 46.005 524.525 ;
        RECT 46.295 524.355 46.465 524.525 ;
        RECT 46.755 524.355 46.925 524.525 ;
        RECT 47.215 524.355 47.385 524.525 ;
        RECT 47.675 524.355 47.845 524.525 ;
        RECT 48.135 524.355 48.305 524.525 ;
        RECT 48.595 524.355 48.765 524.525 ;
        RECT 49.055 524.355 49.225 524.525 ;
        RECT 49.515 524.355 49.685 524.525 ;
        RECT 49.975 524.355 50.145 524.525 ;
        RECT 50.435 524.355 50.605 524.525 ;
        RECT 50.895 524.355 51.065 524.525 ;
        RECT 51.355 524.355 51.525 524.525 ;
        RECT 51.815 524.355 51.985 524.525 ;
        RECT 52.275 524.355 52.445 524.525 ;
        RECT 52.735 524.355 52.905 524.525 ;
        RECT 53.195 524.355 53.365 524.525 ;
        RECT 53.655 524.355 53.825 524.525 ;
        RECT 42.615 521.635 42.785 521.805 ;
        RECT 43.075 521.635 43.245 521.805 ;
        RECT 43.535 521.635 43.705 521.805 ;
        RECT 43.995 521.635 44.165 521.805 ;
        RECT 44.455 521.635 44.625 521.805 ;
        RECT 44.915 521.635 45.085 521.805 ;
        RECT 45.375 521.635 45.545 521.805 ;
        RECT 45.835 521.635 46.005 521.805 ;
        RECT 46.295 521.635 46.465 521.805 ;
        RECT 46.755 521.635 46.925 521.805 ;
        RECT 47.215 521.635 47.385 521.805 ;
        RECT 47.675 521.635 47.845 521.805 ;
        RECT 48.135 521.635 48.305 521.805 ;
        RECT 48.595 521.635 48.765 521.805 ;
        RECT 49.055 521.635 49.225 521.805 ;
        RECT 49.515 521.635 49.685 521.805 ;
        RECT 49.975 521.635 50.145 521.805 ;
        RECT 50.435 521.635 50.605 521.805 ;
        RECT 50.895 521.635 51.065 521.805 ;
        RECT 51.355 521.635 51.525 521.805 ;
        RECT 51.815 521.635 51.985 521.805 ;
        RECT 52.275 521.635 52.445 521.805 ;
        RECT 52.735 521.635 52.905 521.805 ;
        RECT 53.195 521.635 53.365 521.805 ;
        RECT 53.655 521.635 53.825 521.805 ;
        RECT 42.615 518.915 42.785 519.085 ;
        RECT 43.075 518.915 43.245 519.085 ;
        RECT 43.535 518.915 43.705 519.085 ;
        RECT 43.995 518.915 44.165 519.085 ;
        RECT 44.455 518.915 44.625 519.085 ;
        RECT 44.915 518.915 45.085 519.085 ;
        RECT 45.375 518.915 45.545 519.085 ;
        RECT 45.835 518.915 46.005 519.085 ;
        RECT 46.295 518.915 46.465 519.085 ;
        RECT 46.755 518.915 46.925 519.085 ;
        RECT 47.215 518.915 47.385 519.085 ;
        RECT 47.675 518.915 47.845 519.085 ;
        RECT 48.135 518.915 48.305 519.085 ;
        RECT 48.595 518.915 48.765 519.085 ;
        RECT 49.055 518.915 49.225 519.085 ;
        RECT 49.515 518.915 49.685 519.085 ;
        RECT 49.975 518.915 50.145 519.085 ;
        RECT 50.435 518.915 50.605 519.085 ;
        RECT 50.895 518.915 51.065 519.085 ;
        RECT 51.355 518.915 51.525 519.085 ;
        RECT 51.815 518.915 51.985 519.085 ;
        RECT 52.275 518.915 52.445 519.085 ;
        RECT 52.735 518.915 52.905 519.085 ;
        RECT 53.195 518.915 53.365 519.085 ;
        RECT 53.655 518.915 53.825 519.085 ;
        RECT 42.615 516.195 42.785 516.365 ;
        RECT 43.075 516.195 43.245 516.365 ;
        RECT 43.535 516.195 43.705 516.365 ;
        RECT 43.995 516.195 44.165 516.365 ;
        RECT 44.455 516.195 44.625 516.365 ;
        RECT 44.915 516.195 45.085 516.365 ;
        RECT 45.375 516.195 45.545 516.365 ;
        RECT 45.835 516.195 46.005 516.365 ;
        RECT 46.295 516.195 46.465 516.365 ;
        RECT 46.755 516.195 46.925 516.365 ;
        RECT 47.215 516.195 47.385 516.365 ;
        RECT 47.675 516.195 47.845 516.365 ;
        RECT 48.135 516.195 48.305 516.365 ;
        RECT 48.595 516.195 48.765 516.365 ;
        RECT 49.055 516.195 49.225 516.365 ;
        RECT 49.515 516.195 49.685 516.365 ;
        RECT 49.975 516.195 50.145 516.365 ;
        RECT 50.435 516.195 50.605 516.365 ;
        RECT 50.895 516.195 51.065 516.365 ;
        RECT 51.355 516.195 51.525 516.365 ;
        RECT 51.815 516.195 51.985 516.365 ;
        RECT 52.275 516.195 52.445 516.365 ;
        RECT 52.735 516.195 52.905 516.365 ;
        RECT 53.195 516.195 53.365 516.365 ;
        RECT 53.655 516.195 53.825 516.365 ;
        RECT 42.615 513.475 42.785 513.645 ;
        RECT 43.075 513.475 43.245 513.645 ;
        RECT 43.535 513.475 43.705 513.645 ;
        RECT 43.995 513.475 44.165 513.645 ;
        RECT 44.455 513.475 44.625 513.645 ;
        RECT 44.915 513.475 45.085 513.645 ;
        RECT 45.375 513.475 45.545 513.645 ;
        RECT 45.835 513.475 46.005 513.645 ;
        RECT 46.295 513.475 46.465 513.645 ;
        RECT 46.755 513.475 46.925 513.645 ;
        RECT 47.215 513.475 47.385 513.645 ;
        RECT 47.675 513.475 47.845 513.645 ;
        RECT 48.135 513.475 48.305 513.645 ;
        RECT 48.595 513.475 48.765 513.645 ;
        RECT 49.055 513.475 49.225 513.645 ;
        RECT 49.515 513.475 49.685 513.645 ;
        RECT 49.975 513.475 50.145 513.645 ;
        RECT 50.435 513.475 50.605 513.645 ;
        RECT 50.895 513.475 51.065 513.645 ;
        RECT 51.355 513.475 51.525 513.645 ;
        RECT 51.815 513.475 51.985 513.645 ;
        RECT 52.275 513.475 52.445 513.645 ;
        RECT 52.735 513.475 52.905 513.645 ;
        RECT 53.195 513.475 53.365 513.645 ;
        RECT 53.655 513.475 53.825 513.645 ;
        RECT 42.615 510.755 42.785 510.925 ;
        RECT 43.075 510.755 43.245 510.925 ;
        RECT 43.535 510.755 43.705 510.925 ;
        RECT 43.995 510.755 44.165 510.925 ;
        RECT 44.455 510.755 44.625 510.925 ;
        RECT 44.915 510.755 45.085 510.925 ;
        RECT 45.375 510.755 45.545 510.925 ;
        RECT 45.835 510.755 46.005 510.925 ;
        RECT 46.295 510.755 46.465 510.925 ;
        RECT 46.755 510.755 46.925 510.925 ;
        RECT 47.215 510.755 47.385 510.925 ;
        RECT 47.675 510.755 47.845 510.925 ;
        RECT 48.135 510.755 48.305 510.925 ;
        RECT 48.595 510.755 48.765 510.925 ;
        RECT 49.055 510.755 49.225 510.925 ;
        RECT 49.515 510.755 49.685 510.925 ;
        RECT 49.975 510.755 50.145 510.925 ;
        RECT 50.435 510.755 50.605 510.925 ;
        RECT 50.895 510.755 51.065 510.925 ;
        RECT 51.355 510.755 51.525 510.925 ;
        RECT 51.815 510.755 51.985 510.925 ;
        RECT 52.275 510.755 52.445 510.925 ;
        RECT 52.735 510.755 52.905 510.925 ;
        RECT 53.195 510.755 53.365 510.925 ;
        RECT 53.655 510.755 53.825 510.925 ;
        RECT 42.615 508.035 42.785 508.205 ;
        RECT 43.075 508.035 43.245 508.205 ;
        RECT 43.535 508.035 43.705 508.205 ;
        RECT 43.995 508.035 44.165 508.205 ;
        RECT 44.455 508.035 44.625 508.205 ;
        RECT 44.915 508.035 45.085 508.205 ;
        RECT 45.375 508.035 45.545 508.205 ;
        RECT 45.835 508.035 46.005 508.205 ;
        RECT 46.295 508.035 46.465 508.205 ;
        RECT 46.755 508.035 46.925 508.205 ;
        RECT 47.215 508.035 47.385 508.205 ;
        RECT 47.675 508.035 47.845 508.205 ;
        RECT 48.135 508.035 48.305 508.205 ;
        RECT 48.595 508.035 48.765 508.205 ;
        RECT 49.055 508.035 49.225 508.205 ;
        RECT 49.515 508.035 49.685 508.205 ;
        RECT 49.975 508.035 50.145 508.205 ;
        RECT 50.435 508.035 50.605 508.205 ;
        RECT 50.895 508.035 51.065 508.205 ;
        RECT 51.355 508.035 51.525 508.205 ;
        RECT 51.815 508.035 51.985 508.205 ;
        RECT 52.275 508.035 52.445 508.205 ;
        RECT 52.735 508.035 52.905 508.205 ;
        RECT 53.195 508.035 53.365 508.205 ;
        RECT 53.655 508.035 53.825 508.205 ;
        RECT 42.615 505.315 42.785 505.485 ;
        RECT 43.075 505.315 43.245 505.485 ;
        RECT 43.535 505.315 43.705 505.485 ;
        RECT 43.995 505.315 44.165 505.485 ;
        RECT 44.455 505.315 44.625 505.485 ;
        RECT 44.915 505.315 45.085 505.485 ;
        RECT 45.375 505.315 45.545 505.485 ;
        RECT 45.835 505.315 46.005 505.485 ;
        RECT 46.295 505.315 46.465 505.485 ;
        RECT 46.755 505.315 46.925 505.485 ;
        RECT 47.215 505.315 47.385 505.485 ;
        RECT 47.675 505.315 47.845 505.485 ;
        RECT 48.135 505.315 48.305 505.485 ;
        RECT 48.595 505.315 48.765 505.485 ;
        RECT 49.055 505.315 49.225 505.485 ;
        RECT 49.515 505.315 49.685 505.485 ;
        RECT 49.975 505.315 50.145 505.485 ;
        RECT 50.435 505.315 50.605 505.485 ;
        RECT 50.895 505.315 51.065 505.485 ;
        RECT 51.355 505.315 51.525 505.485 ;
        RECT 51.815 505.315 51.985 505.485 ;
        RECT 52.275 505.315 52.445 505.485 ;
        RECT 52.735 505.315 52.905 505.485 ;
        RECT 53.195 505.315 53.365 505.485 ;
        RECT 53.655 505.315 53.825 505.485 ;
        RECT 42.615 502.595 42.785 502.765 ;
        RECT 43.075 502.595 43.245 502.765 ;
        RECT 43.535 502.595 43.705 502.765 ;
        RECT 43.995 502.595 44.165 502.765 ;
        RECT 44.455 502.595 44.625 502.765 ;
        RECT 44.915 502.595 45.085 502.765 ;
        RECT 45.375 502.595 45.545 502.765 ;
        RECT 45.835 502.595 46.005 502.765 ;
        RECT 46.295 502.595 46.465 502.765 ;
        RECT 46.755 502.595 46.925 502.765 ;
        RECT 47.215 502.595 47.385 502.765 ;
        RECT 47.675 502.595 47.845 502.765 ;
        RECT 48.135 502.595 48.305 502.765 ;
        RECT 48.595 502.595 48.765 502.765 ;
        RECT 49.055 502.595 49.225 502.765 ;
        RECT 49.515 502.595 49.685 502.765 ;
        RECT 49.975 502.595 50.145 502.765 ;
        RECT 50.435 502.595 50.605 502.765 ;
        RECT 50.895 502.595 51.065 502.765 ;
        RECT 51.355 502.595 51.525 502.765 ;
        RECT 51.815 502.595 51.985 502.765 ;
        RECT 52.275 502.595 52.445 502.765 ;
        RECT 52.735 502.595 52.905 502.765 ;
        RECT 53.195 502.595 53.365 502.765 ;
        RECT 53.655 502.595 53.825 502.765 ;
        RECT 42.615 499.875 42.785 500.045 ;
        RECT 43.075 499.875 43.245 500.045 ;
        RECT 43.535 499.875 43.705 500.045 ;
        RECT 43.995 499.875 44.165 500.045 ;
        RECT 44.455 499.875 44.625 500.045 ;
        RECT 44.915 499.875 45.085 500.045 ;
        RECT 45.375 499.875 45.545 500.045 ;
        RECT 45.835 499.875 46.005 500.045 ;
        RECT 46.295 499.875 46.465 500.045 ;
        RECT 46.755 499.875 46.925 500.045 ;
        RECT 47.215 499.875 47.385 500.045 ;
        RECT 47.675 499.875 47.845 500.045 ;
        RECT 48.135 499.875 48.305 500.045 ;
        RECT 48.595 499.875 48.765 500.045 ;
        RECT 49.055 499.875 49.225 500.045 ;
        RECT 49.515 499.875 49.685 500.045 ;
        RECT 49.975 499.875 50.145 500.045 ;
        RECT 50.435 499.875 50.605 500.045 ;
        RECT 50.895 499.875 51.065 500.045 ;
        RECT 51.355 499.875 51.525 500.045 ;
        RECT 51.815 499.875 51.985 500.045 ;
        RECT 52.275 499.875 52.445 500.045 ;
        RECT 52.735 499.875 52.905 500.045 ;
        RECT 53.195 499.875 53.365 500.045 ;
        RECT 53.655 499.875 53.825 500.045 ;
        RECT 42.615 497.155 42.785 497.325 ;
        RECT 43.075 497.155 43.245 497.325 ;
        RECT 43.535 497.155 43.705 497.325 ;
        RECT 43.995 497.155 44.165 497.325 ;
        RECT 44.455 497.155 44.625 497.325 ;
        RECT 44.915 497.155 45.085 497.325 ;
        RECT 45.375 497.155 45.545 497.325 ;
        RECT 45.835 497.155 46.005 497.325 ;
        RECT 46.295 497.155 46.465 497.325 ;
        RECT 46.755 497.155 46.925 497.325 ;
        RECT 47.215 497.155 47.385 497.325 ;
        RECT 47.675 497.155 47.845 497.325 ;
        RECT 48.135 497.155 48.305 497.325 ;
        RECT 48.595 497.155 48.765 497.325 ;
        RECT 49.055 497.155 49.225 497.325 ;
        RECT 49.515 497.155 49.685 497.325 ;
        RECT 49.975 497.155 50.145 497.325 ;
        RECT 50.435 497.155 50.605 497.325 ;
        RECT 50.895 497.155 51.065 497.325 ;
        RECT 51.355 497.155 51.525 497.325 ;
        RECT 51.815 497.155 51.985 497.325 ;
        RECT 52.275 497.155 52.445 497.325 ;
        RECT 52.735 497.155 52.905 497.325 ;
        RECT 53.195 497.155 53.365 497.325 ;
        RECT 53.655 497.155 53.825 497.325 ;
        RECT 42.615 494.435 42.785 494.605 ;
        RECT 43.075 494.435 43.245 494.605 ;
        RECT 43.535 494.435 43.705 494.605 ;
        RECT 43.995 494.435 44.165 494.605 ;
        RECT 44.455 494.435 44.625 494.605 ;
        RECT 44.915 494.435 45.085 494.605 ;
        RECT 45.375 494.435 45.545 494.605 ;
        RECT 45.835 494.435 46.005 494.605 ;
        RECT 46.295 494.435 46.465 494.605 ;
        RECT 46.755 494.435 46.925 494.605 ;
        RECT 47.215 494.435 47.385 494.605 ;
        RECT 47.675 494.435 47.845 494.605 ;
        RECT 48.135 494.435 48.305 494.605 ;
        RECT 48.595 494.435 48.765 494.605 ;
        RECT 49.055 494.435 49.225 494.605 ;
        RECT 49.515 494.435 49.685 494.605 ;
        RECT 49.975 494.435 50.145 494.605 ;
        RECT 50.435 494.435 50.605 494.605 ;
        RECT 50.895 494.435 51.065 494.605 ;
        RECT 51.355 494.435 51.525 494.605 ;
        RECT 51.815 494.435 51.985 494.605 ;
        RECT 52.275 494.435 52.445 494.605 ;
        RECT 52.735 494.435 52.905 494.605 ;
        RECT 53.195 494.435 53.365 494.605 ;
        RECT 53.655 494.435 53.825 494.605 ;
        RECT 42.615 491.715 42.785 491.885 ;
        RECT 43.075 491.715 43.245 491.885 ;
        RECT 43.535 491.715 43.705 491.885 ;
        RECT 43.995 491.715 44.165 491.885 ;
        RECT 44.455 491.715 44.625 491.885 ;
        RECT 44.915 491.715 45.085 491.885 ;
        RECT 45.375 491.715 45.545 491.885 ;
        RECT 45.835 491.715 46.005 491.885 ;
        RECT 46.295 491.715 46.465 491.885 ;
        RECT 46.755 491.715 46.925 491.885 ;
        RECT 47.215 491.715 47.385 491.885 ;
        RECT 47.675 491.715 47.845 491.885 ;
        RECT 48.135 491.715 48.305 491.885 ;
        RECT 48.595 491.715 48.765 491.885 ;
        RECT 49.055 491.715 49.225 491.885 ;
        RECT 49.515 491.715 49.685 491.885 ;
        RECT 49.975 491.715 50.145 491.885 ;
        RECT 50.435 491.715 50.605 491.885 ;
        RECT 50.895 491.715 51.065 491.885 ;
        RECT 51.355 491.715 51.525 491.885 ;
        RECT 51.815 491.715 51.985 491.885 ;
        RECT 52.275 491.715 52.445 491.885 ;
        RECT 52.735 491.715 52.905 491.885 ;
        RECT 53.195 491.715 53.365 491.885 ;
        RECT 53.655 491.715 53.825 491.885 ;
        RECT 42.615 488.995 42.785 489.165 ;
        RECT 43.075 488.995 43.245 489.165 ;
        RECT 43.535 488.995 43.705 489.165 ;
        RECT 43.995 488.995 44.165 489.165 ;
        RECT 44.455 488.995 44.625 489.165 ;
        RECT 44.915 488.995 45.085 489.165 ;
        RECT 45.375 488.995 45.545 489.165 ;
        RECT 45.835 488.995 46.005 489.165 ;
        RECT 46.295 488.995 46.465 489.165 ;
        RECT 46.755 488.995 46.925 489.165 ;
        RECT 47.215 488.995 47.385 489.165 ;
        RECT 47.675 488.995 47.845 489.165 ;
        RECT 48.135 488.995 48.305 489.165 ;
        RECT 48.595 488.995 48.765 489.165 ;
        RECT 49.055 488.995 49.225 489.165 ;
        RECT 49.515 488.995 49.685 489.165 ;
        RECT 49.975 488.995 50.145 489.165 ;
        RECT 50.435 488.995 50.605 489.165 ;
        RECT 50.895 488.995 51.065 489.165 ;
        RECT 51.355 488.995 51.525 489.165 ;
        RECT 51.815 488.995 51.985 489.165 ;
        RECT 52.275 488.995 52.445 489.165 ;
        RECT 52.735 488.995 52.905 489.165 ;
        RECT 53.195 488.995 53.365 489.165 ;
        RECT 53.655 488.995 53.825 489.165 ;
        RECT 42.615 486.275 42.785 486.445 ;
        RECT 43.075 486.275 43.245 486.445 ;
        RECT 43.535 486.275 43.705 486.445 ;
        RECT 43.995 486.275 44.165 486.445 ;
        RECT 44.455 486.275 44.625 486.445 ;
        RECT 44.915 486.275 45.085 486.445 ;
        RECT 45.375 486.275 45.545 486.445 ;
        RECT 45.835 486.275 46.005 486.445 ;
        RECT 46.295 486.275 46.465 486.445 ;
        RECT 46.755 486.275 46.925 486.445 ;
        RECT 47.215 486.275 47.385 486.445 ;
        RECT 47.675 486.275 47.845 486.445 ;
        RECT 48.135 486.275 48.305 486.445 ;
        RECT 48.595 486.275 48.765 486.445 ;
        RECT 49.055 486.275 49.225 486.445 ;
        RECT 49.515 486.275 49.685 486.445 ;
        RECT 49.975 486.275 50.145 486.445 ;
        RECT 50.435 486.275 50.605 486.445 ;
        RECT 50.895 486.275 51.065 486.445 ;
        RECT 51.355 486.275 51.525 486.445 ;
        RECT 51.815 486.275 51.985 486.445 ;
        RECT 52.275 486.275 52.445 486.445 ;
        RECT 52.735 486.275 52.905 486.445 ;
        RECT 53.195 486.275 53.365 486.445 ;
        RECT 53.655 486.275 53.825 486.445 ;
        RECT 42.615 483.555 42.785 483.725 ;
        RECT 43.075 483.555 43.245 483.725 ;
        RECT 43.535 483.555 43.705 483.725 ;
        RECT 43.995 483.555 44.165 483.725 ;
        RECT 44.455 483.555 44.625 483.725 ;
        RECT 44.915 483.555 45.085 483.725 ;
        RECT 45.375 483.555 45.545 483.725 ;
        RECT 45.835 483.555 46.005 483.725 ;
        RECT 46.295 483.555 46.465 483.725 ;
        RECT 46.755 483.555 46.925 483.725 ;
        RECT 47.215 483.555 47.385 483.725 ;
        RECT 47.675 483.555 47.845 483.725 ;
        RECT 48.135 483.555 48.305 483.725 ;
        RECT 48.595 483.555 48.765 483.725 ;
        RECT 49.055 483.555 49.225 483.725 ;
        RECT 49.515 483.555 49.685 483.725 ;
        RECT 49.975 483.555 50.145 483.725 ;
        RECT 50.435 483.555 50.605 483.725 ;
        RECT 50.895 483.555 51.065 483.725 ;
        RECT 51.355 483.555 51.525 483.725 ;
        RECT 51.815 483.555 51.985 483.725 ;
        RECT 52.275 483.555 52.445 483.725 ;
        RECT 52.735 483.555 52.905 483.725 ;
        RECT 53.195 483.555 53.365 483.725 ;
        RECT 53.655 483.555 53.825 483.725 ;
        RECT 42.615 480.835 42.785 481.005 ;
        RECT 43.075 480.835 43.245 481.005 ;
        RECT 43.535 480.835 43.705 481.005 ;
        RECT 43.995 480.835 44.165 481.005 ;
        RECT 44.455 480.835 44.625 481.005 ;
        RECT 44.915 480.835 45.085 481.005 ;
        RECT 45.375 480.835 45.545 481.005 ;
        RECT 45.835 480.835 46.005 481.005 ;
        RECT 46.295 480.835 46.465 481.005 ;
        RECT 46.755 480.835 46.925 481.005 ;
        RECT 47.215 480.835 47.385 481.005 ;
        RECT 47.675 480.835 47.845 481.005 ;
        RECT 48.135 480.835 48.305 481.005 ;
        RECT 48.595 480.835 48.765 481.005 ;
        RECT 49.055 480.835 49.225 481.005 ;
        RECT 49.515 480.835 49.685 481.005 ;
        RECT 49.975 480.835 50.145 481.005 ;
        RECT 50.435 480.835 50.605 481.005 ;
        RECT 50.895 480.835 51.065 481.005 ;
        RECT 51.355 480.835 51.525 481.005 ;
        RECT 51.815 480.835 51.985 481.005 ;
        RECT 52.275 480.835 52.445 481.005 ;
        RECT 52.735 480.835 52.905 481.005 ;
        RECT 53.195 480.835 53.365 481.005 ;
        RECT 53.655 480.835 53.825 481.005 ;
        RECT 42.615 478.115 42.785 478.285 ;
        RECT 43.075 478.115 43.245 478.285 ;
        RECT 43.535 478.115 43.705 478.285 ;
        RECT 43.995 478.115 44.165 478.285 ;
        RECT 44.455 478.115 44.625 478.285 ;
        RECT 44.915 478.115 45.085 478.285 ;
        RECT 45.375 478.115 45.545 478.285 ;
        RECT 45.835 478.115 46.005 478.285 ;
        RECT 46.295 478.115 46.465 478.285 ;
        RECT 46.755 478.115 46.925 478.285 ;
        RECT 47.215 478.115 47.385 478.285 ;
        RECT 47.675 478.115 47.845 478.285 ;
        RECT 48.135 478.115 48.305 478.285 ;
        RECT 48.595 478.115 48.765 478.285 ;
        RECT 49.055 478.115 49.225 478.285 ;
        RECT 49.515 478.115 49.685 478.285 ;
        RECT 49.975 478.115 50.145 478.285 ;
        RECT 50.435 478.115 50.605 478.285 ;
        RECT 50.895 478.115 51.065 478.285 ;
        RECT 51.355 478.115 51.525 478.285 ;
        RECT 51.815 478.115 51.985 478.285 ;
        RECT 52.275 478.115 52.445 478.285 ;
        RECT 52.735 478.115 52.905 478.285 ;
        RECT 53.195 478.115 53.365 478.285 ;
        RECT 53.655 478.115 53.825 478.285 ;
        RECT 42.615 475.395 42.785 475.565 ;
        RECT 43.075 475.395 43.245 475.565 ;
        RECT 43.535 475.395 43.705 475.565 ;
        RECT 43.995 475.395 44.165 475.565 ;
        RECT 44.455 475.395 44.625 475.565 ;
        RECT 44.915 475.395 45.085 475.565 ;
        RECT 45.375 475.395 45.545 475.565 ;
        RECT 45.835 475.395 46.005 475.565 ;
        RECT 46.295 475.395 46.465 475.565 ;
        RECT 46.755 475.395 46.925 475.565 ;
        RECT 47.215 475.395 47.385 475.565 ;
        RECT 47.675 475.395 47.845 475.565 ;
        RECT 48.135 475.395 48.305 475.565 ;
        RECT 48.595 475.395 48.765 475.565 ;
        RECT 49.055 475.395 49.225 475.565 ;
        RECT 49.515 475.395 49.685 475.565 ;
        RECT 49.975 475.395 50.145 475.565 ;
        RECT 50.435 475.395 50.605 475.565 ;
        RECT 50.895 475.395 51.065 475.565 ;
        RECT 51.355 475.395 51.525 475.565 ;
        RECT 51.815 475.395 51.985 475.565 ;
        RECT 52.275 475.395 52.445 475.565 ;
        RECT 52.735 475.395 52.905 475.565 ;
        RECT 53.195 475.395 53.365 475.565 ;
        RECT 53.655 475.395 53.825 475.565 ;
        RECT 42.615 472.675 42.785 472.845 ;
        RECT 43.075 472.675 43.245 472.845 ;
        RECT 43.535 472.675 43.705 472.845 ;
        RECT 43.995 472.675 44.165 472.845 ;
        RECT 44.455 472.675 44.625 472.845 ;
        RECT 44.915 472.675 45.085 472.845 ;
        RECT 45.375 472.675 45.545 472.845 ;
        RECT 45.835 472.675 46.005 472.845 ;
        RECT 46.295 472.675 46.465 472.845 ;
        RECT 46.755 472.675 46.925 472.845 ;
        RECT 47.215 472.675 47.385 472.845 ;
        RECT 47.675 472.675 47.845 472.845 ;
        RECT 48.135 472.675 48.305 472.845 ;
        RECT 48.595 472.675 48.765 472.845 ;
        RECT 49.055 472.675 49.225 472.845 ;
        RECT 49.515 472.675 49.685 472.845 ;
        RECT 49.975 472.675 50.145 472.845 ;
        RECT 50.435 472.675 50.605 472.845 ;
        RECT 50.895 472.675 51.065 472.845 ;
        RECT 51.355 472.675 51.525 472.845 ;
        RECT 51.815 472.675 51.985 472.845 ;
        RECT 52.275 472.675 52.445 472.845 ;
        RECT 52.735 472.675 52.905 472.845 ;
        RECT 53.195 472.675 53.365 472.845 ;
        RECT 53.655 472.675 53.825 472.845 ;
        RECT 42.615 469.955 42.785 470.125 ;
        RECT 43.075 469.955 43.245 470.125 ;
        RECT 43.535 469.955 43.705 470.125 ;
        RECT 43.995 469.955 44.165 470.125 ;
        RECT 44.455 469.955 44.625 470.125 ;
        RECT 44.915 469.955 45.085 470.125 ;
        RECT 45.375 469.955 45.545 470.125 ;
        RECT 45.835 469.955 46.005 470.125 ;
        RECT 46.295 469.955 46.465 470.125 ;
        RECT 46.755 469.955 46.925 470.125 ;
        RECT 47.215 469.955 47.385 470.125 ;
        RECT 47.675 469.955 47.845 470.125 ;
        RECT 48.135 469.955 48.305 470.125 ;
        RECT 48.595 469.955 48.765 470.125 ;
        RECT 49.055 469.955 49.225 470.125 ;
        RECT 49.515 469.955 49.685 470.125 ;
        RECT 49.975 469.955 50.145 470.125 ;
        RECT 50.435 469.955 50.605 470.125 ;
        RECT 50.895 469.955 51.065 470.125 ;
        RECT 51.355 469.955 51.525 470.125 ;
        RECT 51.815 469.955 51.985 470.125 ;
        RECT 52.275 469.955 52.445 470.125 ;
        RECT 52.735 469.955 52.905 470.125 ;
        RECT 53.195 469.955 53.365 470.125 ;
        RECT 53.655 469.955 53.825 470.125 ;
        RECT 42.615 467.235 42.785 467.405 ;
        RECT 43.075 467.235 43.245 467.405 ;
        RECT 43.535 467.235 43.705 467.405 ;
        RECT 43.995 467.235 44.165 467.405 ;
        RECT 44.455 467.235 44.625 467.405 ;
        RECT 44.915 467.235 45.085 467.405 ;
        RECT 45.375 467.235 45.545 467.405 ;
        RECT 45.835 467.235 46.005 467.405 ;
        RECT 46.295 467.235 46.465 467.405 ;
        RECT 46.755 467.235 46.925 467.405 ;
        RECT 47.215 467.235 47.385 467.405 ;
        RECT 47.675 467.235 47.845 467.405 ;
        RECT 48.135 467.235 48.305 467.405 ;
        RECT 48.595 467.235 48.765 467.405 ;
        RECT 49.055 467.235 49.225 467.405 ;
        RECT 49.515 467.235 49.685 467.405 ;
        RECT 49.975 467.235 50.145 467.405 ;
        RECT 50.435 467.235 50.605 467.405 ;
        RECT 50.895 467.235 51.065 467.405 ;
        RECT 51.355 467.235 51.525 467.405 ;
        RECT 51.815 467.235 51.985 467.405 ;
        RECT 52.275 467.235 52.445 467.405 ;
        RECT 52.735 467.235 52.905 467.405 ;
        RECT 53.195 467.235 53.365 467.405 ;
        RECT 53.655 467.235 53.825 467.405 ;
        RECT 42.615 464.515 42.785 464.685 ;
        RECT 43.075 464.515 43.245 464.685 ;
        RECT 43.535 464.515 43.705 464.685 ;
        RECT 43.995 464.515 44.165 464.685 ;
        RECT 44.455 464.515 44.625 464.685 ;
        RECT 44.915 464.515 45.085 464.685 ;
        RECT 45.375 464.515 45.545 464.685 ;
        RECT 45.835 464.515 46.005 464.685 ;
        RECT 46.295 464.515 46.465 464.685 ;
        RECT 46.755 464.515 46.925 464.685 ;
        RECT 47.215 464.515 47.385 464.685 ;
        RECT 47.675 464.515 47.845 464.685 ;
        RECT 48.135 464.515 48.305 464.685 ;
        RECT 48.595 464.515 48.765 464.685 ;
        RECT 49.055 464.515 49.225 464.685 ;
        RECT 49.515 464.515 49.685 464.685 ;
        RECT 49.975 464.515 50.145 464.685 ;
        RECT 50.435 464.515 50.605 464.685 ;
        RECT 50.895 464.515 51.065 464.685 ;
        RECT 51.355 464.515 51.525 464.685 ;
        RECT 51.815 464.515 51.985 464.685 ;
        RECT 52.275 464.515 52.445 464.685 ;
        RECT 52.735 464.515 52.905 464.685 ;
        RECT 53.195 464.515 53.365 464.685 ;
        RECT 53.655 464.515 53.825 464.685 ;
        RECT 42.615 461.795 42.785 461.965 ;
        RECT 43.075 461.795 43.245 461.965 ;
        RECT 43.535 461.795 43.705 461.965 ;
        RECT 43.995 461.795 44.165 461.965 ;
        RECT 44.455 461.795 44.625 461.965 ;
        RECT 44.915 461.795 45.085 461.965 ;
        RECT 45.375 461.795 45.545 461.965 ;
        RECT 45.835 461.795 46.005 461.965 ;
        RECT 46.295 461.795 46.465 461.965 ;
        RECT 46.755 461.795 46.925 461.965 ;
        RECT 47.215 461.795 47.385 461.965 ;
        RECT 47.675 461.795 47.845 461.965 ;
        RECT 48.135 461.795 48.305 461.965 ;
        RECT 48.595 461.795 48.765 461.965 ;
        RECT 49.055 461.795 49.225 461.965 ;
        RECT 49.515 461.795 49.685 461.965 ;
        RECT 49.975 461.795 50.145 461.965 ;
        RECT 50.435 461.795 50.605 461.965 ;
        RECT 50.895 461.795 51.065 461.965 ;
        RECT 51.355 461.795 51.525 461.965 ;
        RECT 51.815 461.795 51.985 461.965 ;
        RECT 52.275 461.795 52.445 461.965 ;
        RECT 52.735 461.795 52.905 461.965 ;
        RECT 53.195 461.795 53.365 461.965 ;
        RECT 53.655 461.795 53.825 461.965 ;
        RECT 42.615 459.075 42.785 459.245 ;
        RECT 43.075 459.075 43.245 459.245 ;
        RECT 43.535 459.075 43.705 459.245 ;
        RECT 43.995 459.075 44.165 459.245 ;
        RECT 44.455 459.075 44.625 459.245 ;
        RECT 44.915 459.075 45.085 459.245 ;
        RECT 45.375 459.075 45.545 459.245 ;
        RECT 45.835 459.075 46.005 459.245 ;
        RECT 46.295 459.075 46.465 459.245 ;
        RECT 46.755 459.075 46.925 459.245 ;
        RECT 47.215 459.075 47.385 459.245 ;
        RECT 47.675 459.075 47.845 459.245 ;
        RECT 48.135 459.075 48.305 459.245 ;
        RECT 48.595 459.075 48.765 459.245 ;
        RECT 49.055 459.075 49.225 459.245 ;
        RECT 49.515 459.075 49.685 459.245 ;
        RECT 49.975 459.075 50.145 459.245 ;
        RECT 50.435 459.075 50.605 459.245 ;
        RECT 50.895 459.075 51.065 459.245 ;
        RECT 51.355 459.075 51.525 459.245 ;
        RECT 51.815 459.075 51.985 459.245 ;
        RECT 52.275 459.075 52.445 459.245 ;
        RECT 52.735 459.075 52.905 459.245 ;
        RECT 53.195 459.075 53.365 459.245 ;
        RECT 53.655 459.075 53.825 459.245 ;
        RECT 42.615 456.355 42.785 456.525 ;
        RECT 43.075 456.355 43.245 456.525 ;
        RECT 43.535 456.355 43.705 456.525 ;
        RECT 43.995 456.355 44.165 456.525 ;
        RECT 44.455 456.355 44.625 456.525 ;
        RECT 44.915 456.355 45.085 456.525 ;
        RECT 45.375 456.355 45.545 456.525 ;
        RECT 45.835 456.355 46.005 456.525 ;
        RECT 46.295 456.355 46.465 456.525 ;
        RECT 46.755 456.355 46.925 456.525 ;
        RECT 47.215 456.355 47.385 456.525 ;
        RECT 47.675 456.355 47.845 456.525 ;
        RECT 48.135 456.355 48.305 456.525 ;
        RECT 48.595 456.355 48.765 456.525 ;
        RECT 49.055 456.355 49.225 456.525 ;
        RECT 49.515 456.355 49.685 456.525 ;
        RECT 49.975 456.355 50.145 456.525 ;
        RECT 50.435 456.355 50.605 456.525 ;
        RECT 50.895 456.355 51.065 456.525 ;
        RECT 51.355 456.355 51.525 456.525 ;
        RECT 51.815 456.355 51.985 456.525 ;
        RECT 52.275 456.355 52.445 456.525 ;
        RECT 52.735 456.355 52.905 456.525 ;
        RECT 53.195 456.355 53.365 456.525 ;
        RECT 53.655 456.355 53.825 456.525 ;
        RECT 42.615 453.635 42.785 453.805 ;
        RECT 43.075 453.635 43.245 453.805 ;
        RECT 43.535 453.635 43.705 453.805 ;
        RECT 43.995 453.635 44.165 453.805 ;
        RECT 44.455 453.635 44.625 453.805 ;
        RECT 44.915 453.635 45.085 453.805 ;
        RECT 45.375 453.635 45.545 453.805 ;
        RECT 45.835 453.635 46.005 453.805 ;
        RECT 46.295 453.635 46.465 453.805 ;
        RECT 46.755 453.635 46.925 453.805 ;
        RECT 47.215 453.635 47.385 453.805 ;
        RECT 47.675 453.635 47.845 453.805 ;
        RECT 48.135 453.635 48.305 453.805 ;
        RECT 48.595 453.635 48.765 453.805 ;
        RECT 49.055 453.635 49.225 453.805 ;
        RECT 49.515 453.635 49.685 453.805 ;
        RECT 49.975 453.635 50.145 453.805 ;
        RECT 50.435 453.635 50.605 453.805 ;
        RECT 50.895 453.635 51.065 453.805 ;
        RECT 51.355 453.635 51.525 453.805 ;
        RECT 51.815 453.635 51.985 453.805 ;
        RECT 52.275 453.635 52.445 453.805 ;
        RECT 52.735 453.635 52.905 453.805 ;
        RECT 53.195 453.635 53.365 453.805 ;
        RECT 53.655 453.635 53.825 453.805 ;
        RECT 42.615 450.915 42.785 451.085 ;
        RECT 43.075 450.915 43.245 451.085 ;
        RECT 43.535 450.915 43.705 451.085 ;
        RECT 43.995 450.915 44.165 451.085 ;
        RECT 44.455 450.915 44.625 451.085 ;
        RECT 44.915 450.915 45.085 451.085 ;
        RECT 45.375 450.915 45.545 451.085 ;
        RECT 45.835 450.915 46.005 451.085 ;
        RECT 46.295 450.915 46.465 451.085 ;
        RECT 46.755 450.915 46.925 451.085 ;
        RECT 47.215 450.915 47.385 451.085 ;
        RECT 47.675 450.915 47.845 451.085 ;
        RECT 48.135 450.915 48.305 451.085 ;
        RECT 48.595 450.915 48.765 451.085 ;
        RECT 49.055 450.915 49.225 451.085 ;
        RECT 49.515 450.915 49.685 451.085 ;
        RECT 49.975 450.915 50.145 451.085 ;
        RECT 50.435 450.915 50.605 451.085 ;
        RECT 50.895 450.915 51.065 451.085 ;
        RECT 51.355 450.915 51.525 451.085 ;
        RECT 51.815 450.915 51.985 451.085 ;
        RECT 52.275 450.915 52.445 451.085 ;
        RECT 52.735 450.915 52.905 451.085 ;
        RECT 53.195 450.915 53.365 451.085 ;
        RECT 53.655 450.915 53.825 451.085 ;
        RECT 42.615 448.195 42.785 448.365 ;
        RECT 43.075 448.195 43.245 448.365 ;
        RECT 43.535 448.195 43.705 448.365 ;
        RECT 43.995 448.195 44.165 448.365 ;
        RECT 44.455 448.195 44.625 448.365 ;
        RECT 44.915 448.195 45.085 448.365 ;
        RECT 45.375 448.195 45.545 448.365 ;
        RECT 45.835 448.195 46.005 448.365 ;
        RECT 46.295 448.195 46.465 448.365 ;
        RECT 46.755 448.195 46.925 448.365 ;
        RECT 47.215 448.195 47.385 448.365 ;
        RECT 47.675 448.195 47.845 448.365 ;
        RECT 48.135 448.195 48.305 448.365 ;
        RECT 48.595 448.195 48.765 448.365 ;
        RECT 49.055 448.195 49.225 448.365 ;
        RECT 49.515 448.195 49.685 448.365 ;
        RECT 49.975 448.195 50.145 448.365 ;
        RECT 50.435 448.195 50.605 448.365 ;
        RECT 50.895 448.195 51.065 448.365 ;
        RECT 51.355 448.195 51.525 448.365 ;
        RECT 51.815 448.195 51.985 448.365 ;
        RECT 52.275 448.195 52.445 448.365 ;
        RECT 52.735 448.195 52.905 448.365 ;
        RECT 53.195 448.195 53.365 448.365 ;
        RECT 53.655 448.195 53.825 448.365 ;
        RECT 42.615 445.475 42.785 445.645 ;
        RECT 43.075 445.475 43.245 445.645 ;
        RECT 43.535 445.475 43.705 445.645 ;
        RECT 43.995 445.475 44.165 445.645 ;
        RECT 44.455 445.475 44.625 445.645 ;
        RECT 44.915 445.475 45.085 445.645 ;
        RECT 45.375 445.475 45.545 445.645 ;
        RECT 45.835 445.475 46.005 445.645 ;
        RECT 46.295 445.475 46.465 445.645 ;
        RECT 46.755 445.475 46.925 445.645 ;
        RECT 47.215 445.475 47.385 445.645 ;
        RECT 47.675 445.475 47.845 445.645 ;
        RECT 48.135 445.475 48.305 445.645 ;
        RECT 48.595 445.475 48.765 445.645 ;
        RECT 49.055 445.475 49.225 445.645 ;
        RECT 49.515 445.475 49.685 445.645 ;
        RECT 49.975 445.475 50.145 445.645 ;
        RECT 50.435 445.475 50.605 445.645 ;
        RECT 50.895 445.475 51.065 445.645 ;
        RECT 51.355 445.475 51.525 445.645 ;
        RECT 51.815 445.475 51.985 445.645 ;
        RECT 52.275 445.475 52.445 445.645 ;
        RECT 52.735 445.475 52.905 445.645 ;
        RECT 53.195 445.475 53.365 445.645 ;
        RECT 53.655 445.475 53.825 445.645 ;
        RECT 42.615 442.755 42.785 442.925 ;
        RECT 43.075 442.755 43.245 442.925 ;
        RECT 43.535 442.755 43.705 442.925 ;
        RECT 43.995 442.755 44.165 442.925 ;
        RECT 44.455 442.755 44.625 442.925 ;
        RECT 44.915 442.755 45.085 442.925 ;
        RECT 45.375 442.755 45.545 442.925 ;
        RECT 45.835 442.755 46.005 442.925 ;
        RECT 46.295 442.755 46.465 442.925 ;
        RECT 46.755 442.755 46.925 442.925 ;
        RECT 47.215 442.755 47.385 442.925 ;
        RECT 47.675 442.755 47.845 442.925 ;
        RECT 48.135 442.755 48.305 442.925 ;
        RECT 48.595 442.755 48.765 442.925 ;
        RECT 49.055 442.755 49.225 442.925 ;
        RECT 49.515 442.755 49.685 442.925 ;
        RECT 49.975 442.755 50.145 442.925 ;
        RECT 50.435 442.755 50.605 442.925 ;
        RECT 50.895 442.755 51.065 442.925 ;
        RECT 51.355 442.755 51.525 442.925 ;
        RECT 51.815 442.755 51.985 442.925 ;
        RECT 52.275 442.755 52.445 442.925 ;
        RECT 52.735 442.755 52.905 442.925 ;
        RECT 53.195 442.755 53.365 442.925 ;
        RECT 53.655 442.755 53.825 442.925 ;
        RECT 42.615 440.035 42.785 440.205 ;
        RECT 43.075 440.035 43.245 440.205 ;
        RECT 43.535 440.035 43.705 440.205 ;
        RECT 43.995 440.035 44.165 440.205 ;
        RECT 44.455 440.035 44.625 440.205 ;
        RECT 44.915 440.035 45.085 440.205 ;
        RECT 45.375 440.035 45.545 440.205 ;
        RECT 45.835 440.035 46.005 440.205 ;
        RECT 46.295 440.035 46.465 440.205 ;
        RECT 46.755 440.035 46.925 440.205 ;
        RECT 47.215 440.035 47.385 440.205 ;
        RECT 47.675 440.035 47.845 440.205 ;
        RECT 48.135 440.035 48.305 440.205 ;
        RECT 48.595 440.035 48.765 440.205 ;
        RECT 49.055 440.035 49.225 440.205 ;
        RECT 49.515 440.035 49.685 440.205 ;
        RECT 49.975 440.035 50.145 440.205 ;
        RECT 50.435 440.035 50.605 440.205 ;
        RECT 50.895 440.035 51.065 440.205 ;
        RECT 51.355 440.035 51.525 440.205 ;
        RECT 51.815 440.035 51.985 440.205 ;
        RECT 52.275 440.035 52.445 440.205 ;
        RECT 52.735 440.035 52.905 440.205 ;
        RECT 53.195 440.035 53.365 440.205 ;
        RECT 53.655 440.035 53.825 440.205 ;
        RECT 42.615 437.315 42.785 437.485 ;
        RECT 43.075 437.315 43.245 437.485 ;
        RECT 43.535 437.315 43.705 437.485 ;
        RECT 43.995 437.315 44.165 437.485 ;
        RECT 44.455 437.315 44.625 437.485 ;
        RECT 44.915 437.315 45.085 437.485 ;
        RECT 45.375 437.315 45.545 437.485 ;
        RECT 45.835 437.315 46.005 437.485 ;
        RECT 46.295 437.315 46.465 437.485 ;
        RECT 46.755 437.315 46.925 437.485 ;
        RECT 47.215 437.315 47.385 437.485 ;
        RECT 47.675 437.315 47.845 437.485 ;
        RECT 48.135 437.315 48.305 437.485 ;
        RECT 48.595 437.315 48.765 437.485 ;
        RECT 49.055 437.315 49.225 437.485 ;
        RECT 49.515 437.315 49.685 437.485 ;
        RECT 49.975 437.315 50.145 437.485 ;
        RECT 50.435 437.315 50.605 437.485 ;
        RECT 50.895 437.315 51.065 437.485 ;
        RECT 51.355 437.315 51.525 437.485 ;
        RECT 51.815 437.315 51.985 437.485 ;
        RECT 52.275 437.315 52.445 437.485 ;
        RECT 52.735 437.315 52.905 437.485 ;
        RECT 53.195 437.315 53.365 437.485 ;
        RECT 53.655 437.315 53.825 437.485 ;
        RECT 42.615 434.595 42.785 434.765 ;
        RECT 43.075 434.595 43.245 434.765 ;
        RECT 43.535 434.595 43.705 434.765 ;
        RECT 43.995 434.595 44.165 434.765 ;
        RECT 44.455 434.595 44.625 434.765 ;
        RECT 44.915 434.595 45.085 434.765 ;
        RECT 45.375 434.595 45.545 434.765 ;
        RECT 45.835 434.595 46.005 434.765 ;
        RECT 46.295 434.595 46.465 434.765 ;
        RECT 46.755 434.595 46.925 434.765 ;
        RECT 47.215 434.595 47.385 434.765 ;
        RECT 47.675 434.595 47.845 434.765 ;
        RECT 48.135 434.595 48.305 434.765 ;
        RECT 48.595 434.595 48.765 434.765 ;
        RECT 49.055 434.595 49.225 434.765 ;
        RECT 49.515 434.595 49.685 434.765 ;
        RECT 49.975 434.595 50.145 434.765 ;
        RECT 50.435 434.595 50.605 434.765 ;
        RECT 50.895 434.595 51.065 434.765 ;
        RECT 51.355 434.595 51.525 434.765 ;
        RECT 51.815 434.595 51.985 434.765 ;
        RECT 52.275 434.595 52.445 434.765 ;
        RECT 52.735 434.595 52.905 434.765 ;
        RECT 53.195 434.595 53.365 434.765 ;
        RECT 53.655 434.595 53.825 434.765 ;
        RECT 42.615 431.875 42.785 432.045 ;
        RECT 43.075 431.875 43.245 432.045 ;
        RECT 43.535 431.875 43.705 432.045 ;
        RECT 43.995 431.875 44.165 432.045 ;
        RECT 44.455 431.875 44.625 432.045 ;
        RECT 44.915 431.875 45.085 432.045 ;
        RECT 45.375 431.875 45.545 432.045 ;
        RECT 45.835 431.875 46.005 432.045 ;
        RECT 46.295 431.875 46.465 432.045 ;
        RECT 46.755 431.875 46.925 432.045 ;
        RECT 47.215 431.875 47.385 432.045 ;
        RECT 47.675 431.875 47.845 432.045 ;
        RECT 48.135 431.875 48.305 432.045 ;
        RECT 48.595 431.875 48.765 432.045 ;
        RECT 49.055 431.875 49.225 432.045 ;
        RECT 49.515 431.875 49.685 432.045 ;
        RECT 49.975 431.875 50.145 432.045 ;
        RECT 50.435 431.875 50.605 432.045 ;
        RECT 50.895 431.875 51.065 432.045 ;
        RECT 51.355 431.875 51.525 432.045 ;
        RECT 51.815 431.875 51.985 432.045 ;
        RECT 52.275 431.875 52.445 432.045 ;
        RECT 52.735 431.875 52.905 432.045 ;
        RECT 53.195 431.875 53.365 432.045 ;
        RECT 53.655 431.875 53.825 432.045 ;
        RECT 42.615 429.155 42.785 429.325 ;
        RECT 43.075 429.155 43.245 429.325 ;
        RECT 43.535 429.155 43.705 429.325 ;
        RECT 43.995 429.155 44.165 429.325 ;
        RECT 44.455 429.155 44.625 429.325 ;
        RECT 44.915 429.155 45.085 429.325 ;
        RECT 45.375 429.155 45.545 429.325 ;
        RECT 45.835 429.155 46.005 429.325 ;
        RECT 46.295 429.155 46.465 429.325 ;
        RECT 46.755 429.155 46.925 429.325 ;
        RECT 47.215 429.155 47.385 429.325 ;
        RECT 47.675 429.155 47.845 429.325 ;
        RECT 48.135 429.155 48.305 429.325 ;
        RECT 48.595 429.155 48.765 429.325 ;
        RECT 49.055 429.155 49.225 429.325 ;
        RECT 49.515 429.155 49.685 429.325 ;
        RECT 49.975 429.155 50.145 429.325 ;
        RECT 50.435 429.155 50.605 429.325 ;
        RECT 50.895 429.155 51.065 429.325 ;
        RECT 51.355 429.155 51.525 429.325 ;
        RECT 51.815 429.155 51.985 429.325 ;
        RECT 52.275 429.155 52.445 429.325 ;
        RECT 52.735 429.155 52.905 429.325 ;
        RECT 53.195 429.155 53.365 429.325 ;
        RECT 53.655 429.155 53.825 429.325 ;
        RECT 42.615 426.435 42.785 426.605 ;
        RECT 43.075 426.435 43.245 426.605 ;
        RECT 43.535 426.435 43.705 426.605 ;
        RECT 43.995 426.435 44.165 426.605 ;
        RECT 44.455 426.435 44.625 426.605 ;
        RECT 44.915 426.435 45.085 426.605 ;
        RECT 45.375 426.435 45.545 426.605 ;
        RECT 45.835 426.435 46.005 426.605 ;
        RECT 46.295 426.435 46.465 426.605 ;
        RECT 46.755 426.435 46.925 426.605 ;
        RECT 47.215 426.435 47.385 426.605 ;
        RECT 47.675 426.435 47.845 426.605 ;
        RECT 48.135 426.435 48.305 426.605 ;
        RECT 48.595 426.435 48.765 426.605 ;
        RECT 49.055 426.435 49.225 426.605 ;
        RECT 49.515 426.435 49.685 426.605 ;
        RECT 49.975 426.435 50.145 426.605 ;
        RECT 50.435 426.435 50.605 426.605 ;
        RECT 50.895 426.435 51.065 426.605 ;
        RECT 51.355 426.435 51.525 426.605 ;
        RECT 51.815 426.435 51.985 426.605 ;
        RECT 52.275 426.435 52.445 426.605 ;
        RECT 52.735 426.435 52.905 426.605 ;
        RECT 53.195 426.435 53.365 426.605 ;
        RECT 53.655 426.435 53.825 426.605 ;
        RECT 42.615 423.715 42.785 423.885 ;
        RECT 43.075 423.715 43.245 423.885 ;
        RECT 43.535 423.715 43.705 423.885 ;
        RECT 43.995 423.715 44.165 423.885 ;
        RECT 44.455 423.715 44.625 423.885 ;
        RECT 44.915 423.715 45.085 423.885 ;
        RECT 45.375 423.715 45.545 423.885 ;
        RECT 45.835 423.715 46.005 423.885 ;
        RECT 46.295 423.715 46.465 423.885 ;
        RECT 46.755 423.715 46.925 423.885 ;
        RECT 47.215 423.715 47.385 423.885 ;
        RECT 47.675 423.715 47.845 423.885 ;
        RECT 48.135 423.715 48.305 423.885 ;
        RECT 48.595 423.715 48.765 423.885 ;
        RECT 49.055 423.715 49.225 423.885 ;
        RECT 49.515 423.715 49.685 423.885 ;
        RECT 49.975 423.715 50.145 423.885 ;
        RECT 50.435 423.715 50.605 423.885 ;
        RECT 50.895 423.715 51.065 423.885 ;
        RECT 51.355 423.715 51.525 423.885 ;
        RECT 51.815 423.715 51.985 423.885 ;
        RECT 52.275 423.715 52.445 423.885 ;
        RECT 52.735 423.715 52.905 423.885 ;
        RECT 53.195 423.715 53.365 423.885 ;
        RECT 53.655 423.715 53.825 423.885 ;
        RECT 42.615 420.995 42.785 421.165 ;
        RECT 43.075 420.995 43.245 421.165 ;
        RECT 43.535 420.995 43.705 421.165 ;
        RECT 43.995 420.995 44.165 421.165 ;
        RECT 44.455 420.995 44.625 421.165 ;
        RECT 44.915 420.995 45.085 421.165 ;
        RECT 45.375 420.995 45.545 421.165 ;
        RECT 45.835 420.995 46.005 421.165 ;
        RECT 46.295 420.995 46.465 421.165 ;
        RECT 46.755 420.995 46.925 421.165 ;
        RECT 47.215 420.995 47.385 421.165 ;
        RECT 47.675 420.995 47.845 421.165 ;
        RECT 48.135 420.995 48.305 421.165 ;
        RECT 48.595 420.995 48.765 421.165 ;
        RECT 49.055 420.995 49.225 421.165 ;
        RECT 49.515 420.995 49.685 421.165 ;
        RECT 49.975 420.995 50.145 421.165 ;
        RECT 50.435 420.995 50.605 421.165 ;
        RECT 50.895 420.995 51.065 421.165 ;
        RECT 51.355 420.995 51.525 421.165 ;
        RECT 51.815 420.995 51.985 421.165 ;
        RECT 52.275 420.995 52.445 421.165 ;
        RECT 52.735 420.995 52.905 421.165 ;
        RECT 53.195 420.995 53.365 421.165 ;
        RECT 53.655 420.995 53.825 421.165 ;
        RECT 42.615 418.275 42.785 418.445 ;
        RECT 43.075 418.275 43.245 418.445 ;
        RECT 43.535 418.275 43.705 418.445 ;
        RECT 43.995 418.275 44.165 418.445 ;
        RECT 44.455 418.275 44.625 418.445 ;
        RECT 44.915 418.275 45.085 418.445 ;
        RECT 45.375 418.275 45.545 418.445 ;
        RECT 45.835 418.275 46.005 418.445 ;
        RECT 46.295 418.275 46.465 418.445 ;
        RECT 46.755 418.275 46.925 418.445 ;
        RECT 47.215 418.275 47.385 418.445 ;
        RECT 47.675 418.275 47.845 418.445 ;
        RECT 48.135 418.275 48.305 418.445 ;
        RECT 48.595 418.275 48.765 418.445 ;
        RECT 49.055 418.275 49.225 418.445 ;
        RECT 49.515 418.275 49.685 418.445 ;
        RECT 49.975 418.275 50.145 418.445 ;
        RECT 50.435 418.275 50.605 418.445 ;
        RECT 50.895 418.275 51.065 418.445 ;
        RECT 51.355 418.275 51.525 418.445 ;
        RECT 51.815 418.275 51.985 418.445 ;
        RECT 52.275 418.275 52.445 418.445 ;
        RECT 52.735 418.275 52.905 418.445 ;
        RECT 53.195 418.275 53.365 418.445 ;
        RECT 53.655 418.275 53.825 418.445 ;
        RECT 42.615 415.555 42.785 415.725 ;
        RECT 43.075 415.555 43.245 415.725 ;
        RECT 43.535 415.555 43.705 415.725 ;
        RECT 43.995 415.555 44.165 415.725 ;
        RECT 44.455 415.555 44.625 415.725 ;
        RECT 44.915 415.555 45.085 415.725 ;
        RECT 45.375 415.555 45.545 415.725 ;
        RECT 45.835 415.555 46.005 415.725 ;
        RECT 46.295 415.555 46.465 415.725 ;
        RECT 46.755 415.555 46.925 415.725 ;
        RECT 47.215 415.555 47.385 415.725 ;
        RECT 47.675 415.555 47.845 415.725 ;
        RECT 48.135 415.555 48.305 415.725 ;
        RECT 48.595 415.555 48.765 415.725 ;
        RECT 49.055 415.555 49.225 415.725 ;
        RECT 49.515 415.555 49.685 415.725 ;
        RECT 49.975 415.555 50.145 415.725 ;
        RECT 50.435 415.555 50.605 415.725 ;
        RECT 50.895 415.555 51.065 415.725 ;
        RECT 51.355 415.555 51.525 415.725 ;
        RECT 51.815 415.555 51.985 415.725 ;
        RECT 52.275 415.555 52.445 415.725 ;
        RECT 52.735 415.555 52.905 415.725 ;
        RECT 53.195 415.555 53.365 415.725 ;
        RECT 53.655 415.555 53.825 415.725 ;
        RECT 42.615 412.835 42.785 413.005 ;
        RECT 43.075 412.835 43.245 413.005 ;
        RECT 43.535 412.835 43.705 413.005 ;
        RECT 43.995 412.835 44.165 413.005 ;
        RECT 44.455 412.835 44.625 413.005 ;
        RECT 44.915 412.835 45.085 413.005 ;
        RECT 45.375 412.835 45.545 413.005 ;
        RECT 45.835 412.835 46.005 413.005 ;
        RECT 46.295 412.835 46.465 413.005 ;
        RECT 46.755 412.835 46.925 413.005 ;
        RECT 47.215 412.835 47.385 413.005 ;
        RECT 47.675 412.835 47.845 413.005 ;
        RECT 48.135 412.835 48.305 413.005 ;
        RECT 48.595 412.835 48.765 413.005 ;
        RECT 49.055 412.835 49.225 413.005 ;
        RECT 49.515 412.835 49.685 413.005 ;
        RECT 49.975 412.835 50.145 413.005 ;
        RECT 50.435 412.835 50.605 413.005 ;
        RECT 50.895 412.835 51.065 413.005 ;
        RECT 51.355 412.835 51.525 413.005 ;
        RECT 51.815 412.835 51.985 413.005 ;
        RECT 52.275 412.835 52.445 413.005 ;
        RECT 52.735 412.835 52.905 413.005 ;
        RECT 53.195 412.835 53.365 413.005 ;
        RECT 53.655 412.835 53.825 413.005 ;
        RECT 42.615 410.115 42.785 410.285 ;
        RECT 43.075 410.115 43.245 410.285 ;
        RECT 43.535 410.115 43.705 410.285 ;
        RECT 43.995 410.115 44.165 410.285 ;
        RECT 44.455 410.115 44.625 410.285 ;
        RECT 44.915 410.115 45.085 410.285 ;
        RECT 45.375 410.115 45.545 410.285 ;
        RECT 45.835 410.115 46.005 410.285 ;
        RECT 46.295 410.115 46.465 410.285 ;
        RECT 46.755 410.115 46.925 410.285 ;
        RECT 47.215 410.115 47.385 410.285 ;
        RECT 47.675 410.115 47.845 410.285 ;
        RECT 48.135 410.115 48.305 410.285 ;
        RECT 48.595 410.115 48.765 410.285 ;
        RECT 49.055 410.115 49.225 410.285 ;
        RECT 49.515 410.115 49.685 410.285 ;
        RECT 49.975 410.115 50.145 410.285 ;
        RECT 50.435 410.115 50.605 410.285 ;
        RECT 50.895 410.115 51.065 410.285 ;
        RECT 51.355 410.115 51.525 410.285 ;
        RECT 51.815 410.115 51.985 410.285 ;
        RECT 52.275 410.115 52.445 410.285 ;
        RECT 52.735 410.115 52.905 410.285 ;
        RECT 53.195 410.115 53.365 410.285 ;
        RECT 53.655 410.115 53.825 410.285 ;
        RECT 42.615 407.395 42.785 407.565 ;
        RECT 43.075 407.395 43.245 407.565 ;
        RECT 43.535 407.395 43.705 407.565 ;
        RECT 43.995 407.395 44.165 407.565 ;
        RECT 44.455 407.395 44.625 407.565 ;
        RECT 44.915 407.395 45.085 407.565 ;
        RECT 45.375 407.395 45.545 407.565 ;
        RECT 45.835 407.395 46.005 407.565 ;
        RECT 46.295 407.395 46.465 407.565 ;
        RECT 46.755 407.395 46.925 407.565 ;
        RECT 47.215 407.395 47.385 407.565 ;
        RECT 47.675 407.395 47.845 407.565 ;
        RECT 48.135 407.395 48.305 407.565 ;
        RECT 48.595 407.395 48.765 407.565 ;
        RECT 49.055 407.395 49.225 407.565 ;
        RECT 49.515 407.395 49.685 407.565 ;
        RECT 49.975 407.395 50.145 407.565 ;
        RECT 50.435 407.395 50.605 407.565 ;
        RECT 50.895 407.395 51.065 407.565 ;
        RECT 51.355 407.395 51.525 407.565 ;
        RECT 51.815 407.395 51.985 407.565 ;
        RECT 52.275 407.395 52.445 407.565 ;
        RECT 52.735 407.395 52.905 407.565 ;
        RECT 53.195 407.395 53.365 407.565 ;
        RECT 53.655 407.395 53.825 407.565 ;
        RECT 42.615 404.675 42.785 404.845 ;
        RECT 43.075 404.675 43.245 404.845 ;
        RECT 43.535 404.675 43.705 404.845 ;
        RECT 43.995 404.675 44.165 404.845 ;
        RECT 44.455 404.675 44.625 404.845 ;
        RECT 44.915 404.675 45.085 404.845 ;
        RECT 45.375 404.675 45.545 404.845 ;
        RECT 45.835 404.675 46.005 404.845 ;
        RECT 46.295 404.675 46.465 404.845 ;
        RECT 46.755 404.675 46.925 404.845 ;
        RECT 47.215 404.675 47.385 404.845 ;
        RECT 47.675 404.675 47.845 404.845 ;
        RECT 48.135 404.675 48.305 404.845 ;
        RECT 48.595 404.675 48.765 404.845 ;
        RECT 49.055 404.675 49.225 404.845 ;
        RECT 49.515 404.675 49.685 404.845 ;
        RECT 49.975 404.675 50.145 404.845 ;
        RECT 50.435 404.675 50.605 404.845 ;
        RECT 50.895 404.675 51.065 404.845 ;
        RECT 51.355 404.675 51.525 404.845 ;
        RECT 51.815 404.675 51.985 404.845 ;
        RECT 52.275 404.675 52.445 404.845 ;
        RECT 52.735 404.675 52.905 404.845 ;
        RECT 53.195 404.675 53.365 404.845 ;
        RECT 53.655 404.675 53.825 404.845 ;
        RECT 42.615 401.955 42.785 402.125 ;
        RECT 43.075 401.955 43.245 402.125 ;
        RECT 43.535 401.955 43.705 402.125 ;
        RECT 43.995 401.955 44.165 402.125 ;
        RECT 44.455 401.955 44.625 402.125 ;
        RECT 44.915 401.955 45.085 402.125 ;
        RECT 45.375 401.955 45.545 402.125 ;
        RECT 45.835 401.955 46.005 402.125 ;
        RECT 46.295 401.955 46.465 402.125 ;
        RECT 46.755 401.955 46.925 402.125 ;
        RECT 47.215 401.955 47.385 402.125 ;
        RECT 47.675 401.955 47.845 402.125 ;
        RECT 48.135 401.955 48.305 402.125 ;
        RECT 48.595 401.955 48.765 402.125 ;
        RECT 49.055 401.955 49.225 402.125 ;
        RECT 49.515 401.955 49.685 402.125 ;
        RECT 49.975 401.955 50.145 402.125 ;
        RECT 50.435 401.955 50.605 402.125 ;
        RECT 50.895 401.955 51.065 402.125 ;
        RECT 51.355 401.955 51.525 402.125 ;
        RECT 51.815 401.955 51.985 402.125 ;
        RECT 52.275 401.955 52.445 402.125 ;
        RECT 52.735 401.955 52.905 402.125 ;
        RECT 53.195 401.955 53.365 402.125 ;
        RECT 53.655 401.955 53.825 402.125 ;
        RECT 42.615 399.235 42.785 399.405 ;
        RECT 43.075 399.235 43.245 399.405 ;
        RECT 43.535 399.235 43.705 399.405 ;
        RECT 43.995 399.235 44.165 399.405 ;
        RECT 44.455 399.235 44.625 399.405 ;
        RECT 44.915 399.235 45.085 399.405 ;
        RECT 45.375 399.235 45.545 399.405 ;
        RECT 45.835 399.235 46.005 399.405 ;
        RECT 46.295 399.235 46.465 399.405 ;
        RECT 46.755 399.235 46.925 399.405 ;
        RECT 47.215 399.235 47.385 399.405 ;
        RECT 47.675 399.235 47.845 399.405 ;
        RECT 48.135 399.235 48.305 399.405 ;
        RECT 48.595 399.235 48.765 399.405 ;
        RECT 49.055 399.235 49.225 399.405 ;
        RECT 49.515 399.235 49.685 399.405 ;
        RECT 49.975 399.235 50.145 399.405 ;
        RECT 50.435 399.235 50.605 399.405 ;
        RECT 50.895 399.235 51.065 399.405 ;
        RECT 51.355 399.235 51.525 399.405 ;
        RECT 51.815 399.235 51.985 399.405 ;
        RECT 52.275 399.235 52.445 399.405 ;
        RECT 52.735 399.235 52.905 399.405 ;
        RECT 53.195 399.235 53.365 399.405 ;
        RECT 53.655 399.235 53.825 399.405 ;
        RECT 42.615 396.515 42.785 396.685 ;
        RECT 43.075 396.515 43.245 396.685 ;
        RECT 43.535 396.515 43.705 396.685 ;
        RECT 43.995 396.515 44.165 396.685 ;
        RECT 44.455 396.515 44.625 396.685 ;
        RECT 44.915 396.515 45.085 396.685 ;
        RECT 45.375 396.515 45.545 396.685 ;
        RECT 45.835 396.515 46.005 396.685 ;
        RECT 46.295 396.515 46.465 396.685 ;
        RECT 46.755 396.515 46.925 396.685 ;
        RECT 47.215 396.515 47.385 396.685 ;
        RECT 47.675 396.515 47.845 396.685 ;
        RECT 48.135 396.515 48.305 396.685 ;
        RECT 48.595 396.515 48.765 396.685 ;
        RECT 49.055 396.515 49.225 396.685 ;
        RECT 49.515 396.515 49.685 396.685 ;
        RECT 49.975 396.515 50.145 396.685 ;
        RECT 50.435 396.515 50.605 396.685 ;
        RECT 50.895 396.515 51.065 396.685 ;
        RECT 51.355 396.515 51.525 396.685 ;
        RECT 51.815 396.515 51.985 396.685 ;
        RECT 52.275 396.515 52.445 396.685 ;
        RECT 52.735 396.515 52.905 396.685 ;
        RECT 53.195 396.515 53.365 396.685 ;
        RECT 53.655 396.515 53.825 396.685 ;
        RECT 42.615 393.795 42.785 393.965 ;
        RECT 43.075 393.795 43.245 393.965 ;
        RECT 43.535 393.795 43.705 393.965 ;
        RECT 43.995 393.795 44.165 393.965 ;
        RECT 44.455 393.795 44.625 393.965 ;
        RECT 44.915 393.795 45.085 393.965 ;
        RECT 45.375 393.795 45.545 393.965 ;
        RECT 45.835 393.795 46.005 393.965 ;
        RECT 46.295 393.795 46.465 393.965 ;
        RECT 46.755 393.795 46.925 393.965 ;
        RECT 47.215 393.795 47.385 393.965 ;
        RECT 47.675 393.795 47.845 393.965 ;
        RECT 48.135 393.795 48.305 393.965 ;
        RECT 48.595 393.795 48.765 393.965 ;
        RECT 49.055 393.795 49.225 393.965 ;
        RECT 49.515 393.795 49.685 393.965 ;
        RECT 49.975 393.795 50.145 393.965 ;
        RECT 50.435 393.795 50.605 393.965 ;
        RECT 50.895 393.795 51.065 393.965 ;
        RECT 51.355 393.795 51.525 393.965 ;
        RECT 51.815 393.795 51.985 393.965 ;
        RECT 52.275 393.795 52.445 393.965 ;
        RECT 52.735 393.795 52.905 393.965 ;
        RECT 53.195 393.795 53.365 393.965 ;
        RECT 53.655 393.795 53.825 393.965 ;
        RECT 42.615 391.075 42.785 391.245 ;
        RECT 43.075 391.075 43.245 391.245 ;
        RECT 43.535 391.075 43.705 391.245 ;
        RECT 43.995 391.075 44.165 391.245 ;
        RECT 44.455 391.075 44.625 391.245 ;
        RECT 44.915 391.075 45.085 391.245 ;
        RECT 45.375 391.075 45.545 391.245 ;
        RECT 45.835 391.075 46.005 391.245 ;
        RECT 46.295 391.075 46.465 391.245 ;
        RECT 46.755 391.075 46.925 391.245 ;
        RECT 47.215 391.075 47.385 391.245 ;
        RECT 47.675 391.075 47.845 391.245 ;
        RECT 48.135 391.075 48.305 391.245 ;
        RECT 48.595 391.075 48.765 391.245 ;
        RECT 49.055 391.075 49.225 391.245 ;
        RECT 49.515 391.075 49.685 391.245 ;
        RECT 49.975 391.075 50.145 391.245 ;
        RECT 50.435 391.075 50.605 391.245 ;
        RECT 50.895 391.075 51.065 391.245 ;
        RECT 51.355 391.075 51.525 391.245 ;
        RECT 51.815 391.075 51.985 391.245 ;
        RECT 52.275 391.075 52.445 391.245 ;
        RECT 52.735 391.075 52.905 391.245 ;
        RECT 53.195 391.075 53.365 391.245 ;
        RECT 53.655 391.075 53.825 391.245 ;
        RECT 42.615 388.355 42.785 388.525 ;
        RECT 43.075 388.355 43.245 388.525 ;
        RECT 43.535 388.355 43.705 388.525 ;
        RECT 43.995 388.355 44.165 388.525 ;
        RECT 44.455 388.355 44.625 388.525 ;
        RECT 44.915 388.355 45.085 388.525 ;
        RECT 45.375 388.355 45.545 388.525 ;
        RECT 45.835 388.355 46.005 388.525 ;
        RECT 46.295 388.355 46.465 388.525 ;
        RECT 46.755 388.355 46.925 388.525 ;
        RECT 47.215 388.355 47.385 388.525 ;
        RECT 47.675 388.355 47.845 388.525 ;
        RECT 48.135 388.355 48.305 388.525 ;
        RECT 48.595 388.355 48.765 388.525 ;
        RECT 49.055 388.355 49.225 388.525 ;
        RECT 49.515 388.355 49.685 388.525 ;
        RECT 49.975 388.355 50.145 388.525 ;
        RECT 50.435 388.355 50.605 388.525 ;
        RECT 50.895 388.355 51.065 388.525 ;
        RECT 51.355 388.355 51.525 388.525 ;
        RECT 51.815 388.355 51.985 388.525 ;
        RECT 52.275 388.355 52.445 388.525 ;
        RECT 52.735 388.355 52.905 388.525 ;
        RECT 53.195 388.355 53.365 388.525 ;
        RECT 53.655 388.355 53.825 388.525 ;
        RECT 42.615 385.635 42.785 385.805 ;
        RECT 43.075 385.635 43.245 385.805 ;
        RECT 43.535 385.635 43.705 385.805 ;
        RECT 43.995 385.635 44.165 385.805 ;
        RECT 44.455 385.635 44.625 385.805 ;
        RECT 44.915 385.635 45.085 385.805 ;
        RECT 45.375 385.635 45.545 385.805 ;
        RECT 45.835 385.635 46.005 385.805 ;
        RECT 46.295 385.635 46.465 385.805 ;
        RECT 46.755 385.635 46.925 385.805 ;
        RECT 47.215 385.635 47.385 385.805 ;
        RECT 47.675 385.635 47.845 385.805 ;
        RECT 48.135 385.635 48.305 385.805 ;
        RECT 48.595 385.635 48.765 385.805 ;
        RECT 49.055 385.635 49.225 385.805 ;
        RECT 49.515 385.635 49.685 385.805 ;
        RECT 49.975 385.635 50.145 385.805 ;
        RECT 50.435 385.635 50.605 385.805 ;
        RECT 50.895 385.635 51.065 385.805 ;
        RECT 51.355 385.635 51.525 385.805 ;
        RECT 51.815 385.635 51.985 385.805 ;
        RECT 52.275 385.635 52.445 385.805 ;
        RECT 52.735 385.635 52.905 385.805 ;
        RECT 53.195 385.635 53.365 385.805 ;
        RECT 53.655 385.635 53.825 385.805 ;
        RECT 42.615 382.915 42.785 383.085 ;
        RECT 43.075 382.915 43.245 383.085 ;
        RECT 43.535 382.915 43.705 383.085 ;
        RECT 43.995 382.915 44.165 383.085 ;
        RECT 44.455 382.915 44.625 383.085 ;
        RECT 44.915 382.915 45.085 383.085 ;
        RECT 45.375 382.915 45.545 383.085 ;
        RECT 45.835 382.915 46.005 383.085 ;
        RECT 46.295 382.915 46.465 383.085 ;
        RECT 46.755 382.915 46.925 383.085 ;
        RECT 47.215 382.915 47.385 383.085 ;
        RECT 47.675 382.915 47.845 383.085 ;
        RECT 48.135 382.915 48.305 383.085 ;
        RECT 48.595 382.915 48.765 383.085 ;
        RECT 49.055 382.915 49.225 383.085 ;
        RECT 49.515 382.915 49.685 383.085 ;
        RECT 49.975 382.915 50.145 383.085 ;
        RECT 50.435 382.915 50.605 383.085 ;
        RECT 50.895 382.915 51.065 383.085 ;
        RECT 51.355 382.915 51.525 383.085 ;
        RECT 51.815 382.915 51.985 383.085 ;
        RECT 52.275 382.915 52.445 383.085 ;
        RECT 52.735 382.915 52.905 383.085 ;
        RECT 53.195 382.915 53.365 383.085 ;
        RECT 53.655 382.915 53.825 383.085 ;
        RECT 42.615 380.195 42.785 380.365 ;
        RECT 43.075 380.195 43.245 380.365 ;
        RECT 43.535 380.195 43.705 380.365 ;
        RECT 43.995 380.195 44.165 380.365 ;
        RECT 44.455 380.195 44.625 380.365 ;
        RECT 44.915 380.195 45.085 380.365 ;
        RECT 45.375 380.195 45.545 380.365 ;
        RECT 45.835 380.195 46.005 380.365 ;
        RECT 46.295 380.195 46.465 380.365 ;
        RECT 46.755 380.195 46.925 380.365 ;
        RECT 47.215 380.195 47.385 380.365 ;
        RECT 47.675 380.195 47.845 380.365 ;
        RECT 48.135 380.195 48.305 380.365 ;
        RECT 48.595 380.195 48.765 380.365 ;
        RECT 49.055 380.195 49.225 380.365 ;
        RECT 49.515 380.195 49.685 380.365 ;
        RECT 49.975 380.195 50.145 380.365 ;
        RECT 50.435 380.195 50.605 380.365 ;
        RECT 50.895 380.195 51.065 380.365 ;
        RECT 51.355 380.195 51.525 380.365 ;
        RECT 51.815 380.195 51.985 380.365 ;
        RECT 52.275 380.195 52.445 380.365 ;
        RECT 52.735 380.195 52.905 380.365 ;
        RECT 53.195 380.195 53.365 380.365 ;
        RECT 53.655 380.195 53.825 380.365 ;
        RECT 42.615 377.475 42.785 377.645 ;
        RECT 43.075 377.475 43.245 377.645 ;
        RECT 43.535 377.475 43.705 377.645 ;
        RECT 43.995 377.475 44.165 377.645 ;
        RECT 44.455 377.475 44.625 377.645 ;
        RECT 44.915 377.475 45.085 377.645 ;
        RECT 45.375 377.475 45.545 377.645 ;
        RECT 45.835 377.475 46.005 377.645 ;
        RECT 46.295 377.475 46.465 377.645 ;
        RECT 46.755 377.475 46.925 377.645 ;
        RECT 47.215 377.475 47.385 377.645 ;
        RECT 47.675 377.475 47.845 377.645 ;
        RECT 48.135 377.475 48.305 377.645 ;
        RECT 48.595 377.475 48.765 377.645 ;
        RECT 49.055 377.475 49.225 377.645 ;
        RECT 49.515 377.475 49.685 377.645 ;
        RECT 49.975 377.475 50.145 377.645 ;
        RECT 50.435 377.475 50.605 377.645 ;
        RECT 50.895 377.475 51.065 377.645 ;
        RECT 51.355 377.475 51.525 377.645 ;
        RECT 51.815 377.475 51.985 377.645 ;
        RECT 52.275 377.475 52.445 377.645 ;
        RECT 52.735 377.475 52.905 377.645 ;
        RECT 53.195 377.475 53.365 377.645 ;
        RECT 53.655 377.475 53.825 377.645 ;
        RECT 42.615 374.755 42.785 374.925 ;
        RECT 43.075 374.755 43.245 374.925 ;
        RECT 43.535 374.755 43.705 374.925 ;
        RECT 43.995 374.755 44.165 374.925 ;
        RECT 44.455 374.755 44.625 374.925 ;
        RECT 44.915 374.755 45.085 374.925 ;
        RECT 45.375 374.755 45.545 374.925 ;
        RECT 45.835 374.755 46.005 374.925 ;
        RECT 46.295 374.755 46.465 374.925 ;
        RECT 46.755 374.755 46.925 374.925 ;
        RECT 47.215 374.755 47.385 374.925 ;
        RECT 47.675 374.755 47.845 374.925 ;
        RECT 48.135 374.755 48.305 374.925 ;
        RECT 48.595 374.755 48.765 374.925 ;
        RECT 49.055 374.755 49.225 374.925 ;
        RECT 49.515 374.755 49.685 374.925 ;
        RECT 49.975 374.755 50.145 374.925 ;
        RECT 50.435 374.755 50.605 374.925 ;
        RECT 50.895 374.755 51.065 374.925 ;
        RECT 51.355 374.755 51.525 374.925 ;
        RECT 51.815 374.755 51.985 374.925 ;
        RECT 52.275 374.755 52.445 374.925 ;
        RECT 52.735 374.755 52.905 374.925 ;
        RECT 53.195 374.755 53.365 374.925 ;
        RECT 53.655 374.755 53.825 374.925 ;
        RECT 42.615 372.035 42.785 372.205 ;
        RECT 43.075 372.035 43.245 372.205 ;
        RECT 43.535 372.035 43.705 372.205 ;
        RECT 43.995 372.035 44.165 372.205 ;
        RECT 44.455 372.035 44.625 372.205 ;
        RECT 44.915 372.035 45.085 372.205 ;
        RECT 45.375 372.035 45.545 372.205 ;
        RECT 45.835 372.035 46.005 372.205 ;
        RECT 46.295 372.035 46.465 372.205 ;
        RECT 46.755 372.035 46.925 372.205 ;
        RECT 47.215 372.035 47.385 372.205 ;
        RECT 47.675 372.035 47.845 372.205 ;
        RECT 48.135 372.035 48.305 372.205 ;
        RECT 48.595 372.035 48.765 372.205 ;
        RECT 49.055 372.035 49.225 372.205 ;
        RECT 49.515 372.035 49.685 372.205 ;
        RECT 49.975 372.035 50.145 372.205 ;
        RECT 50.435 372.035 50.605 372.205 ;
        RECT 50.895 372.035 51.065 372.205 ;
        RECT 51.355 372.035 51.525 372.205 ;
        RECT 51.815 372.035 51.985 372.205 ;
        RECT 52.275 372.035 52.445 372.205 ;
        RECT 52.735 372.035 52.905 372.205 ;
        RECT 53.195 372.035 53.365 372.205 ;
        RECT 53.655 372.035 53.825 372.205 ;
        RECT 42.615 369.315 42.785 369.485 ;
        RECT 43.075 369.315 43.245 369.485 ;
        RECT 43.535 369.315 43.705 369.485 ;
        RECT 43.995 369.315 44.165 369.485 ;
        RECT 44.455 369.315 44.625 369.485 ;
        RECT 44.915 369.315 45.085 369.485 ;
        RECT 45.375 369.315 45.545 369.485 ;
        RECT 45.835 369.315 46.005 369.485 ;
        RECT 46.295 369.315 46.465 369.485 ;
        RECT 46.755 369.315 46.925 369.485 ;
        RECT 47.215 369.315 47.385 369.485 ;
        RECT 47.675 369.315 47.845 369.485 ;
        RECT 48.135 369.315 48.305 369.485 ;
        RECT 48.595 369.315 48.765 369.485 ;
        RECT 49.055 369.315 49.225 369.485 ;
        RECT 49.515 369.315 49.685 369.485 ;
        RECT 49.975 369.315 50.145 369.485 ;
        RECT 50.435 369.315 50.605 369.485 ;
        RECT 50.895 369.315 51.065 369.485 ;
        RECT 51.355 369.315 51.525 369.485 ;
        RECT 51.815 369.315 51.985 369.485 ;
        RECT 52.275 369.315 52.445 369.485 ;
        RECT 52.735 369.315 52.905 369.485 ;
        RECT 53.195 369.315 53.365 369.485 ;
        RECT 53.655 369.315 53.825 369.485 ;
        RECT 42.615 366.595 42.785 366.765 ;
        RECT 43.075 366.595 43.245 366.765 ;
        RECT 43.535 366.595 43.705 366.765 ;
        RECT 43.995 366.595 44.165 366.765 ;
        RECT 44.455 366.595 44.625 366.765 ;
        RECT 44.915 366.595 45.085 366.765 ;
        RECT 45.375 366.595 45.545 366.765 ;
        RECT 45.835 366.595 46.005 366.765 ;
        RECT 46.295 366.595 46.465 366.765 ;
        RECT 46.755 366.595 46.925 366.765 ;
        RECT 47.215 366.595 47.385 366.765 ;
        RECT 47.675 366.595 47.845 366.765 ;
        RECT 48.135 366.595 48.305 366.765 ;
        RECT 48.595 366.595 48.765 366.765 ;
        RECT 49.055 366.595 49.225 366.765 ;
        RECT 49.515 366.595 49.685 366.765 ;
        RECT 49.975 366.595 50.145 366.765 ;
        RECT 50.435 366.595 50.605 366.765 ;
        RECT 50.895 366.595 51.065 366.765 ;
        RECT 51.355 366.595 51.525 366.765 ;
        RECT 51.815 366.595 51.985 366.765 ;
        RECT 52.275 366.595 52.445 366.765 ;
        RECT 52.735 366.595 52.905 366.765 ;
        RECT 53.195 366.595 53.365 366.765 ;
        RECT 53.655 366.595 53.825 366.765 ;
        RECT 42.615 363.875 42.785 364.045 ;
        RECT 43.075 363.875 43.245 364.045 ;
        RECT 43.535 363.875 43.705 364.045 ;
        RECT 43.995 363.875 44.165 364.045 ;
        RECT 44.455 363.875 44.625 364.045 ;
        RECT 44.915 363.875 45.085 364.045 ;
        RECT 45.375 363.875 45.545 364.045 ;
        RECT 45.835 363.875 46.005 364.045 ;
        RECT 46.295 363.875 46.465 364.045 ;
        RECT 46.755 363.875 46.925 364.045 ;
        RECT 47.215 363.875 47.385 364.045 ;
        RECT 47.675 363.875 47.845 364.045 ;
        RECT 48.135 363.875 48.305 364.045 ;
        RECT 48.595 363.875 48.765 364.045 ;
        RECT 49.055 363.875 49.225 364.045 ;
        RECT 49.515 363.875 49.685 364.045 ;
        RECT 49.975 363.875 50.145 364.045 ;
        RECT 50.435 363.875 50.605 364.045 ;
        RECT 50.895 363.875 51.065 364.045 ;
        RECT 51.355 363.875 51.525 364.045 ;
        RECT 51.815 363.875 51.985 364.045 ;
        RECT 52.275 363.875 52.445 364.045 ;
        RECT 52.735 363.875 52.905 364.045 ;
        RECT 53.195 363.875 53.365 364.045 ;
        RECT 53.655 363.875 53.825 364.045 ;
        RECT 42.615 361.155 42.785 361.325 ;
        RECT 43.075 361.155 43.245 361.325 ;
        RECT 43.535 361.155 43.705 361.325 ;
        RECT 43.995 361.155 44.165 361.325 ;
        RECT 44.455 361.155 44.625 361.325 ;
        RECT 44.915 361.155 45.085 361.325 ;
        RECT 45.375 361.155 45.545 361.325 ;
        RECT 45.835 361.155 46.005 361.325 ;
        RECT 46.295 361.155 46.465 361.325 ;
        RECT 46.755 361.155 46.925 361.325 ;
        RECT 47.215 361.155 47.385 361.325 ;
        RECT 47.675 361.155 47.845 361.325 ;
        RECT 48.135 361.155 48.305 361.325 ;
        RECT 48.595 361.155 48.765 361.325 ;
        RECT 49.055 361.155 49.225 361.325 ;
        RECT 49.515 361.155 49.685 361.325 ;
        RECT 49.975 361.155 50.145 361.325 ;
        RECT 50.435 361.155 50.605 361.325 ;
        RECT 50.895 361.155 51.065 361.325 ;
        RECT 51.355 361.155 51.525 361.325 ;
        RECT 51.815 361.155 51.985 361.325 ;
        RECT 52.275 361.155 52.445 361.325 ;
        RECT 52.735 361.155 52.905 361.325 ;
        RECT 53.195 361.155 53.365 361.325 ;
        RECT 53.655 361.155 53.825 361.325 ;
        RECT 42.615 358.435 42.785 358.605 ;
        RECT 43.075 358.435 43.245 358.605 ;
        RECT 43.535 358.435 43.705 358.605 ;
        RECT 43.995 358.435 44.165 358.605 ;
        RECT 44.455 358.435 44.625 358.605 ;
        RECT 44.915 358.435 45.085 358.605 ;
        RECT 45.375 358.435 45.545 358.605 ;
        RECT 45.835 358.435 46.005 358.605 ;
        RECT 46.295 358.435 46.465 358.605 ;
        RECT 46.755 358.435 46.925 358.605 ;
        RECT 47.215 358.435 47.385 358.605 ;
        RECT 47.675 358.435 47.845 358.605 ;
        RECT 48.135 358.435 48.305 358.605 ;
        RECT 48.595 358.435 48.765 358.605 ;
        RECT 49.055 358.435 49.225 358.605 ;
        RECT 49.515 358.435 49.685 358.605 ;
        RECT 49.975 358.435 50.145 358.605 ;
        RECT 50.435 358.435 50.605 358.605 ;
        RECT 50.895 358.435 51.065 358.605 ;
        RECT 51.355 358.435 51.525 358.605 ;
        RECT 51.815 358.435 51.985 358.605 ;
        RECT 52.275 358.435 52.445 358.605 ;
        RECT 52.735 358.435 52.905 358.605 ;
        RECT 53.195 358.435 53.365 358.605 ;
        RECT 53.655 358.435 53.825 358.605 ;
        RECT 42.615 355.715 42.785 355.885 ;
        RECT 43.075 355.715 43.245 355.885 ;
        RECT 43.535 355.715 43.705 355.885 ;
        RECT 43.995 355.715 44.165 355.885 ;
        RECT 44.455 355.715 44.625 355.885 ;
        RECT 44.915 355.715 45.085 355.885 ;
        RECT 45.375 355.715 45.545 355.885 ;
        RECT 45.835 355.715 46.005 355.885 ;
        RECT 46.295 355.715 46.465 355.885 ;
        RECT 46.755 355.715 46.925 355.885 ;
        RECT 47.215 355.715 47.385 355.885 ;
        RECT 47.675 355.715 47.845 355.885 ;
        RECT 48.135 355.715 48.305 355.885 ;
        RECT 48.595 355.715 48.765 355.885 ;
        RECT 49.055 355.715 49.225 355.885 ;
        RECT 49.515 355.715 49.685 355.885 ;
        RECT 49.975 355.715 50.145 355.885 ;
        RECT 50.435 355.715 50.605 355.885 ;
        RECT 50.895 355.715 51.065 355.885 ;
        RECT 51.355 355.715 51.525 355.885 ;
        RECT 51.815 355.715 51.985 355.885 ;
        RECT 52.275 355.715 52.445 355.885 ;
        RECT 52.735 355.715 52.905 355.885 ;
        RECT 53.195 355.715 53.365 355.885 ;
        RECT 53.655 355.715 53.825 355.885 ;
        RECT 42.615 352.995 42.785 353.165 ;
        RECT 43.075 352.995 43.245 353.165 ;
        RECT 43.535 352.995 43.705 353.165 ;
        RECT 43.995 352.995 44.165 353.165 ;
        RECT 44.455 352.995 44.625 353.165 ;
        RECT 44.915 352.995 45.085 353.165 ;
        RECT 45.375 352.995 45.545 353.165 ;
        RECT 45.835 352.995 46.005 353.165 ;
        RECT 46.295 352.995 46.465 353.165 ;
        RECT 46.755 352.995 46.925 353.165 ;
        RECT 47.215 352.995 47.385 353.165 ;
        RECT 47.675 352.995 47.845 353.165 ;
        RECT 48.135 352.995 48.305 353.165 ;
        RECT 48.595 352.995 48.765 353.165 ;
        RECT 49.055 352.995 49.225 353.165 ;
        RECT 49.515 352.995 49.685 353.165 ;
        RECT 49.975 352.995 50.145 353.165 ;
        RECT 50.435 352.995 50.605 353.165 ;
        RECT 50.895 352.995 51.065 353.165 ;
        RECT 51.355 352.995 51.525 353.165 ;
        RECT 51.815 352.995 51.985 353.165 ;
        RECT 52.275 352.995 52.445 353.165 ;
        RECT 52.735 352.995 52.905 353.165 ;
        RECT 53.195 352.995 53.365 353.165 ;
        RECT 53.655 352.995 53.825 353.165 ;
        RECT 42.615 350.275 42.785 350.445 ;
        RECT 43.075 350.275 43.245 350.445 ;
        RECT 43.535 350.275 43.705 350.445 ;
        RECT 43.995 350.275 44.165 350.445 ;
        RECT 44.455 350.275 44.625 350.445 ;
        RECT 44.915 350.275 45.085 350.445 ;
        RECT 45.375 350.275 45.545 350.445 ;
        RECT 45.835 350.275 46.005 350.445 ;
        RECT 46.295 350.275 46.465 350.445 ;
        RECT 46.755 350.275 46.925 350.445 ;
        RECT 47.215 350.275 47.385 350.445 ;
        RECT 47.675 350.275 47.845 350.445 ;
        RECT 48.135 350.275 48.305 350.445 ;
        RECT 48.595 350.275 48.765 350.445 ;
        RECT 49.055 350.275 49.225 350.445 ;
        RECT 49.515 350.275 49.685 350.445 ;
        RECT 49.975 350.275 50.145 350.445 ;
        RECT 50.435 350.275 50.605 350.445 ;
        RECT 50.895 350.275 51.065 350.445 ;
        RECT 51.355 350.275 51.525 350.445 ;
        RECT 51.815 350.275 51.985 350.445 ;
        RECT 52.275 350.275 52.445 350.445 ;
        RECT 52.735 350.275 52.905 350.445 ;
        RECT 53.195 350.275 53.365 350.445 ;
        RECT 53.655 350.275 53.825 350.445 ;
        RECT 42.615 347.555 42.785 347.725 ;
        RECT 43.075 347.555 43.245 347.725 ;
        RECT 43.535 347.555 43.705 347.725 ;
        RECT 43.995 347.555 44.165 347.725 ;
        RECT 44.455 347.555 44.625 347.725 ;
        RECT 44.915 347.555 45.085 347.725 ;
        RECT 45.375 347.555 45.545 347.725 ;
        RECT 45.835 347.555 46.005 347.725 ;
        RECT 46.295 347.555 46.465 347.725 ;
        RECT 46.755 347.555 46.925 347.725 ;
        RECT 47.215 347.555 47.385 347.725 ;
        RECT 47.675 347.555 47.845 347.725 ;
        RECT 48.135 347.555 48.305 347.725 ;
        RECT 48.595 347.555 48.765 347.725 ;
        RECT 49.055 347.555 49.225 347.725 ;
        RECT 49.515 347.555 49.685 347.725 ;
        RECT 49.975 347.555 50.145 347.725 ;
        RECT 50.435 347.555 50.605 347.725 ;
        RECT 50.895 347.555 51.065 347.725 ;
        RECT 51.355 347.555 51.525 347.725 ;
        RECT 51.815 347.555 51.985 347.725 ;
        RECT 52.275 347.555 52.445 347.725 ;
        RECT 52.735 347.555 52.905 347.725 ;
        RECT 53.195 347.555 53.365 347.725 ;
        RECT 53.655 347.555 53.825 347.725 ;
        RECT 42.615 344.835 42.785 345.005 ;
        RECT 43.075 344.835 43.245 345.005 ;
        RECT 43.535 344.835 43.705 345.005 ;
        RECT 43.995 344.835 44.165 345.005 ;
        RECT 44.455 344.835 44.625 345.005 ;
        RECT 44.915 344.835 45.085 345.005 ;
        RECT 45.375 344.835 45.545 345.005 ;
        RECT 45.835 344.835 46.005 345.005 ;
        RECT 46.295 344.835 46.465 345.005 ;
        RECT 46.755 344.835 46.925 345.005 ;
        RECT 47.215 344.835 47.385 345.005 ;
        RECT 47.675 344.835 47.845 345.005 ;
        RECT 48.135 344.835 48.305 345.005 ;
        RECT 48.595 344.835 48.765 345.005 ;
        RECT 49.055 344.835 49.225 345.005 ;
        RECT 49.515 344.835 49.685 345.005 ;
        RECT 49.975 344.835 50.145 345.005 ;
        RECT 50.435 344.835 50.605 345.005 ;
        RECT 50.895 344.835 51.065 345.005 ;
        RECT 51.355 344.835 51.525 345.005 ;
        RECT 51.815 344.835 51.985 345.005 ;
        RECT 52.275 344.835 52.445 345.005 ;
        RECT 52.735 344.835 52.905 345.005 ;
        RECT 53.195 344.835 53.365 345.005 ;
        RECT 53.655 344.835 53.825 345.005 ;
        RECT 42.615 342.115 42.785 342.285 ;
        RECT 43.075 342.115 43.245 342.285 ;
        RECT 43.535 342.115 43.705 342.285 ;
        RECT 43.995 342.115 44.165 342.285 ;
        RECT 44.455 342.115 44.625 342.285 ;
        RECT 44.915 342.115 45.085 342.285 ;
        RECT 45.375 342.115 45.545 342.285 ;
        RECT 45.835 342.115 46.005 342.285 ;
        RECT 46.295 342.115 46.465 342.285 ;
        RECT 46.755 342.115 46.925 342.285 ;
        RECT 47.215 342.115 47.385 342.285 ;
        RECT 47.675 342.115 47.845 342.285 ;
        RECT 48.135 342.115 48.305 342.285 ;
        RECT 48.595 342.115 48.765 342.285 ;
        RECT 49.055 342.115 49.225 342.285 ;
        RECT 49.515 342.115 49.685 342.285 ;
        RECT 49.975 342.115 50.145 342.285 ;
        RECT 50.435 342.115 50.605 342.285 ;
        RECT 50.895 342.115 51.065 342.285 ;
        RECT 51.355 342.115 51.525 342.285 ;
        RECT 51.815 342.115 51.985 342.285 ;
        RECT 52.275 342.115 52.445 342.285 ;
        RECT 52.735 342.115 52.905 342.285 ;
        RECT 53.195 342.115 53.365 342.285 ;
        RECT 53.655 342.115 53.825 342.285 ;
        RECT 42.615 339.395 42.785 339.565 ;
        RECT 43.075 339.395 43.245 339.565 ;
        RECT 43.535 339.395 43.705 339.565 ;
        RECT 43.995 339.395 44.165 339.565 ;
        RECT 44.455 339.395 44.625 339.565 ;
        RECT 44.915 339.395 45.085 339.565 ;
        RECT 45.375 339.395 45.545 339.565 ;
        RECT 45.835 339.395 46.005 339.565 ;
        RECT 46.295 339.395 46.465 339.565 ;
        RECT 46.755 339.395 46.925 339.565 ;
        RECT 47.215 339.395 47.385 339.565 ;
        RECT 47.675 339.395 47.845 339.565 ;
        RECT 48.135 339.395 48.305 339.565 ;
        RECT 48.595 339.395 48.765 339.565 ;
        RECT 49.055 339.395 49.225 339.565 ;
        RECT 49.515 339.395 49.685 339.565 ;
        RECT 49.975 339.395 50.145 339.565 ;
        RECT 50.435 339.395 50.605 339.565 ;
        RECT 50.895 339.395 51.065 339.565 ;
        RECT 51.355 339.395 51.525 339.565 ;
        RECT 51.815 339.395 51.985 339.565 ;
        RECT 52.275 339.395 52.445 339.565 ;
        RECT 52.735 339.395 52.905 339.565 ;
        RECT 53.195 339.395 53.365 339.565 ;
        RECT 53.655 339.395 53.825 339.565 ;
        RECT 42.615 336.675 42.785 336.845 ;
        RECT 43.075 336.675 43.245 336.845 ;
        RECT 43.535 336.675 43.705 336.845 ;
        RECT 43.995 336.675 44.165 336.845 ;
        RECT 44.455 336.675 44.625 336.845 ;
        RECT 44.915 336.675 45.085 336.845 ;
        RECT 45.375 336.675 45.545 336.845 ;
        RECT 45.835 336.675 46.005 336.845 ;
        RECT 46.295 336.675 46.465 336.845 ;
        RECT 46.755 336.675 46.925 336.845 ;
        RECT 47.215 336.675 47.385 336.845 ;
        RECT 47.675 336.675 47.845 336.845 ;
        RECT 48.135 336.675 48.305 336.845 ;
        RECT 48.595 336.675 48.765 336.845 ;
        RECT 49.055 336.675 49.225 336.845 ;
        RECT 49.515 336.675 49.685 336.845 ;
        RECT 49.975 336.675 50.145 336.845 ;
        RECT 50.435 336.675 50.605 336.845 ;
        RECT 50.895 336.675 51.065 336.845 ;
        RECT 51.355 336.675 51.525 336.845 ;
        RECT 51.815 336.675 51.985 336.845 ;
        RECT 52.275 336.675 52.445 336.845 ;
        RECT 52.735 336.675 52.905 336.845 ;
        RECT 53.195 336.675 53.365 336.845 ;
        RECT 53.655 336.675 53.825 336.845 ;
        RECT 42.615 333.955 42.785 334.125 ;
        RECT 43.075 333.955 43.245 334.125 ;
        RECT 43.535 333.955 43.705 334.125 ;
        RECT 43.995 333.955 44.165 334.125 ;
        RECT 44.455 333.955 44.625 334.125 ;
        RECT 44.915 333.955 45.085 334.125 ;
        RECT 45.375 333.955 45.545 334.125 ;
        RECT 45.835 333.955 46.005 334.125 ;
        RECT 46.295 333.955 46.465 334.125 ;
        RECT 46.755 333.955 46.925 334.125 ;
        RECT 47.215 333.955 47.385 334.125 ;
        RECT 47.675 333.955 47.845 334.125 ;
        RECT 48.135 333.955 48.305 334.125 ;
        RECT 48.595 333.955 48.765 334.125 ;
        RECT 49.055 333.955 49.225 334.125 ;
        RECT 49.515 333.955 49.685 334.125 ;
        RECT 49.975 333.955 50.145 334.125 ;
        RECT 50.435 333.955 50.605 334.125 ;
        RECT 50.895 333.955 51.065 334.125 ;
        RECT 51.355 333.955 51.525 334.125 ;
        RECT 51.815 333.955 51.985 334.125 ;
        RECT 52.275 333.955 52.445 334.125 ;
        RECT 52.735 333.955 52.905 334.125 ;
        RECT 53.195 333.955 53.365 334.125 ;
        RECT 53.655 333.955 53.825 334.125 ;
        RECT 42.615 331.235 42.785 331.405 ;
        RECT 43.075 331.235 43.245 331.405 ;
        RECT 43.535 331.235 43.705 331.405 ;
        RECT 43.995 331.235 44.165 331.405 ;
        RECT 44.455 331.235 44.625 331.405 ;
        RECT 44.915 331.235 45.085 331.405 ;
        RECT 45.375 331.235 45.545 331.405 ;
        RECT 45.835 331.235 46.005 331.405 ;
        RECT 46.295 331.235 46.465 331.405 ;
        RECT 46.755 331.235 46.925 331.405 ;
        RECT 47.215 331.235 47.385 331.405 ;
        RECT 47.675 331.235 47.845 331.405 ;
        RECT 48.135 331.235 48.305 331.405 ;
        RECT 48.595 331.235 48.765 331.405 ;
        RECT 49.055 331.235 49.225 331.405 ;
        RECT 49.515 331.235 49.685 331.405 ;
        RECT 49.975 331.235 50.145 331.405 ;
        RECT 50.435 331.235 50.605 331.405 ;
        RECT 50.895 331.235 51.065 331.405 ;
        RECT 51.355 331.235 51.525 331.405 ;
        RECT 51.815 331.235 51.985 331.405 ;
        RECT 52.275 331.235 52.445 331.405 ;
        RECT 52.735 331.235 52.905 331.405 ;
        RECT 53.195 331.235 53.365 331.405 ;
        RECT 53.655 331.235 53.825 331.405 ;
        RECT 42.615 328.515 42.785 328.685 ;
        RECT 43.075 328.515 43.245 328.685 ;
        RECT 43.535 328.515 43.705 328.685 ;
        RECT 43.995 328.515 44.165 328.685 ;
        RECT 44.455 328.515 44.625 328.685 ;
        RECT 44.915 328.515 45.085 328.685 ;
        RECT 45.375 328.515 45.545 328.685 ;
        RECT 45.835 328.515 46.005 328.685 ;
        RECT 46.295 328.515 46.465 328.685 ;
        RECT 46.755 328.515 46.925 328.685 ;
        RECT 47.215 328.515 47.385 328.685 ;
        RECT 47.675 328.515 47.845 328.685 ;
        RECT 48.135 328.515 48.305 328.685 ;
        RECT 48.595 328.515 48.765 328.685 ;
        RECT 49.055 328.515 49.225 328.685 ;
        RECT 49.515 328.515 49.685 328.685 ;
        RECT 49.975 328.515 50.145 328.685 ;
        RECT 50.435 328.515 50.605 328.685 ;
        RECT 50.895 328.515 51.065 328.685 ;
        RECT 51.355 328.515 51.525 328.685 ;
        RECT 51.815 328.515 51.985 328.685 ;
        RECT 52.275 328.515 52.445 328.685 ;
        RECT 52.735 328.515 52.905 328.685 ;
        RECT 53.195 328.515 53.365 328.685 ;
        RECT 53.655 328.515 53.825 328.685 ;
        RECT 42.615 325.795 42.785 325.965 ;
        RECT 43.075 325.795 43.245 325.965 ;
        RECT 43.535 325.795 43.705 325.965 ;
        RECT 43.995 325.795 44.165 325.965 ;
        RECT 44.455 325.795 44.625 325.965 ;
        RECT 44.915 325.795 45.085 325.965 ;
        RECT 45.375 325.795 45.545 325.965 ;
        RECT 45.835 325.795 46.005 325.965 ;
        RECT 46.295 325.795 46.465 325.965 ;
        RECT 46.755 325.795 46.925 325.965 ;
        RECT 47.215 325.795 47.385 325.965 ;
        RECT 47.675 325.795 47.845 325.965 ;
        RECT 48.135 325.795 48.305 325.965 ;
        RECT 48.595 325.795 48.765 325.965 ;
        RECT 49.055 325.795 49.225 325.965 ;
        RECT 49.515 325.795 49.685 325.965 ;
        RECT 49.975 325.795 50.145 325.965 ;
        RECT 50.435 325.795 50.605 325.965 ;
        RECT 50.895 325.795 51.065 325.965 ;
        RECT 51.355 325.795 51.525 325.965 ;
        RECT 51.815 325.795 51.985 325.965 ;
        RECT 52.275 325.795 52.445 325.965 ;
        RECT 52.735 325.795 52.905 325.965 ;
        RECT 53.195 325.795 53.365 325.965 ;
        RECT 53.655 325.795 53.825 325.965 ;
        RECT 42.615 323.075 42.785 323.245 ;
        RECT 43.075 323.075 43.245 323.245 ;
        RECT 43.535 323.075 43.705 323.245 ;
        RECT 43.995 323.075 44.165 323.245 ;
        RECT 44.455 323.075 44.625 323.245 ;
        RECT 44.915 323.075 45.085 323.245 ;
        RECT 45.375 323.075 45.545 323.245 ;
        RECT 45.835 323.075 46.005 323.245 ;
        RECT 46.295 323.075 46.465 323.245 ;
        RECT 46.755 323.075 46.925 323.245 ;
        RECT 47.215 323.075 47.385 323.245 ;
        RECT 47.675 323.075 47.845 323.245 ;
        RECT 48.135 323.075 48.305 323.245 ;
        RECT 48.595 323.075 48.765 323.245 ;
        RECT 49.055 323.075 49.225 323.245 ;
        RECT 49.515 323.075 49.685 323.245 ;
        RECT 49.975 323.075 50.145 323.245 ;
        RECT 50.435 323.075 50.605 323.245 ;
        RECT 50.895 323.075 51.065 323.245 ;
        RECT 51.355 323.075 51.525 323.245 ;
        RECT 51.815 323.075 51.985 323.245 ;
        RECT 52.275 323.075 52.445 323.245 ;
        RECT 52.735 323.075 52.905 323.245 ;
        RECT 53.195 323.075 53.365 323.245 ;
        RECT 53.655 323.075 53.825 323.245 ;
        RECT 42.615 320.355 42.785 320.525 ;
        RECT 43.075 320.355 43.245 320.525 ;
        RECT 43.535 320.355 43.705 320.525 ;
        RECT 43.995 320.355 44.165 320.525 ;
        RECT 44.455 320.355 44.625 320.525 ;
        RECT 44.915 320.355 45.085 320.525 ;
        RECT 45.375 320.355 45.545 320.525 ;
        RECT 45.835 320.355 46.005 320.525 ;
        RECT 46.295 320.355 46.465 320.525 ;
        RECT 46.755 320.355 46.925 320.525 ;
        RECT 47.215 320.355 47.385 320.525 ;
        RECT 47.675 320.355 47.845 320.525 ;
        RECT 48.135 320.355 48.305 320.525 ;
        RECT 48.595 320.355 48.765 320.525 ;
        RECT 49.055 320.355 49.225 320.525 ;
        RECT 49.515 320.355 49.685 320.525 ;
        RECT 49.975 320.355 50.145 320.525 ;
        RECT 50.435 320.355 50.605 320.525 ;
        RECT 50.895 320.355 51.065 320.525 ;
        RECT 51.355 320.355 51.525 320.525 ;
        RECT 51.815 320.355 51.985 320.525 ;
        RECT 52.275 320.355 52.445 320.525 ;
        RECT 52.735 320.355 52.905 320.525 ;
        RECT 53.195 320.355 53.365 320.525 ;
        RECT 53.655 320.355 53.825 320.525 ;
        RECT 42.615 317.635 42.785 317.805 ;
        RECT 43.075 317.635 43.245 317.805 ;
        RECT 43.535 317.635 43.705 317.805 ;
        RECT 43.995 317.635 44.165 317.805 ;
        RECT 44.455 317.635 44.625 317.805 ;
        RECT 44.915 317.635 45.085 317.805 ;
        RECT 45.375 317.635 45.545 317.805 ;
        RECT 45.835 317.635 46.005 317.805 ;
        RECT 46.295 317.635 46.465 317.805 ;
        RECT 46.755 317.635 46.925 317.805 ;
        RECT 47.215 317.635 47.385 317.805 ;
        RECT 47.675 317.635 47.845 317.805 ;
        RECT 48.135 317.635 48.305 317.805 ;
        RECT 48.595 317.635 48.765 317.805 ;
        RECT 49.055 317.635 49.225 317.805 ;
        RECT 49.515 317.635 49.685 317.805 ;
        RECT 49.975 317.635 50.145 317.805 ;
        RECT 50.435 317.635 50.605 317.805 ;
        RECT 50.895 317.635 51.065 317.805 ;
        RECT 51.355 317.635 51.525 317.805 ;
        RECT 51.815 317.635 51.985 317.805 ;
        RECT 52.275 317.635 52.445 317.805 ;
        RECT 52.735 317.635 52.905 317.805 ;
        RECT 53.195 317.635 53.365 317.805 ;
        RECT 53.655 317.635 53.825 317.805 ;
        RECT 42.615 314.915 42.785 315.085 ;
        RECT 43.075 314.915 43.245 315.085 ;
        RECT 43.535 314.915 43.705 315.085 ;
        RECT 43.995 314.915 44.165 315.085 ;
        RECT 44.455 314.915 44.625 315.085 ;
        RECT 44.915 314.915 45.085 315.085 ;
        RECT 45.375 314.915 45.545 315.085 ;
        RECT 45.835 314.915 46.005 315.085 ;
        RECT 46.295 314.915 46.465 315.085 ;
        RECT 46.755 314.915 46.925 315.085 ;
        RECT 47.215 314.915 47.385 315.085 ;
        RECT 47.675 314.915 47.845 315.085 ;
        RECT 48.135 314.915 48.305 315.085 ;
        RECT 48.595 314.915 48.765 315.085 ;
        RECT 49.055 314.915 49.225 315.085 ;
        RECT 49.515 314.915 49.685 315.085 ;
        RECT 49.975 314.915 50.145 315.085 ;
        RECT 50.435 314.915 50.605 315.085 ;
        RECT 50.895 314.915 51.065 315.085 ;
        RECT 51.355 314.915 51.525 315.085 ;
        RECT 51.815 314.915 51.985 315.085 ;
        RECT 52.275 314.915 52.445 315.085 ;
        RECT 52.735 314.915 52.905 315.085 ;
        RECT 53.195 314.915 53.365 315.085 ;
        RECT 53.655 314.915 53.825 315.085 ;
        RECT 42.615 312.195 42.785 312.365 ;
        RECT 43.075 312.195 43.245 312.365 ;
        RECT 43.535 312.195 43.705 312.365 ;
        RECT 43.995 312.195 44.165 312.365 ;
        RECT 44.455 312.195 44.625 312.365 ;
        RECT 44.915 312.195 45.085 312.365 ;
        RECT 45.375 312.195 45.545 312.365 ;
        RECT 45.835 312.195 46.005 312.365 ;
        RECT 46.295 312.195 46.465 312.365 ;
        RECT 46.755 312.195 46.925 312.365 ;
        RECT 47.215 312.195 47.385 312.365 ;
        RECT 47.675 312.195 47.845 312.365 ;
        RECT 48.135 312.195 48.305 312.365 ;
        RECT 48.595 312.195 48.765 312.365 ;
        RECT 49.055 312.195 49.225 312.365 ;
        RECT 49.515 312.195 49.685 312.365 ;
        RECT 49.975 312.195 50.145 312.365 ;
        RECT 50.435 312.195 50.605 312.365 ;
        RECT 50.895 312.195 51.065 312.365 ;
        RECT 51.355 312.195 51.525 312.365 ;
        RECT 51.815 312.195 51.985 312.365 ;
        RECT 52.275 312.195 52.445 312.365 ;
        RECT 52.735 312.195 52.905 312.365 ;
        RECT 53.195 312.195 53.365 312.365 ;
        RECT 53.655 312.195 53.825 312.365 ;
        RECT 42.615 309.475 42.785 309.645 ;
        RECT 43.075 309.475 43.245 309.645 ;
        RECT 43.535 309.475 43.705 309.645 ;
        RECT 43.995 309.475 44.165 309.645 ;
        RECT 44.455 309.475 44.625 309.645 ;
        RECT 44.915 309.475 45.085 309.645 ;
        RECT 45.375 309.475 45.545 309.645 ;
        RECT 45.835 309.475 46.005 309.645 ;
        RECT 46.295 309.475 46.465 309.645 ;
        RECT 46.755 309.475 46.925 309.645 ;
        RECT 47.215 309.475 47.385 309.645 ;
        RECT 47.675 309.475 47.845 309.645 ;
        RECT 48.135 309.475 48.305 309.645 ;
        RECT 48.595 309.475 48.765 309.645 ;
        RECT 49.055 309.475 49.225 309.645 ;
        RECT 49.515 309.475 49.685 309.645 ;
        RECT 49.975 309.475 50.145 309.645 ;
        RECT 50.435 309.475 50.605 309.645 ;
        RECT 50.895 309.475 51.065 309.645 ;
        RECT 51.355 309.475 51.525 309.645 ;
        RECT 51.815 309.475 51.985 309.645 ;
        RECT 52.275 309.475 52.445 309.645 ;
        RECT 52.735 309.475 52.905 309.645 ;
        RECT 53.195 309.475 53.365 309.645 ;
        RECT 53.655 309.475 53.825 309.645 ;
        RECT 42.615 306.755 42.785 306.925 ;
        RECT 43.075 306.755 43.245 306.925 ;
        RECT 43.535 306.755 43.705 306.925 ;
        RECT 43.995 306.755 44.165 306.925 ;
        RECT 44.455 306.755 44.625 306.925 ;
        RECT 44.915 306.755 45.085 306.925 ;
        RECT 45.375 306.755 45.545 306.925 ;
        RECT 45.835 306.755 46.005 306.925 ;
        RECT 46.295 306.755 46.465 306.925 ;
        RECT 46.755 306.755 46.925 306.925 ;
        RECT 47.215 306.755 47.385 306.925 ;
        RECT 47.675 306.755 47.845 306.925 ;
        RECT 48.135 306.755 48.305 306.925 ;
        RECT 48.595 306.755 48.765 306.925 ;
        RECT 49.055 306.755 49.225 306.925 ;
        RECT 49.515 306.755 49.685 306.925 ;
        RECT 49.975 306.755 50.145 306.925 ;
        RECT 50.435 306.755 50.605 306.925 ;
        RECT 50.895 306.755 51.065 306.925 ;
        RECT 51.355 306.755 51.525 306.925 ;
        RECT 51.815 306.755 51.985 306.925 ;
        RECT 52.275 306.755 52.445 306.925 ;
        RECT 52.735 306.755 52.905 306.925 ;
        RECT 53.195 306.755 53.365 306.925 ;
        RECT 53.655 306.755 53.825 306.925 ;
        RECT 42.615 304.035 42.785 304.205 ;
        RECT 43.075 304.035 43.245 304.205 ;
        RECT 43.535 304.035 43.705 304.205 ;
        RECT 43.995 304.035 44.165 304.205 ;
        RECT 44.455 304.035 44.625 304.205 ;
        RECT 44.915 304.035 45.085 304.205 ;
        RECT 45.375 304.035 45.545 304.205 ;
        RECT 45.835 304.035 46.005 304.205 ;
        RECT 46.295 304.035 46.465 304.205 ;
        RECT 46.755 304.035 46.925 304.205 ;
        RECT 47.215 304.035 47.385 304.205 ;
        RECT 47.675 304.035 47.845 304.205 ;
        RECT 48.135 304.035 48.305 304.205 ;
        RECT 48.595 304.035 48.765 304.205 ;
        RECT 49.055 304.035 49.225 304.205 ;
        RECT 49.515 304.035 49.685 304.205 ;
        RECT 49.975 304.035 50.145 304.205 ;
        RECT 50.435 304.035 50.605 304.205 ;
        RECT 50.895 304.035 51.065 304.205 ;
        RECT 51.355 304.035 51.525 304.205 ;
        RECT 51.815 304.035 51.985 304.205 ;
        RECT 52.275 304.035 52.445 304.205 ;
        RECT 52.735 304.035 52.905 304.205 ;
        RECT 53.195 304.035 53.365 304.205 ;
        RECT 53.655 304.035 53.825 304.205 ;
        RECT 42.615 301.315 42.785 301.485 ;
        RECT 43.075 301.315 43.245 301.485 ;
        RECT 43.535 301.315 43.705 301.485 ;
        RECT 43.995 301.315 44.165 301.485 ;
        RECT 44.455 301.315 44.625 301.485 ;
        RECT 44.915 301.315 45.085 301.485 ;
        RECT 45.375 301.315 45.545 301.485 ;
        RECT 45.835 301.315 46.005 301.485 ;
        RECT 46.295 301.315 46.465 301.485 ;
        RECT 46.755 301.315 46.925 301.485 ;
        RECT 47.215 301.315 47.385 301.485 ;
        RECT 47.675 301.315 47.845 301.485 ;
        RECT 48.135 301.315 48.305 301.485 ;
        RECT 48.595 301.315 48.765 301.485 ;
        RECT 49.055 301.315 49.225 301.485 ;
        RECT 49.515 301.315 49.685 301.485 ;
        RECT 49.975 301.315 50.145 301.485 ;
        RECT 50.435 301.315 50.605 301.485 ;
        RECT 50.895 301.315 51.065 301.485 ;
        RECT 51.355 301.315 51.525 301.485 ;
        RECT 51.815 301.315 51.985 301.485 ;
        RECT 52.275 301.315 52.445 301.485 ;
        RECT 52.735 301.315 52.905 301.485 ;
        RECT 53.195 301.315 53.365 301.485 ;
        RECT 53.655 301.315 53.825 301.485 ;
        RECT 42.615 298.595 42.785 298.765 ;
        RECT 43.075 298.595 43.245 298.765 ;
        RECT 43.535 298.595 43.705 298.765 ;
        RECT 43.995 298.595 44.165 298.765 ;
        RECT 44.455 298.595 44.625 298.765 ;
        RECT 44.915 298.595 45.085 298.765 ;
        RECT 45.375 298.595 45.545 298.765 ;
        RECT 45.835 298.595 46.005 298.765 ;
        RECT 46.295 298.595 46.465 298.765 ;
        RECT 46.755 298.595 46.925 298.765 ;
        RECT 47.215 298.595 47.385 298.765 ;
        RECT 47.675 298.595 47.845 298.765 ;
        RECT 48.135 298.595 48.305 298.765 ;
        RECT 48.595 298.595 48.765 298.765 ;
        RECT 49.055 298.595 49.225 298.765 ;
        RECT 49.515 298.595 49.685 298.765 ;
        RECT 49.975 298.595 50.145 298.765 ;
        RECT 50.435 298.595 50.605 298.765 ;
        RECT 50.895 298.595 51.065 298.765 ;
        RECT 51.355 298.595 51.525 298.765 ;
        RECT 51.815 298.595 51.985 298.765 ;
        RECT 52.275 298.595 52.445 298.765 ;
        RECT 52.735 298.595 52.905 298.765 ;
        RECT 53.195 298.595 53.365 298.765 ;
        RECT 53.655 298.595 53.825 298.765 ;
        RECT 42.615 295.875 42.785 296.045 ;
        RECT 43.075 295.875 43.245 296.045 ;
        RECT 43.535 295.875 43.705 296.045 ;
        RECT 43.995 295.875 44.165 296.045 ;
        RECT 44.455 295.875 44.625 296.045 ;
        RECT 44.915 295.875 45.085 296.045 ;
        RECT 45.375 295.875 45.545 296.045 ;
        RECT 45.835 295.875 46.005 296.045 ;
        RECT 46.295 295.875 46.465 296.045 ;
        RECT 46.755 295.875 46.925 296.045 ;
        RECT 47.215 295.875 47.385 296.045 ;
        RECT 47.675 295.875 47.845 296.045 ;
        RECT 48.135 295.875 48.305 296.045 ;
        RECT 48.595 295.875 48.765 296.045 ;
        RECT 49.055 295.875 49.225 296.045 ;
        RECT 49.515 295.875 49.685 296.045 ;
        RECT 49.975 295.875 50.145 296.045 ;
        RECT 50.435 295.875 50.605 296.045 ;
        RECT 50.895 295.875 51.065 296.045 ;
        RECT 51.355 295.875 51.525 296.045 ;
        RECT 51.815 295.875 51.985 296.045 ;
        RECT 52.275 295.875 52.445 296.045 ;
        RECT 52.735 295.875 52.905 296.045 ;
        RECT 53.195 295.875 53.365 296.045 ;
        RECT 53.655 295.875 53.825 296.045 ;
        RECT 42.615 293.155 42.785 293.325 ;
        RECT 43.075 293.155 43.245 293.325 ;
        RECT 43.535 293.155 43.705 293.325 ;
        RECT 43.995 293.155 44.165 293.325 ;
        RECT 44.455 293.155 44.625 293.325 ;
        RECT 44.915 293.155 45.085 293.325 ;
        RECT 45.375 293.155 45.545 293.325 ;
        RECT 45.835 293.155 46.005 293.325 ;
        RECT 46.295 293.155 46.465 293.325 ;
        RECT 46.755 293.155 46.925 293.325 ;
        RECT 47.215 293.155 47.385 293.325 ;
        RECT 47.675 293.155 47.845 293.325 ;
        RECT 48.135 293.155 48.305 293.325 ;
        RECT 48.595 293.155 48.765 293.325 ;
        RECT 49.055 293.155 49.225 293.325 ;
        RECT 49.515 293.155 49.685 293.325 ;
        RECT 49.975 293.155 50.145 293.325 ;
        RECT 50.435 293.155 50.605 293.325 ;
        RECT 50.895 293.155 51.065 293.325 ;
        RECT 51.355 293.155 51.525 293.325 ;
        RECT 51.815 293.155 51.985 293.325 ;
        RECT 52.275 293.155 52.445 293.325 ;
        RECT 52.735 293.155 52.905 293.325 ;
        RECT 53.195 293.155 53.365 293.325 ;
        RECT 53.655 293.155 53.825 293.325 ;
        RECT 42.615 290.435 42.785 290.605 ;
        RECT 43.075 290.435 43.245 290.605 ;
        RECT 43.535 290.435 43.705 290.605 ;
        RECT 43.995 290.435 44.165 290.605 ;
        RECT 44.455 290.435 44.625 290.605 ;
        RECT 44.915 290.435 45.085 290.605 ;
        RECT 45.375 290.435 45.545 290.605 ;
        RECT 45.835 290.435 46.005 290.605 ;
        RECT 46.295 290.435 46.465 290.605 ;
        RECT 46.755 290.435 46.925 290.605 ;
        RECT 47.215 290.435 47.385 290.605 ;
        RECT 47.675 290.435 47.845 290.605 ;
        RECT 48.135 290.435 48.305 290.605 ;
        RECT 48.595 290.435 48.765 290.605 ;
        RECT 49.055 290.435 49.225 290.605 ;
        RECT 49.515 290.435 49.685 290.605 ;
        RECT 49.975 290.435 50.145 290.605 ;
        RECT 50.435 290.435 50.605 290.605 ;
        RECT 50.895 290.435 51.065 290.605 ;
        RECT 51.355 290.435 51.525 290.605 ;
        RECT 51.815 290.435 51.985 290.605 ;
        RECT 52.275 290.435 52.445 290.605 ;
        RECT 52.735 290.435 52.905 290.605 ;
        RECT 53.195 290.435 53.365 290.605 ;
        RECT 53.655 290.435 53.825 290.605 ;
        RECT 42.615 287.715 42.785 287.885 ;
        RECT 43.075 287.715 43.245 287.885 ;
        RECT 43.535 287.715 43.705 287.885 ;
        RECT 43.995 287.715 44.165 287.885 ;
        RECT 44.455 287.715 44.625 287.885 ;
        RECT 44.915 287.715 45.085 287.885 ;
        RECT 45.375 287.715 45.545 287.885 ;
        RECT 45.835 287.715 46.005 287.885 ;
        RECT 46.295 287.715 46.465 287.885 ;
        RECT 46.755 287.715 46.925 287.885 ;
        RECT 47.215 287.715 47.385 287.885 ;
        RECT 47.675 287.715 47.845 287.885 ;
        RECT 48.135 287.715 48.305 287.885 ;
        RECT 48.595 287.715 48.765 287.885 ;
        RECT 49.055 287.715 49.225 287.885 ;
        RECT 49.515 287.715 49.685 287.885 ;
        RECT 49.975 287.715 50.145 287.885 ;
        RECT 50.435 287.715 50.605 287.885 ;
        RECT 50.895 287.715 51.065 287.885 ;
        RECT 51.355 287.715 51.525 287.885 ;
        RECT 51.815 287.715 51.985 287.885 ;
        RECT 52.275 287.715 52.445 287.885 ;
        RECT 52.735 287.715 52.905 287.885 ;
        RECT 53.195 287.715 53.365 287.885 ;
        RECT 53.655 287.715 53.825 287.885 ;
        RECT 42.615 284.995 42.785 285.165 ;
        RECT 43.075 284.995 43.245 285.165 ;
        RECT 43.535 284.995 43.705 285.165 ;
        RECT 43.995 284.995 44.165 285.165 ;
        RECT 44.455 284.995 44.625 285.165 ;
        RECT 44.915 284.995 45.085 285.165 ;
        RECT 45.375 284.995 45.545 285.165 ;
        RECT 45.835 284.995 46.005 285.165 ;
        RECT 46.295 284.995 46.465 285.165 ;
        RECT 46.755 284.995 46.925 285.165 ;
        RECT 47.215 284.995 47.385 285.165 ;
        RECT 47.675 284.995 47.845 285.165 ;
        RECT 48.135 284.995 48.305 285.165 ;
        RECT 48.595 284.995 48.765 285.165 ;
        RECT 49.055 284.995 49.225 285.165 ;
        RECT 49.515 284.995 49.685 285.165 ;
        RECT 49.975 284.995 50.145 285.165 ;
        RECT 50.435 284.995 50.605 285.165 ;
        RECT 50.895 284.995 51.065 285.165 ;
        RECT 51.355 284.995 51.525 285.165 ;
        RECT 51.815 284.995 51.985 285.165 ;
        RECT 52.275 284.995 52.445 285.165 ;
        RECT 52.735 284.995 52.905 285.165 ;
        RECT 53.195 284.995 53.365 285.165 ;
        RECT 53.655 284.995 53.825 285.165 ;
        RECT 42.615 282.275 42.785 282.445 ;
        RECT 43.075 282.275 43.245 282.445 ;
        RECT 43.535 282.275 43.705 282.445 ;
        RECT 43.995 282.275 44.165 282.445 ;
        RECT 44.455 282.275 44.625 282.445 ;
        RECT 44.915 282.275 45.085 282.445 ;
        RECT 45.375 282.275 45.545 282.445 ;
        RECT 45.835 282.275 46.005 282.445 ;
        RECT 46.295 282.275 46.465 282.445 ;
        RECT 46.755 282.275 46.925 282.445 ;
        RECT 47.215 282.275 47.385 282.445 ;
        RECT 47.675 282.275 47.845 282.445 ;
        RECT 48.135 282.275 48.305 282.445 ;
        RECT 48.595 282.275 48.765 282.445 ;
        RECT 49.055 282.275 49.225 282.445 ;
        RECT 49.515 282.275 49.685 282.445 ;
        RECT 49.975 282.275 50.145 282.445 ;
        RECT 50.435 282.275 50.605 282.445 ;
        RECT 50.895 282.275 51.065 282.445 ;
        RECT 51.355 282.275 51.525 282.445 ;
        RECT 51.815 282.275 51.985 282.445 ;
        RECT 52.275 282.275 52.445 282.445 ;
        RECT 52.735 282.275 52.905 282.445 ;
        RECT 53.195 282.275 53.365 282.445 ;
        RECT 53.655 282.275 53.825 282.445 ;
        RECT 42.615 279.555 42.785 279.725 ;
        RECT 43.075 279.555 43.245 279.725 ;
        RECT 43.535 279.555 43.705 279.725 ;
        RECT 43.995 279.555 44.165 279.725 ;
        RECT 44.455 279.555 44.625 279.725 ;
        RECT 44.915 279.555 45.085 279.725 ;
        RECT 45.375 279.555 45.545 279.725 ;
        RECT 45.835 279.555 46.005 279.725 ;
        RECT 46.295 279.555 46.465 279.725 ;
        RECT 46.755 279.555 46.925 279.725 ;
        RECT 47.215 279.555 47.385 279.725 ;
        RECT 47.675 279.555 47.845 279.725 ;
        RECT 48.135 279.555 48.305 279.725 ;
        RECT 48.595 279.555 48.765 279.725 ;
        RECT 49.055 279.555 49.225 279.725 ;
        RECT 49.515 279.555 49.685 279.725 ;
        RECT 49.975 279.555 50.145 279.725 ;
        RECT 50.435 279.555 50.605 279.725 ;
        RECT 50.895 279.555 51.065 279.725 ;
        RECT 51.355 279.555 51.525 279.725 ;
        RECT 51.815 279.555 51.985 279.725 ;
        RECT 52.275 279.555 52.445 279.725 ;
        RECT 52.735 279.555 52.905 279.725 ;
        RECT 53.195 279.555 53.365 279.725 ;
        RECT 53.655 279.555 53.825 279.725 ;
        RECT 42.615 276.835 42.785 277.005 ;
        RECT 43.075 276.835 43.245 277.005 ;
        RECT 43.535 276.835 43.705 277.005 ;
        RECT 43.995 276.835 44.165 277.005 ;
        RECT 44.455 276.835 44.625 277.005 ;
        RECT 44.915 276.835 45.085 277.005 ;
        RECT 45.375 276.835 45.545 277.005 ;
        RECT 45.835 276.835 46.005 277.005 ;
        RECT 46.295 276.835 46.465 277.005 ;
        RECT 46.755 276.835 46.925 277.005 ;
        RECT 47.215 276.835 47.385 277.005 ;
        RECT 47.675 276.835 47.845 277.005 ;
        RECT 48.135 276.835 48.305 277.005 ;
        RECT 48.595 276.835 48.765 277.005 ;
        RECT 49.055 276.835 49.225 277.005 ;
        RECT 49.515 276.835 49.685 277.005 ;
        RECT 49.975 276.835 50.145 277.005 ;
        RECT 50.435 276.835 50.605 277.005 ;
        RECT 50.895 276.835 51.065 277.005 ;
        RECT 51.355 276.835 51.525 277.005 ;
        RECT 51.815 276.835 51.985 277.005 ;
        RECT 52.275 276.835 52.445 277.005 ;
        RECT 52.735 276.835 52.905 277.005 ;
        RECT 53.195 276.835 53.365 277.005 ;
        RECT 53.655 276.835 53.825 277.005 ;
        RECT 42.615 274.115 42.785 274.285 ;
        RECT 43.075 274.115 43.245 274.285 ;
        RECT 43.535 274.115 43.705 274.285 ;
        RECT 43.995 274.115 44.165 274.285 ;
        RECT 44.455 274.115 44.625 274.285 ;
        RECT 44.915 274.115 45.085 274.285 ;
        RECT 45.375 274.115 45.545 274.285 ;
        RECT 45.835 274.115 46.005 274.285 ;
        RECT 46.295 274.115 46.465 274.285 ;
        RECT 46.755 274.115 46.925 274.285 ;
        RECT 47.215 274.115 47.385 274.285 ;
        RECT 47.675 274.115 47.845 274.285 ;
        RECT 48.135 274.115 48.305 274.285 ;
        RECT 48.595 274.115 48.765 274.285 ;
        RECT 49.055 274.115 49.225 274.285 ;
        RECT 49.515 274.115 49.685 274.285 ;
        RECT 49.975 274.115 50.145 274.285 ;
        RECT 50.435 274.115 50.605 274.285 ;
        RECT 50.895 274.115 51.065 274.285 ;
        RECT 51.355 274.115 51.525 274.285 ;
        RECT 51.815 274.115 51.985 274.285 ;
        RECT 52.275 274.115 52.445 274.285 ;
        RECT 52.735 274.115 52.905 274.285 ;
        RECT 53.195 274.115 53.365 274.285 ;
        RECT 53.655 274.115 53.825 274.285 ;
        RECT 42.615 271.395 42.785 271.565 ;
        RECT 43.075 271.395 43.245 271.565 ;
        RECT 43.535 271.395 43.705 271.565 ;
        RECT 43.995 271.395 44.165 271.565 ;
        RECT 44.455 271.395 44.625 271.565 ;
        RECT 44.915 271.395 45.085 271.565 ;
        RECT 45.375 271.395 45.545 271.565 ;
        RECT 45.835 271.395 46.005 271.565 ;
        RECT 46.295 271.395 46.465 271.565 ;
        RECT 46.755 271.395 46.925 271.565 ;
        RECT 47.215 271.395 47.385 271.565 ;
        RECT 47.675 271.395 47.845 271.565 ;
        RECT 48.135 271.395 48.305 271.565 ;
        RECT 48.595 271.395 48.765 271.565 ;
        RECT 49.055 271.395 49.225 271.565 ;
        RECT 49.515 271.395 49.685 271.565 ;
        RECT 49.975 271.395 50.145 271.565 ;
        RECT 50.435 271.395 50.605 271.565 ;
        RECT 50.895 271.395 51.065 271.565 ;
        RECT 51.355 271.395 51.525 271.565 ;
        RECT 51.815 271.395 51.985 271.565 ;
        RECT 52.275 271.395 52.445 271.565 ;
        RECT 52.735 271.395 52.905 271.565 ;
        RECT 53.195 271.395 53.365 271.565 ;
        RECT 53.655 271.395 53.825 271.565 ;
        RECT 42.615 268.675 42.785 268.845 ;
        RECT 43.075 268.675 43.245 268.845 ;
        RECT 43.535 268.675 43.705 268.845 ;
        RECT 43.995 268.675 44.165 268.845 ;
        RECT 44.455 268.675 44.625 268.845 ;
        RECT 44.915 268.675 45.085 268.845 ;
        RECT 45.375 268.675 45.545 268.845 ;
        RECT 45.835 268.675 46.005 268.845 ;
        RECT 46.295 268.675 46.465 268.845 ;
        RECT 46.755 268.675 46.925 268.845 ;
        RECT 47.215 268.675 47.385 268.845 ;
        RECT 47.675 268.675 47.845 268.845 ;
        RECT 48.135 268.675 48.305 268.845 ;
        RECT 48.595 268.675 48.765 268.845 ;
        RECT 49.055 268.675 49.225 268.845 ;
        RECT 49.515 268.675 49.685 268.845 ;
        RECT 49.975 268.675 50.145 268.845 ;
        RECT 50.435 268.675 50.605 268.845 ;
        RECT 50.895 268.675 51.065 268.845 ;
        RECT 51.355 268.675 51.525 268.845 ;
        RECT 51.815 268.675 51.985 268.845 ;
        RECT 52.275 268.675 52.445 268.845 ;
        RECT 52.735 268.675 52.905 268.845 ;
        RECT 53.195 268.675 53.365 268.845 ;
        RECT 53.655 268.675 53.825 268.845 ;
        RECT 42.615 265.955 42.785 266.125 ;
        RECT 43.075 265.955 43.245 266.125 ;
        RECT 43.535 265.955 43.705 266.125 ;
        RECT 43.995 265.955 44.165 266.125 ;
        RECT 44.455 265.955 44.625 266.125 ;
        RECT 44.915 265.955 45.085 266.125 ;
        RECT 45.375 265.955 45.545 266.125 ;
        RECT 45.835 265.955 46.005 266.125 ;
        RECT 46.295 265.955 46.465 266.125 ;
        RECT 46.755 265.955 46.925 266.125 ;
        RECT 47.215 265.955 47.385 266.125 ;
        RECT 47.675 265.955 47.845 266.125 ;
        RECT 48.135 265.955 48.305 266.125 ;
        RECT 48.595 265.955 48.765 266.125 ;
        RECT 49.055 265.955 49.225 266.125 ;
        RECT 49.515 265.955 49.685 266.125 ;
        RECT 49.975 265.955 50.145 266.125 ;
        RECT 50.435 265.955 50.605 266.125 ;
        RECT 50.895 265.955 51.065 266.125 ;
        RECT 51.355 265.955 51.525 266.125 ;
        RECT 51.815 265.955 51.985 266.125 ;
        RECT 52.275 265.955 52.445 266.125 ;
        RECT 52.735 265.955 52.905 266.125 ;
        RECT 53.195 265.955 53.365 266.125 ;
        RECT 53.655 265.955 53.825 266.125 ;
        RECT 42.615 263.235 42.785 263.405 ;
        RECT 43.075 263.235 43.245 263.405 ;
        RECT 43.535 263.235 43.705 263.405 ;
        RECT 43.995 263.235 44.165 263.405 ;
        RECT 44.455 263.235 44.625 263.405 ;
        RECT 44.915 263.235 45.085 263.405 ;
        RECT 45.375 263.235 45.545 263.405 ;
        RECT 45.835 263.235 46.005 263.405 ;
        RECT 46.295 263.235 46.465 263.405 ;
        RECT 46.755 263.235 46.925 263.405 ;
        RECT 47.215 263.235 47.385 263.405 ;
        RECT 47.675 263.235 47.845 263.405 ;
        RECT 48.135 263.235 48.305 263.405 ;
        RECT 48.595 263.235 48.765 263.405 ;
        RECT 49.055 263.235 49.225 263.405 ;
        RECT 49.515 263.235 49.685 263.405 ;
        RECT 49.975 263.235 50.145 263.405 ;
        RECT 50.435 263.235 50.605 263.405 ;
        RECT 50.895 263.235 51.065 263.405 ;
        RECT 51.355 263.235 51.525 263.405 ;
        RECT 51.815 263.235 51.985 263.405 ;
        RECT 52.275 263.235 52.445 263.405 ;
        RECT 52.735 263.235 52.905 263.405 ;
        RECT 53.195 263.235 53.365 263.405 ;
        RECT 53.655 263.235 53.825 263.405 ;
        RECT 42.615 260.515 42.785 260.685 ;
        RECT 43.075 260.515 43.245 260.685 ;
        RECT 43.535 260.515 43.705 260.685 ;
        RECT 43.995 260.515 44.165 260.685 ;
        RECT 44.455 260.515 44.625 260.685 ;
        RECT 44.915 260.515 45.085 260.685 ;
        RECT 45.375 260.515 45.545 260.685 ;
        RECT 45.835 260.515 46.005 260.685 ;
        RECT 46.295 260.515 46.465 260.685 ;
        RECT 46.755 260.515 46.925 260.685 ;
        RECT 47.215 260.515 47.385 260.685 ;
        RECT 47.675 260.515 47.845 260.685 ;
        RECT 48.135 260.515 48.305 260.685 ;
        RECT 48.595 260.515 48.765 260.685 ;
        RECT 49.055 260.515 49.225 260.685 ;
        RECT 49.515 260.515 49.685 260.685 ;
        RECT 49.975 260.515 50.145 260.685 ;
        RECT 50.435 260.515 50.605 260.685 ;
        RECT 50.895 260.515 51.065 260.685 ;
        RECT 51.355 260.515 51.525 260.685 ;
        RECT 51.815 260.515 51.985 260.685 ;
        RECT 52.275 260.515 52.445 260.685 ;
        RECT 52.735 260.515 52.905 260.685 ;
        RECT 53.195 260.515 53.365 260.685 ;
        RECT 53.655 260.515 53.825 260.685 ;
        RECT 42.615 257.795 42.785 257.965 ;
        RECT 43.075 257.795 43.245 257.965 ;
        RECT 43.535 257.795 43.705 257.965 ;
        RECT 43.995 257.795 44.165 257.965 ;
        RECT 44.455 257.795 44.625 257.965 ;
        RECT 44.915 257.795 45.085 257.965 ;
        RECT 45.375 257.795 45.545 257.965 ;
        RECT 45.835 257.795 46.005 257.965 ;
        RECT 46.295 257.795 46.465 257.965 ;
        RECT 46.755 257.795 46.925 257.965 ;
        RECT 47.215 257.795 47.385 257.965 ;
        RECT 47.675 257.795 47.845 257.965 ;
        RECT 48.135 257.795 48.305 257.965 ;
        RECT 48.595 257.795 48.765 257.965 ;
        RECT 49.055 257.795 49.225 257.965 ;
        RECT 49.515 257.795 49.685 257.965 ;
        RECT 49.975 257.795 50.145 257.965 ;
        RECT 50.435 257.795 50.605 257.965 ;
        RECT 50.895 257.795 51.065 257.965 ;
        RECT 51.355 257.795 51.525 257.965 ;
        RECT 51.815 257.795 51.985 257.965 ;
        RECT 52.275 257.795 52.445 257.965 ;
        RECT 52.735 257.795 52.905 257.965 ;
        RECT 53.195 257.795 53.365 257.965 ;
        RECT 53.655 257.795 53.825 257.965 ;
        RECT 42.615 255.075 42.785 255.245 ;
        RECT 43.075 255.075 43.245 255.245 ;
        RECT 43.535 255.075 43.705 255.245 ;
        RECT 43.995 255.075 44.165 255.245 ;
        RECT 44.455 255.075 44.625 255.245 ;
        RECT 44.915 255.075 45.085 255.245 ;
        RECT 45.375 255.075 45.545 255.245 ;
        RECT 45.835 255.075 46.005 255.245 ;
        RECT 46.295 255.075 46.465 255.245 ;
        RECT 46.755 255.075 46.925 255.245 ;
        RECT 47.215 255.075 47.385 255.245 ;
        RECT 47.675 255.075 47.845 255.245 ;
        RECT 48.135 255.075 48.305 255.245 ;
        RECT 48.595 255.075 48.765 255.245 ;
        RECT 49.055 255.075 49.225 255.245 ;
        RECT 49.515 255.075 49.685 255.245 ;
        RECT 49.975 255.075 50.145 255.245 ;
        RECT 50.435 255.075 50.605 255.245 ;
        RECT 50.895 255.075 51.065 255.245 ;
        RECT 51.355 255.075 51.525 255.245 ;
        RECT 51.815 255.075 51.985 255.245 ;
        RECT 52.275 255.075 52.445 255.245 ;
        RECT 52.735 255.075 52.905 255.245 ;
        RECT 53.195 255.075 53.365 255.245 ;
        RECT 53.655 255.075 53.825 255.245 ;
        RECT 42.615 252.355 42.785 252.525 ;
        RECT 43.075 252.355 43.245 252.525 ;
        RECT 43.535 252.355 43.705 252.525 ;
        RECT 43.995 252.355 44.165 252.525 ;
        RECT 44.455 252.355 44.625 252.525 ;
        RECT 44.915 252.355 45.085 252.525 ;
        RECT 45.375 252.355 45.545 252.525 ;
        RECT 45.835 252.355 46.005 252.525 ;
        RECT 46.295 252.355 46.465 252.525 ;
        RECT 46.755 252.355 46.925 252.525 ;
        RECT 47.215 252.355 47.385 252.525 ;
        RECT 47.675 252.355 47.845 252.525 ;
        RECT 48.135 252.355 48.305 252.525 ;
        RECT 48.595 252.355 48.765 252.525 ;
        RECT 49.055 252.355 49.225 252.525 ;
        RECT 49.515 252.355 49.685 252.525 ;
        RECT 49.975 252.355 50.145 252.525 ;
        RECT 50.435 252.355 50.605 252.525 ;
        RECT 50.895 252.355 51.065 252.525 ;
        RECT 51.355 252.355 51.525 252.525 ;
        RECT 51.815 252.355 51.985 252.525 ;
        RECT 52.275 252.355 52.445 252.525 ;
        RECT 52.735 252.355 52.905 252.525 ;
        RECT 53.195 252.355 53.365 252.525 ;
        RECT 53.655 252.355 53.825 252.525 ;
        RECT 42.615 249.635 42.785 249.805 ;
        RECT 43.075 249.635 43.245 249.805 ;
        RECT 43.535 249.635 43.705 249.805 ;
        RECT 43.995 249.635 44.165 249.805 ;
        RECT 44.455 249.635 44.625 249.805 ;
        RECT 44.915 249.635 45.085 249.805 ;
        RECT 45.375 249.635 45.545 249.805 ;
        RECT 45.835 249.635 46.005 249.805 ;
        RECT 46.295 249.635 46.465 249.805 ;
        RECT 46.755 249.635 46.925 249.805 ;
        RECT 47.215 249.635 47.385 249.805 ;
        RECT 47.675 249.635 47.845 249.805 ;
        RECT 48.135 249.635 48.305 249.805 ;
        RECT 48.595 249.635 48.765 249.805 ;
        RECT 49.055 249.635 49.225 249.805 ;
        RECT 49.515 249.635 49.685 249.805 ;
        RECT 49.975 249.635 50.145 249.805 ;
        RECT 50.435 249.635 50.605 249.805 ;
        RECT 50.895 249.635 51.065 249.805 ;
        RECT 51.355 249.635 51.525 249.805 ;
        RECT 51.815 249.635 51.985 249.805 ;
        RECT 52.275 249.635 52.445 249.805 ;
        RECT 52.735 249.635 52.905 249.805 ;
        RECT 53.195 249.635 53.365 249.805 ;
        RECT 53.655 249.635 53.825 249.805 ;
        RECT 42.615 246.915 42.785 247.085 ;
        RECT 43.075 246.915 43.245 247.085 ;
        RECT 43.535 246.915 43.705 247.085 ;
        RECT 43.995 246.915 44.165 247.085 ;
        RECT 44.455 246.915 44.625 247.085 ;
        RECT 44.915 246.915 45.085 247.085 ;
        RECT 45.375 246.915 45.545 247.085 ;
        RECT 45.835 246.915 46.005 247.085 ;
        RECT 46.295 246.915 46.465 247.085 ;
        RECT 46.755 246.915 46.925 247.085 ;
        RECT 47.215 246.915 47.385 247.085 ;
        RECT 47.675 246.915 47.845 247.085 ;
        RECT 48.135 246.915 48.305 247.085 ;
        RECT 48.595 246.915 48.765 247.085 ;
        RECT 49.055 246.915 49.225 247.085 ;
        RECT 49.515 246.915 49.685 247.085 ;
        RECT 49.975 246.915 50.145 247.085 ;
        RECT 50.435 246.915 50.605 247.085 ;
        RECT 50.895 246.915 51.065 247.085 ;
        RECT 51.355 246.915 51.525 247.085 ;
        RECT 51.815 246.915 51.985 247.085 ;
        RECT 52.275 246.915 52.445 247.085 ;
        RECT 52.735 246.915 52.905 247.085 ;
        RECT 53.195 246.915 53.365 247.085 ;
        RECT 53.655 246.915 53.825 247.085 ;
        RECT 42.615 244.195 42.785 244.365 ;
        RECT 43.075 244.195 43.245 244.365 ;
        RECT 43.535 244.195 43.705 244.365 ;
        RECT 43.995 244.195 44.165 244.365 ;
        RECT 44.455 244.195 44.625 244.365 ;
        RECT 44.915 244.195 45.085 244.365 ;
        RECT 45.375 244.195 45.545 244.365 ;
        RECT 45.835 244.195 46.005 244.365 ;
        RECT 46.295 244.195 46.465 244.365 ;
        RECT 46.755 244.195 46.925 244.365 ;
        RECT 47.215 244.195 47.385 244.365 ;
        RECT 47.675 244.195 47.845 244.365 ;
        RECT 48.135 244.195 48.305 244.365 ;
        RECT 48.595 244.195 48.765 244.365 ;
        RECT 49.055 244.195 49.225 244.365 ;
        RECT 49.515 244.195 49.685 244.365 ;
        RECT 49.975 244.195 50.145 244.365 ;
        RECT 50.435 244.195 50.605 244.365 ;
        RECT 50.895 244.195 51.065 244.365 ;
        RECT 51.355 244.195 51.525 244.365 ;
        RECT 51.815 244.195 51.985 244.365 ;
        RECT 52.275 244.195 52.445 244.365 ;
        RECT 52.735 244.195 52.905 244.365 ;
        RECT 53.195 244.195 53.365 244.365 ;
        RECT 53.655 244.195 53.825 244.365 ;
        RECT 42.615 241.475 42.785 241.645 ;
        RECT 43.075 241.475 43.245 241.645 ;
        RECT 43.535 241.475 43.705 241.645 ;
        RECT 43.995 241.475 44.165 241.645 ;
        RECT 44.455 241.475 44.625 241.645 ;
        RECT 44.915 241.475 45.085 241.645 ;
        RECT 45.375 241.475 45.545 241.645 ;
        RECT 45.835 241.475 46.005 241.645 ;
        RECT 46.295 241.475 46.465 241.645 ;
        RECT 46.755 241.475 46.925 241.645 ;
        RECT 47.215 241.475 47.385 241.645 ;
        RECT 47.675 241.475 47.845 241.645 ;
        RECT 48.135 241.475 48.305 241.645 ;
        RECT 48.595 241.475 48.765 241.645 ;
        RECT 49.055 241.475 49.225 241.645 ;
        RECT 49.515 241.475 49.685 241.645 ;
        RECT 49.975 241.475 50.145 241.645 ;
        RECT 50.435 241.475 50.605 241.645 ;
        RECT 50.895 241.475 51.065 241.645 ;
        RECT 51.355 241.475 51.525 241.645 ;
        RECT 51.815 241.475 51.985 241.645 ;
        RECT 52.275 241.475 52.445 241.645 ;
        RECT 52.735 241.475 52.905 241.645 ;
        RECT 53.195 241.475 53.365 241.645 ;
        RECT 53.655 241.475 53.825 241.645 ;
        RECT 42.615 238.755 42.785 238.925 ;
        RECT 43.075 238.755 43.245 238.925 ;
        RECT 43.535 238.755 43.705 238.925 ;
        RECT 43.995 238.755 44.165 238.925 ;
        RECT 44.455 238.755 44.625 238.925 ;
        RECT 44.915 238.755 45.085 238.925 ;
        RECT 45.375 238.755 45.545 238.925 ;
        RECT 45.835 238.755 46.005 238.925 ;
        RECT 46.295 238.755 46.465 238.925 ;
        RECT 46.755 238.755 46.925 238.925 ;
        RECT 47.215 238.755 47.385 238.925 ;
        RECT 47.675 238.755 47.845 238.925 ;
        RECT 48.135 238.755 48.305 238.925 ;
        RECT 48.595 238.755 48.765 238.925 ;
        RECT 49.055 238.755 49.225 238.925 ;
        RECT 49.515 238.755 49.685 238.925 ;
        RECT 49.975 238.755 50.145 238.925 ;
        RECT 50.435 238.755 50.605 238.925 ;
        RECT 50.895 238.755 51.065 238.925 ;
        RECT 51.355 238.755 51.525 238.925 ;
        RECT 51.815 238.755 51.985 238.925 ;
        RECT 52.275 238.755 52.445 238.925 ;
        RECT 52.735 238.755 52.905 238.925 ;
        RECT 53.195 238.755 53.365 238.925 ;
        RECT 53.655 238.755 53.825 238.925 ;
        RECT 42.615 236.035 42.785 236.205 ;
        RECT 43.075 236.035 43.245 236.205 ;
        RECT 43.535 236.035 43.705 236.205 ;
        RECT 43.995 236.035 44.165 236.205 ;
        RECT 44.455 236.035 44.625 236.205 ;
        RECT 44.915 236.035 45.085 236.205 ;
        RECT 45.375 236.035 45.545 236.205 ;
        RECT 45.835 236.035 46.005 236.205 ;
        RECT 46.295 236.035 46.465 236.205 ;
        RECT 46.755 236.035 46.925 236.205 ;
        RECT 47.215 236.035 47.385 236.205 ;
        RECT 47.675 236.035 47.845 236.205 ;
        RECT 48.135 236.035 48.305 236.205 ;
        RECT 48.595 236.035 48.765 236.205 ;
        RECT 49.055 236.035 49.225 236.205 ;
        RECT 49.515 236.035 49.685 236.205 ;
        RECT 49.975 236.035 50.145 236.205 ;
        RECT 50.435 236.035 50.605 236.205 ;
        RECT 50.895 236.035 51.065 236.205 ;
        RECT 51.355 236.035 51.525 236.205 ;
        RECT 51.815 236.035 51.985 236.205 ;
        RECT 52.275 236.035 52.445 236.205 ;
        RECT 52.735 236.035 52.905 236.205 ;
        RECT 53.195 236.035 53.365 236.205 ;
        RECT 53.655 236.035 53.825 236.205 ;
        RECT 42.615 233.315 42.785 233.485 ;
        RECT 43.075 233.315 43.245 233.485 ;
        RECT 43.535 233.315 43.705 233.485 ;
        RECT 43.995 233.315 44.165 233.485 ;
        RECT 44.455 233.315 44.625 233.485 ;
        RECT 44.915 233.315 45.085 233.485 ;
        RECT 45.375 233.315 45.545 233.485 ;
        RECT 45.835 233.315 46.005 233.485 ;
        RECT 46.295 233.315 46.465 233.485 ;
        RECT 46.755 233.315 46.925 233.485 ;
        RECT 47.215 233.315 47.385 233.485 ;
        RECT 47.675 233.315 47.845 233.485 ;
        RECT 48.135 233.315 48.305 233.485 ;
        RECT 48.595 233.315 48.765 233.485 ;
        RECT 49.055 233.315 49.225 233.485 ;
        RECT 49.515 233.315 49.685 233.485 ;
        RECT 49.975 233.315 50.145 233.485 ;
        RECT 50.435 233.315 50.605 233.485 ;
        RECT 50.895 233.315 51.065 233.485 ;
        RECT 51.355 233.315 51.525 233.485 ;
        RECT 51.815 233.315 51.985 233.485 ;
        RECT 52.275 233.315 52.445 233.485 ;
        RECT 52.735 233.315 52.905 233.485 ;
        RECT 53.195 233.315 53.365 233.485 ;
        RECT 53.655 233.315 53.825 233.485 ;
        RECT 42.615 230.595 42.785 230.765 ;
        RECT 43.075 230.595 43.245 230.765 ;
        RECT 43.535 230.595 43.705 230.765 ;
        RECT 43.995 230.595 44.165 230.765 ;
        RECT 44.455 230.595 44.625 230.765 ;
        RECT 44.915 230.595 45.085 230.765 ;
        RECT 45.375 230.595 45.545 230.765 ;
        RECT 45.835 230.595 46.005 230.765 ;
        RECT 46.295 230.595 46.465 230.765 ;
        RECT 46.755 230.595 46.925 230.765 ;
        RECT 47.215 230.595 47.385 230.765 ;
        RECT 47.675 230.595 47.845 230.765 ;
        RECT 48.135 230.595 48.305 230.765 ;
        RECT 48.595 230.595 48.765 230.765 ;
        RECT 49.055 230.595 49.225 230.765 ;
        RECT 49.515 230.595 49.685 230.765 ;
        RECT 49.975 230.595 50.145 230.765 ;
        RECT 50.435 230.595 50.605 230.765 ;
        RECT 50.895 230.595 51.065 230.765 ;
        RECT 51.355 230.595 51.525 230.765 ;
        RECT 51.815 230.595 51.985 230.765 ;
        RECT 52.275 230.595 52.445 230.765 ;
        RECT 52.735 230.595 52.905 230.765 ;
        RECT 53.195 230.595 53.365 230.765 ;
        RECT 53.655 230.595 53.825 230.765 ;
        RECT 42.615 227.875 42.785 228.045 ;
        RECT 43.075 227.875 43.245 228.045 ;
        RECT 43.535 227.875 43.705 228.045 ;
        RECT 43.995 227.875 44.165 228.045 ;
        RECT 44.455 227.875 44.625 228.045 ;
        RECT 44.915 227.875 45.085 228.045 ;
        RECT 45.375 227.875 45.545 228.045 ;
        RECT 45.835 227.875 46.005 228.045 ;
        RECT 46.295 227.875 46.465 228.045 ;
        RECT 46.755 227.875 46.925 228.045 ;
        RECT 47.215 227.875 47.385 228.045 ;
        RECT 47.675 227.875 47.845 228.045 ;
        RECT 48.135 227.875 48.305 228.045 ;
        RECT 48.595 227.875 48.765 228.045 ;
        RECT 49.055 227.875 49.225 228.045 ;
        RECT 49.515 227.875 49.685 228.045 ;
        RECT 49.975 227.875 50.145 228.045 ;
        RECT 50.435 227.875 50.605 228.045 ;
        RECT 50.895 227.875 51.065 228.045 ;
        RECT 51.355 227.875 51.525 228.045 ;
        RECT 51.815 227.875 51.985 228.045 ;
        RECT 52.275 227.875 52.445 228.045 ;
        RECT 52.735 227.875 52.905 228.045 ;
        RECT 53.195 227.875 53.365 228.045 ;
        RECT 53.655 227.875 53.825 228.045 ;
        RECT 42.615 225.155 42.785 225.325 ;
        RECT 43.075 225.155 43.245 225.325 ;
        RECT 43.535 225.155 43.705 225.325 ;
        RECT 43.995 225.155 44.165 225.325 ;
        RECT 44.455 225.155 44.625 225.325 ;
        RECT 44.915 225.155 45.085 225.325 ;
        RECT 45.375 225.155 45.545 225.325 ;
        RECT 45.835 225.155 46.005 225.325 ;
        RECT 46.295 225.155 46.465 225.325 ;
        RECT 46.755 225.155 46.925 225.325 ;
        RECT 47.215 225.155 47.385 225.325 ;
        RECT 47.675 225.155 47.845 225.325 ;
        RECT 48.135 225.155 48.305 225.325 ;
        RECT 48.595 225.155 48.765 225.325 ;
        RECT 49.055 225.155 49.225 225.325 ;
        RECT 49.515 225.155 49.685 225.325 ;
        RECT 49.975 225.155 50.145 225.325 ;
        RECT 50.435 225.155 50.605 225.325 ;
        RECT 50.895 225.155 51.065 225.325 ;
        RECT 51.355 225.155 51.525 225.325 ;
        RECT 51.815 225.155 51.985 225.325 ;
        RECT 52.275 225.155 52.445 225.325 ;
        RECT 52.735 225.155 52.905 225.325 ;
        RECT 53.195 225.155 53.365 225.325 ;
        RECT 53.655 225.155 53.825 225.325 ;
        RECT 42.615 222.435 42.785 222.605 ;
        RECT 43.075 222.435 43.245 222.605 ;
        RECT 43.535 222.435 43.705 222.605 ;
        RECT 43.995 222.435 44.165 222.605 ;
        RECT 44.455 222.435 44.625 222.605 ;
        RECT 44.915 222.435 45.085 222.605 ;
        RECT 45.375 222.435 45.545 222.605 ;
        RECT 45.835 222.435 46.005 222.605 ;
        RECT 46.295 222.435 46.465 222.605 ;
        RECT 46.755 222.435 46.925 222.605 ;
        RECT 47.215 222.435 47.385 222.605 ;
        RECT 47.675 222.435 47.845 222.605 ;
        RECT 48.135 222.435 48.305 222.605 ;
        RECT 48.595 222.435 48.765 222.605 ;
        RECT 49.055 222.435 49.225 222.605 ;
        RECT 49.515 222.435 49.685 222.605 ;
        RECT 49.975 222.435 50.145 222.605 ;
        RECT 50.435 222.435 50.605 222.605 ;
        RECT 50.895 222.435 51.065 222.605 ;
        RECT 51.355 222.435 51.525 222.605 ;
        RECT 51.815 222.435 51.985 222.605 ;
        RECT 52.275 222.435 52.445 222.605 ;
        RECT 52.735 222.435 52.905 222.605 ;
        RECT 53.195 222.435 53.365 222.605 ;
        RECT 53.655 222.435 53.825 222.605 ;
        RECT 42.615 219.715 42.785 219.885 ;
        RECT 43.075 219.715 43.245 219.885 ;
        RECT 43.535 219.715 43.705 219.885 ;
        RECT 43.995 219.715 44.165 219.885 ;
        RECT 44.455 219.715 44.625 219.885 ;
        RECT 44.915 219.715 45.085 219.885 ;
        RECT 45.375 219.715 45.545 219.885 ;
        RECT 45.835 219.715 46.005 219.885 ;
        RECT 46.295 219.715 46.465 219.885 ;
        RECT 46.755 219.715 46.925 219.885 ;
        RECT 47.215 219.715 47.385 219.885 ;
        RECT 47.675 219.715 47.845 219.885 ;
        RECT 48.135 219.715 48.305 219.885 ;
        RECT 48.595 219.715 48.765 219.885 ;
        RECT 49.055 219.715 49.225 219.885 ;
        RECT 49.515 219.715 49.685 219.885 ;
        RECT 49.975 219.715 50.145 219.885 ;
        RECT 50.435 219.715 50.605 219.885 ;
        RECT 50.895 219.715 51.065 219.885 ;
        RECT 51.355 219.715 51.525 219.885 ;
        RECT 51.815 219.715 51.985 219.885 ;
        RECT 52.275 219.715 52.445 219.885 ;
        RECT 52.735 219.715 52.905 219.885 ;
        RECT 53.195 219.715 53.365 219.885 ;
        RECT 53.655 219.715 53.825 219.885 ;
        RECT 42.615 216.995 42.785 217.165 ;
        RECT 43.075 216.995 43.245 217.165 ;
        RECT 43.535 216.995 43.705 217.165 ;
        RECT 43.995 216.995 44.165 217.165 ;
        RECT 44.455 216.995 44.625 217.165 ;
        RECT 44.915 216.995 45.085 217.165 ;
        RECT 45.375 216.995 45.545 217.165 ;
        RECT 45.835 216.995 46.005 217.165 ;
        RECT 46.295 216.995 46.465 217.165 ;
        RECT 46.755 216.995 46.925 217.165 ;
        RECT 47.215 216.995 47.385 217.165 ;
        RECT 47.675 216.995 47.845 217.165 ;
        RECT 48.135 216.995 48.305 217.165 ;
        RECT 48.595 216.995 48.765 217.165 ;
        RECT 49.055 216.995 49.225 217.165 ;
        RECT 49.515 216.995 49.685 217.165 ;
        RECT 49.975 216.995 50.145 217.165 ;
        RECT 50.435 216.995 50.605 217.165 ;
        RECT 50.895 216.995 51.065 217.165 ;
        RECT 51.355 216.995 51.525 217.165 ;
        RECT 51.815 216.995 51.985 217.165 ;
        RECT 52.275 216.995 52.445 217.165 ;
        RECT 52.735 216.995 52.905 217.165 ;
        RECT 53.195 216.995 53.365 217.165 ;
        RECT 53.655 216.995 53.825 217.165 ;
        RECT 42.615 214.275 42.785 214.445 ;
        RECT 43.075 214.275 43.245 214.445 ;
        RECT 43.535 214.275 43.705 214.445 ;
        RECT 43.995 214.275 44.165 214.445 ;
        RECT 44.455 214.275 44.625 214.445 ;
        RECT 44.915 214.275 45.085 214.445 ;
        RECT 45.375 214.275 45.545 214.445 ;
        RECT 45.835 214.275 46.005 214.445 ;
        RECT 46.295 214.275 46.465 214.445 ;
        RECT 46.755 214.275 46.925 214.445 ;
        RECT 47.215 214.275 47.385 214.445 ;
        RECT 47.675 214.275 47.845 214.445 ;
        RECT 48.135 214.275 48.305 214.445 ;
        RECT 48.595 214.275 48.765 214.445 ;
        RECT 49.055 214.275 49.225 214.445 ;
        RECT 49.515 214.275 49.685 214.445 ;
        RECT 49.975 214.275 50.145 214.445 ;
        RECT 50.435 214.275 50.605 214.445 ;
        RECT 50.895 214.275 51.065 214.445 ;
        RECT 51.355 214.275 51.525 214.445 ;
        RECT 51.815 214.275 51.985 214.445 ;
        RECT 52.275 214.275 52.445 214.445 ;
        RECT 52.735 214.275 52.905 214.445 ;
        RECT 53.195 214.275 53.365 214.445 ;
        RECT 53.655 214.275 53.825 214.445 ;
        RECT 42.615 211.555 42.785 211.725 ;
        RECT 43.075 211.555 43.245 211.725 ;
        RECT 43.535 211.555 43.705 211.725 ;
        RECT 43.995 211.555 44.165 211.725 ;
        RECT 44.455 211.555 44.625 211.725 ;
        RECT 44.915 211.555 45.085 211.725 ;
        RECT 45.375 211.555 45.545 211.725 ;
        RECT 45.835 211.555 46.005 211.725 ;
        RECT 46.295 211.555 46.465 211.725 ;
        RECT 46.755 211.555 46.925 211.725 ;
        RECT 47.215 211.555 47.385 211.725 ;
        RECT 47.675 211.555 47.845 211.725 ;
        RECT 48.135 211.555 48.305 211.725 ;
        RECT 48.595 211.555 48.765 211.725 ;
        RECT 49.055 211.555 49.225 211.725 ;
        RECT 49.515 211.555 49.685 211.725 ;
        RECT 49.975 211.555 50.145 211.725 ;
        RECT 50.435 211.555 50.605 211.725 ;
        RECT 50.895 211.555 51.065 211.725 ;
        RECT 51.355 211.555 51.525 211.725 ;
        RECT 51.815 211.555 51.985 211.725 ;
        RECT 52.275 211.555 52.445 211.725 ;
        RECT 52.735 211.555 52.905 211.725 ;
        RECT 53.195 211.555 53.365 211.725 ;
        RECT 53.655 211.555 53.825 211.725 ;
        RECT 42.615 208.835 42.785 209.005 ;
        RECT 43.075 208.835 43.245 209.005 ;
        RECT 43.535 208.835 43.705 209.005 ;
        RECT 43.995 208.835 44.165 209.005 ;
        RECT 44.455 208.835 44.625 209.005 ;
        RECT 44.915 208.835 45.085 209.005 ;
        RECT 45.375 208.835 45.545 209.005 ;
        RECT 45.835 208.835 46.005 209.005 ;
        RECT 46.295 208.835 46.465 209.005 ;
        RECT 46.755 208.835 46.925 209.005 ;
        RECT 47.215 208.835 47.385 209.005 ;
        RECT 47.675 208.835 47.845 209.005 ;
        RECT 48.135 208.835 48.305 209.005 ;
        RECT 48.595 208.835 48.765 209.005 ;
        RECT 49.055 208.835 49.225 209.005 ;
        RECT 49.515 208.835 49.685 209.005 ;
        RECT 49.975 208.835 50.145 209.005 ;
        RECT 50.435 208.835 50.605 209.005 ;
        RECT 50.895 208.835 51.065 209.005 ;
        RECT 51.355 208.835 51.525 209.005 ;
        RECT 51.815 208.835 51.985 209.005 ;
        RECT 52.275 208.835 52.445 209.005 ;
        RECT 52.735 208.835 52.905 209.005 ;
        RECT 53.195 208.835 53.365 209.005 ;
        RECT 53.655 208.835 53.825 209.005 ;
        RECT 42.615 206.115 42.785 206.285 ;
        RECT 43.075 206.115 43.245 206.285 ;
        RECT 43.535 206.115 43.705 206.285 ;
        RECT 43.995 206.115 44.165 206.285 ;
        RECT 44.455 206.115 44.625 206.285 ;
        RECT 44.915 206.115 45.085 206.285 ;
        RECT 45.375 206.115 45.545 206.285 ;
        RECT 45.835 206.115 46.005 206.285 ;
        RECT 46.295 206.115 46.465 206.285 ;
        RECT 46.755 206.115 46.925 206.285 ;
        RECT 47.215 206.115 47.385 206.285 ;
        RECT 47.675 206.115 47.845 206.285 ;
        RECT 48.135 206.115 48.305 206.285 ;
        RECT 48.595 206.115 48.765 206.285 ;
        RECT 49.055 206.115 49.225 206.285 ;
        RECT 49.515 206.115 49.685 206.285 ;
        RECT 49.975 206.115 50.145 206.285 ;
        RECT 50.435 206.115 50.605 206.285 ;
        RECT 50.895 206.115 51.065 206.285 ;
        RECT 51.355 206.115 51.525 206.285 ;
        RECT 51.815 206.115 51.985 206.285 ;
        RECT 52.275 206.115 52.445 206.285 ;
        RECT 52.735 206.115 52.905 206.285 ;
        RECT 53.195 206.115 53.365 206.285 ;
        RECT 53.655 206.115 53.825 206.285 ;
        RECT 42.615 203.395 42.785 203.565 ;
        RECT 43.075 203.395 43.245 203.565 ;
        RECT 43.535 203.395 43.705 203.565 ;
        RECT 43.995 203.395 44.165 203.565 ;
        RECT 44.455 203.395 44.625 203.565 ;
        RECT 44.915 203.395 45.085 203.565 ;
        RECT 45.375 203.395 45.545 203.565 ;
        RECT 45.835 203.395 46.005 203.565 ;
        RECT 46.295 203.395 46.465 203.565 ;
        RECT 46.755 203.395 46.925 203.565 ;
        RECT 47.215 203.395 47.385 203.565 ;
        RECT 47.675 203.395 47.845 203.565 ;
        RECT 48.135 203.395 48.305 203.565 ;
        RECT 48.595 203.395 48.765 203.565 ;
        RECT 49.055 203.395 49.225 203.565 ;
        RECT 49.515 203.395 49.685 203.565 ;
        RECT 49.975 203.395 50.145 203.565 ;
        RECT 50.435 203.395 50.605 203.565 ;
        RECT 50.895 203.395 51.065 203.565 ;
        RECT 51.355 203.395 51.525 203.565 ;
        RECT 51.815 203.395 51.985 203.565 ;
        RECT 52.275 203.395 52.445 203.565 ;
        RECT 52.735 203.395 52.905 203.565 ;
        RECT 53.195 203.395 53.365 203.565 ;
        RECT 53.655 203.395 53.825 203.565 ;
        RECT 42.615 200.675 42.785 200.845 ;
        RECT 43.075 200.675 43.245 200.845 ;
        RECT 43.535 200.675 43.705 200.845 ;
        RECT 43.995 200.675 44.165 200.845 ;
        RECT 44.455 200.675 44.625 200.845 ;
        RECT 44.915 200.675 45.085 200.845 ;
        RECT 45.375 200.675 45.545 200.845 ;
        RECT 45.835 200.675 46.005 200.845 ;
        RECT 46.295 200.675 46.465 200.845 ;
        RECT 46.755 200.675 46.925 200.845 ;
        RECT 47.215 200.675 47.385 200.845 ;
        RECT 47.675 200.675 47.845 200.845 ;
        RECT 48.135 200.675 48.305 200.845 ;
        RECT 48.595 200.675 48.765 200.845 ;
        RECT 49.055 200.675 49.225 200.845 ;
        RECT 49.515 200.675 49.685 200.845 ;
        RECT 49.975 200.675 50.145 200.845 ;
        RECT 50.435 200.675 50.605 200.845 ;
        RECT 50.895 200.675 51.065 200.845 ;
        RECT 51.355 200.675 51.525 200.845 ;
        RECT 51.815 200.675 51.985 200.845 ;
        RECT 52.275 200.675 52.445 200.845 ;
        RECT 52.735 200.675 52.905 200.845 ;
        RECT 53.195 200.675 53.365 200.845 ;
        RECT 53.655 200.675 53.825 200.845 ;
        RECT 42.615 197.955 42.785 198.125 ;
        RECT 43.075 197.955 43.245 198.125 ;
        RECT 43.535 197.955 43.705 198.125 ;
        RECT 43.995 197.955 44.165 198.125 ;
        RECT 44.455 197.955 44.625 198.125 ;
        RECT 44.915 197.955 45.085 198.125 ;
        RECT 45.375 197.955 45.545 198.125 ;
        RECT 45.835 197.955 46.005 198.125 ;
        RECT 46.295 197.955 46.465 198.125 ;
        RECT 46.755 197.955 46.925 198.125 ;
        RECT 47.215 197.955 47.385 198.125 ;
        RECT 47.675 197.955 47.845 198.125 ;
        RECT 48.135 197.955 48.305 198.125 ;
        RECT 48.595 197.955 48.765 198.125 ;
        RECT 49.055 197.955 49.225 198.125 ;
        RECT 49.515 197.955 49.685 198.125 ;
        RECT 49.975 197.955 50.145 198.125 ;
        RECT 50.435 197.955 50.605 198.125 ;
        RECT 50.895 197.955 51.065 198.125 ;
        RECT 51.355 197.955 51.525 198.125 ;
        RECT 51.815 197.955 51.985 198.125 ;
        RECT 52.275 197.955 52.445 198.125 ;
        RECT 52.735 197.955 52.905 198.125 ;
        RECT 53.195 197.955 53.365 198.125 ;
        RECT 53.655 197.955 53.825 198.125 ;
        RECT 42.615 195.235 42.785 195.405 ;
        RECT 43.075 195.235 43.245 195.405 ;
        RECT 43.535 195.235 43.705 195.405 ;
        RECT 43.995 195.235 44.165 195.405 ;
        RECT 44.455 195.235 44.625 195.405 ;
        RECT 44.915 195.235 45.085 195.405 ;
        RECT 45.375 195.235 45.545 195.405 ;
        RECT 45.835 195.235 46.005 195.405 ;
        RECT 46.295 195.235 46.465 195.405 ;
        RECT 46.755 195.235 46.925 195.405 ;
        RECT 47.215 195.235 47.385 195.405 ;
        RECT 47.675 195.235 47.845 195.405 ;
        RECT 48.135 195.235 48.305 195.405 ;
        RECT 48.595 195.235 48.765 195.405 ;
        RECT 49.055 195.235 49.225 195.405 ;
        RECT 49.515 195.235 49.685 195.405 ;
        RECT 49.975 195.235 50.145 195.405 ;
        RECT 50.435 195.235 50.605 195.405 ;
        RECT 50.895 195.235 51.065 195.405 ;
        RECT 51.355 195.235 51.525 195.405 ;
        RECT 51.815 195.235 51.985 195.405 ;
        RECT 52.275 195.235 52.445 195.405 ;
        RECT 52.735 195.235 52.905 195.405 ;
        RECT 53.195 195.235 53.365 195.405 ;
        RECT 53.655 195.235 53.825 195.405 ;
        RECT 42.615 192.515 42.785 192.685 ;
        RECT 43.075 192.515 43.245 192.685 ;
        RECT 43.535 192.515 43.705 192.685 ;
        RECT 43.995 192.515 44.165 192.685 ;
        RECT 44.455 192.515 44.625 192.685 ;
        RECT 44.915 192.515 45.085 192.685 ;
        RECT 45.375 192.515 45.545 192.685 ;
        RECT 45.835 192.515 46.005 192.685 ;
        RECT 46.295 192.515 46.465 192.685 ;
        RECT 46.755 192.515 46.925 192.685 ;
        RECT 47.215 192.515 47.385 192.685 ;
        RECT 47.675 192.515 47.845 192.685 ;
        RECT 48.135 192.515 48.305 192.685 ;
        RECT 48.595 192.515 48.765 192.685 ;
        RECT 49.055 192.515 49.225 192.685 ;
        RECT 49.515 192.515 49.685 192.685 ;
        RECT 49.975 192.515 50.145 192.685 ;
        RECT 50.435 192.515 50.605 192.685 ;
        RECT 50.895 192.515 51.065 192.685 ;
        RECT 51.355 192.515 51.525 192.685 ;
        RECT 51.815 192.515 51.985 192.685 ;
        RECT 52.275 192.515 52.445 192.685 ;
        RECT 52.735 192.515 52.905 192.685 ;
        RECT 53.195 192.515 53.365 192.685 ;
        RECT 53.655 192.515 53.825 192.685 ;
        RECT 42.615 189.795 42.785 189.965 ;
        RECT 43.075 189.795 43.245 189.965 ;
        RECT 43.535 189.795 43.705 189.965 ;
        RECT 43.995 189.795 44.165 189.965 ;
        RECT 44.455 189.795 44.625 189.965 ;
        RECT 44.915 189.795 45.085 189.965 ;
        RECT 45.375 189.795 45.545 189.965 ;
        RECT 45.835 189.795 46.005 189.965 ;
        RECT 46.295 189.795 46.465 189.965 ;
        RECT 46.755 189.795 46.925 189.965 ;
        RECT 47.215 189.795 47.385 189.965 ;
        RECT 47.675 189.795 47.845 189.965 ;
        RECT 48.135 189.795 48.305 189.965 ;
        RECT 48.595 189.795 48.765 189.965 ;
        RECT 49.055 189.795 49.225 189.965 ;
        RECT 49.515 189.795 49.685 189.965 ;
        RECT 49.975 189.795 50.145 189.965 ;
        RECT 50.435 189.795 50.605 189.965 ;
        RECT 50.895 189.795 51.065 189.965 ;
        RECT 51.355 189.795 51.525 189.965 ;
        RECT 51.815 189.795 51.985 189.965 ;
        RECT 52.275 189.795 52.445 189.965 ;
        RECT 52.735 189.795 52.905 189.965 ;
        RECT 53.195 189.795 53.365 189.965 ;
        RECT 53.655 189.795 53.825 189.965 ;
        RECT 42.615 187.075 42.785 187.245 ;
        RECT 43.075 187.075 43.245 187.245 ;
        RECT 43.535 187.075 43.705 187.245 ;
        RECT 43.995 187.075 44.165 187.245 ;
        RECT 44.455 187.075 44.625 187.245 ;
        RECT 44.915 187.075 45.085 187.245 ;
        RECT 45.375 187.075 45.545 187.245 ;
        RECT 45.835 187.075 46.005 187.245 ;
        RECT 46.295 187.075 46.465 187.245 ;
        RECT 46.755 187.075 46.925 187.245 ;
        RECT 47.215 187.075 47.385 187.245 ;
        RECT 47.675 187.075 47.845 187.245 ;
        RECT 48.135 187.075 48.305 187.245 ;
        RECT 48.595 187.075 48.765 187.245 ;
        RECT 49.055 187.075 49.225 187.245 ;
        RECT 49.515 187.075 49.685 187.245 ;
        RECT 49.975 187.075 50.145 187.245 ;
        RECT 50.435 187.075 50.605 187.245 ;
        RECT 50.895 187.075 51.065 187.245 ;
        RECT 51.355 187.075 51.525 187.245 ;
        RECT 51.815 187.075 51.985 187.245 ;
        RECT 52.275 187.075 52.445 187.245 ;
        RECT 52.735 187.075 52.905 187.245 ;
        RECT 53.195 187.075 53.365 187.245 ;
        RECT 53.655 187.075 53.825 187.245 ;
        RECT 42.615 184.355 42.785 184.525 ;
        RECT 43.075 184.355 43.245 184.525 ;
        RECT 43.535 184.355 43.705 184.525 ;
        RECT 43.995 184.355 44.165 184.525 ;
        RECT 44.455 184.355 44.625 184.525 ;
        RECT 44.915 184.355 45.085 184.525 ;
        RECT 45.375 184.355 45.545 184.525 ;
        RECT 45.835 184.355 46.005 184.525 ;
        RECT 46.295 184.355 46.465 184.525 ;
        RECT 46.755 184.355 46.925 184.525 ;
        RECT 47.215 184.355 47.385 184.525 ;
        RECT 47.675 184.355 47.845 184.525 ;
        RECT 48.135 184.355 48.305 184.525 ;
        RECT 48.595 184.355 48.765 184.525 ;
        RECT 49.055 184.355 49.225 184.525 ;
        RECT 49.515 184.355 49.685 184.525 ;
        RECT 49.975 184.355 50.145 184.525 ;
        RECT 50.435 184.355 50.605 184.525 ;
        RECT 50.895 184.355 51.065 184.525 ;
        RECT 51.355 184.355 51.525 184.525 ;
        RECT 51.815 184.355 51.985 184.525 ;
        RECT 52.275 184.355 52.445 184.525 ;
        RECT 52.735 184.355 52.905 184.525 ;
        RECT 53.195 184.355 53.365 184.525 ;
        RECT 53.655 184.355 53.825 184.525 ;
        RECT 42.615 181.635 42.785 181.805 ;
        RECT 43.075 181.635 43.245 181.805 ;
        RECT 43.535 181.635 43.705 181.805 ;
        RECT 43.995 181.635 44.165 181.805 ;
        RECT 44.455 181.635 44.625 181.805 ;
        RECT 44.915 181.635 45.085 181.805 ;
        RECT 45.375 181.635 45.545 181.805 ;
        RECT 45.835 181.635 46.005 181.805 ;
        RECT 46.295 181.635 46.465 181.805 ;
        RECT 46.755 181.635 46.925 181.805 ;
        RECT 47.215 181.635 47.385 181.805 ;
        RECT 47.675 181.635 47.845 181.805 ;
        RECT 48.135 181.635 48.305 181.805 ;
        RECT 48.595 181.635 48.765 181.805 ;
        RECT 49.055 181.635 49.225 181.805 ;
        RECT 49.515 181.635 49.685 181.805 ;
        RECT 49.975 181.635 50.145 181.805 ;
        RECT 50.435 181.635 50.605 181.805 ;
        RECT 50.895 181.635 51.065 181.805 ;
        RECT 51.355 181.635 51.525 181.805 ;
        RECT 51.815 181.635 51.985 181.805 ;
        RECT 52.275 181.635 52.445 181.805 ;
        RECT 52.735 181.635 52.905 181.805 ;
        RECT 53.195 181.635 53.365 181.805 ;
        RECT 53.655 181.635 53.825 181.805 ;
        RECT 42.615 178.915 42.785 179.085 ;
        RECT 43.075 178.915 43.245 179.085 ;
        RECT 43.535 178.915 43.705 179.085 ;
        RECT 43.995 178.915 44.165 179.085 ;
        RECT 44.455 178.915 44.625 179.085 ;
        RECT 44.915 178.915 45.085 179.085 ;
        RECT 45.375 178.915 45.545 179.085 ;
        RECT 45.835 178.915 46.005 179.085 ;
        RECT 46.295 178.915 46.465 179.085 ;
        RECT 46.755 178.915 46.925 179.085 ;
        RECT 47.215 178.915 47.385 179.085 ;
        RECT 47.675 178.915 47.845 179.085 ;
        RECT 48.135 178.915 48.305 179.085 ;
        RECT 48.595 178.915 48.765 179.085 ;
        RECT 49.055 178.915 49.225 179.085 ;
        RECT 49.515 178.915 49.685 179.085 ;
        RECT 49.975 178.915 50.145 179.085 ;
        RECT 50.435 178.915 50.605 179.085 ;
        RECT 50.895 178.915 51.065 179.085 ;
        RECT 51.355 178.915 51.525 179.085 ;
        RECT 51.815 178.915 51.985 179.085 ;
        RECT 52.275 178.915 52.445 179.085 ;
        RECT 52.735 178.915 52.905 179.085 ;
        RECT 53.195 178.915 53.365 179.085 ;
        RECT 53.655 178.915 53.825 179.085 ;
        RECT 42.615 176.195 42.785 176.365 ;
        RECT 43.075 176.195 43.245 176.365 ;
        RECT 43.535 176.195 43.705 176.365 ;
        RECT 43.995 176.195 44.165 176.365 ;
        RECT 44.455 176.195 44.625 176.365 ;
        RECT 44.915 176.195 45.085 176.365 ;
        RECT 45.375 176.195 45.545 176.365 ;
        RECT 45.835 176.195 46.005 176.365 ;
        RECT 46.295 176.195 46.465 176.365 ;
        RECT 46.755 176.195 46.925 176.365 ;
        RECT 47.215 176.195 47.385 176.365 ;
        RECT 47.675 176.195 47.845 176.365 ;
        RECT 48.135 176.195 48.305 176.365 ;
        RECT 48.595 176.195 48.765 176.365 ;
        RECT 49.055 176.195 49.225 176.365 ;
        RECT 49.515 176.195 49.685 176.365 ;
        RECT 49.975 176.195 50.145 176.365 ;
        RECT 50.435 176.195 50.605 176.365 ;
        RECT 50.895 176.195 51.065 176.365 ;
        RECT 51.355 176.195 51.525 176.365 ;
        RECT 51.815 176.195 51.985 176.365 ;
        RECT 52.275 176.195 52.445 176.365 ;
        RECT 52.735 176.195 52.905 176.365 ;
        RECT 53.195 176.195 53.365 176.365 ;
        RECT 53.655 176.195 53.825 176.365 ;
        RECT 42.615 173.475 42.785 173.645 ;
        RECT 43.075 173.475 43.245 173.645 ;
        RECT 43.535 173.475 43.705 173.645 ;
        RECT 43.995 173.475 44.165 173.645 ;
        RECT 44.455 173.475 44.625 173.645 ;
        RECT 44.915 173.475 45.085 173.645 ;
        RECT 45.375 173.475 45.545 173.645 ;
        RECT 45.835 173.475 46.005 173.645 ;
        RECT 46.295 173.475 46.465 173.645 ;
        RECT 46.755 173.475 46.925 173.645 ;
        RECT 47.215 173.475 47.385 173.645 ;
        RECT 47.675 173.475 47.845 173.645 ;
        RECT 48.135 173.475 48.305 173.645 ;
        RECT 48.595 173.475 48.765 173.645 ;
        RECT 49.055 173.475 49.225 173.645 ;
        RECT 49.515 173.475 49.685 173.645 ;
        RECT 49.975 173.475 50.145 173.645 ;
        RECT 50.435 173.475 50.605 173.645 ;
        RECT 50.895 173.475 51.065 173.645 ;
        RECT 51.355 173.475 51.525 173.645 ;
        RECT 51.815 173.475 51.985 173.645 ;
        RECT 52.275 173.475 52.445 173.645 ;
        RECT 52.735 173.475 52.905 173.645 ;
        RECT 53.195 173.475 53.365 173.645 ;
        RECT 53.655 173.475 53.825 173.645 ;
        RECT 42.615 170.755 42.785 170.925 ;
        RECT 43.075 170.755 43.245 170.925 ;
        RECT 43.535 170.755 43.705 170.925 ;
        RECT 43.995 170.755 44.165 170.925 ;
        RECT 44.455 170.755 44.625 170.925 ;
        RECT 44.915 170.755 45.085 170.925 ;
        RECT 45.375 170.755 45.545 170.925 ;
        RECT 45.835 170.755 46.005 170.925 ;
        RECT 46.295 170.755 46.465 170.925 ;
        RECT 46.755 170.755 46.925 170.925 ;
        RECT 47.215 170.755 47.385 170.925 ;
        RECT 47.675 170.755 47.845 170.925 ;
        RECT 48.135 170.755 48.305 170.925 ;
        RECT 48.595 170.755 48.765 170.925 ;
        RECT 49.055 170.755 49.225 170.925 ;
        RECT 49.515 170.755 49.685 170.925 ;
        RECT 49.975 170.755 50.145 170.925 ;
        RECT 50.435 170.755 50.605 170.925 ;
        RECT 50.895 170.755 51.065 170.925 ;
        RECT 51.355 170.755 51.525 170.925 ;
        RECT 51.815 170.755 51.985 170.925 ;
        RECT 52.275 170.755 52.445 170.925 ;
        RECT 52.735 170.755 52.905 170.925 ;
        RECT 53.195 170.755 53.365 170.925 ;
        RECT 53.655 170.755 53.825 170.925 ;
        RECT 42.615 168.035 42.785 168.205 ;
        RECT 43.075 168.035 43.245 168.205 ;
        RECT 43.535 168.035 43.705 168.205 ;
        RECT 43.995 168.035 44.165 168.205 ;
        RECT 44.455 168.035 44.625 168.205 ;
        RECT 44.915 168.035 45.085 168.205 ;
        RECT 45.375 168.035 45.545 168.205 ;
        RECT 45.835 168.035 46.005 168.205 ;
        RECT 46.295 168.035 46.465 168.205 ;
        RECT 46.755 168.035 46.925 168.205 ;
        RECT 47.215 168.035 47.385 168.205 ;
        RECT 47.675 168.035 47.845 168.205 ;
        RECT 48.135 168.035 48.305 168.205 ;
        RECT 48.595 168.035 48.765 168.205 ;
        RECT 49.055 168.035 49.225 168.205 ;
        RECT 49.515 168.035 49.685 168.205 ;
        RECT 49.975 168.035 50.145 168.205 ;
        RECT 50.435 168.035 50.605 168.205 ;
        RECT 50.895 168.035 51.065 168.205 ;
        RECT 51.355 168.035 51.525 168.205 ;
        RECT 51.815 168.035 51.985 168.205 ;
        RECT 52.275 168.035 52.445 168.205 ;
        RECT 52.735 168.035 52.905 168.205 ;
        RECT 53.195 168.035 53.365 168.205 ;
        RECT 53.655 168.035 53.825 168.205 ;
        RECT 42.615 165.315 42.785 165.485 ;
        RECT 43.075 165.315 43.245 165.485 ;
        RECT 43.535 165.315 43.705 165.485 ;
        RECT 43.995 165.315 44.165 165.485 ;
        RECT 44.455 165.315 44.625 165.485 ;
        RECT 44.915 165.315 45.085 165.485 ;
        RECT 45.375 165.315 45.545 165.485 ;
        RECT 45.835 165.315 46.005 165.485 ;
        RECT 46.295 165.315 46.465 165.485 ;
        RECT 46.755 165.315 46.925 165.485 ;
        RECT 47.215 165.315 47.385 165.485 ;
        RECT 47.675 165.315 47.845 165.485 ;
        RECT 48.135 165.315 48.305 165.485 ;
        RECT 48.595 165.315 48.765 165.485 ;
        RECT 49.055 165.315 49.225 165.485 ;
        RECT 49.515 165.315 49.685 165.485 ;
        RECT 49.975 165.315 50.145 165.485 ;
        RECT 50.435 165.315 50.605 165.485 ;
        RECT 50.895 165.315 51.065 165.485 ;
        RECT 51.355 165.315 51.525 165.485 ;
        RECT 51.815 165.315 51.985 165.485 ;
        RECT 52.275 165.315 52.445 165.485 ;
        RECT 52.735 165.315 52.905 165.485 ;
        RECT 53.195 165.315 53.365 165.485 ;
        RECT 53.655 165.315 53.825 165.485 ;
        RECT 42.615 162.595 42.785 162.765 ;
        RECT 43.075 162.595 43.245 162.765 ;
        RECT 43.535 162.595 43.705 162.765 ;
        RECT 43.995 162.595 44.165 162.765 ;
        RECT 44.455 162.595 44.625 162.765 ;
        RECT 44.915 162.595 45.085 162.765 ;
        RECT 45.375 162.595 45.545 162.765 ;
        RECT 45.835 162.595 46.005 162.765 ;
        RECT 46.295 162.595 46.465 162.765 ;
        RECT 46.755 162.595 46.925 162.765 ;
        RECT 47.215 162.595 47.385 162.765 ;
        RECT 47.675 162.595 47.845 162.765 ;
        RECT 48.135 162.595 48.305 162.765 ;
        RECT 48.595 162.595 48.765 162.765 ;
        RECT 49.055 162.595 49.225 162.765 ;
        RECT 49.515 162.595 49.685 162.765 ;
        RECT 49.975 162.595 50.145 162.765 ;
        RECT 50.435 162.595 50.605 162.765 ;
        RECT 50.895 162.595 51.065 162.765 ;
        RECT 51.355 162.595 51.525 162.765 ;
        RECT 51.815 162.595 51.985 162.765 ;
        RECT 52.275 162.595 52.445 162.765 ;
        RECT 52.735 162.595 52.905 162.765 ;
        RECT 53.195 162.595 53.365 162.765 ;
        RECT 53.655 162.595 53.825 162.765 ;
        RECT 42.615 159.875 42.785 160.045 ;
        RECT 43.075 159.875 43.245 160.045 ;
        RECT 43.535 159.875 43.705 160.045 ;
        RECT 43.995 159.875 44.165 160.045 ;
        RECT 44.455 159.875 44.625 160.045 ;
        RECT 44.915 159.875 45.085 160.045 ;
        RECT 45.375 159.875 45.545 160.045 ;
        RECT 45.835 159.875 46.005 160.045 ;
        RECT 46.295 159.875 46.465 160.045 ;
        RECT 46.755 159.875 46.925 160.045 ;
        RECT 47.215 159.875 47.385 160.045 ;
        RECT 47.675 159.875 47.845 160.045 ;
        RECT 48.135 159.875 48.305 160.045 ;
        RECT 48.595 159.875 48.765 160.045 ;
        RECT 49.055 159.875 49.225 160.045 ;
        RECT 49.515 159.875 49.685 160.045 ;
        RECT 49.975 159.875 50.145 160.045 ;
        RECT 50.435 159.875 50.605 160.045 ;
        RECT 50.895 159.875 51.065 160.045 ;
        RECT 51.355 159.875 51.525 160.045 ;
        RECT 51.815 159.875 51.985 160.045 ;
        RECT 52.275 159.875 52.445 160.045 ;
        RECT 52.735 159.875 52.905 160.045 ;
        RECT 53.195 159.875 53.365 160.045 ;
        RECT 53.655 159.875 53.825 160.045 ;
        RECT 42.615 157.155 42.785 157.325 ;
        RECT 43.075 157.155 43.245 157.325 ;
        RECT 43.535 157.155 43.705 157.325 ;
        RECT 43.995 157.155 44.165 157.325 ;
        RECT 44.455 157.155 44.625 157.325 ;
        RECT 44.915 157.155 45.085 157.325 ;
        RECT 45.375 157.155 45.545 157.325 ;
        RECT 45.835 157.155 46.005 157.325 ;
        RECT 46.295 157.155 46.465 157.325 ;
        RECT 46.755 157.155 46.925 157.325 ;
        RECT 47.215 157.155 47.385 157.325 ;
        RECT 47.675 157.155 47.845 157.325 ;
        RECT 48.135 157.155 48.305 157.325 ;
        RECT 48.595 157.155 48.765 157.325 ;
        RECT 49.055 157.155 49.225 157.325 ;
        RECT 49.515 157.155 49.685 157.325 ;
        RECT 49.975 157.155 50.145 157.325 ;
        RECT 50.435 157.155 50.605 157.325 ;
        RECT 50.895 157.155 51.065 157.325 ;
        RECT 51.355 157.155 51.525 157.325 ;
        RECT 51.815 157.155 51.985 157.325 ;
        RECT 52.275 157.155 52.445 157.325 ;
        RECT 52.735 157.155 52.905 157.325 ;
        RECT 53.195 157.155 53.365 157.325 ;
        RECT 53.655 157.155 53.825 157.325 ;
        RECT 42.615 154.435 42.785 154.605 ;
        RECT 43.075 154.435 43.245 154.605 ;
        RECT 43.535 154.435 43.705 154.605 ;
        RECT 43.995 154.435 44.165 154.605 ;
        RECT 44.455 154.435 44.625 154.605 ;
        RECT 44.915 154.435 45.085 154.605 ;
        RECT 45.375 154.435 45.545 154.605 ;
        RECT 45.835 154.435 46.005 154.605 ;
        RECT 46.295 154.435 46.465 154.605 ;
        RECT 46.755 154.435 46.925 154.605 ;
        RECT 47.215 154.435 47.385 154.605 ;
        RECT 47.675 154.435 47.845 154.605 ;
        RECT 48.135 154.435 48.305 154.605 ;
        RECT 48.595 154.435 48.765 154.605 ;
        RECT 49.055 154.435 49.225 154.605 ;
        RECT 49.515 154.435 49.685 154.605 ;
        RECT 49.975 154.435 50.145 154.605 ;
        RECT 50.435 154.435 50.605 154.605 ;
        RECT 50.895 154.435 51.065 154.605 ;
        RECT 51.355 154.435 51.525 154.605 ;
        RECT 51.815 154.435 51.985 154.605 ;
        RECT 52.275 154.435 52.445 154.605 ;
        RECT 52.735 154.435 52.905 154.605 ;
        RECT 53.195 154.435 53.365 154.605 ;
        RECT 53.655 154.435 53.825 154.605 ;
        RECT 42.615 151.715 42.785 151.885 ;
        RECT 43.075 151.715 43.245 151.885 ;
        RECT 43.535 151.715 43.705 151.885 ;
        RECT 43.995 151.715 44.165 151.885 ;
        RECT 44.455 151.715 44.625 151.885 ;
        RECT 44.915 151.715 45.085 151.885 ;
        RECT 45.375 151.715 45.545 151.885 ;
        RECT 45.835 151.715 46.005 151.885 ;
        RECT 46.295 151.715 46.465 151.885 ;
        RECT 46.755 151.715 46.925 151.885 ;
        RECT 47.215 151.715 47.385 151.885 ;
        RECT 47.675 151.715 47.845 151.885 ;
        RECT 48.135 151.715 48.305 151.885 ;
        RECT 48.595 151.715 48.765 151.885 ;
        RECT 49.055 151.715 49.225 151.885 ;
        RECT 49.515 151.715 49.685 151.885 ;
        RECT 49.975 151.715 50.145 151.885 ;
        RECT 50.435 151.715 50.605 151.885 ;
        RECT 50.895 151.715 51.065 151.885 ;
        RECT 51.355 151.715 51.525 151.885 ;
        RECT 51.815 151.715 51.985 151.885 ;
        RECT 52.275 151.715 52.445 151.885 ;
        RECT 52.735 151.715 52.905 151.885 ;
        RECT 53.195 151.715 53.365 151.885 ;
        RECT 53.655 151.715 53.825 151.885 ;
        RECT 42.615 148.995 42.785 149.165 ;
        RECT 43.075 148.995 43.245 149.165 ;
        RECT 43.535 148.995 43.705 149.165 ;
        RECT 43.995 148.995 44.165 149.165 ;
        RECT 44.455 148.995 44.625 149.165 ;
        RECT 44.915 148.995 45.085 149.165 ;
        RECT 45.375 148.995 45.545 149.165 ;
        RECT 45.835 148.995 46.005 149.165 ;
        RECT 46.295 148.995 46.465 149.165 ;
        RECT 46.755 148.995 46.925 149.165 ;
        RECT 47.215 148.995 47.385 149.165 ;
        RECT 47.675 148.995 47.845 149.165 ;
        RECT 48.135 148.995 48.305 149.165 ;
        RECT 48.595 148.995 48.765 149.165 ;
        RECT 49.055 148.995 49.225 149.165 ;
        RECT 49.515 148.995 49.685 149.165 ;
        RECT 49.975 148.995 50.145 149.165 ;
        RECT 50.435 148.995 50.605 149.165 ;
        RECT 50.895 148.995 51.065 149.165 ;
        RECT 51.355 148.995 51.525 149.165 ;
        RECT 51.815 148.995 51.985 149.165 ;
        RECT 52.275 148.995 52.445 149.165 ;
        RECT 52.735 148.995 52.905 149.165 ;
        RECT 53.195 148.995 53.365 149.165 ;
        RECT 53.655 148.995 53.825 149.165 ;
        RECT 42.615 146.275 42.785 146.445 ;
        RECT 43.075 146.275 43.245 146.445 ;
        RECT 43.535 146.275 43.705 146.445 ;
        RECT 43.995 146.275 44.165 146.445 ;
        RECT 44.455 146.275 44.625 146.445 ;
        RECT 44.915 146.275 45.085 146.445 ;
        RECT 45.375 146.275 45.545 146.445 ;
        RECT 45.835 146.275 46.005 146.445 ;
        RECT 46.295 146.275 46.465 146.445 ;
        RECT 46.755 146.275 46.925 146.445 ;
        RECT 47.215 146.275 47.385 146.445 ;
        RECT 47.675 146.275 47.845 146.445 ;
        RECT 48.135 146.275 48.305 146.445 ;
        RECT 48.595 146.275 48.765 146.445 ;
        RECT 49.055 146.275 49.225 146.445 ;
        RECT 49.515 146.275 49.685 146.445 ;
        RECT 49.975 146.275 50.145 146.445 ;
        RECT 50.435 146.275 50.605 146.445 ;
        RECT 50.895 146.275 51.065 146.445 ;
        RECT 51.355 146.275 51.525 146.445 ;
        RECT 51.815 146.275 51.985 146.445 ;
        RECT 52.275 146.275 52.445 146.445 ;
        RECT 52.735 146.275 52.905 146.445 ;
        RECT 53.195 146.275 53.365 146.445 ;
        RECT 53.655 146.275 53.825 146.445 ;
        RECT 42.615 143.555 42.785 143.725 ;
        RECT 43.075 143.555 43.245 143.725 ;
        RECT 43.535 143.555 43.705 143.725 ;
        RECT 43.995 143.555 44.165 143.725 ;
        RECT 44.455 143.555 44.625 143.725 ;
        RECT 44.915 143.555 45.085 143.725 ;
        RECT 45.375 143.555 45.545 143.725 ;
        RECT 45.835 143.555 46.005 143.725 ;
        RECT 46.295 143.555 46.465 143.725 ;
        RECT 46.755 143.555 46.925 143.725 ;
        RECT 47.215 143.555 47.385 143.725 ;
        RECT 47.675 143.555 47.845 143.725 ;
        RECT 48.135 143.555 48.305 143.725 ;
        RECT 48.595 143.555 48.765 143.725 ;
        RECT 49.055 143.555 49.225 143.725 ;
        RECT 49.515 143.555 49.685 143.725 ;
        RECT 49.975 143.555 50.145 143.725 ;
        RECT 50.435 143.555 50.605 143.725 ;
        RECT 50.895 143.555 51.065 143.725 ;
        RECT 51.355 143.555 51.525 143.725 ;
        RECT 51.815 143.555 51.985 143.725 ;
        RECT 52.275 143.555 52.445 143.725 ;
        RECT 52.735 143.555 52.905 143.725 ;
        RECT 53.195 143.555 53.365 143.725 ;
        RECT 53.655 143.555 53.825 143.725 ;
        RECT 42.615 140.835 42.785 141.005 ;
        RECT 43.075 140.835 43.245 141.005 ;
        RECT 43.535 140.835 43.705 141.005 ;
        RECT 43.995 140.835 44.165 141.005 ;
        RECT 44.455 140.835 44.625 141.005 ;
        RECT 44.915 140.835 45.085 141.005 ;
        RECT 45.375 140.835 45.545 141.005 ;
        RECT 45.835 140.835 46.005 141.005 ;
        RECT 46.295 140.835 46.465 141.005 ;
        RECT 46.755 140.835 46.925 141.005 ;
        RECT 47.215 140.835 47.385 141.005 ;
        RECT 47.675 140.835 47.845 141.005 ;
        RECT 48.135 140.835 48.305 141.005 ;
        RECT 48.595 140.835 48.765 141.005 ;
        RECT 49.055 140.835 49.225 141.005 ;
        RECT 49.515 140.835 49.685 141.005 ;
        RECT 49.975 140.835 50.145 141.005 ;
        RECT 50.435 140.835 50.605 141.005 ;
        RECT 50.895 140.835 51.065 141.005 ;
        RECT 51.355 140.835 51.525 141.005 ;
        RECT 51.815 140.835 51.985 141.005 ;
        RECT 52.275 140.835 52.445 141.005 ;
        RECT 52.735 140.835 52.905 141.005 ;
        RECT 53.195 140.835 53.365 141.005 ;
        RECT 53.655 140.835 53.825 141.005 ;
        RECT 42.615 138.115 42.785 138.285 ;
        RECT 43.075 138.115 43.245 138.285 ;
        RECT 43.535 138.115 43.705 138.285 ;
        RECT 43.995 138.115 44.165 138.285 ;
        RECT 44.455 138.115 44.625 138.285 ;
        RECT 44.915 138.115 45.085 138.285 ;
        RECT 45.375 138.115 45.545 138.285 ;
        RECT 45.835 138.115 46.005 138.285 ;
        RECT 46.295 138.115 46.465 138.285 ;
        RECT 46.755 138.115 46.925 138.285 ;
        RECT 47.215 138.115 47.385 138.285 ;
        RECT 47.675 138.115 47.845 138.285 ;
        RECT 48.135 138.115 48.305 138.285 ;
        RECT 48.595 138.115 48.765 138.285 ;
        RECT 49.055 138.115 49.225 138.285 ;
        RECT 49.515 138.115 49.685 138.285 ;
        RECT 49.975 138.115 50.145 138.285 ;
        RECT 50.435 138.115 50.605 138.285 ;
        RECT 50.895 138.115 51.065 138.285 ;
        RECT 51.355 138.115 51.525 138.285 ;
        RECT 51.815 138.115 51.985 138.285 ;
        RECT 52.275 138.115 52.445 138.285 ;
        RECT 52.735 138.115 52.905 138.285 ;
        RECT 53.195 138.115 53.365 138.285 ;
        RECT 53.655 138.115 53.825 138.285 ;
        RECT 42.615 135.395 42.785 135.565 ;
        RECT 43.075 135.395 43.245 135.565 ;
        RECT 43.535 135.395 43.705 135.565 ;
        RECT 43.995 135.395 44.165 135.565 ;
        RECT 44.455 135.395 44.625 135.565 ;
        RECT 44.915 135.395 45.085 135.565 ;
        RECT 45.375 135.395 45.545 135.565 ;
        RECT 45.835 135.395 46.005 135.565 ;
        RECT 46.295 135.395 46.465 135.565 ;
        RECT 46.755 135.395 46.925 135.565 ;
        RECT 47.215 135.395 47.385 135.565 ;
        RECT 47.675 135.395 47.845 135.565 ;
        RECT 48.135 135.395 48.305 135.565 ;
        RECT 48.595 135.395 48.765 135.565 ;
        RECT 49.055 135.395 49.225 135.565 ;
        RECT 49.515 135.395 49.685 135.565 ;
        RECT 49.975 135.395 50.145 135.565 ;
        RECT 50.435 135.395 50.605 135.565 ;
        RECT 50.895 135.395 51.065 135.565 ;
        RECT 51.355 135.395 51.525 135.565 ;
        RECT 51.815 135.395 51.985 135.565 ;
        RECT 52.275 135.395 52.445 135.565 ;
        RECT 52.735 135.395 52.905 135.565 ;
        RECT 53.195 135.395 53.365 135.565 ;
        RECT 53.655 135.395 53.825 135.565 ;
        RECT 42.615 132.675 42.785 132.845 ;
        RECT 43.075 132.675 43.245 132.845 ;
        RECT 43.535 132.675 43.705 132.845 ;
        RECT 43.995 132.675 44.165 132.845 ;
        RECT 44.455 132.675 44.625 132.845 ;
        RECT 44.915 132.675 45.085 132.845 ;
        RECT 45.375 132.675 45.545 132.845 ;
        RECT 45.835 132.675 46.005 132.845 ;
        RECT 46.295 132.675 46.465 132.845 ;
        RECT 46.755 132.675 46.925 132.845 ;
        RECT 47.215 132.675 47.385 132.845 ;
        RECT 47.675 132.675 47.845 132.845 ;
        RECT 48.135 132.675 48.305 132.845 ;
        RECT 48.595 132.675 48.765 132.845 ;
        RECT 49.055 132.675 49.225 132.845 ;
        RECT 49.515 132.675 49.685 132.845 ;
        RECT 49.975 132.675 50.145 132.845 ;
        RECT 50.435 132.675 50.605 132.845 ;
        RECT 50.895 132.675 51.065 132.845 ;
        RECT 51.355 132.675 51.525 132.845 ;
        RECT 51.815 132.675 51.985 132.845 ;
        RECT 52.275 132.675 52.445 132.845 ;
        RECT 52.735 132.675 52.905 132.845 ;
        RECT 53.195 132.675 53.365 132.845 ;
        RECT 53.655 132.675 53.825 132.845 ;
        RECT 42.615 129.955 42.785 130.125 ;
        RECT 43.075 129.955 43.245 130.125 ;
        RECT 43.535 129.955 43.705 130.125 ;
        RECT 43.995 129.955 44.165 130.125 ;
        RECT 44.455 129.955 44.625 130.125 ;
        RECT 44.915 129.955 45.085 130.125 ;
        RECT 45.375 129.955 45.545 130.125 ;
        RECT 45.835 129.955 46.005 130.125 ;
        RECT 46.295 129.955 46.465 130.125 ;
        RECT 46.755 129.955 46.925 130.125 ;
        RECT 47.215 129.955 47.385 130.125 ;
        RECT 47.675 129.955 47.845 130.125 ;
        RECT 48.135 129.955 48.305 130.125 ;
        RECT 48.595 129.955 48.765 130.125 ;
        RECT 49.055 129.955 49.225 130.125 ;
        RECT 49.515 129.955 49.685 130.125 ;
        RECT 49.975 129.955 50.145 130.125 ;
        RECT 50.435 129.955 50.605 130.125 ;
        RECT 50.895 129.955 51.065 130.125 ;
        RECT 51.355 129.955 51.525 130.125 ;
        RECT 51.815 129.955 51.985 130.125 ;
        RECT 52.275 129.955 52.445 130.125 ;
        RECT 52.735 129.955 52.905 130.125 ;
        RECT 53.195 129.955 53.365 130.125 ;
        RECT 53.655 129.955 53.825 130.125 ;
        RECT 42.615 127.235 42.785 127.405 ;
        RECT 43.075 127.235 43.245 127.405 ;
        RECT 43.535 127.235 43.705 127.405 ;
        RECT 43.995 127.235 44.165 127.405 ;
        RECT 44.455 127.235 44.625 127.405 ;
        RECT 44.915 127.235 45.085 127.405 ;
        RECT 45.375 127.235 45.545 127.405 ;
        RECT 45.835 127.235 46.005 127.405 ;
        RECT 46.295 127.235 46.465 127.405 ;
        RECT 46.755 127.235 46.925 127.405 ;
        RECT 47.215 127.235 47.385 127.405 ;
        RECT 47.675 127.235 47.845 127.405 ;
        RECT 48.135 127.235 48.305 127.405 ;
        RECT 48.595 127.235 48.765 127.405 ;
        RECT 49.055 127.235 49.225 127.405 ;
        RECT 49.515 127.235 49.685 127.405 ;
        RECT 49.975 127.235 50.145 127.405 ;
        RECT 50.435 127.235 50.605 127.405 ;
        RECT 50.895 127.235 51.065 127.405 ;
        RECT 51.355 127.235 51.525 127.405 ;
        RECT 51.815 127.235 51.985 127.405 ;
        RECT 52.275 127.235 52.445 127.405 ;
        RECT 52.735 127.235 52.905 127.405 ;
        RECT 53.195 127.235 53.365 127.405 ;
        RECT 53.655 127.235 53.825 127.405 ;
        RECT 42.615 124.515 42.785 124.685 ;
        RECT 43.075 124.515 43.245 124.685 ;
        RECT 43.535 124.515 43.705 124.685 ;
        RECT 43.995 124.515 44.165 124.685 ;
        RECT 44.455 124.515 44.625 124.685 ;
        RECT 44.915 124.515 45.085 124.685 ;
        RECT 45.375 124.515 45.545 124.685 ;
        RECT 45.835 124.515 46.005 124.685 ;
        RECT 46.295 124.515 46.465 124.685 ;
        RECT 46.755 124.515 46.925 124.685 ;
        RECT 47.215 124.515 47.385 124.685 ;
        RECT 47.675 124.515 47.845 124.685 ;
        RECT 48.135 124.515 48.305 124.685 ;
        RECT 48.595 124.515 48.765 124.685 ;
        RECT 49.055 124.515 49.225 124.685 ;
        RECT 49.515 124.515 49.685 124.685 ;
        RECT 49.975 124.515 50.145 124.685 ;
        RECT 50.435 124.515 50.605 124.685 ;
        RECT 50.895 124.515 51.065 124.685 ;
        RECT 51.355 124.515 51.525 124.685 ;
        RECT 51.815 124.515 51.985 124.685 ;
        RECT 52.275 124.515 52.445 124.685 ;
        RECT 52.735 124.515 52.905 124.685 ;
        RECT 53.195 124.515 53.365 124.685 ;
        RECT 53.655 124.515 53.825 124.685 ;
        RECT 42.615 121.795 42.785 121.965 ;
        RECT 43.075 121.795 43.245 121.965 ;
        RECT 43.535 121.795 43.705 121.965 ;
        RECT 43.995 121.795 44.165 121.965 ;
        RECT 44.455 121.795 44.625 121.965 ;
        RECT 44.915 121.795 45.085 121.965 ;
        RECT 45.375 121.795 45.545 121.965 ;
        RECT 45.835 121.795 46.005 121.965 ;
        RECT 46.295 121.795 46.465 121.965 ;
        RECT 46.755 121.795 46.925 121.965 ;
        RECT 47.215 121.795 47.385 121.965 ;
        RECT 47.675 121.795 47.845 121.965 ;
        RECT 48.135 121.795 48.305 121.965 ;
        RECT 48.595 121.795 48.765 121.965 ;
        RECT 49.055 121.795 49.225 121.965 ;
        RECT 49.515 121.795 49.685 121.965 ;
        RECT 49.975 121.795 50.145 121.965 ;
        RECT 50.435 121.795 50.605 121.965 ;
        RECT 50.895 121.795 51.065 121.965 ;
        RECT 51.355 121.795 51.525 121.965 ;
        RECT 51.815 121.795 51.985 121.965 ;
        RECT 52.275 121.795 52.445 121.965 ;
        RECT 52.735 121.795 52.905 121.965 ;
        RECT 53.195 121.795 53.365 121.965 ;
        RECT 53.655 121.795 53.825 121.965 ;
        RECT 42.615 119.075 42.785 119.245 ;
        RECT 43.075 119.075 43.245 119.245 ;
        RECT 43.535 119.075 43.705 119.245 ;
        RECT 43.995 119.075 44.165 119.245 ;
        RECT 44.455 119.075 44.625 119.245 ;
        RECT 44.915 119.075 45.085 119.245 ;
        RECT 45.375 119.075 45.545 119.245 ;
        RECT 45.835 119.075 46.005 119.245 ;
        RECT 46.295 119.075 46.465 119.245 ;
        RECT 46.755 119.075 46.925 119.245 ;
        RECT 47.215 119.075 47.385 119.245 ;
        RECT 47.675 119.075 47.845 119.245 ;
        RECT 48.135 119.075 48.305 119.245 ;
        RECT 48.595 119.075 48.765 119.245 ;
        RECT 49.055 119.075 49.225 119.245 ;
        RECT 49.515 119.075 49.685 119.245 ;
        RECT 49.975 119.075 50.145 119.245 ;
        RECT 50.435 119.075 50.605 119.245 ;
        RECT 50.895 119.075 51.065 119.245 ;
        RECT 51.355 119.075 51.525 119.245 ;
        RECT 51.815 119.075 51.985 119.245 ;
        RECT 52.275 119.075 52.445 119.245 ;
        RECT 52.735 119.075 52.905 119.245 ;
        RECT 53.195 119.075 53.365 119.245 ;
        RECT 53.655 119.075 53.825 119.245 ;
        RECT 42.615 116.355 42.785 116.525 ;
        RECT 43.075 116.355 43.245 116.525 ;
        RECT 43.535 116.355 43.705 116.525 ;
        RECT 43.995 116.355 44.165 116.525 ;
        RECT 44.455 116.355 44.625 116.525 ;
        RECT 44.915 116.355 45.085 116.525 ;
        RECT 45.375 116.355 45.545 116.525 ;
        RECT 45.835 116.355 46.005 116.525 ;
        RECT 46.295 116.355 46.465 116.525 ;
        RECT 46.755 116.355 46.925 116.525 ;
        RECT 47.215 116.355 47.385 116.525 ;
        RECT 47.675 116.355 47.845 116.525 ;
        RECT 48.135 116.355 48.305 116.525 ;
        RECT 48.595 116.355 48.765 116.525 ;
        RECT 49.055 116.355 49.225 116.525 ;
        RECT 49.515 116.355 49.685 116.525 ;
        RECT 49.975 116.355 50.145 116.525 ;
        RECT 50.435 116.355 50.605 116.525 ;
        RECT 50.895 116.355 51.065 116.525 ;
        RECT 51.355 116.355 51.525 116.525 ;
        RECT 51.815 116.355 51.985 116.525 ;
        RECT 52.275 116.355 52.445 116.525 ;
        RECT 52.735 116.355 52.905 116.525 ;
        RECT 53.195 116.355 53.365 116.525 ;
        RECT 53.655 116.355 53.825 116.525 ;
        RECT 42.615 113.635 42.785 113.805 ;
        RECT 43.075 113.635 43.245 113.805 ;
        RECT 43.535 113.635 43.705 113.805 ;
        RECT 43.995 113.635 44.165 113.805 ;
        RECT 44.455 113.635 44.625 113.805 ;
        RECT 44.915 113.635 45.085 113.805 ;
        RECT 45.375 113.635 45.545 113.805 ;
        RECT 45.835 113.635 46.005 113.805 ;
        RECT 46.295 113.635 46.465 113.805 ;
        RECT 46.755 113.635 46.925 113.805 ;
        RECT 47.215 113.635 47.385 113.805 ;
        RECT 47.675 113.635 47.845 113.805 ;
        RECT 48.135 113.635 48.305 113.805 ;
        RECT 48.595 113.635 48.765 113.805 ;
        RECT 49.055 113.635 49.225 113.805 ;
        RECT 49.515 113.635 49.685 113.805 ;
        RECT 49.975 113.635 50.145 113.805 ;
        RECT 50.435 113.635 50.605 113.805 ;
        RECT 50.895 113.635 51.065 113.805 ;
        RECT 51.355 113.635 51.525 113.805 ;
        RECT 51.815 113.635 51.985 113.805 ;
        RECT 52.275 113.635 52.445 113.805 ;
        RECT 52.735 113.635 52.905 113.805 ;
        RECT 53.195 113.635 53.365 113.805 ;
        RECT 53.655 113.635 53.825 113.805 ;
        RECT 42.615 110.915 42.785 111.085 ;
        RECT 43.075 110.915 43.245 111.085 ;
        RECT 43.535 110.915 43.705 111.085 ;
        RECT 43.995 110.915 44.165 111.085 ;
        RECT 44.455 110.915 44.625 111.085 ;
        RECT 44.915 110.915 45.085 111.085 ;
        RECT 45.375 110.915 45.545 111.085 ;
        RECT 45.835 110.915 46.005 111.085 ;
        RECT 46.295 110.915 46.465 111.085 ;
        RECT 46.755 110.915 46.925 111.085 ;
        RECT 47.215 110.915 47.385 111.085 ;
        RECT 47.675 110.915 47.845 111.085 ;
        RECT 48.135 110.915 48.305 111.085 ;
        RECT 48.595 110.915 48.765 111.085 ;
        RECT 49.055 110.915 49.225 111.085 ;
        RECT 49.515 110.915 49.685 111.085 ;
        RECT 49.975 110.915 50.145 111.085 ;
        RECT 50.435 110.915 50.605 111.085 ;
        RECT 50.895 110.915 51.065 111.085 ;
        RECT 51.355 110.915 51.525 111.085 ;
        RECT 51.815 110.915 51.985 111.085 ;
        RECT 52.275 110.915 52.445 111.085 ;
        RECT 52.735 110.915 52.905 111.085 ;
        RECT 53.195 110.915 53.365 111.085 ;
        RECT 53.655 110.915 53.825 111.085 ;
        RECT 42.615 108.195 42.785 108.365 ;
        RECT 43.075 108.195 43.245 108.365 ;
        RECT 43.535 108.195 43.705 108.365 ;
        RECT 43.995 108.195 44.165 108.365 ;
        RECT 44.455 108.195 44.625 108.365 ;
        RECT 44.915 108.195 45.085 108.365 ;
        RECT 45.375 108.195 45.545 108.365 ;
        RECT 45.835 108.195 46.005 108.365 ;
        RECT 46.295 108.195 46.465 108.365 ;
        RECT 46.755 108.195 46.925 108.365 ;
        RECT 47.215 108.195 47.385 108.365 ;
        RECT 47.675 108.195 47.845 108.365 ;
        RECT 48.135 108.195 48.305 108.365 ;
        RECT 48.595 108.195 48.765 108.365 ;
        RECT 49.055 108.195 49.225 108.365 ;
        RECT 49.515 108.195 49.685 108.365 ;
        RECT 49.975 108.195 50.145 108.365 ;
        RECT 50.435 108.195 50.605 108.365 ;
        RECT 50.895 108.195 51.065 108.365 ;
        RECT 51.355 108.195 51.525 108.365 ;
        RECT 51.815 108.195 51.985 108.365 ;
        RECT 52.275 108.195 52.445 108.365 ;
        RECT 52.735 108.195 52.905 108.365 ;
        RECT 53.195 108.195 53.365 108.365 ;
        RECT 53.655 108.195 53.825 108.365 ;
        RECT 42.615 105.475 42.785 105.645 ;
        RECT 43.075 105.475 43.245 105.645 ;
        RECT 43.535 105.475 43.705 105.645 ;
        RECT 43.995 105.475 44.165 105.645 ;
        RECT 44.455 105.475 44.625 105.645 ;
        RECT 44.915 105.475 45.085 105.645 ;
        RECT 45.375 105.475 45.545 105.645 ;
        RECT 45.835 105.475 46.005 105.645 ;
        RECT 46.295 105.475 46.465 105.645 ;
        RECT 46.755 105.475 46.925 105.645 ;
        RECT 47.215 105.475 47.385 105.645 ;
        RECT 47.675 105.475 47.845 105.645 ;
        RECT 48.135 105.475 48.305 105.645 ;
        RECT 48.595 105.475 48.765 105.645 ;
        RECT 49.055 105.475 49.225 105.645 ;
        RECT 49.515 105.475 49.685 105.645 ;
        RECT 49.975 105.475 50.145 105.645 ;
        RECT 50.435 105.475 50.605 105.645 ;
        RECT 50.895 105.475 51.065 105.645 ;
        RECT 51.355 105.475 51.525 105.645 ;
        RECT 51.815 105.475 51.985 105.645 ;
        RECT 52.275 105.475 52.445 105.645 ;
        RECT 52.735 105.475 52.905 105.645 ;
        RECT 53.195 105.475 53.365 105.645 ;
        RECT 53.655 105.475 53.825 105.645 ;
        RECT 42.615 102.755 42.785 102.925 ;
        RECT 43.075 102.755 43.245 102.925 ;
        RECT 43.535 102.755 43.705 102.925 ;
        RECT 43.995 102.755 44.165 102.925 ;
        RECT 44.455 102.755 44.625 102.925 ;
        RECT 44.915 102.755 45.085 102.925 ;
        RECT 45.375 102.755 45.545 102.925 ;
        RECT 45.835 102.755 46.005 102.925 ;
        RECT 46.295 102.755 46.465 102.925 ;
        RECT 46.755 102.755 46.925 102.925 ;
        RECT 47.215 102.755 47.385 102.925 ;
        RECT 47.675 102.755 47.845 102.925 ;
        RECT 48.135 102.755 48.305 102.925 ;
        RECT 48.595 102.755 48.765 102.925 ;
        RECT 49.055 102.755 49.225 102.925 ;
        RECT 49.515 102.755 49.685 102.925 ;
        RECT 49.975 102.755 50.145 102.925 ;
        RECT 50.435 102.755 50.605 102.925 ;
        RECT 50.895 102.755 51.065 102.925 ;
        RECT 51.355 102.755 51.525 102.925 ;
        RECT 51.815 102.755 51.985 102.925 ;
        RECT 52.275 102.755 52.445 102.925 ;
        RECT 52.735 102.755 52.905 102.925 ;
        RECT 53.195 102.755 53.365 102.925 ;
        RECT 53.655 102.755 53.825 102.925 ;
        RECT 42.615 100.035 42.785 100.205 ;
        RECT 43.075 100.035 43.245 100.205 ;
        RECT 43.535 100.035 43.705 100.205 ;
        RECT 43.995 100.035 44.165 100.205 ;
        RECT 44.455 100.035 44.625 100.205 ;
        RECT 44.915 100.035 45.085 100.205 ;
        RECT 45.375 100.035 45.545 100.205 ;
        RECT 45.835 100.035 46.005 100.205 ;
        RECT 46.295 100.035 46.465 100.205 ;
        RECT 46.755 100.035 46.925 100.205 ;
        RECT 47.215 100.035 47.385 100.205 ;
        RECT 47.675 100.035 47.845 100.205 ;
        RECT 48.135 100.035 48.305 100.205 ;
        RECT 48.595 100.035 48.765 100.205 ;
        RECT 49.055 100.035 49.225 100.205 ;
        RECT 49.515 100.035 49.685 100.205 ;
        RECT 49.975 100.035 50.145 100.205 ;
        RECT 50.435 100.035 50.605 100.205 ;
        RECT 50.895 100.035 51.065 100.205 ;
        RECT 51.355 100.035 51.525 100.205 ;
        RECT 51.815 100.035 51.985 100.205 ;
        RECT 52.275 100.035 52.445 100.205 ;
        RECT 52.735 100.035 52.905 100.205 ;
        RECT 53.195 100.035 53.365 100.205 ;
        RECT 53.655 100.035 53.825 100.205 ;
        RECT 42.615 97.315 42.785 97.485 ;
        RECT 43.075 97.315 43.245 97.485 ;
        RECT 43.535 97.315 43.705 97.485 ;
        RECT 43.995 97.315 44.165 97.485 ;
        RECT 44.455 97.315 44.625 97.485 ;
        RECT 44.915 97.315 45.085 97.485 ;
        RECT 45.375 97.315 45.545 97.485 ;
        RECT 45.835 97.315 46.005 97.485 ;
        RECT 46.295 97.315 46.465 97.485 ;
        RECT 46.755 97.315 46.925 97.485 ;
        RECT 47.215 97.315 47.385 97.485 ;
        RECT 47.675 97.315 47.845 97.485 ;
        RECT 48.135 97.315 48.305 97.485 ;
        RECT 48.595 97.315 48.765 97.485 ;
        RECT 49.055 97.315 49.225 97.485 ;
        RECT 49.515 97.315 49.685 97.485 ;
        RECT 49.975 97.315 50.145 97.485 ;
        RECT 50.435 97.315 50.605 97.485 ;
        RECT 50.895 97.315 51.065 97.485 ;
        RECT 51.355 97.315 51.525 97.485 ;
        RECT 51.815 97.315 51.985 97.485 ;
        RECT 52.275 97.315 52.445 97.485 ;
        RECT 52.735 97.315 52.905 97.485 ;
        RECT 53.195 97.315 53.365 97.485 ;
        RECT 53.655 97.315 53.825 97.485 ;
        RECT 42.615 94.595 42.785 94.765 ;
        RECT 43.075 94.595 43.245 94.765 ;
        RECT 43.535 94.595 43.705 94.765 ;
        RECT 43.995 94.595 44.165 94.765 ;
        RECT 44.455 94.595 44.625 94.765 ;
        RECT 44.915 94.595 45.085 94.765 ;
        RECT 45.375 94.595 45.545 94.765 ;
        RECT 45.835 94.595 46.005 94.765 ;
        RECT 46.295 94.595 46.465 94.765 ;
        RECT 46.755 94.595 46.925 94.765 ;
        RECT 47.215 94.595 47.385 94.765 ;
        RECT 47.675 94.595 47.845 94.765 ;
        RECT 48.135 94.595 48.305 94.765 ;
        RECT 48.595 94.595 48.765 94.765 ;
        RECT 49.055 94.595 49.225 94.765 ;
        RECT 49.515 94.595 49.685 94.765 ;
        RECT 49.975 94.595 50.145 94.765 ;
        RECT 50.435 94.595 50.605 94.765 ;
        RECT 50.895 94.595 51.065 94.765 ;
        RECT 51.355 94.595 51.525 94.765 ;
        RECT 51.815 94.595 51.985 94.765 ;
        RECT 52.275 94.595 52.445 94.765 ;
        RECT 52.735 94.595 52.905 94.765 ;
        RECT 53.195 94.595 53.365 94.765 ;
        RECT 53.655 94.595 53.825 94.765 ;
        RECT 42.615 91.875 42.785 92.045 ;
        RECT 43.075 91.875 43.245 92.045 ;
        RECT 43.535 91.875 43.705 92.045 ;
        RECT 43.995 91.875 44.165 92.045 ;
        RECT 44.455 91.875 44.625 92.045 ;
        RECT 44.915 91.875 45.085 92.045 ;
        RECT 45.375 91.875 45.545 92.045 ;
        RECT 45.835 91.875 46.005 92.045 ;
        RECT 46.295 91.875 46.465 92.045 ;
        RECT 46.755 91.875 46.925 92.045 ;
        RECT 47.215 91.875 47.385 92.045 ;
        RECT 47.675 91.875 47.845 92.045 ;
        RECT 48.135 91.875 48.305 92.045 ;
        RECT 48.595 91.875 48.765 92.045 ;
        RECT 49.055 91.875 49.225 92.045 ;
        RECT 49.515 91.875 49.685 92.045 ;
        RECT 49.975 91.875 50.145 92.045 ;
        RECT 50.435 91.875 50.605 92.045 ;
        RECT 50.895 91.875 51.065 92.045 ;
        RECT 51.355 91.875 51.525 92.045 ;
        RECT 51.815 91.875 51.985 92.045 ;
        RECT 52.275 91.875 52.445 92.045 ;
        RECT 52.735 91.875 52.905 92.045 ;
        RECT 53.195 91.875 53.365 92.045 ;
        RECT 53.655 91.875 53.825 92.045 ;
        RECT 42.615 89.155 42.785 89.325 ;
        RECT 43.075 89.155 43.245 89.325 ;
        RECT 43.535 89.155 43.705 89.325 ;
        RECT 43.995 89.155 44.165 89.325 ;
        RECT 44.455 89.155 44.625 89.325 ;
        RECT 44.915 89.155 45.085 89.325 ;
        RECT 45.375 89.155 45.545 89.325 ;
        RECT 45.835 89.155 46.005 89.325 ;
        RECT 46.295 89.155 46.465 89.325 ;
        RECT 46.755 89.155 46.925 89.325 ;
        RECT 47.215 89.155 47.385 89.325 ;
        RECT 47.675 89.155 47.845 89.325 ;
        RECT 48.135 89.155 48.305 89.325 ;
        RECT 48.595 89.155 48.765 89.325 ;
        RECT 49.055 89.155 49.225 89.325 ;
        RECT 49.515 89.155 49.685 89.325 ;
        RECT 49.975 89.155 50.145 89.325 ;
        RECT 50.435 89.155 50.605 89.325 ;
        RECT 50.895 89.155 51.065 89.325 ;
        RECT 51.355 89.155 51.525 89.325 ;
        RECT 51.815 89.155 51.985 89.325 ;
        RECT 52.275 89.155 52.445 89.325 ;
        RECT 52.735 89.155 52.905 89.325 ;
        RECT 53.195 89.155 53.365 89.325 ;
        RECT 53.655 89.155 53.825 89.325 ;
        RECT 42.615 86.435 42.785 86.605 ;
        RECT 43.075 86.435 43.245 86.605 ;
        RECT 43.535 86.435 43.705 86.605 ;
        RECT 43.995 86.435 44.165 86.605 ;
        RECT 44.455 86.435 44.625 86.605 ;
        RECT 44.915 86.435 45.085 86.605 ;
        RECT 45.375 86.435 45.545 86.605 ;
        RECT 45.835 86.435 46.005 86.605 ;
        RECT 46.295 86.435 46.465 86.605 ;
        RECT 46.755 86.435 46.925 86.605 ;
        RECT 47.215 86.435 47.385 86.605 ;
        RECT 47.675 86.435 47.845 86.605 ;
        RECT 48.135 86.435 48.305 86.605 ;
        RECT 48.595 86.435 48.765 86.605 ;
        RECT 49.055 86.435 49.225 86.605 ;
        RECT 49.515 86.435 49.685 86.605 ;
        RECT 49.975 86.435 50.145 86.605 ;
        RECT 50.435 86.435 50.605 86.605 ;
        RECT 50.895 86.435 51.065 86.605 ;
        RECT 51.355 86.435 51.525 86.605 ;
        RECT 51.815 86.435 51.985 86.605 ;
        RECT 52.275 86.435 52.445 86.605 ;
        RECT 52.735 86.435 52.905 86.605 ;
        RECT 53.195 86.435 53.365 86.605 ;
        RECT 53.655 86.435 53.825 86.605 ;
        RECT 42.615 83.715 42.785 83.885 ;
        RECT 43.075 83.715 43.245 83.885 ;
        RECT 43.535 83.715 43.705 83.885 ;
        RECT 43.995 83.715 44.165 83.885 ;
        RECT 44.455 83.715 44.625 83.885 ;
        RECT 44.915 83.715 45.085 83.885 ;
        RECT 45.375 83.715 45.545 83.885 ;
        RECT 45.835 83.715 46.005 83.885 ;
        RECT 46.295 83.715 46.465 83.885 ;
        RECT 46.755 83.715 46.925 83.885 ;
        RECT 47.215 83.715 47.385 83.885 ;
        RECT 47.675 83.715 47.845 83.885 ;
        RECT 48.135 83.715 48.305 83.885 ;
        RECT 48.595 83.715 48.765 83.885 ;
        RECT 49.055 83.715 49.225 83.885 ;
        RECT 49.515 83.715 49.685 83.885 ;
        RECT 49.975 83.715 50.145 83.885 ;
        RECT 50.435 83.715 50.605 83.885 ;
        RECT 50.895 83.715 51.065 83.885 ;
        RECT 51.355 83.715 51.525 83.885 ;
        RECT 51.815 83.715 51.985 83.885 ;
        RECT 52.275 83.715 52.445 83.885 ;
        RECT 52.735 83.715 52.905 83.885 ;
        RECT 53.195 83.715 53.365 83.885 ;
        RECT 53.655 83.715 53.825 83.885 ;
        RECT 42.615 80.995 42.785 81.165 ;
        RECT 43.075 80.995 43.245 81.165 ;
        RECT 43.535 80.995 43.705 81.165 ;
        RECT 43.995 80.995 44.165 81.165 ;
        RECT 44.455 80.995 44.625 81.165 ;
        RECT 44.915 80.995 45.085 81.165 ;
        RECT 45.375 80.995 45.545 81.165 ;
        RECT 45.835 80.995 46.005 81.165 ;
        RECT 46.295 80.995 46.465 81.165 ;
        RECT 46.755 80.995 46.925 81.165 ;
        RECT 47.215 80.995 47.385 81.165 ;
        RECT 47.675 80.995 47.845 81.165 ;
        RECT 48.135 80.995 48.305 81.165 ;
        RECT 48.595 80.995 48.765 81.165 ;
        RECT 49.055 80.995 49.225 81.165 ;
        RECT 49.515 80.995 49.685 81.165 ;
        RECT 49.975 80.995 50.145 81.165 ;
        RECT 50.435 80.995 50.605 81.165 ;
        RECT 50.895 80.995 51.065 81.165 ;
        RECT 51.355 80.995 51.525 81.165 ;
        RECT 51.815 80.995 51.985 81.165 ;
        RECT 52.275 80.995 52.445 81.165 ;
        RECT 52.735 80.995 52.905 81.165 ;
        RECT 53.195 80.995 53.365 81.165 ;
        RECT 53.655 80.995 53.825 81.165 ;
        RECT 42.615 78.275 42.785 78.445 ;
        RECT 43.075 78.275 43.245 78.445 ;
        RECT 43.535 78.275 43.705 78.445 ;
        RECT 43.995 78.275 44.165 78.445 ;
        RECT 44.455 78.275 44.625 78.445 ;
        RECT 44.915 78.275 45.085 78.445 ;
        RECT 45.375 78.275 45.545 78.445 ;
        RECT 45.835 78.275 46.005 78.445 ;
        RECT 46.295 78.275 46.465 78.445 ;
        RECT 46.755 78.275 46.925 78.445 ;
        RECT 47.215 78.275 47.385 78.445 ;
        RECT 47.675 78.275 47.845 78.445 ;
        RECT 48.135 78.275 48.305 78.445 ;
        RECT 48.595 78.275 48.765 78.445 ;
        RECT 49.055 78.275 49.225 78.445 ;
        RECT 49.515 78.275 49.685 78.445 ;
        RECT 49.975 78.275 50.145 78.445 ;
        RECT 50.435 78.275 50.605 78.445 ;
        RECT 50.895 78.275 51.065 78.445 ;
        RECT 51.355 78.275 51.525 78.445 ;
        RECT 51.815 78.275 51.985 78.445 ;
        RECT 52.275 78.275 52.445 78.445 ;
        RECT 52.735 78.275 52.905 78.445 ;
        RECT 53.195 78.275 53.365 78.445 ;
        RECT 53.655 78.275 53.825 78.445 ;
        RECT 42.615 75.555 42.785 75.725 ;
        RECT 43.075 75.555 43.245 75.725 ;
        RECT 43.535 75.555 43.705 75.725 ;
        RECT 43.995 75.555 44.165 75.725 ;
        RECT 44.455 75.555 44.625 75.725 ;
        RECT 44.915 75.555 45.085 75.725 ;
        RECT 45.375 75.555 45.545 75.725 ;
        RECT 45.835 75.555 46.005 75.725 ;
        RECT 46.295 75.555 46.465 75.725 ;
        RECT 46.755 75.555 46.925 75.725 ;
        RECT 47.215 75.555 47.385 75.725 ;
        RECT 47.675 75.555 47.845 75.725 ;
        RECT 48.135 75.555 48.305 75.725 ;
        RECT 48.595 75.555 48.765 75.725 ;
        RECT 49.055 75.555 49.225 75.725 ;
        RECT 49.515 75.555 49.685 75.725 ;
        RECT 49.975 75.555 50.145 75.725 ;
        RECT 50.435 75.555 50.605 75.725 ;
        RECT 50.895 75.555 51.065 75.725 ;
        RECT 51.355 75.555 51.525 75.725 ;
        RECT 51.815 75.555 51.985 75.725 ;
        RECT 52.275 75.555 52.445 75.725 ;
        RECT 52.735 75.555 52.905 75.725 ;
        RECT 53.195 75.555 53.365 75.725 ;
        RECT 53.655 75.555 53.825 75.725 ;
        RECT 42.615 72.835 42.785 73.005 ;
        RECT 43.075 72.835 43.245 73.005 ;
        RECT 43.535 72.835 43.705 73.005 ;
        RECT 43.995 72.835 44.165 73.005 ;
        RECT 44.455 72.835 44.625 73.005 ;
        RECT 44.915 72.835 45.085 73.005 ;
        RECT 45.375 72.835 45.545 73.005 ;
        RECT 45.835 72.835 46.005 73.005 ;
        RECT 46.295 72.835 46.465 73.005 ;
        RECT 46.755 72.835 46.925 73.005 ;
        RECT 47.215 72.835 47.385 73.005 ;
        RECT 47.675 72.835 47.845 73.005 ;
        RECT 48.135 72.835 48.305 73.005 ;
        RECT 48.595 72.835 48.765 73.005 ;
        RECT 49.055 72.835 49.225 73.005 ;
        RECT 49.515 72.835 49.685 73.005 ;
        RECT 49.975 72.835 50.145 73.005 ;
        RECT 50.435 72.835 50.605 73.005 ;
        RECT 50.895 72.835 51.065 73.005 ;
        RECT 51.355 72.835 51.525 73.005 ;
        RECT 51.815 72.835 51.985 73.005 ;
        RECT 52.275 72.835 52.445 73.005 ;
        RECT 52.735 72.835 52.905 73.005 ;
        RECT 53.195 72.835 53.365 73.005 ;
        RECT 53.655 72.835 53.825 73.005 ;
        RECT 42.615 70.115 42.785 70.285 ;
        RECT 43.075 70.115 43.245 70.285 ;
        RECT 43.535 70.115 43.705 70.285 ;
        RECT 43.995 70.115 44.165 70.285 ;
        RECT 44.455 70.115 44.625 70.285 ;
        RECT 44.915 70.115 45.085 70.285 ;
        RECT 45.375 70.115 45.545 70.285 ;
        RECT 45.835 70.115 46.005 70.285 ;
        RECT 46.295 70.115 46.465 70.285 ;
        RECT 46.755 70.115 46.925 70.285 ;
        RECT 47.215 70.115 47.385 70.285 ;
        RECT 47.675 70.115 47.845 70.285 ;
        RECT 48.135 70.115 48.305 70.285 ;
        RECT 48.595 70.115 48.765 70.285 ;
        RECT 49.055 70.115 49.225 70.285 ;
        RECT 49.515 70.115 49.685 70.285 ;
        RECT 49.975 70.115 50.145 70.285 ;
        RECT 50.435 70.115 50.605 70.285 ;
        RECT 50.895 70.115 51.065 70.285 ;
        RECT 51.355 70.115 51.525 70.285 ;
        RECT 51.815 70.115 51.985 70.285 ;
        RECT 52.275 70.115 52.445 70.285 ;
        RECT 52.735 70.115 52.905 70.285 ;
        RECT 53.195 70.115 53.365 70.285 ;
        RECT 53.655 70.115 53.825 70.285 ;
        RECT 42.615 67.395 42.785 67.565 ;
        RECT 43.075 67.395 43.245 67.565 ;
        RECT 43.535 67.395 43.705 67.565 ;
        RECT 43.995 67.395 44.165 67.565 ;
        RECT 44.455 67.395 44.625 67.565 ;
        RECT 44.915 67.395 45.085 67.565 ;
        RECT 45.375 67.395 45.545 67.565 ;
        RECT 45.835 67.395 46.005 67.565 ;
        RECT 46.295 67.395 46.465 67.565 ;
        RECT 46.755 67.395 46.925 67.565 ;
        RECT 47.215 67.395 47.385 67.565 ;
        RECT 47.675 67.395 47.845 67.565 ;
        RECT 48.135 67.395 48.305 67.565 ;
        RECT 48.595 67.395 48.765 67.565 ;
        RECT 49.055 67.395 49.225 67.565 ;
        RECT 49.515 67.395 49.685 67.565 ;
        RECT 49.975 67.395 50.145 67.565 ;
        RECT 50.435 67.395 50.605 67.565 ;
        RECT 50.895 67.395 51.065 67.565 ;
        RECT 51.355 67.395 51.525 67.565 ;
        RECT 51.815 67.395 51.985 67.565 ;
        RECT 52.275 67.395 52.445 67.565 ;
        RECT 52.735 67.395 52.905 67.565 ;
        RECT 53.195 67.395 53.365 67.565 ;
        RECT 53.655 67.395 53.825 67.565 ;
        RECT 42.615 64.675 42.785 64.845 ;
        RECT 43.075 64.675 43.245 64.845 ;
        RECT 43.535 64.675 43.705 64.845 ;
        RECT 43.995 64.675 44.165 64.845 ;
        RECT 44.455 64.675 44.625 64.845 ;
        RECT 44.915 64.675 45.085 64.845 ;
        RECT 45.375 64.675 45.545 64.845 ;
        RECT 45.835 64.675 46.005 64.845 ;
        RECT 46.295 64.675 46.465 64.845 ;
        RECT 46.755 64.675 46.925 64.845 ;
        RECT 47.215 64.675 47.385 64.845 ;
        RECT 47.675 64.675 47.845 64.845 ;
        RECT 48.135 64.675 48.305 64.845 ;
        RECT 48.595 64.675 48.765 64.845 ;
        RECT 49.055 64.675 49.225 64.845 ;
        RECT 49.515 64.675 49.685 64.845 ;
        RECT 49.975 64.675 50.145 64.845 ;
        RECT 50.435 64.675 50.605 64.845 ;
        RECT 50.895 64.675 51.065 64.845 ;
        RECT 51.355 64.675 51.525 64.845 ;
        RECT 51.815 64.675 51.985 64.845 ;
        RECT 52.275 64.675 52.445 64.845 ;
        RECT 52.735 64.675 52.905 64.845 ;
        RECT 53.195 64.675 53.365 64.845 ;
        RECT 53.655 64.675 53.825 64.845 ;
        RECT 42.615 61.955 42.785 62.125 ;
        RECT 43.075 61.955 43.245 62.125 ;
        RECT 43.535 61.955 43.705 62.125 ;
        RECT 43.995 61.955 44.165 62.125 ;
        RECT 44.455 61.955 44.625 62.125 ;
        RECT 44.915 61.955 45.085 62.125 ;
        RECT 45.375 61.955 45.545 62.125 ;
        RECT 45.835 61.955 46.005 62.125 ;
        RECT 46.295 61.955 46.465 62.125 ;
        RECT 46.755 61.955 46.925 62.125 ;
        RECT 47.215 61.955 47.385 62.125 ;
        RECT 47.675 61.955 47.845 62.125 ;
        RECT 48.135 61.955 48.305 62.125 ;
        RECT 48.595 61.955 48.765 62.125 ;
        RECT 49.055 61.955 49.225 62.125 ;
        RECT 49.515 61.955 49.685 62.125 ;
        RECT 49.975 61.955 50.145 62.125 ;
        RECT 50.435 61.955 50.605 62.125 ;
        RECT 50.895 61.955 51.065 62.125 ;
        RECT 51.355 61.955 51.525 62.125 ;
        RECT 51.815 61.955 51.985 62.125 ;
        RECT 52.275 61.955 52.445 62.125 ;
        RECT 52.735 61.955 52.905 62.125 ;
        RECT 53.195 61.955 53.365 62.125 ;
        RECT 53.655 61.955 53.825 62.125 ;
        RECT 42.615 59.235 42.785 59.405 ;
        RECT 43.075 59.235 43.245 59.405 ;
        RECT 43.535 59.235 43.705 59.405 ;
        RECT 43.995 59.235 44.165 59.405 ;
        RECT 44.455 59.235 44.625 59.405 ;
        RECT 44.915 59.235 45.085 59.405 ;
        RECT 45.375 59.235 45.545 59.405 ;
        RECT 45.835 59.235 46.005 59.405 ;
        RECT 46.295 59.235 46.465 59.405 ;
        RECT 46.755 59.235 46.925 59.405 ;
        RECT 47.215 59.235 47.385 59.405 ;
        RECT 47.675 59.235 47.845 59.405 ;
        RECT 48.135 59.235 48.305 59.405 ;
        RECT 48.595 59.235 48.765 59.405 ;
        RECT 49.055 59.235 49.225 59.405 ;
        RECT 49.515 59.235 49.685 59.405 ;
        RECT 49.975 59.235 50.145 59.405 ;
        RECT 50.435 59.235 50.605 59.405 ;
        RECT 50.895 59.235 51.065 59.405 ;
        RECT 51.355 59.235 51.525 59.405 ;
        RECT 51.815 59.235 51.985 59.405 ;
        RECT 52.275 59.235 52.445 59.405 ;
        RECT 52.735 59.235 52.905 59.405 ;
        RECT 53.195 59.235 53.365 59.405 ;
        RECT 53.655 59.235 53.825 59.405 ;
        RECT 42.615 56.515 42.785 56.685 ;
        RECT 43.075 56.515 43.245 56.685 ;
        RECT 43.535 56.515 43.705 56.685 ;
        RECT 43.995 56.515 44.165 56.685 ;
        RECT 44.455 56.515 44.625 56.685 ;
        RECT 44.915 56.515 45.085 56.685 ;
        RECT 45.375 56.515 45.545 56.685 ;
        RECT 45.835 56.515 46.005 56.685 ;
        RECT 46.295 56.515 46.465 56.685 ;
        RECT 46.755 56.515 46.925 56.685 ;
        RECT 47.215 56.515 47.385 56.685 ;
        RECT 47.675 56.515 47.845 56.685 ;
        RECT 48.135 56.515 48.305 56.685 ;
        RECT 48.595 56.515 48.765 56.685 ;
        RECT 49.055 56.515 49.225 56.685 ;
        RECT 49.515 56.515 49.685 56.685 ;
        RECT 49.975 56.515 50.145 56.685 ;
        RECT 50.435 56.515 50.605 56.685 ;
        RECT 50.895 56.515 51.065 56.685 ;
        RECT 51.355 56.515 51.525 56.685 ;
        RECT 51.815 56.515 51.985 56.685 ;
        RECT 52.275 56.515 52.445 56.685 ;
        RECT 52.735 56.515 52.905 56.685 ;
        RECT 53.195 56.515 53.365 56.685 ;
        RECT 53.655 56.515 53.825 56.685 ;
      LAYER met1 ;
        RECT 42.470 619.400 633.960 619.880 ;
        RECT 54.000 617.160 633.960 619.400 ;
        RECT 42.470 616.680 633.960 617.160 ;
        RECT 54.000 614.440 633.960 616.680 ;
        RECT 42.470 613.960 633.960 614.440 ;
        RECT 54.000 611.720 633.960 613.960 ;
        RECT 42.470 611.240 633.960 611.720 ;
        RECT 44.380 611.040 44.700 611.100 ;
        RECT 54.000 611.040 633.960 611.240 ;
        RECT 44.380 610.900 633.960 611.040 ;
        RECT 44.380 610.840 44.700 610.900 ;
        RECT 49.440 609.340 49.760 609.400 ;
        RECT 54.000 609.340 633.960 610.900 ;
        RECT 49.440 609.200 633.960 609.340 ;
        RECT 49.440 609.140 49.760 609.200 ;
        RECT 54.000 609.000 633.960 609.200 ;
        RECT 42.470 608.520 633.960 609.000 ;
        RECT 54.000 606.280 633.960 608.520 ;
        RECT 42.470 605.800 633.960 606.280 ;
        RECT 54.000 603.560 633.960 605.800 ;
        RECT 42.470 603.080 633.960 603.560 ;
        RECT 54.000 600.840 633.960 603.080 ;
        RECT 42.470 600.360 633.960 600.840 ;
        RECT 54.000 598.120 633.960 600.360 ;
        RECT 42.470 597.640 633.960 598.120 ;
        RECT 54.000 595.400 633.960 597.640 ;
        RECT 42.470 594.920 633.960 595.400 ;
        RECT 54.000 592.680 633.960 594.920 ;
        RECT 42.470 592.200 633.960 592.680 ;
        RECT 54.000 589.960 633.960 592.200 ;
        RECT 42.470 589.480 633.960 589.960 ;
        RECT 54.000 587.240 633.960 589.480 ;
        RECT 42.470 586.760 633.960 587.240 ;
        RECT 54.000 584.520 633.960 586.760 ;
        RECT 42.470 584.040 633.960 584.520 ;
        RECT 54.000 581.800 633.960 584.040 ;
        RECT 42.470 581.320 633.960 581.800 ;
        RECT 54.000 579.080 633.960 581.320 ;
        RECT 42.470 578.600 633.960 579.080 ;
        RECT 54.000 576.360 633.960 578.600 ;
        RECT 42.470 575.880 633.960 576.360 ;
        RECT 54.000 573.640 633.960 575.880 ;
        RECT 42.470 573.160 633.960 573.640 ;
        RECT 54.000 570.920 633.960 573.160 ;
        RECT 42.470 570.440 633.960 570.920 ;
        RECT 54.000 568.200 633.960 570.440 ;
        RECT 42.470 567.720 633.960 568.200 ;
        RECT 54.000 565.480 633.960 567.720 ;
        RECT 42.470 565.000 633.960 565.480 ;
        RECT 54.000 562.760 633.960 565.000 ;
        RECT 42.470 562.280 633.960 562.760 ;
        RECT 54.000 560.040 633.960 562.280 ;
        RECT 42.470 559.560 633.960 560.040 ;
        RECT 54.000 557.320 633.960 559.560 ;
        RECT 42.470 556.840 633.960 557.320 ;
        RECT 54.000 554.600 633.960 556.840 ;
        RECT 42.470 554.120 633.960 554.600 ;
        RECT 54.000 551.880 633.960 554.120 ;
        RECT 42.470 551.400 633.960 551.880 ;
        RECT 54.000 549.160 633.960 551.400 ;
        RECT 42.470 548.680 633.960 549.160 ;
        RECT 54.000 546.440 633.960 548.680 ;
        RECT 42.470 545.960 633.960 546.440 ;
        RECT 54.000 543.720 633.960 545.960 ;
        RECT 42.470 543.240 633.960 543.720 ;
        RECT 54.000 541.000 633.960 543.240 ;
        RECT 42.470 540.520 633.960 541.000 ;
        RECT 54.000 538.280 633.960 540.520 ;
        RECT 42.470 537.800 633.960 538.280 ;
        RECT 54.000 535.560 633.960 537.800 ;
        RECT 42.470 535.080 633.960 535.560 ;
        RECT 54.000 532.840 633.960 535.080 ;
        RECT 42.470 532.360 633.960 532.840 ;
        RECT 54.000 530.120 633.960 532.360 ;
        RECT 42.470 529.640 633.960 530.120 ;
        RECT 54.000 527.400 633.960 529.640 ;
        RECT 42.470 526.920 633.960 527.400 ;
        RECT 54.000 524.680 633.960 526.920 ;
        RECT 42.470 524.200 633.960 524.680 ;
        RECT 54.000 521.960 633.960 524.200 ;
        RECT 42.470 521.480 633.960 521.960 ;
        RECT 54.000 519.240 633.960 521.480 ;
        RECT 42.470 518.760 633.960 519.240 ;
        RECT 54.000 516.520 633.960 518.760 ;
        RECT 42.470 516.040 633.960 516.520 ;
        RECT 54.000 513.800 633.960 516.040 ;
        RECT 42.470 513.320 633.960 513.800 ;
        RECT 54.000 511.080 633.960 513.320 ;
        RECT 42.470 510.600 633.960 511.080 ;
        RECT 54.000 508.360 633.960 510.600 ;
        RECT 42.470 507.880 633.960 508.360 ;
        RECT 54.000 505.640 633.960 507.880 ;
        RECT 42.470 505.160 633.960 505.640 ;
        RECT 54.000 502.920 633.960 505.160 ;
        RECT 42.470 502.440 633.960 502.920 ;
        RECT 54.000 500.200 633.960 502.440 ;
        RECT 42.470 499.720 633.960 500.200 ;
        RECT 54.000 497.480 633.960 499.720 ;
        RECT 42.470 497.000 633.960 497.480 ;
        RECT 54.000 494.760 633.960 497.000 ;
        RECT 42.470 494.280 633.960 494.760 ;
        RECT 54.000 492.040 633.960 494.280 ;
        RECT 42.470 491.560 633.960 492.040 ;
        RECT 54.000 489.320 633.960 491.560 ;
        RECT 42.470 488.840 633.960 489.320 ;
        RECT 54.000 486.600 633.960 488.840 ;
        RECT 42.470 486.120 633.960 486.600 ;
        RECT 54.000 483.880 633.960 486.120 ;
        RECT 42.470 483.400 633.960 483.880 ;
        RECT 54.000 481.160 633.960 483.400 ;
        RECT 42.470 480.680 633.960 481.160 ;
        RECT 54.000 478.440 633.960 480.680 ;
        RECT 42.470 477.960 633.960 478.440 ;
        RECT 54.000 475.720 633.960 477.960 ;
        RECT 42.470 475.240 633.960 475.720 ;
        RECT 54.000 473.000 633.960 475.240 ;
        RECT 42.470 472.520 633.960 473.000 ;
        RECT 54.000 470.280 633.960 472.520 ;
        RECT 42.470 469.800 633.960 470.280 ;
        RECT 54.000 467.560 633.960 469.800 ;
        RECT 42.470 467.080 633.960 467.560 ;
        RECT 54.000 464.840 633.960 467.080 ;
        RECT 42.470 464.360 633.960 464.840 ;
        RECT 54.000 462.120 633.960 464.360 ;
        RECT 42.470 461.640 633.960 462.120 ;
        RECT 54.000 459.400 633.960 461.640 ;
        RECT 42.470 458.920 633.960 459.400 ;
        RECT 54.000 456.680 633.960 458.920 ;
        RECT 42.470 456.200 633.960 456.680 ;
        RECT 54.000 453.960 633.960 456.200 ;
        RECT 42.470 453.480 633.960 453.960 ;
        RECT 54.000 451.240 633.960 453.480 ;
        RECT 42.470 450.760 633.960 451.240 ;
        RECT 54.000 448.520 633.960 450.760 ;
        RECT 42.470 448.040 633.960 448.520 ;
        RECT 54.000 445.800 633.960 448.040 ;
        RECT 42.470 445.320 633.960 445.800 ;
        RECT 54.000 443.080 633.960 445.320 ;
        RECT 42.470 442.600 633.960 443.080 ;
        RECT 54.000 440.360 633.960 442.600 ;
        RECT 42.470 439.880 633.960 440.360 ;
        RECT 54.000 437.640 633.960 439.880 ;
        RECT 42.470 437.160 633.960 437.640 ;
        RECT 54.000 434.920 633.960 437.160 ;
        RECT 42.470 434.440 633.960 434.920 ;
        RECT 54.000 432.200 633.960 434.440 ;
        RECT 42.470 431.720 633.960 432.200 ;
        RECT 54.000 429.480 633.960 431.720 ;
        RECT 42.470 429.000 633.960 429.480 ;
        RECT 54.000 426.760 633.960 429.000 ;
        RECT 42.470 426.280 633.960 426.760 ;
        RECT 54.000 424.040 633.960 426.280 ;
        RECT 42.470 423.560 633.960 424.040 ;
        RECT 54.000 421.320 633.960 423.560 ;
        RECT 42.470 420.840 633.960 421.320 ;
        RECT 54.000 418.600 633.960 420.840 ;
        RECT 42.470 418.120 633.960 418.600 ;
        RECT 54.000 415.880 633.960 418.120 ;
        RECT 42.470 415.400 633.960 415.880 ;
        RECT 54.000 413.160 633.960 415.400 ;
        RECT 42.470 412.680 633.960 413.160 ;
        RECT 54.000 410.440 633.960 412.680 ;
        RECT 42.470 409.960 633.960 410.440 ;
        RECT 54.000 407.720 633.960 409.960 ;
        RECT 42.470 407.240 633.960 407.720 ;
        RECT 54.000 405.000 633.960 407.240 ;
        RECT 42.470 404.520 633.960 405.000 ;
        RECT 54.000 402.280 633.960 404.520 ;
        RECT 42.470 401.800 633.960 402.280 ;
        RECT 54.000 399.560 633.960 401.800 ;
        RECT 42.470 399.080 633.960 399.560 ;
        RECT 54.000 396.840 633.960 399.080 ;
        RECT 42.470 396.360 633.960 396.840 ;
        RECT 54.000 394.120 633.960 396.360 ;
        RECT 42.470 393.640 633.960 394.120 ;
        RECT 54.000 391.400 633.960 393.640 ;
        RECT 42.470 390.920 633.960 391.400 ;
        RECT 54.000 388.680 633.960 390.920 ;
        RECT 42.470 388.200 633.960 388.680 ;
        RECT 54.000 385.960 633.960 388.200 ;
        RECT 42.470 385.480 633.960 385.960 ;
        RECT 54.000 383.240 633.960 385.480 ;
        RECT 42.470 382.760 633.960 383.240 ;
        RECT 54.000 380.520 633.960 382.760 ;
        RECT 42.470 380.040 633.960 380.520 ;
        RECT 54.000 377.800 633.960 380.040 ;
        RECT 42.470 377.320 633.960 377.800 ;
        RECT 54.000 375.080 633.960 377.320 ;
        RECT 42.470 374.600 633.960 375.080 ;
        RECT 54.000 372.360 633.960 374.600 ;
        RECT 42.470 371.880 633.960 372.360 ;
        RECT 54.000 369.640 633.960 371.880 ;
        RECT 42.470 369.160 633.960 369.640 ;
        RECT 54.000 366.920 633.960 369.160 ;
        RECT 42.470 366.440 633.960 366.920 ;
        RECT 54.000 364.200 633.960 366.440 ;
        RECT 42.470 363.720 633.960 364.200 ;
        RECT 54.000 361.480 633.960 363.720 ;
        RECT 42.470 361.000 633.960 361.480 ;
        RECT 54.000 358.760 633.960 361.000 ;
        RECT 42.470 358.280 633.960 358.760 ;
        RECT 54.000 356.040 633.960 358.280 ;
        RECT 42.470 355.560 633.960 356.040 ;
        RECT 54.000 353.320 633.960 355.560 ;
        RECT 42.470 352.840 633.960 353.320 ;
        RECT 54.000 350.600 633.960 352.840 ;
        RECT 42.470 350.120 633.960 350.600 ;
        RECT 54.000 347.880 633.960 350.120 ;
        RECT 42.470 347.400 633.960 347.880 ;
        RECT 54.000 345.160 633.960 347.400 ;
        RECT 42.470 344.680 633.960 345.160 ;
        RECT 54.000 342.440 633.960 344.680 ;
        RECT 42.470 341.960 633.960 342.440 ;
        RECT 54.000 339.720 633.960 341.960 ;
        RECT 42.470 339.240 633.960 339.720 ;
        RECT 54.000 337.000 633.960 339.240 ;
        RECT 42.470 336.520 633.960 337.000 ;
        RECT 54.000 334.280 633.960 336.520 ;
        RECT 42.470 333.800 633.960 334.280 ;
        RECT 54.000 331.560 633.960 333.800 ;
        RECT 42.470 331.080 633.960 331.560 ;
        RECT 54.000 328.840 633.960 331.080 ;
        RECT 42.470 328.360 633.960 328.840 ;
        RECT 54.000 326.120 633.960 328.360 ;
        RECT 42.470 325.640 633.960 326.120 ;
        RECT 54.000 323.400 633.960 325.640 ;
        RECT 42.470 322.920 633.960 323.400 ;
        RECT 54.000 320.680 633.960 322.920 ;
        RECT 42.470 320.200 633.960 320.680 ;
        RECT 54.000 317.960 633.960 320.200 ;
        RECT 42.470 317.480 633.960 317.960 ;
        RECT 54.000 315.240 633.960 317.480 ;
        RECT 42.470 314.760 633.960 315.240 ;
        RECT 54.000 312.520 633.960 314.760 ;
        RECT 42.470 312.040 633.960 312.520 ;
        RECT 54.000 309.800 633.960 312.040 ;
        RECT 42.470 309.320 633.960 309.800 ;
        RECT 54.000 307.080 633.960 309.320 ;
        RECT 42.470 306.600 633.960 307.080 ;
        RECT 54.000 304.360 633.960 306.600 ;
        RECT 42.470 303.880 633.960 304.360 ;
        RECT 54.000 301.640 633.960 303.880 ;
        RECT 42.470 301.160 633.960 301.640 ;
        RECT 54.000 298.920 633.960 301.160 ;
        RECT 42.470 298.440 633.960 298.920 ;
        RECT 54.000 296.200 633.960 298.440 ;
        RECT 42.470 295.720 633.960 296.200 ;
        RECT 54.000 293.480 633.960 295.720 ;
        RECT 42.470 293.000 633.960 293.480 ;
        RECT 54.000 290.760 633.960 293.000 ;
        RECT 42.470 290.280 633.960 290.760 ;
        RECT 54.000 288.040 633.960 290.280 ;
        RECT 42.470 287.560 633.960 288.040 ;
        RECT 54.000 285.320 633.960 287.560 ;
        RECT 42.470 284.840 633.960 285.320 ;
        RECT 54.000 282.600 633.960 284.840 ;
        RECT 42.470 282.120 633.960 282.600 ;
        RECT 54.000 279.880 633.960 282.120 ;
        RECT 42.470 279.400 633.960 279.880 ;
        RECT 54.000 277.160 633.960 279.400 ;
        RECT 42.470 276.680 633.960 277.160 ;
        RECT 54.000 274.440 633.960 276.680 ;
        RECT 42.470 273.960 633.960 274.440 ;
        RECT 54.000 271.720 633.960 273.960 ;
        RECT 42.470 271.240 633.960 271.720 ;
        RECT 54.000 269.000 633.960 271.240 ;
        RECT 42.470 268.520 633.960 269.000 ;
        RECT 54.000 266.280 633.960 268.520 ;
        RECT 42.470 265.800 633.960 266.280 ;
        RECT 54.000 263.560 633.960 265.800 ;
        RECT 42.470 263.080 633.960 263.560 ;
        RECT 54.000 260.840 633.960 263.080 ;
        RECT 42.470 260.360 633.960 260.840 ;
        RECT 54.000 258.120 633.960 260.360 ;
        RECT 42.470 257.640 633.960 258.120 ;
        RECT 54.000 255.400 633.960 257.640 ;
        RECT 42.470 254.920 633.960 255.400 ;
        RECT 54.000 252.680 633.960 254.920 ;
        RECT 42.470 252.200 633.960 252.680 ;
        RECT 54.000 249.960 633.960 252.200 ;
        RECT 42.470 249.480 633.960 249.960 ;
        RECT 54.000 247.240 633.960 249.480 ;
        RECT 42.470 246.760 633.960 247.240 ;
        RECT 54.000 244.520 633.960 246.760 ;
        RECT 42.470 244.040 633.960 244.520 ;
        RECT 54.000 241.800 633.960 244.040 ;
        RECT 42.470 241.320 633.960 241.800 ;
        RECT 54.000 239.080 633.960 241.320 ;
        RECT 42.470 238.600 633.960 239.080 ;
        RECT 54.000 236.360 633.960 238.600 ;
        RECT 42.470 235.880 633.960 236.360 ;
        RECT 54.000 233.640 633.960 235.880 ;
        RECT 42.470 233.160 633.960 233.640 ;
        RECT 54.000 230.920 633.960 233.160 ;
        RECT 42.470 230.440 633.960 230.920 ;
        RECT 54.000 228.200 633.960 230.440 ;
        RECT 42.470 227.720 633.960 228.200 ;
        RECT 54.000 225.480 633.960 227.720 ;
        RECT 42.470 225.000 633.960 225.480 ;
        RECT 54.000 222.760 633.960 225.000 ;
        RECT 42.470 222.280 633.960 222.760 ;
        RECT 54.000 220.040 633.960 222.280 ;
        RECT 42.470 219.560 633.960 220.040 ;
        RECT 54.000 217.320 633.960 219.560 ;
        RECT 42.470 216.840 633.960 217.320 ;
        RECT 54.000 214.600 633.960 216.840 ;
        RECT 42.470 214.120 633.960 214.600 ;
        RECT 54.000 211.880 633.960 214.120 ;
        RECT 42.470 211.400 633.960 211.880 ;
        RECT 54.000 209.160 633.960 211.400 ;
        RECT 42.470 208.680 633.960 209.160 ;
        RECT 54.000 206.440 633.960 208.680 ;
        RECT 42.470 205.960 633.960 206.440 ;
        RECT 54.000 203.720 633.960 205.960 ;
        RECT 42.470 203.240 633.960 203.720 ;
        RECT 54.000 201.000 633.960 203.240 ;
        RECT 42.470 200.520 633.960 201.000 ;
        RECT 54.000 198.280 633.960 200.520 ;
        RECT 42.470 197.800 633.960 198.280 ;
        RECT 54.000 195.560 633.960 197.800 ;
        RECT 42.470 195.080 633.960 195.560 ;
        RECT 54.000 192.840 633.960 195.080 ;
        RECT 42.470 192.360 633.960 192.840 ;
        RECT 54.000 190.120 633.960 192.360 ;
        RECT 42.470 189.640 633.960 190.120 ;
        RECT 54.000 187.400 633.960 189.640 ;
        RECT 42.470 186.920 633.960 187.400 ;
        RECT 54.000 184.680 633.960 186.920 ;
        RECT 42.470 184.200 633.960 184.680 ;
        RECT 54.000 181.960 633.960 184.200 ;
        RECT 42.470 181.480 633.960 181.960 ;
        RECT 54.000 179.240 633.960 181.480 ;
        RECT 42.470 178.760 633.960 179.240 ;
        RECT 54.000 176.520 633.960 178.760 ;
        RECT 42.470 176.040 633.960 176.520 ;
        RECT 54.000 173.800 633.960 176.040 ;
        RECT 42.470 173.320 633.960 173.800 ;
        RECT 54.000 171.080 633.960 173.320 ;
        RECT 42.470 170.600 633.960 171.080 ;
        RECT 54.000 168.360 633.960 170.600 ;
        RECT 42.470 167.880 633.960 168.360 ;
        RECT 54.000 165.640 633.960 167.880 ;
        RECT 42.470 165.160 633.960 165.640 ;
        RECT 54.000 162.920 633.960 165.160 ;
        RECT 42.470 162.440 633.960 162.920 ;
        RECT 54.000 160.200 633.960 162.440 ;
        RECT 42.470 159.720 633.960 160.200 ;
        RECT 54.000 157.480 633.960 159.720 ;
        RECT 42.470 157.000 633.960 157.480 ;
        RECT 54.000 154.760 633.960 157.000 ;
        RECT 42.470 154.280 633.960 154.760 ;
        RECT 54.000 152.040 633.960 154.280 ;
        RECT 42.470 151.560 633.960 152.040 ;
        RECT 54.000 149.320 633.960 151.560 ;
        RECT 42.470 148.840 633.960 149.320 ;
        RECT 54.000 146.600 633.960 148.840 ;
        RECT 42.470 146.120 633.960 146.600 ;
        RECT 54.000 143.880 633.960 146.120 ;
        RECT 42.470 143.400 633.960 143.880 ;
        RECT 54.000 141.160 633.960 143.400 ;
        RECT 42.470 140.680 633.960 141.160 ;
        RECT 54.000 138.440 633.960 140.680 ;
        RECT 42.470 137.960 633.960 138.440 ;
        RECT 54.000 135.720 633.960 137.960 ;
        RECT 42.470 135.240 633.960 135.720 ;
        RECT 54.000 133.000 633.960 135.240 ;
        RECT 42.470 132.520 633.960 133.000 ;
        RECT 54.000 130.280 633.960 132.520 ;
        RECT 42.470 129.800 633.960 130.280 ;
        RECT 54.000 127.560 633.960 129.800 ;
        RECT 42.470 127.080 633.960 127.560 ;
        RECT 54.000 124.840 633.960 127.080 ;
        RECT 42.470 124.360 633.960 124.840 ;
        RECT 54.000 122.120 633.960 124.360 ;
        RECT 42.470 121.640 633.960 122.120 ;
        RECT 54.000 119.400 633.960 121.640 ;
        RECT 42.470 118.920 633.960 119.400 ;
        RECT 54.000 116.680 633.960 118.920 ;
        RECT 42.470 116.200 633.960 116.680 ;
        RECT 54.000 113.960 633.960 116.200 ;
        RECT 42.470 113.480 633.960 113.960 ;
        RECT 54.000 111.240 633.960 113.480 ;
        RECT 42.470 110.760 633.960 111.240 ;
        RECT 54.000 108.520 633.960 110.760 ;
        RECT 42.470 108.040 633.960 108.520 ;
        RECT 54.000 105.800 633.960 108.040 ;
        RECT 42.470 105.320 633.960 105.800 ;
        RECT 54.000 103.080 633.960 105.320 ;
        RECT 42.470 102.600 633.960 103.080 ;
        RECT 54.000 100.360 633.960 102.600 ;
        RECT 42.470 99.880 633.960 100.360 ;
        RECT 54.000 97.640 633.960 99.880 ;
        RECT 42.470 97.160 633.960 97.640 ;
        RECT 54.000 94.920 633.960 97.160 ;
        RECT 42.470 94.440 633.960 94.920 ;
        RECT 54.000 92.200 633.960 94.440 ;
        RECT 42.470 91.720 633.960 92.200 ;
        RECT 54.000 89.480 633.960 91.720 ;
        RECT 42.470 89.000 633.960 89.480 ;
        RECT 54.000 86.760 633.960 89.000 ;
        RECT 42.470 86.280 633.960 86.760 ;
        RECT 54.000 84.040 633.960 86.280 ;
        RECT 42.470 83.560 633.960 84.040 ;
        RECT 54.000 81.320 633.960 83.560 ;
        RECT 42.470 80.840 633.960 81.320 ;
        RECT 54.000 78.600 633.960 80.840 ;
        RECT 42.470 78.120 633.960 78.600 ;
        RECT 54.000 75.880 633.960 78.120 ;
        RECT 42.470 75.400 633.960 75.880 ;
        RECT 54.000 73.160 633.960 75.400 ;
        RECT 42.470 72.680 633.960 73.160 ;
        RECT 54.000 70.440 633.960 72.680 ;
        RECT 42.470 69.960 633.960 70.440 ;
        RECT 54.000 67.720 633.960 69.960 ;
        RECT 42.470 67.240 633.960 67.720 ;
        RECT 54.000 65.000 633.960 67.240 ;
        RECT 42.470 64.520 633.960 65.000 ;
        RECT 54.000 62.280 633.960 64.520 ;
        RECT 42.470 61.800 633.960 62.280 ;
        RECT 54.000 59.560 633.960 61.800 ;
        RECT 42.470 59.080 633.960 59.560 ;
        RECT 54.000 56.840 633.960 59.080 ;
        RECT 42.470 56.360 633.960 56.840 ;
        RECT 54.000 54.120 633.960 56.360 ;
        RECT 42.470 54.000 633.960 54.120 ;
        RECT 42.470 53.640 631.270 54.000 ;
        RECT 92.680 53.440 93.000 53.500 ;
        RECT 138.680 53.440 139.000 53.500 ;
        RECT 145.120 53.440 145.440 53.500 ;
        RECT 152.020 53.440 152.340 53.500 ;
        RECT 82.190 53.300 93.000 53.440 ;
        RECT 50.820 52.760 51.140 52.820 ;
        RECT 65.080 52.760 65.400 52.820 ;
        RECT 50.820 52.620 65.400 52.760 ;
        RECT 50.820 52.560 51.140 52.620 ;
        RECT 65.080 52.560 65.400 52.620 ;
        RECT 72.900 52.760 73.220 52.820 ;
        RECT 82.190 52.760 82.330 53.300 ;
        RECT 92.680 53.240 93.000 53.300 ;
        RECT 93.230 53.300 139.000 53.440 ;
        RECT 83.040 53.100 83.330 53.145 ;
        RECT 85.360 53.100 85.650 53.145 ;
        RECT 86.740 53.100 87.030 53.145 ;
        RECT 83.040 52.960 87.030 53.100 ;
        RECT 83.040 52.915 83.330 52.960 ;
        RECT 85.360 52.915 85.650 52.960 ;
        RECT 86.740 52.915 87.030 52.960 ;
        RECT 88.080 53.100 88.400 53.160 ;
        RECT 93.230 53.100 93.370 53.300 ;
        RECT 138.680 53.240 139.000 53.300 ;
        RECT 139.690 53.300 144.430 53.440 ;
        RECT 99.120 53.100 99.440 53.160 ;
        RECT 88.080 52.960 93.370 53.100 ;
        RECT 98.290 52.960 99.440 53.100 ;
        RECT 88.080 52.900 88.400 52.960 ;
        RECT 72.900 52.620 82.330 52.760 ;
        RECT 82.575 52.760 82.865 52.805 ;
        RECT 91.760 52.760 92.080 52.820 ;
        RECT 98.290 52.760 98.430 52.960 ;
        RECT 99.120 52.900 99.440 52.960 ;
        RECT 99.600 53.100 99.890 53.145 ;
        RECT 101.920 53.100 102.210 53.145 ;
        RECT 103.300 53.100 103.590 53.145 ;
        RECT 99.600 52.960 103.590 53.100 ;
        RECT 99.600 52.915 99.890 52.960 ;
        RECT 101.920 52.915 102.210 52.960 ;
        RECT 103.300 52.915 103.590 52.960 ;
        RECT 112.020 53.100 112.310 53.145 ;
        RECT 114.340 53.100 114.630 53.145 ;
        RECT 115.720 53.100 116.010 53.145 ;
        RECT 112.020 52.960 116.010 53.100 ;
        RECT 112.020 52.915 112.310 52.960 ;
        RECT 114.340 52.915 114.630 52.960 ;
        RECT 115.720 52.915 116.010 52.960 ;
        RECT 127.660 53.100 127.950 53.145 ;
        RECT 129.980 53.100 130.270 53.145 ;
        RECT 131.360 53.100 131.650 53.145 ;
        RECT 127.660 52.960 131.650 53.100 ;
        RECT 127.660 52.915 127.950 52.960 ;
        RECT 129.980 52.915 130.270 52.960 ;
        RECT 131.360 52.915 131.650 52.960 ;
        RECT 133.160 53.100 133.480 53.160 ;
        RECT 139.140 53.100 139.460 53.160 ;
        RECT 139.690 53.100 139.830 53.300 ;
        RECT 133.160 52.960 139.830 53.100 ;
        RECT 140.080 53.100 140.370 53.145 ;
        RECT 142.400 53.100 142.690 53.145 ;
        RECT 143.780 53.100 144.070 53.145 ;
        RECT 140.080 52.960 144.070 53.100 ;
        RECT 144.290 53.100 144.430 53.300 ;
        RECT 145.120 53.300 152.340 53.440 ;
        RECT 145.120 53.240 145.440 53.300 ;
        RECT 152.020 53.240 152.340 53.300 ;
        RECT 152.480 53.440 152.800 53.500 ;
        RECT 162.155 53.440 162.445 53.485 ;
        RECT 152.480 53.300 162.445 53.440 ;
        RECT 152.480 53.240 152.800 53.300 ;
        RECT 162.155 53.255 162.445 53.300 ;
        RECT 163.520 53.440 163.840 53.500 ;
        RECT 184.220 53.440 184.540 53.500 ;
        RECT 186.520 53.440 186.840 53.500 ;
        RECT 163.520 53.300 186.840 53.440 ;
        RECT 163.520 53.240 163.840 53.300 ;
        RECT 184.220 53.240 184.540 53.300 ;
        RECT 186.520 53.240 186.840 53.300 ;
        RECT 188.360 53.440 188.680 53.500 ;
        RECT 210.900 53.440 211.220 53.500 ;
        RECT 219.180 53.440 219.500 53.500 ;
        RECT 248.160 53.440 248.480 53.500 ;
        RECT 188.360 53.300 209.290 53.440 ;
        RECT 188.360 53.240 188.680 53.300 ;
        RECT 148.340 53.100 148.660 53.160 ;
        RECT 144.290 52.960 148.660 53.100 ;
        RECT 133.160 52.900 133.480 52.960 ;
        RECT 139.140 52.900 139.460 52.960 ;
        RECT 140.080 52.915 140.370 52.960 ;
        RECT 142.400 52.915 142.690 52.960 ;
        RECT 143.780 52.915 144.070 52.960 ;
        RECT 148.340 52.900 148.660 52.960 ;
        RECT 155.720 53.100 156.010 53.145 ;
        RECT 158.040 53.100 158.330 53.145 ;
        RECT 159.420 53.100 159.710 53.145 ;
        RECT 155.720 52.960 159.710 53.100 ;
        RECT 155.720 52.915 156.010 52.960 ;
        RECT 158.040 52.915 158.330 52.960 ;
        RECT 159.420 52.915 159.710 52.960 ;
        RECT 170.900 53.100 171.190 53.145 ;
        RECT 173.220 53.100 173.510 53.145 ;
        RECT 174.600 53.100 174.890 53.145 ;
        RECT 170.900 52.960 174.890 53.100 ;
        RECT 170.900 52.915 171.190 52.960 ;
        RECT 173.220 52.915 173.510 52.960 ;
        RECT 174.600 52.915 174.890 52.960 ;
        RECT 185.620 53.100 185.910 53.145 ;
        RECT 187.940 53.100 188.230 53.145 ;
        RECT 189.320 53.100 189.610 53.145 ;
        RECT 185.620 52.960 189.610 53.100 ;
        RECT 185.620 52.915 185.910 52.960 ;
        RECT 187.940 52.915 188.230 52.960 ;
        RECT 189.320 52.915 189.610 52.960 ;
        RECT 198.500 53.100 198.790 53.145 ;
        RECT 200.820 53.100 201.110 53.145 ;
        RECT 202.200 53.100 202.490 53.145 ;
        RECT 198.500 52.960 202.490 53.100 ;
        RECT 209.150 53.100 209.290 53.300 ;
        RECT 210.900 53.300 218.950 53.440 ;
        RECT 210.900 53.240 211.220 53.300 ;
        RECT 218.810 53.100 218.950 53.300 ;
        RECT 219.180 53.300 248.480 53.440 ;
        RECT 219.180 53.240 219.500 53.300 ;
        RECT 248.160 53.240 248.480 53.300 ;
        RECT 249.080 53.440 249.400 53.500 ;
        RECT 260.120 53.440 260.440 53.500 ;
        RECT 261.960 53.440 262.280 53.500 ;
        RECT 279.440 53.440 279.760 53.500 ;
        RECT 249.080 53.300 260.440 53.440 ;
        RECT 249.080 53.240 249.400 53.300 ;
        RECT 260.120 53.240 260.440 53.300 ;
        RECT 260.670 53.300 261.730 53.440 ;
        RECT 228.840 53.100 229.160 53.160 ;
        RECT 238.040 53.100 238.360 53.160 ;
        RECT 209.150 52.960 218.030 53.100 ;
        RECT 218.810 52.960 227.690 53.100 ;
        RECT 198.500 52.915 198.790 52.960 ;
        RECT 200.820 52.915 201.110 52.960 ;
        RECT 202.200 52.915 202.490 52.960 ;
        RECT 82.575 52.620 86.010 52.760 ;
        RECT 72.900 52.560 73.220 52.620 ;
        RECT 82.575 52.575 82.865 52.620 ;
        RECT 53.120 52.420 53.440 52.480 ;
        RECT 77.515 52.420 77.805 52.465 ;
        RECT 53.120 52.280 77.805 52.420 ;
        RECT 53.120 52.220 53.440 52.280 ;
        RECT 77.515 52.235 77.805 52.280 ;
        RECT 83.955 52.420 84.245 52.465 ;
        RECT 85.320 52.420 85.640 52.480 ;
        RECT 83.955 52.280 85.640 52.420 ;
        RECT 85.870 52.420 86.010 52.620 ;
        RECT 91.760 52.620 98.430 52.760 ;
        RECT 98.660 52.760 98.980 52.820 ;
        RECT 100.040 52.760 100.360 52.820 ;
        RECT 98.660 52.620 100.360 52.760 ;
        RECT 91.760 52.560 92.080 52.620 ;
        RECT 98.660 52.560 98.980 52.620 ;
        RECT 100.040 52.560 100.360 52.620 ;
        RECT 100.515 52.760 100.805 52.805 ;
        RECT 107.400 52.760 107.720 52.820 ;
        RECT 100.515 52.620 107.720 52.760 ;
        RECT 100.515 52.575 100.805 52.620 ;
        RECT 107.400 52.560 107.720 52.620 ;
        RECT 112.935 52.760 113.225 52.805 ;
        RECT 121.660 52.760 121.980 52.820 ;
        RECT 134.095 52.760 134.385 52.805 ;
        RECT 112.935 52.620 121.980 52.760 ;
        RECT 112.935 52.575 113.225 52.620 ;
        RECT 121.660 52.560 121.980 52.620 ;
        RECT 122.210 52.620 134.385 52.760 ;
        RECT 99.135 52.420 99.425 52.465 ;
        RECT 111.555 52.420 111.845 52.465 ;
        RECT 113.380 52.420 113.700 52.480 ;
        RECT 85.870 52.280 113.700 52.420 ;
        RECT 83.955 52.235 84.245 52.280 ;
        RECT 85.320 52.220 85.640 52.280 ;
        RECT 99.135 52.235 99.425 52.280 ;
        RECT 111.555 52.235 111.845 52.280 ;
        RECT 113.380 52.220 113.700 52.280 ;
        RECT 114.300 52.420 114.620 52.480 ;
        RECT 122.210 52.420 122.350 52.620 ;
        RECT 134.095 52.575 134.385 52.620 ;
        RECT 141.900 52.760 142.220 52.820 ;
        RECT 146.515 52.760 146.805 52.805 ;
        RECT 141.900 52.620 146.805 52.760 ;
        RECT 141.900 52.560 142.220 52.620 ;
        RECT 146.515 52.575 146.805 52.620 ;
        RECT 153.860 52.760 154.180 52.820 ;
        RECT 155.255 52.760 155.545 52.805 ;
        RECT 156.620 52.760 156.940 52.820 ;
        RECT 153.860 52.620 155.545 52.760 ;
        RECT 156.425 52.620 156.940 52.760 ;
        RECT 153.860 52.560 154.180 52.620 ;
        RECT 155.255 52.575 155.545 52.620 ;
        RECT 114.300 52.280 122.350 52.420 ;
        RECT 125.800 52.420 126.120 52.480 ;
        RECT 127.195 52.420 127.485 52.465 ;
        RECT 128.560 52.420 128.880 52.480 ;
        RECT 125.800 52.280 127.485 52.420 ;
        RECT 128.365 52.280 128.880 52.420 ;
        RECT 114.300 52.220 114.620 52.280 ;
        RECT 125.800 52.220 126.120 52.280 ;
        RECT 127.195 52.235 127.485 52.280 ;
        RECT 128.560 52.220 128.880 52.280 ;
        RECT 132.240 52.420 132.560 52.480 ;
        RECT 139.600 52.420 139.920 52.480 ;
        RECT 132.240 52.280 139.920 52.420 ;
        RECT 132.240 52.220 132.560 52.280 ;
        RECT 139.600 52.220 139.920 52.280 ;
        RECT 140.995 52.420 141.285 52.465 ;
        RECT 149.720 52.420 150.040 52.480 ;
        RECT 140.995 52.280 150.040 52.420 ;
        RECT 155.330 52.420 155.470 52.575 ;
        RECT 156.620 52.560 156.940 52.620 ;
        RECT 158.920 52.760 159.240 52.820 ;
        RECT 171.800 52.760 172.120 52.820 ;
        RECT 158.920 52.620 171.110 52.760 ;
        RECT 171.605 52.620 172.120 52.760 ;
        RECT 158.920 52.560 159.240 52.620 ;
        RECT 170.420 52.420 170.740 52.480 ;
        RECT 155.330 52.280 170.740 52.420 ;
        RECT 170.970 52.420 171.110 52.620 ;
        RECT 171.800 52.560 172.120 52.620 ;
        RECT 177.335 52.575 177.625 52.805 ;
        RECT 178.700 52.760 179.020 52.820 ;
        RECT 186.535 52.760 186.825 52.805 ;
        RECT 190.660 52.760 190.980 52.820 ;
        RECT 210.455 52.760 210.745 52.805 ;
        RECT 212.280 52.760 212.600 52.820 ;
        RECT 214.600 52.760 214.890 52.805 ;
        RECT 217.380 52.760 217.670 52.805 ;
        RECT 178.700 52.620 186.290 52.760 ;
        RECT 177.410 52.420 177.550 52.575 ;
        RECT 178.700 52.560 179.020 52.620 ;
        RECT 170.970 52.280 177.550 52.420 ;
        RECT 181.920 52.420 182.240 52.480 ;
        RECT 183.760 52.420 184.080 52.480 ;
        RECT 185.155 52.420 185.445 52.465 ;
        RECT 181.920 52.280 185.445 52.420 ;
        RECT 186.150 52.420 186.290 52.620 ;
        RECT 186.535 52.620 190.980 52.760 ;
        RECT 186.535 52.575 186.825 52.620 ;
        RECT 190.660 52.560 190.980 52.620 ;
        RECT 191.210 52.620 210.745 52.760 ;
        RECT 212.085 52.620 212.600 52.760 ;
        RECT 191.210 52.420 191.350 52.620 ;
        RECT 210.455 52.575 210.745 52.620 ;
        RECT 212.280 52.560 212.600 52.620 ;
        RECT 212.830 52.620 214.350 52.760 ;
        RECT 186.150 52.280 191.350 52.420 ;
        RECT 197.560 52.420 197.880 52.480 ;
        RECT 198.035 52.420 198.325 52.465 ;
        RECT 197.560 52.280 198.325 52.420 ;
        RECT 140.995 52.235 141.285 52.280 ;
        RECT 149.720 52.220 150.040 52.280 ;
        RECT 170.420 52.220 170.740 52.280 ;
        RECT 181.920 52.220 182.240 52.280 ;
        RECT 183.760 52.220 184.080 52.280 ;
        RECT 185.155 52.235 185.445 52.280 ;
        RECT 197.560 52.220 197.880 52.280 ;
        RECT 198.035 52.235 198.325 52.280 ;
        RECT 199.415 52.420 199.705 52.465 ;
        RECT 202.620 52.420 202.940 52.480 ;
        RECT 212.830 52.420 212.970 52.620 ;
        RECT 199.415 52.280 202.940 52.420 ;
        RECT 199.415 52.235 199.705 52.280 ;
        RECT 202.620 52.220 202.940 52.280 ;
        RECT 203.170 52.280 212.970 52.420 ;
        RECT 213.200 52.420 213.520 52.480 ;
        RECT 214.210 52.420 214.350 52.620 ;
        RECT 214.600 52.620 217.670 52.760 ;
        RECT 217.890 52.760 218.030 52.960 ;
        RECT 217.890 52.620 225.850 52.760 ;
        RECT 214.600 52.575 214.890 52.620 ;
        RECT 217.380 52.575 217.670 52.620 ;
        RECT 215.515 52.420 215.805 52.465 ;
        RECT 213.200 52.280 213.715 52.420 ;
        RECT 214.210 52.280 215.805 52.420 ;
        RECT 81.640 52.080 81.960 52.140 ;
        RECT 51.370 51.940 81.960 52.080 ;
        RECT 47.140 51.740 47.460 51.800 ;
        RECT 51.370 51.740 51.510 51.940 ;
        RECT 81.640 51.880 81.960 51.940 ;
        RECT 83.500 52.080 83.790 52.125 ;
        RECT 84.900 52.080 85.190 52.125 ;
        RECT 86.740 52.080 87.030 52.125 ;
        RECT 83.500 51.940 87.030 52.080 ;
        RECT 83.500 51.895 83.790 51.940 ;
        RECT 84.900 51.895 85.190 51.940 ;
        RECT 86.740 51.895 87.030 51.940 ;
        RECT 100.060 52.080 100.350 52.125 ;
        RECT 101.460 52.080 101.750 52.125 ;
        RECT 103.300 52.080 103.590 52.125 ;
        RECT 100.060 51.940 103.590 52.080 ;
        RECT 100.060 51.895 100.350 51.940 ;
        RECT 101.460 51.895 101.750 51.940 ;
        RECT 103.300 51.895 103.590 51.940 ;
        RECT 112.480 52.080 112.770 52.125 ;
        RECT 113.880 52.080 114.170 52.125 ;
        RECT 115.720 52.080 116.010 52.125 ;
        RECT 112.480 51.940 116.010 52.080 ;
        RECT 112.480 51.895 112.770 51.940 ;
        RECT 113.880 51.895 114.170 51.940 ;
        RECT 115.720 51.895 116.010 51.940 ;
        RECT 125.340 52.080 125.660 52.140 ;
        RECT 127.640 52.080 127.960 52.140 ;
        RECT 125.340 51.940 127.960 52.080 ;
        RECT 125.340 51.880 125.660 51.940 ;
        RECT 127.640 51.880 127.960 51.940 ;
        RECT 128.120 52.080 128.410 52.125 ;
        RECT 129.520 52.080 129.810 52.125 ;
        RECT 131.360 52.080 131.650 52.125 ;
        RECT 128.120 51.940 131.650 52.080 ;
        RECT 128.120 51.895 128.410 51.940 ;
        RECT 129.520 51.895 129.810 51.940 ;
        RECT 131.360 51.895 131.650 51.940 ;
        RECT 136.840 52.080 137.160 52.140 ;
        RECT 140.060 52.080 140.380 52.140 ;
        RECT 136.840 51.940 140.380 52.080 ;
        RECT 136.840 51.880 137.160 51.940 ;
        RECT 140.060 51.880 140.380 51.940 ;
        RECT 140.540 52.080 140.830 52.125 ;
        RECT 141.940 52.080 142.230 52.125 ;
        RECT 143.780 52.080 144.070 52.125 ;
        RECT 154.780 52.080 155.100 52.140 ;
        RECT 140.540 51.940 144.070 52.080 ;
        RECT 140.540 51.895 140.830 51.940 ;
        RECT 141.940 51.895 142.230 51.940 ;
        RECT 143.780 51.895 144.070 51.940 ;
        RECT 144.290 51.940 155.100 52.080 ;
        RECT 47.140 51.600 51.510 51.740 ;
        RECT 77.500 51.740 77.820 51.800 ;
        RECT 77.975 51.740 78.265 51.785 ;
        RECT 77.500 51.600 78.265 51.740 ;
        RECT 81.730 51.740 81.870 51.880 ;
        RECT 89.475 51.740 89.765 51.785 ;
        RECT 81.730 51.600 89.765 51.740 ;
        RECT 47.140 51.540 47.460 51.600 ;
        RECT 77.500 51.540 77.820 51.600 ;
        RECT 77.975 51.555 78.265 51.600 ;
        RECT 89.475 51.555 89.765 51.600 ;
        RECT 89.920 51.740 90.240 51.800 ;
        RECT 106.035 51.740 106.325 51.785 ;
        RECT 89.920 51.600 106.325 51.740 ;
        RECT 89.920 51.540 90.240 51.600 ;
        RECT 106.035 51.555 106.325 51.600 ;
        RECT 108.320 51.740 108.640 51.800 ;
        RECT 118.455 51.740 118.745 51.785 ;
        RECT 108.320 51.600 118.745 51.740 ;
        RECT 108.320 51.540 108.640 51.600 ;
        RECT 118.455 51.555 118.745 51.600 ;
        RECT 119.360 51.740 119.680 51.800 ;
        RECT 133.160 51.740 133.480 51.800 ;
        RECT 119.360 51.600 133.480 51.740 ;
        RECT 119.360 51.540 119.680 51.600 ;
        RECT 133.160 51.540 133.480 51.600 ;
        RECT 138.680 51.740 139.000 51.800 ;
        RECT 144.290 51.740 144.430 51.940 ;
        RECT 154.780 51.880 155.100 51.940 ;
        RECT 156.180 52.080 156.470 52.125 ;
        RECT 157.580 52.080 157.870 52.125 ;
        RECT 159.420 52.080 159.710 52.125 ;
        RECT 156.180 51.940 159.710 52.080 ;
        RECT 156.180 51.895 156.470 51.940 ;
        RECT 157.580 51.895 157.870 51.940 ;
        RECT 159.420 51.895 159.710 51.940 ;
        RECT 171.360 52.080 171.650 52.125 ;
        RECT 172.760 52.080 173.050 52.125 ;
        RECT 174.600 52.080 174.890 52.125 ;
        RECT 171.360 51.940 174.890 52.080 ;
        RECT 171.360 51.895 171.650 51.940 ;
        RECT 172.760 51.895 173.050 51.940 ;
        RECT 174.600 51.895 174.890 51.940 ;
        RECT 178.240 52.080 178.560 52.140 ;
        RECT 186.080 52.080 186.370 52.125 ;
        RECT 187.480 52.080 187.770 52.125 ;
        RECT 189.320 52.080 189.610 52.125 ;
        RECT 178.240 51.940 185.830 52.080 ;
        RECT 178.240 51.880 178.560 51.940 ;
        RECT 138.680 51.600 144.430 51.740 ;
        RECT 185.690 51.740 185.830 51.940 ;
        RECT 186.080 51.940 189.610 52.080 ;
        RECT 186.080 51.895 186.370 51.940 ;
        RECT 187.480 51.895 187.770 51.940 ;
        RECT 189.320 51.895 189.610 51.940 ;
        RECT 190.660 52.080 190.980 52.140 ;
        RECT 198.960 52.080 199.250 52.125 ;
        RECT 200.360 52.080 200.650 52.125 ;
        RECT 202.200 52.080 202.490 52.125 ;
        RECT 190.660 51.940 192.270 52.080 ;
        RECT 190.660 51.880 190.980 51.940 ;
        RECT 191.580 51.740 191.900 51.800 ;
        RECT 192.130 51.785 192.270 51.940 ;
        RECT 198.960 51.940 202.490 52.080 ;
        RECT 198.960 51.895 199.250 51.940 ;
        RECT 200.360 51.895 200.650 51.940 ;
        RECT 202.200 51.895 202.490 51.940 ;
        RECT 185.690 51.600 191.900 51.740 ;
        RECT 138.680 51.540 139.000 51.600 ;
        RECT 191.580 51.540 191.900 51.600 ;
        RECT 192.055 51.555 192.345 51.785 ;
        RECT 197.100 51.740 197.420 51.800 ;
        RECT 203.170 51.740 203.310 52.280 ;
        RECT 213.200 52.220 213.520 52.280 ;
        RECT 215.515 52.235 215.805 52.280 ;
        RECT 215.975 52.420 216.265 52.465 ;
        RECT 220.100 52.420 220.420 52.480 ;
        RECT 225.710 52.465 225.850 52.620 ;
        RECT 226.095 52.575 226.385 52.805 ;
        RECT 227.550 52.760 227.690 52.960 ;
        RECT 228.840 52.960 238.360 53.100 ;
        RECT 228.840 52.900 229.160 52.960 ;
        RECT 238.040 52.900 238.360 52.960 ;
        RECT 238.960 53.100 239.280 53.160 ;
        RECT 252.760 53.100 253.080 53.160 ;
        RECT 260.670 53.100 260.810 53.300 ;
        RECT 238.960 52.960 253.080 53.100 ;
        RECT 238.960 52.900 239.280 52.960 ;
        RECT 252.760 52.900 253.080 52.960 ;
        RECT 257.910 52.960 260.810 53.100 ;
        RECT 234.835 52.760 235.125 52.805 ;
        RECT 243.100 52.760 243.420 52.820 ;
        RECT 227.550 52.620 232.290 52.760 ;
        RECT 215.975 52.280 220.420 52.420 ;
        RECT 215.975 52.235 216.265 52.280 ;
        RECT 220.100 52.220 220.420 52.280 ;
        RECT 223.335 52.235 223.625 52.465 ;
        RECT 225.635 52.235 225.925 52.465 ;
        RECT 210.455 52.080 210.745 52.125 ;
        RECT 223.410 52.080 223.550 52.235 ;
        RECT 210.455 51.940 223.550 52.080 ;
        RECT 210.455 51.895 210.745 51.940 ;
        RECT 197.100 51.600 203.310 51.740 ;
        RECT 204.000 51.740 204.320 51.800 ;
        RECT 204.935 51.740 205.225 51.785 ;
        RECT 204.000 51.600 205.225 51.740 ;
        RECT 197.100 51.540 197.420 51.600 ;
        RECT 204.000 51.540 204.320 51.600 ;
        RECT 204.935 51.555 205.225 51.600 ;
        RECT 205.380 51.740 205.700 51.800 ;
        RECT 218.275 51.740 218.565 51.785 ;
        RECT 205.380 51.600 218.565 51.740 ;
        RECT 205.380 51.540 205.700 51.600 ;
        RECT 218.275 51.555 218.565 51.600 ;
        RECT 225.160 51.740 225.480 51.800 ;
        RECT 226.170 51.740 226.310 52.575 ;
        RECT 226.540 52.420 226.860 52.480 ;
        RECT 228.840 52.420 229.160 52.480 ;
        RECT 232.150 52.465 232.290 52.620 ;
        RECT 234.835 52.620 243.420 52.760 ;
        RECT 234.835 52.575 235.125 52.620 ;
        RECT 243.100 52.560 243.420 52.620 ;
        RECT 247.260 52.760 247.550 52.805 ;
        RECT 250.040 52.760 250.330 52.805 ;
        RECT 247.260 52.620 250.330 52.760 ;
        RECT 247.260 52.575 247.550 52.620 ;
        RECT 250.040 52.575 250.330 52.620 ;
        RECT 256.440 52.760 256.760 52.820 ;
        RECT 256.440 52.620 256.955 52.760 ;
        RECT 256.440 52.560 256.760 52.620 ;
        RECT 231.155 52.420 231.445 52.465 ;
        RECT 226.540 52.280 231.445 52.420 ;
        RECT 226.540 52.220 226.860 52.280 ;
        RECT 228.840 52.220 229.160 52.280 ;
        RECT 231.155 52.235 231.445 52.280 ;
        RECT 232.075 52.235 232.365 52.465 ;
        RECT 232.535 52.420 232.825 52.465 ;
        RECT 235.280 52.420 235.600 52.480 ;
        RECT 232.535 52.280 235.600 52.420 ;
        RECT 232.535 52.235 232.825 52.280 ;
        RECT 235.280 52.220 235.600 52.280 ;
        RECT 238.040 52.420 238.360 52.480 ;
        RECT 239.435 52.420 239.725 52.465 ;
        RECT 238.040 52.280 239.725 52.420 ;
        RECT 238.040 52.220 238.360 52.280 ;
        RECT 239.435 52.235 239.725 52.280 ;
        RECT 244.955 52.235 245.245 52.465 ;
        RECT 245.875 52.420 246.165 52.465 ;
        RECT 248.635 52.420 248.925 52.465 ;
        RECT 249.080 52.420 249.400 52.480 ;
        RECT 245.875 52.280 249.400 52.420 ;
        RECT 245.875 52.235 246.165 52.280 ;
        RECT 248.635 52.235 248.925 52.280 ;
        RECT 230.220 52.080 230.540 52.140 ;
        RECT 235.740 52.080 236.060 52.140 ;
        RECT 230.220 51.940 236.060 52.080 ;
        RECT 245.030 52.080 245.170 52.235 ;
        RECT 249.080 52.220 249.400 52.280 ;
        RECT 249.540 52.420 249.860 52.480 ;
        RECT 256.915 52.420 257.205 52.465 ;
        RECT 257.910 52.420 258.050 52.960 ;
        RECT 258.300 52.760 258.590 52.805 ;
        RECT 261.080 52.760 261.370 52.805 ;
        RECT 258.300 52.620 261.370 52.760 ;
        RECT 258.300 52.575 258.590 52.620 ;
        RECT 261.080 52.575 261.370 52.620 ;
        RECT 249.540 52.280 250.055 52.420 ;
        RECT 256.915 52.280 258.050 52.420 ;
        RECT 258.740 52.420 259.060 52.480 ;
        RECT 259.215 52.420 259.505 52.465 ;
        RECT 258.740 52.280 259.505 52.420 ;
        RECT 249.540 52.220 249.860 52.280 ;
        RECT 256.915 52.235 257.205 52.280 ;
        RECT 258.740 52.220 259.060 52.280 ;
        RECT 259.215 52.235 259.505 52.280 ;
        RECT 259.675 52.420 259.965 52.465 ;
        RECT 261.590 52.420 261.730 53.300 ;
        RECT 261.960 53.300 279.760 53.440 ;
        RECT 261.960 53.240 262.280 53.300 ;
        RECT 279.440 53.240 279.760 53.300 ;
        RECT 279.900 53.440 280.220 53.500 ;
        RECT 290.480 53.440 290.800 53.500 ;
        RECT 279.900 53.300 290.800 53.440 ;
        RECT 279.900 53.240 280.220 53.300 ;
        RECT 290.480 53.240 290.800 53.300 ;
        RECT 328.660 53.440 328.980 53.500 ;
        RECT 350.280 53.440 350.600 53.500 ;
        RECT 371.900 53.440 372.220 53.500 ;
        RECT 382.020 53.440 382.340 53.500 ;
        RECT 328.660 53.300 350.600 53.440 ;
        RECT 328.660 53.240 328.980 53.300 ;
        RECT 350.280 53.240 350.600 53.300 ;
        RECT 352.210 53.300 371.670 53.440 ;
        RECT 268.400 53.100 268.720 53.160 ;
        RECT 302.900 53.100 303.220 53.160 ;
        RECT 327.740 53.100 328.060 53.160 ;
        RECT 342.920 53.100 343.240 53.160 ;
        RECT 268.400 52.960 303.220 53.100 ;
        RECT 268.400 52.900 268.720 52.960 ;
        RECT 302.900 52.900 303.220 52.960 ;
        RECT 305.750 52.960 328.060 53.100 ;
        RECT 261.960 52.760 262.280 52.820 ;
        RECT 273.000 52.760 273.320 52.820 ;
        RECT 261.960 52.620 262.475 52.760 ;
        RECT 267.110 52.620 273.320 52.760 ;
        RECT 261.960 52.560 262.280 52.620 ;
        RECT 267.110 52.420 267.250 52.620 ;
        RECT 273.000 52.560 273.320 52.620 ;
        RECT 273.480 52.760 273.770 52.805 ;
        RECT 276.260 52.760 276.550 52.805 ;
        RECT 277.140 52.760 277.460 52.820 ;
        RECT 273.480 52.620 276.550 52.760 ;
        RECT 276.945 52.620 277.460 52.760 ;
        RECT 273.480 52.575 273.770 52.620 ;
        RECT 276.260 52.575 276.550 52.620 ;
        RECT 277.140 52.560 277.460 52.620 ;
        RECT 277.600 52.760 277.920 52.820 ;
        RECT 284.040 52.760 284.360 52.820 ;
        RECT 277.600 52.620 284.360 52.760 ;
        RECT 277.600 52.560 277.920 52.620 ;
        RECT 284.040 52.560 284.360 52.620 ;
        RECT 284.520 52.760 284.810 52.805 ;
        RECT 287.300 52.760 287.590 52.805 ;
        RECT 288.180 52.760 288.500 52.820 ;
        RECT 305.750 52.760 305.890 52.960 ;
        RECT 327.740 52.900 328.060 52.960 ;
        RECT 342.090 52.960 343.240 53.100 ;
        RECT 308.440 52.760 308.730 52.805 ;
        RECT 311.220 52.760 311.510 52.805 ;
        RECT 284.520 52.620 287.590 52.760 ;
        RECT 287.985 52.620 288.500 52.760 ;
        RECT 284.520 52.575 284.810 52.620 ;
        RECT 287.300 52.575 287.590 52.620 ;
        RECT 288.180 52.560 288.500 52.620 ;
        RECT 296.550 52.620 305.890 52.760 ;
        RECT 307.130 52.620 308.190 52.760 ;
        RECT 259.675 52.280 267.250 52.420 ;
        RECT 270.240 52.420 270.560 52.480 ;
        RECT 272.095 52.420 272.385 52.465 ;
        RECT 270.240 52.280 272.385 52.420 ;
        RECT 259.675 52.235 259.965 52.280 ;
        RECT 270.240 52.220 270.560 52.280 ;
        RECT 272.095 52.235 272.385 52.280 ;
        RECT 272.540 52.420 272.860 52.480 ;
        RECT 274.380 52.420 274.700 52.480 ;
        RECT 272.540 52.280 273.055 52.420 ;
        RECT 274.185 52.280 274.700 52.420 ;
        RECT 272.540 52.220 272.860 52.280 ;
        RECT 274.380 52.220 274.700 52.280 ;
        RECT 274.855 52.420 275.145 52.465 ;
        RECT 275.300 52.420 275.620 52.480 ;
        RECT 282.660 52.420 282.980 52.480 ;
        RECT 274.855 52.280 282.980 52.420 ;
        RECT 274.855 52.235 275.145 52.280 ;
        RECT 275.300 52.220 275.620 52.280 ;
        RECT 282.660 52.220 282.980 52.280 ;
        RECT 283.135 52.235 283.425 52.465 ;
        RECT 283.580 52.420 283.900 52.480 ;
        RECT 285.420 52.420 285.740 52.480 ;
        RECT 283.580 52.280 284.095 52.420 ;
        RECT 285.225 52.280 285.740 52.420 ;
        RECT 281.740 52.080 282.060 52.140 ;
        RECT 245.030 51.940 258.050 52.080 ;
        RECT 230.220 51.880 230.540 51.940 ;
        RECT 235.740 51.880 236.060 51.940 ;
        RECT 225.160 51.600 226.310 51.740 ;
        RECT 227.000 51.740 227.320 51.800 ;
        RECT 240.355 51.740 240.645 51.785 ;
        RECT 227.000 51.600 240.645 51.740 ;
        RECT 225.160 51.540 225.480 51.600 ;
        RECT 227.000 51.540 227.320 51.600 ;
        RECT 240.355 51.555 240.645 51.600 ;
        RECT 241.720 51.740 242.040 51.800 ;
        RECT 244.940 51.740 245.260 51.800 ;
        RECT 241.720 51.600 245.260 51.740 ;
        RECT 241.720 51.540 242.040 51.600 ;
        RECT 244.940 51.540 245.260 51.600 ;
        RECT 250.935 51.740 251.225 51.785 ;
        RECT 251.380 51.740 251.700 51.800 ;
        RECT 250.935 51.600 251.700 51.740 ;
        RECT 250.935 51.555 251.225 51.600 ;
        RECT 251.380 51.540 251.700 51.600 ;
        RECT 251.840 51.740 252.160 51.800 ;
        RECT 253.680 51.740 254.000 51.800 ;
        RECT 256.440 51.740 256.760 51.800 ;
        RECT 251.840 51.600 256.760 51.740 ;
        RECT 257.910 51.740 258.050 51.940 ;
        RECT 262.510 51.940 282.060 52.080 ;
        RECT 283.210 52.080 283.350 52.235 ;
        RECT 283.580 52.220 283.900 52.280 ;
        RECT 285.420 52.220 285.740 52.280 ;
        RECT 285.895 52.420 286.185 52.465 ;
        RECT 295.540 52.420 295.860 52.480 ;
        RECT 285.895 52.280 295.860 52.420 ;
        RECT 285.895 52.235 286.185 52.280 ;
        RECT 285.970 52.080 286.110 52.235 ;
        RECT 295.540 52.220 295.860 52.280 ;
        RECT 283.210 51.940 286.110 52.080 ;
        RECT 286.340 52.080 286.660 52.140 ;
        RECT 296.550 52.080 296.690 52.620 ;
        RECT 296.935 52.235 297.225 52.465 ;
        RECT 298.300 52.420 298.620 52.480 ;
        RECT 307.130 52.465 307.270 52.620 ;
        RECT 298.105 52.280 298.620 52.420 ;
        RECT 286.340 51.940 296.690 52.080 ;
        RECT 262.510 51.740 262.650 51.940 ;
        RECT 281.740 51.880 282.060 51.940 ;
        RECT 286.340 51.880 286.660 51.940 ;
        RECT 257.910 51.600 262.650 51.740 ;
        RECT 274.840 51.740 275.160 51.800 ;
        RECT 280.360 51.740 280.680 51.800 ;
        RECT 274.840 51.600 280.680 51.740 ;
        RECT 251.840 51.540 252.160 51.600 ;
        RECT 253.680 51.540 254.000 51.600 ;
        RECT 256.440 51.540 256.760 51.600 ;
        RECT 274.840 51.540 275.160 51.600 ;
        RECT 280.360 51.540 280.680 51.600 ;
        RECT 287.720 51.740 288.040 51.800 ;
        RECT 296.015 51.740 296.305 51.785 ;
        RECT 287.720 51.600 296.305 51.740 ;
        RECT 297.010 51.740 297.150 52.235 ;
        RECT 298.300 52.220 298.620 52.280 ;
        RECT 307.055 52.235 307.345 52.465 ;
        RECT 307.515 52.235 307.805 52.465 ;
        RECT 308.050 52.420 308.190 52.620 ;
        RECT 308.440 52.620 311.510 52.760 ;
        RECT 308.440 52.575 308.730 52.620 ;
        RECT 311.220 52.575 311.510 52.620 ;
        RECT 315.320 52.760 315.640 52.820 ;
        RECT 320.840 52.760 321.160 52.820 ;
        RECT 326.820 52.760 327.140 52.820 ;
        RECT 329.580 52.760 329.900 52.820 ;
        RECT 315.320 52.620 321.160 52.760 ;
        RECT 315.320 52.560 315.640 52.620 ;
        RECT 320.840 52.560 321.160 52.620 ;
        RECT 321.390 52.620 324.290 52.760 ;
        RECT 308.880 52.420 309.200 52.480 ;
        RECT 308.050 52.280 309.200 52.420 ;
        RECT 307.590 52.080 307.730 52.235 ;
        RECT 308.880 52.220 309.200 52.280 ;
        RECT 309.800 52.420 310.120 52.480 ;
        RECT 310.735 52.420 311.025 52.465 ;
        RECT 311.640 52.420 311.960 52.480 ;
        RECT 317.160 52.420 317.480 52.480 ;
        RECT 309.800 52.280 310.315 52.420 ;
        RECT 310.735 52.280 311.960 52.420 ;
        RECT 316.965 52.280 317.480 52.420 ;
        RECT 309.800 52.220 310.120 52.280 ;
        RECT 310.735 52.235 311.025 52.280 ;
        RECT 311.640 52.220 311.960 52.280 ;
        RECT 317.160 52.220 317.480 52.280 ;
        RECT 318.080 52.420 318.400 52.480 ;
        RECT 321.390 52.420 321.530 52.620 ;
        RECT 323.600 52.420 323.920 52.480 ;
        RECT 318.080 52.280 321.530 52.420 ;
        RECT 323.405 52.280 323.920 52.420 ;
        RECT 324.150 52.420 324.290 52.620 ;
        RECT 326.820 52.620 329.900 52.760 ;
        RECT 326.820 52.560 327.140 52.620 ;
        RECT 329.580 52.560 329.900 52.620 ;
        RECT 331.440 52.760 331.730 52.805 ;
        RECT 334.220 52.760 334.510 52.805 ;
        RECT 335.100 52.760 335.420 52.820 ;
        RECT 331.440 52.620 334.510 52.760 ;
        RECT 334.905 52.620 335.420 52.760 ;
        RECT 331.440 52.575 331.730 52.620 ;
        RECT 334.220 52.575 334.510 52.620 ;
        RECT 335.100 52.560 335.420 52.620 ;
        RECT 340.635 52.760 340.925 52.805 ;
        RECT 342.090 52.760 342.230 52.960 ;
        RECT 342.920 52.900 343.240 52.960 ;
        RECT 340.635 52.620 342.230 52.760 ;
        RECT 342.480 52.760 342.770 52.805 ;
        RECT 345.260 52.760 345.550 52.805 ;
        RECT 346.140 52.760 346.460 52.820 ;
        RECT 352.210 52.805 352.350 53.300 ;
        RECT 352.580 53.100 352.900 53.160 ;
        RECT 371.530 53.100 371.670 53.300 ;
        RECT 371.900 53.300 382.340 53.440 ;
        RECT 371.900 53.240 372.220 53.300 ;
        RECT 382.020 53.240 382.340 53.300 ;
        RECT 377.420 53.100 377.740 53.160 ;
        RECT 385.715 53.100 386.005 53.145 ;
        RECT 352.580 52.960 365.690 53.100 ;
        RECT 371.530 52.960 373.510 53.100 ;
        RECT 352.580 52.900 352.900 52.960 ;
        RECT 342.480 52.620 345.550 52.760 ;
        RECT 345.945 52.620 346.460 52.760 ;
        RECT 340.635 52.575 340.925 52.620 ;
        RECT 342.480 52.575 342.770 52.620 ;
        RECT 345.260 52.575 345.550 52.620 ;
        RECT 346.140 52.560 346.460 52.620 ;
        RECT 352.135 52.575 352.425 52.805 ;
        RECT 353.980 52.760 354.270 52.805 ;
        RECT 356.760 52.760 357.050 52.805 ;
        RECT 357.640 52.760 357.960 52.820 ;
        RECT 353.980 52.620 357.050 52.760 ;
        RECT 357.445 52.620 357.960 52.760 ;
        RECT 353.980 52.575 354.270 52.620 ;
        RECT 356.760 52.575 357.050 52.620 ;
        RECT 357.640 52.560 357.960 52.620 ;
        RECT 358.560 52.760 358.880 52.820 ;
        RECT 365.550 52.805 365.690 52.960 ;
        RECT 358.560 52.620 365.230 52.760 ;
        RECT 358.560 52.560 358.880 52.620 ;
        RECT 327.740 52.420 328.060 52.480 ;
        RECT 329.120 52.420 329.440 52.480 ;
        RECT 330.040 52.420 330.360 52.480 ;
        RECT 332.340 52.420 332.660 52.480 ;
        RECT 324.150 52.280 328.060 52.420 ;
        RECT 328.925 52.280 329.440 52.420 ;
        RECT 329.845 52.280 330.360 52.420 ;
        RECT 332.145 52.280 332.660 52.420 ;
        RECT 318.080 52.220 318.400 52.280 ;
        RECT 323.600 52.220 323.920 52.280 ;
        RECT 327.740 52.220 328.060 52.280 ;
        RECT 329.120 52.220 329.440 52.280 ;
        RECT 330.040 52.220 330.360 52.280 ;
        RECT 332.340 52.220 332.660 52.280 ;
        RECT 332.800 52.420 333.120 52.480 ;
        RECT 341.020 52.420 341.310 52.465 ;
        RECT 343.380 52.420 343.700 52.480 ;
        RECT 332.800 52.280 333.315 52.420 ;
        RECT 341.020 52.280 342.690 52.420 ;
        RECT 343.185 52.280 343.700 52.420 ;
        RECT 332.800 52.220 333.120 52.280 ;
        RECT 341.020 52.235 341.310 52.280 ;
        RECT 334.180 52.080 334.500 52.140 ;
        RECT 307.590 51.940 334.500 52.080 ;
        RECT 342.550 52.080 342.690 52.280 ;
        RECT 343.380 52.220 343.700 52.280 ;
        RECT 343.855 52.420 344.145 52.465 ;
        RECT 351.660 52.420 351.980 52.480 ;
        RECT 343.855 52.280 351.980 52.420 ;
        RECT 343.855 52.235 344.145 52.280 ;
        RECT 343.930 52.080 344.070 52.235 ;
        RECT 351.660 52.220 351.980 52.280 ;
        RECT 352.595 52.235 352.885 52.465 ;
        RECT 353.500 52.420 353.820 52.480 ;
        RECT 354.895 52.420 355.185 52.465 ;
        RECT 353.500 52.280 355.185 52.420 ;
        RECT 342.550 51.940 344.070 52.080 ;
        RECT 352.670 52.080 352.810 52.235 ;
        RECT 353.500 52.220 353.820 52.280 ;
        RECT 354.895 52.235 355.185 52.280 ;
        RECT 355.355 52.420 355.645 52.465 ;
        RECT 358.100 52.420 358.420 52.480 ;
        RECT 365.090 52.465 365.230 52.620 ;
        RECT 365.475 52.575 365.765 52.805 ;
        RECT 355.355 52.280 358.420 52.420 ;
        RECT 355.355 52.235 355.645 52.280 ;
        RECT 355.430 52.080 355.570 52.235 ;
        RECT 358.100 52.220 358.420 52.280 ;
        RECT 364.095 52.235 364.385 52.465 ;
        RECT 365.015 52.420 365.305 52.465 ;
        RECT 368.680 52.420 369.000 52.480 ;
        RECT 365.015 52.280 369.000 52.420 ;
        RECT 365.015 52.235 365.305 52.280 ;
        RECT 352.670 51.940 355.570 52.080 ;
        RECT 359.480 52.080 359.800 52.140 ;
        RECT 364.170 52.080 364.310 52.235 ;
        RECT 368.680 52.220 369.000 52.280 ;
        RECT 371.915 52.235 372.205 52.465 ;
        RECT 372.820 52.420 373.140 52.480 ;
        RECT 372.625 52.280 373.140 52.420 ;
        RECT 373.370 52.420 373.510 52.960 ;
        RECT 377.420 52.960 386.005 53.100 ;
        RECT 377.420 52.900 377.740 52.960 ;
        RECT 385.715 52.915 386.005 52.960 ;
        RECT 375.120 52.760 375.440 52.820 ;
        RECT 380.655 52.760 380.945 52.805 ;
        RECT 375.120 52.620 380.945 52.760 ;
        RECT 375.120 52.560 375.440 52.620 ;
        RECT 380.655 52.575 380.945 52.620 ;
        RECT 387.540 52.420 387.860 52.480 ;
        RECT 373.370 52.280 387.860 52.420 ;
        RECT 371.990 52.080 372.130 52.235 ;
        RECT 372.820 52.220 373.140 52.280 ;
        RECT 387.540 52.220 387.860 52.280 ;
        RECT 388.460 52.420 388.780 52.480 ;
        RECT 390.775 52.420 391.065 52.465 ;
        RECT 388.460 52.280 391.065 52.420 ;
        RECT 388.460 52.220 388.780 52.280 ;
        RECT 390.775 52.235 391.065 52.280 ;
        RECT 624.915 52.420 625.205 52.465 ;
        RECT 630.880 52.420 631.200 52.480 ;
        RECT 624.915 52.280 631.200 52.420 ;
        RECT 624.915 52.235 625.205 52.280 ;
        RECT 630.880 52.220 631.200 52.280 ;
        RECT 393.520 52.080 393.840 52.140 ;
        RECT 359.480 51.940 363.850 52.080 ;
        RECT 364.170 51.940 371.670 52.080 ;
        RECT 371.990 51.940 393.840 52.080 ;
        RECT 334.180 51.880 334.500 51.940 ;
        RECT 359.480 51.880 359.800 51.940 ;
        RECT 308.880 51.740 309.200 51.800 ;
        RECT 312.100 51.740 312.420 51.800 ;
        RECT 318.080 51.740 318.400 51.800 ;
        RECT 297.010 51.600 309.200 51.740 ;
        RECT 311.905 51.600 312.420 51.740 ;
        RECT 317.885 51.600 318.400 51.740 ;
        RECT 287.720 51.540 288.040 51.600 ;
        RECT 296.015 51.555 296.305 51.600 ;
        RECT 308.880 51.540 309.200 51.600 ;
        RECT 312.100 51.540 312.420 51.600 ;
        RECT 318.080 51.540 318.400 51.600 ;
        RECT 318.540 51.740 318.860 51.800 ;
        RECT 324.535 51.740 324.825 51.785 ;
        RECT 318.540 51.600 324.825 51.740 ;
        RECT 318.540 51.540 318.860 51.600 ;
        RECT 324.535 51.555 324.825 51.600 ;
        RECT 327.280 51.740 327.600 51.800 ;
        RECT 328.200 51.740 328.520 51.800 ;
        RECT 327.280 51.600 328.520 51.740 ;
        RECT 327.280 51.540 327.600 51.600 ;
        RECT 328.200 51.540 328.520 51.600 ;
        RECT 330.040 51.740 330.360 51.800 ;
        RECT 332.800 51.740 333.120 51.800 ;
        RECT 330.040 51.600 333.120 51.740 ;
        RECT 330.040 51.540 330.360 51.600 ;
        RECT 332.800 51.540 333.120 51.600 ;
        RECT 336.020 51.740 336.340 51.800 ;
        RECT 354.880 51.740 355.200 51.800 ;
        RECT 336.020 51.600 355.200 51.740 ;
        RECT 363.710 51.740 363.850 51.940 ;
        RECT 370.995 51.740 371.285 51.785 ;
        RECT 363.710 51.600 371.285 51.740 ;
        RECT 371.530 51.740 371.670 51.940 ;
        RECT 393.520 51.880 393.840 51.940 ;
        RECT 385.700 51.740 386.020 51.800 ;
        RECT 371.530 51.600 386.020 51.740 ;
        RECT 336.020 51.540 336.340 51.600 ;
        RECT 354.880 51.540 355.200 51.600 ;
        RECT 370.995 51.555 371.285 51.600 ;
        RECT 385.700 51.540 386.020 51.600 ;
        RECT 42.470 50.920 631.270 51.400 ;
        RECT 56.800 50.720 57.120 50.780 ;
        RECT 72.440 50.720 72.760 50.780 ;
        RECT 56.800 50.580 72.760 50.720 ;
        RECT 56.800 50.520 57.120 50.580 ;
        RECT 72.440 50.520 72.760 50.580 ;
        RECT 73.375 50.720 73.665 50.765 ;
        RECT 98.660 50.720 98.980 50.780 ;
        RECT 73.375 50.580 98.980 50.720 ;
        RECT 73.375 50.535 73.665 50.580 ;
        RECT 98.660 50.520 98.980 50.580 ;
        RECT 100.500 50.720 100.820 50.780 ;
        RECT 133.160 50.720 133.480 50.780 ;
        RECT 133.635 50.720 133.925 50.765 ;
        RECT 100.500 50.580 113.150 50.720 ;
        RECT 100.500 50.520 100.820 50.580 ;
        RECT 60.020 50.380 60.340 50.440 ;
        RECT 86.700 50.380 87.020 50.440 ;
        RECT 60.020 50.240 87.020 50.380 ;
        RECT 60.020 50.180 60.340 50.240 ;
        RECT 86.700 50.180 87.020 50.240 ;
        RECT 92.240 50.380 92.530 50.425 ;
        RECT 93.640 50.380 93.930 50.425 ;
        RECT 95.480 50.380 95.770 50.425 ;
        RECT 106.020 50.380 106.340 50.440 ;
        RECT 92.240 50.240 95.770 50.380 ;
        RECT 92.240 50.195 92.530 50.240 ;
        RECT 93.640 50.195 93.930 50.240 ;
        RECT 95.480 50.195 95.770 50.240 ;
        RECT 95.990 50.240 106.340 50.380 ;
        RECT 72.915 49.855 73.205 50.085 ;
        RECT 77.960 50.040 78.280 50.100 ;
        RECT 78.880 50.040 79.200 50.100 ;
        RECT 80.720 50.040 81.040 50.100 ;
        RECT 77.960 49.900 78.475 50.040 ;
        RECT 78.880 49.900 79.395 50.040 ;
        RECT 80.525 49.900 81.040 50.040 ;
        RECT 61.860 49.700 62.180 49.760 ;
        RECT 72.990 49.700 73.130 49.855 ;
        RECT 77.960 49.840 78.280 49.900 ;
        RECT 78.880 49.840 79.200 49.900 ;
        RECT 80.720 49.840 81.040 49.900 ;
        RECT 85.795 50.040 86.085 50.085 ;
        RECT 91.760 50.040 92.080 50.100 ;
        RECT 85.795 49.900 92.080 50.040 ;
        RECT 85.795 49.855 86.085 49.900 ;
        RECT 91.760 49.840 92.080 49.900 ;
        RECT 92.695 50.040 92.985 50.085 ;
        RECT 95.990 50.040 96.130 50.240 ;
        RECT 106.020 50.180 106.340 50.240 ;
        RECT 92.695 49.900 96.130 50.040 ;
        RECT 99.580 50.040 99.900 50.100 ;
        RECT 105.115 50.040 105.405 50.085 ;
        RECT 99.580 49.900 105.405 50.040 ;
        RECT 92.695 49.855 92.985 49.900 ;
        RECT 99.580 49.840 99.900 49.900 ;
        RECT 105.115 49.855 105.405 49.900 ;
        RECT 107.875 49.855 108.165 50.085 ;
        RECT 108.795 50.040 109.085 50.085 ;
        RECT 112.000 50.040 112.320 50.100 ;
        RECT 108.795 49.900 112.320 50.040 ;
        RECT 113.010 50.040 113.150 50.580 ;
        RECT 133.160 50.580 133.925 50.720 ;
        RECT 133.160 50.520 133.480 50.580 ;
        RECT 133.635 50.535 133.925 50.580 ;
        RECT 157.080 50.720 157.400 50.780 ;
        RECT 162.600 50.720 162.920 50.780 ;
        RECT 194.800 50.720 195.120 50.780 ;
        RECT 213.660 50.720 213.980 50.780 ;
        RECT 249.540 50.720 249.860 50.780 ;
        RECT 157.080 50.580 162.920 50.720 ;
        RECT 157.080 50.520 157.400 50.580 ;
        RECT 162.600 50.520 162.920 50.580 ;
        RECT 163.150 50.580 195.120 50.720 ;
        RECT 114.320 50.380 114.610 50.425 ;
        RECT 115.720 50.380 116.010 50.425 ;
        RECT 117.560 50.380 117.850 50.425 ;
        RECT 114.320 50.240 117.850 50.380 ;
        RECT 114.320 50.195 114.610 50.240 ;
        RECT 115.720 50.195 116.010 50.240 ;
        RECT 117.560 50.195 117.850 50.240 ;
        RECT 126.740 50.380 127.030 50.425 ;
        RECT 128.140 50.380 128.430 50.425 ;
        RECT 129.980 50.380 130.270 50.425 ;
        RECT 126.740 50.240 130.270 50.380 ;
        RECT 126.740 50.195 127.030 50.240 ;
        RECT 128.140 50.195 128.430 50.240 ;
        RECT 129.980 50.195 130.270 50.240 ;
        RECT 130.860 50.380 131.180 50.440 ;
        RECT 141.900 50.380 142.220 50.440 ;
        RECT 130.860 50.240 142.220 50.380 ;
        RECT 130.860 50.180 131.180 50.240 ;
        RECT 141.900 50.180 142.220 50.240 ;
        RECT 142.380 50.380 142.670 50.425 ;
        RECT 143.780 50.380 144.070 50.425 ;
        RECT 145.620 50.380 145.910 50.425 ;
        RECT 148.800 50.380 149.120 50.440 ;
        RECT 142.380 50.240 145.910 50.380 ;
        RECT 142.380 50.195 142.670 50.240 ;
        RECT 143.780 50.195 144.070 50.240 ;
        RECT 145.620 50.195 145.910 50.240 ;
        RECT 146.130 50.240 149.120 50.380 ;
        RECT 113.395 50.040 113.685 50.085 ;
        RECT 113.010 49.900 113.685 50.040 ;
        RECT 108.795 49.855 109.085 49.900 ;
        RECT 89.920 49.700 90.240 49.760 ;
        RECT 91.300 49.700 91.620 49.760 ;
        RECT 61.860 49.560 90.240 49.700 ;
        RECT 91.105 49.560 91.620 49.700 ;
        RECT 61.860 49.500 62.180 49.560 ;
        RECT 89.920 49.500 90.240 49.560 ;
        RECT 91.300 49.500 91.620 49.560 ;
        RECT 106.020 49.700 106.340 49.760 ;
        RECT 107.950 49.700 108.090 49.855 ;
        RECT 112.000 49.840 112.320 49.900 ;
        RECT 113.395 49.855 113.685 49.900 ;
        RECT 114.775 50.040 115.065 50.085 ;
        RECT 120.280 50.040 120.600 50.100 ;
        RECT 114.775 49.900 120.600 50.040 ;
        RECT 114.775 49.855 115.065 49.900 ;
        RECT 112.460 49.700 112.780 49.760 ;
        RECT 106.020 49.560 112.780 49.700 ;
        RECT 113.470 49.700 113.610 49.855 ;
        RECT 120.280 49.840 120.600 49.900 ;
        RECT 126.260 49.840 126.580 50.100 ;
        RECT 127.195 50.040 127.485 50.085 ;
        RECT 133.620 50.040 133.940 50.100 ;
        RECT 127.195 49.900 133.940 50.040 ;
        RECT 127.195 49.855 127.485 49.900 ;
        RECT 133.620 49.840 133.940 49.900 ;
        RECT 139.600 50.040 139.920 50.100 ;
        RECT 141.455 50.040 141.745 50.085 ;
        RECT 139.600 49.900 141.745 50.040 ;
        RECT 139.600 49.840 139.920 49.900 ;
        RECT 141.455 49.855 141.745 49.900 ;
        RECT 142.835 50.040 143.125 50.085 ;
        RECT 146.130 50.040 146.270 50.240 ;
        RECT 148.800 50.180 149.120 50.240 ;
        RECT 154.800 50.380 155.090 50.425 ;
        RECT 156.200 50.380 156.490 50.425 ;
        RECT 158.040 50.380 158.330 50.425 ;
        RECT 154.800 50.240 158.330 50.380 ;
        RECT 154.800 50.195 155.090 50.240 ;
        RECT 156.200 50.195 156.490 50.240 ;
        RECT 158.040 50.195 158.330 50.240 ;
        RECT 162.140 50.380 162.460 50.440 ;
        RECT 163.150 50.380 163.290 50.580 ;
        RECT 194.800 50.520 195.120 50.580 ;
        RECT 195.350 50.580 202.850 50.720 ;
        RECT 162.140 50.240 163.290 50.380 ;
        RECT 170.440 50.380 170.730 50.425 ;
        RECT 171.840 50.380 172.130 50.425 ;
        RECT 173.680 50.380 173.970 50.425 ;
        RECT 170.440 50.240 173.970 50.380 ;
        RECT 162.140 50.180 162.460 50.240 ;
        RECT 170.440 50.195 170.730 50.240 ;
        RECT 171.840 50.195 172.130 50.240 ;
        RECT 173.680 50.195 173.970 50.240 ;
        RECT 182.860 50.380 183.150 50.425 ;
        RECT 184.260 50.380 184.550 50.425 ;
        RECT 186.100 50.380 186.390 50.425 ;
        RECT 182.860 50.240 186.390 50.380 ;
        RECT 182.860 50.195 183.150 50.240 ;
        RECT 184.260 50.195 184.550 50.240 ;
        RECT 186.100 50.195 186.390 50.240 ;
        RECT 191.580 50.380 191.900 50.440 ;
        RECT 195.350 50.380 195.490 50.580 ;
        RECT 191.580 50.240 195.490 50.380 ;
        RECT 198.500 50.380 198.790 50.425 ;
        RECT 199.900 50.380 200.190 50.425 ;
        RECT 201.740 50.380 202.030 50.425 ;
        RECT 198.500 50.240 202.030 50.380 ;
        RECT 202.710 50.380 202.850 50.580 ;
        RECT 213.660 50.580 249.860 50.720 ;
        RECT 213.660 50.520 213.980 50.580 ;
        RECT 249.540 50.520 249.860 50.580 ;
        RECT 250.000 50.720 250.320 50.780 ;
        RECT 256.900 50.720 257.220 50.780 ;
        RECT 259.660 50.720 259.980 50.780 ;
        RECT 250.000 50.580 257.220 50.720 ;
        RECT 259.465 50.580 259.980 50.720 ;
        RECT 250.000 50.520 250.320 50.580 ;
        RECT 256.900 50.520 257.220 50.580 ;
        RECT 259.660 50.520 259.980 50.580 ;
        RECT 272.540 50.720 272.860 50.780 ;
        RECT 282.660 50.720 282.980 50.780 ;
        RECT 291.860 50.720 292.180 50.780 ;
        RECT 272.540 50.580 282.980 50.720 ;
        RECT 272.540 50.520 272.860 50.580 ;
        RECT 282.660 50.520 282.980 50.580 ;
        RECT 291.490 50.580 292.180 50.720 ;
        RECT 230.680 50.380 231.000 50.440 ;
        RECT 238.960 50.380 239.280 50.440 ;
        RECT 257.820 50.380 258.140 50.440 ;
        RECT 258.740 50.380 259.060 50.440 ;
        RECT 275.760 50.380 276.080 50.440 ;
        RECT 291.490 50.380 291.630 50.580 ;
        RECT 291.860 50.520 292.180 50.580 ;
        RECT 292.320 50.720 292.640 50.780 ;
        RECT 314.875 50.720 315.165 50.765 ;
        RECT 318.080 50.720 318.400 50.780 ;
        RECT 331.880 50.720 332.200 50.780 ;
        RECT 347.980 50.720 348.300 50.780 ;
        RECT 349.375 50.720 349.665 50.765 ;
        RECT 354.880 50.720 355.200 50.780 ;
        RECT 374.660 50.720 374.980 50.780 ;
        RECT 292.320 50.580 315.165 50.720 ;
        RECT 292.320 50.520 292.640 50.580 ;
        RECT 314.875 50.535 315.165 50.580 ;
        RECT 317.250 50.580 332.200 50.720 ;
        RECT 202.710 50.240 225.390 50.380 ;
        RECT 230.485 50.240 231.000 50.380 ;
        RECT 191.580 50.180 191.900 50.240 ;
        RECT 198.500 50.195 198.790 50.240 ;
        RECT 199.900 50.195 200.190 50.240 ;
        RECT 201.740 50.195 202.030 50.240 ;
        RECT 142.835 49.900 146.270 50.040 ;
        RECT 147.880 50.040 148.200 50.100 ;
        RECT 155.240 50.040 155.560 50.100 ;
        RECT 147.880 49.900 154.550 50.040 ;
        RECT 155.045 49.900 155.560 50.040 ;
        RECT 142.835 49.855 143.125 49.900 ;
        RECT 147.880 49.840 148.200 49.900 ;
        RECT 125.800 49.700 126.120 49.760 ;
        RECT 113.470 49.560 126.120 49.700 ;
        RECT 126.350 49.700 126.490 49.840 ;
        RECT 130.400 49.700 130.720 49.760 ;
        RECT 134.540 49.700 134.860 49.760 ;
        RECT 153.860 49.700 154.180 49.760 ;
        RECT 126.350 49.560 134.860 49.700 ;
        RECT 153.665 49.560 154.180 49.700 ;
        RECT 154.410 49.700 154.550 49.900 ;
        RECT 155.240 49.840 155.560 49.900 ;
        RECT 163.060 50.040 163.380 50.100 ;
        RECT 169.515 50.040 169.805 50.085 ;
        RECT 170.880 50.040 171.200 50.100 ;
        RECT 181.920 50.040 182.240 50.100 ;
        RECT 183.315 50.040 183.605 50.085 ;
        RECT 192.040 50.040 192.360 50.100 ;
        RECT 163.060 49.900 169.805 50.040 ;
        RECT 170.685 49.900 171.200 50.040 ;
        RECT 163.060 49.840 163.380 49.900 ;
        RECT 169.515 49.855 169.805 49.900 ;
        RECT 169.590 49.700 169.730 49.855 ;
        RECT 170.880 49.840 171.200 49.900 ;
        RECT 171.430 49.900 182.435 50.040 ;
        RECT 183.315 49.900 192.360 50.040 ;
        RECT 171.430 49.700 171.570 49.900 ;
        RECT 181.920 49.840 182.240 49.900 ;
        RECT 183.315 49.855 183.605 49.900 ;
        RECT 192.040 49.840 192.360 49.900 ;
        RECT 194.340 50.040 194.660 50.100 ;
        RECT 195.275 50.040 195.565 50.085 ;
        RECT 194.340 49.900 195.565 50.040 ;
        RECT 194.340 49.840 194.660 49.900 ;
        RECT 195.275 49.855 195.565 49.900 ;
        RECT 198.955 50.040 199.245 50.085 ;
        RECT 205.380 50.040 205.700 50.100 ;
        RECT 198.955 49.900 205.700 50.040 ;
        RECT 198.955 49.855 199.245 49.900 ;
        RECT 205.380 49.840 205.700 49.900 ;
        RECT 210.915 50.040 211.205 50.085 ;
        RECT 213.200 50.040 213.520 50.100 ;
        RECT 213.675 50.040 213.965 50.085 ;
        RECT 214.580 50.040 214.900 50.100 ;
        RECT 210.915 49.900 213.965 50.040 ;
        RECT 214.385 49.900 214.900 50.040 ;
        RECT 210.915 49.855 211.205 49.900 ;
        RECT 213.200 49.840 213.520 49.900 ;
        RECT 213.675 49.855 213.965 49.900 ;
        RECT 214.580 49.840 214.900 49.900 ;
        RECT 219.640 50.040 219.960 50.100 ;
        RECT 224.700 50.040 225.020 50.100 ;
        RECT 219.640 49.900 225.020 50.040 ;
        RECT 219.640 49.840 219.960 49.900 ;
        RECT 224.700 49.840 225.020 49.900 ;
        RECT 154.410 49.560 161.450 49.700 ;
        RECT 169.590 49.560 171.570 49.700 ;
        RECT 175.940 49.700 176.260 49.760 ;
        RECT 191.120 49.700 191.440 49.760 ;
        RECT 197.560 49.700 197.880 49.760 ;
        RECT 210.440 49.700 210.760 49.760 ;
        RECT 175.940 49.560 191.440 49.700 ;
        RECT 106.020 49.500 106.340 49.560 ;
        RECT 112.460 49.500 112.780 49.560 ;
        RECT 125.800 49.500 126.120 49.560 ;
        RECT 130.400 49.500 130.720 49.560 ;
        RECT 134.540 49.500 134.860 49.560 ;
        RECT 153.860 49.500 154.180 49.560 ;
        RECT 66.460 49.360 66.780 49.420 ;
        RECT 90.840 49.360 91.160 49.420 ;
        RECT 66.460 49.220 91.160 49.360 ;
        RECT 66.460 49.160 66.780 49.220 ;
        RECT 90.840 49.160 91.160 49.220 ;
        RECT 91.780 49.360 92.070 49.405 ;
        RECT 94.100 49.360 94.390 49.405 ;
        RECT 95.480 49.360 95.770 49.405 ;
        RECT 91.780 49.220 95.770 49.360 ;
        RECT 91.780 49.175 92.070 49.220 ;
        RECT 94.100 49.175 94.390 49.220 ;
        RECT 95.480 49.175 95.770 49.220 ;
        RECT 113.860 49.360 114.150 49.405 ;
        RECT 116.180 49.360 116.470 49.405 ;
        RECT 117.560 49.360 117.850 49.405 ;
        RECT 113.860 49.220 117.850 49.360 ;
        RECT 113.860 49.175 114.150 49.220 ;
        RECT 116.180 49.175 116.470 49.220 ;
        RECT 117.560 49.175 117.850 49.220 ;
        RECT 126.280 49.360 126.570 49.405 ;
        RECT 128.600 49.360 128.890 49.405 ;
        RECT 129.980 49.360 130.270 49.405 ;
        RECT 126.280 49.220 130.270 49.360 ;
        RECT 126.280 49.175 126.570 49.220 ;
        RECT 128.600 49.175 128.890 49.220 ;
        RECT 129.980 49.175 130.270 49.220 ;
        RECT 141.920 49.360 142.210 49.405 ;
        RECT 144.240 49.360 144.530 49.405 ;
        RECT 145.620 49.360 145.910 49.405 ;
        RECT 141.920 49.220 145.910 49.360 ;
        RECT 141.920 49.175 142.210 49.220 ;
        RECT 144.240 49.175 144.530 49.220 ;
        RECT 145.620 49.175 145.910 49.220 ;
        RECT 154.340 49.360 154.630 49.405 ;
        RECT 156.660 49.360 156.950 49.405 ;
        RECT 158.040 49.360 158.330 49.405 ;
        RECT 154.340 49.220 158.330 49.360 ;
        RECT 154.340 49.175 154.630 49.220 ;
        RECT 156.660 49.175 156.950 49.220 ;
        RECT 158.040 49.175 158.330 49.220 ;
        RECT 70.140 49.020 70.460 49.080 ;
        RECT 86.240 49.020 86.560 49.080 ;
        RECT 70.140 48.880 86.560 49.020 ;
        RECT 70.140 48.820 70.460 48.880 ;
        RECT 86.240 48.820 86.560 48.880 ;
        RECT 86.715 49.020 87.005 49.065 ;
        RECT 87.160 49.020 87.480 49.080 ;
        RECT 86.715 48.880 87.480 49.020 ;
        RECT 86.715 48.835 87.005 48.880 ;
        RECT 87.160 48.820 87.480 48.880 ;
        RECT 96.820 49.020 97.140 49.080 ;
        RECT 99.135 49.020 99.425 49.065 ;
        RECT 96.820 48.880 99.425 49.020 ;
        RECT 96.820 48.820 97.140 48.880 ;
        RECT 99.135 48.835 99.425 48.880 ;
        RECT 108.780 49.020 109.100 49.080 ;
        RECT 120.295 49.020 120.585 49.065 ;
        RECT 108.780 48.880 120.585 49.020 ;
        RECT 108.780 48.820 109.100 48.880 ;
        RECT 120.295 48.835 120.585 48.880 ;
        RECT 150.640 49.020 150.960 49.080 ;
        RECT 160.775 49.020 161.065 49.065 ;
        RECT 150.640 48.880 161.065 49.020 ;
        RECT 161.310 49.020 161.450 49.560 ;
        RECT 175.940 49.500 176.260 49.560 ;
        RECT 191.120 49.500 191.440 49.560 ;
        RECT 196.730 49.560 197.880 49.700 ;
        RECT 210.245 49.560 210.760 49.700 ;
        RECT 169.980 49.360 170.270 49.405 ;
        RECT 172.300 49.360 172.590 49.405 ;
        RECT 173.680 49.360 173.970 49.405 ;
        RECT 169.980 49.220 173.970 49.360 ;
        RECT 169.980 49.175 170.270 49.220 ;
        RECT 172.300 49.175 172.590 49.220 ;
        RECT 173.680 49.175 173.970 49.220 ;
        RECT 182.400 49.360 182.690 49.405 ;
        RECT 184.720 49.360 185.010 49.405 ;
        RECT 186.100 49.360 186.390 49.405 ;
        RECT 193.420 49.360 193.740 49.420 ;
        RECT 194.355 49.360 194.645 49.405 ;
        RECT 182.400 49.220 186.390 49.360 ;
        RECT 182.400 49.175 182.690 49.220 ;
        RECT 184.720 49.175 185.010 49.220 ;
        RECT 186.100 49.175 186.390 49.220 ;
        RECT 187.070 49.220 194.645 49.360 ;
        RECT 176.415 49.020 176.705 49.065 ;
        RECT 161.310 48.880 176.705 49.020 ;
        RECT 150.640 48.820 150.960 48.880 ;
        RECT 160.775 48.835 161.065 48.880 ;
        RECT 176.415 48.835 176.705 48.880 ;
        RECT 185.140 49.020 185.460 49.080 ;
        RECT 187.070 49.020 187.210 49.220 ;
        RECT 193.420 49.160 193.740 49.220 ;
        RECT 194.355 49.175 194.645 49.220 ;
        RECT 188.820 49.020 189.140 49.080 ;
        RECT 185.140 48.880 187.210 49.020 ;
        RECT 188.625 48.880 189.140 49.020 ;
        RECT 194.430 49.020 194.570 49.175 ;
        RECT 196.730 49.020 196.870 49.560 ;
        RECT 197.560 49.500 197.880 49.560 ;
        RECT 210.440 49.500 210.760 49.560 ;
        RECT 212.300 49.700 212.590 49.745 ;
        RECT 215.080 49.700 215.370 49.745 ;
        RECT 212.300 49.560 215.370 49.700 ;
        RECT 212.300 49.515 212.590 49.560 ;
        RECT 215.080 49.515 215.370 49.560 ;
        RECT 198.040 49.360 198.330 49.405 ;
        RECT 200.360 49.360 200.650 49.405 ;
        RECT 201.740 49.360 202.030 49.405 ;
        RECT 198.040 49.220 202.030 49.360 ;
        RECT 198.040 49.175 198.330 49.220 ;
        RECT 200.360 49.175 200.650 49.220 ;
        RECT 201.740 49.175 202.030 49.220 ;
        RECT 202.620 49.360 202.940 49.420 ;
        RECT 223.320 49.360 223.640 49.420 ;
        RECT 202.620 49.220 223.640 49.360 ;
        RECT 225.250 49.360 225.390 50.240 ;
        RECT 230.680 50.180 231.000 50.240 ;
        RECT 231.230 50.240 239.280 50.380 ;
        RECT 228.840 50.040 229.160 50.100 ;
        RECT 231.230 50.085 231.370 50.240 ;
        RECT 238.960 50.180 239.280 50.240 ;
        RECT 254.690 50.240 257.590 50.380 ;
        RECT 230.235 50.040 230.525 50.085 ;
        RECT 228.840 49.900 230.525 50.040 ;
        RECT 228.840 49.840 229.160 49.900 ;
        RECT 230.235 49.855 230.525 49.900 ;
        RECT 231.155 49.855 231.445 50.085 ;
        RECT 238.515 50.040 238.805 50.085 ;
        RECT 241.260 50.040 241.580 50.100 ;
        RECT 242.180 50.040 242.500 50.100 ;
        RECT 238.515 49.900 241.580 50.040 ;
        RECT 241.985 49.900 242.500 50.040 ;
        RECT 238.515 49.855 238.805 49.900 ;
        RECT 241.260 49.840 241.580 49.900 ;
        RECT 242.180 49.840 242.500 49.900 ;
        RECT 252.760 50.040 253.080 50.100 ;
        RECT 254.690 50.085 254.830 50.240 ;
        RECT 253.695 50.040 253.985 50.085 ;
        RECT 252.760 49.900 253.985 50.040 ;
        RECT 252.760 49.840 253.080 49.900 ;
        RECT 253.695 49.855 253.985 49.900 ;
        RECT 254.615 49.855 254.905 50.085 ;
        RECT 256.900 50.040 257.220 50.100 ;
        RECT 257.450 50.085 257.590 50.240 ;
        RECT 257.820 50.240 259.060 50.380 ;
        RECT 257.820 50.180 258.140 50.240 ;
        RECT 258.740 50.180 259.060 50.240 ;
        RECT 271.250 50.240 274.150 50.380 ;
        RECT 256.705 49.900 257.220 50.040 ;
        RECT 256.900 49.840 257.220 49.900 ;
        RECT 257.375 50.040 257.665 50.085 ;
        RECT 260.580 50.040 260.900 50.100 ;
        RECT 257.375 49.900 260.900 50.040 ;
        RECT 257.375 49.855 257.665 49.900 ;
        RECT 260.580 49.840 260.900 49.900 ;
        RECT 264.735 50.040 265.025 50.085 ;
        RECT 265.640 50.040 265.960 50.100 ;
        RECT 271.250 50.085 271.390 50.240 ;
        RECT 264.735 49.900 265.960 50.040 ;
        RECT 264.735 49.855 265.025 49.900 ;
        RECT 265.640 49.840 265.960 49.900 ;
        RECT 271.175 49.855 271.465 50.085 ;
        RECT 272.080 50.040 272.400 50.100 ;
        RECT 274.010 50.085 274.150 50.240 ;
        RECT 275.760 50.240 291.630 50.380 ;
        RECT 295.080 50.380 295.400 50.440 ;
        RECT 296.015 50.380 296.305 50.425 ;
        RECT 295.080 50.240 296.305 50.380 ;
        RECT 275.760 50.180 276.080 50.240 ;
        RECT 273.475 50.040 273.765 50.085 ;
        RECT 272.080 49.900 273.765 50.040 ;
        RECT 272.080 49.840 272.400 49.900 ;
        RECT 273.475 49.855 273.765 49.900 ;
        RECT 273.935 50.040 274.225 50.085 ;
        RECT 280.360 50.040 280.680 50.100 ;
        RECT 282.200 50.040 282.520 50.100 ;
        RECT 283.120 50.040 283.440 50.100 ;
        RECT 284.130 50.085 284.270 50.240 ;
        RECT 295.080 50.180 295.400 50.240 ;
        RECT 296.015 50.195 296.305 50.240 ;
        RECT 273.935 49.900 282.520 50.040 ;
        RECT 282.925 49.900 283.440 50.040 ;
        RECT 273.935 49.855 274.225 49.900 ;
        RECT 280.360 49.840 280.680 49.900 ;
        RECT 282.200 49.840 282.520 49.900 ;
        RECT 283.120 49.840 283.440 49.900 ;
        RECT 284.055 49.855 284.345 50.085 ;
        RECT 284.960 50.040 285.280 50.100 ;
        RECT 287.720 50.040 288.040 50.100 ;
        RECT 284.960 49.900 288.040 50.040 ;
        RECT 284.960 49.840 285.280 49.900 ;
        RECT 287.720 49.840 288.040 49.900 ;
        RECT 290.495 50.040 290.785 50.085 ;
        RECT 292.780 50.040 293.100 50.100 ;
        RECT 293.255 50.040 293.545 50.085 ;
        RECT 294.160 50.040 294.480 50.100 ;
        RECT 290.495 49.900 293.545 50.040 ;
        RECT 293.965 49.900 294.480 50.040 ;
        RECT 290.495 49.855 290.785 49.900 ;
        RECT 292.780 49.840 293.100 49.900 ;
        RECT 293.255 49.855 293.545 49.900 ;
        RECT 294.160 49.840 294.480 49.900 ;
        RECT 299.220 50.040 299.540 50.100 ;
        RECT 300.615 50.040 300.905 50.085 ;
        RECT 303.360 50.040 303.680 50.100 ;
        RECT 317.250 50.085 317.390 50.580 ;
        RECT 318.080 50.520 318.400 50.580 ;
        RECT 331.880 50.520 332.200 50.580 ;
        RECT 344.390 50.580 347.290 50.720 ;
        RECT 319.000 50.380 319.320 50.440 ;
        RECT 325.440 50.380 325.760 50.440 ;
        RECT 319.000 50.240 325.760 50.380 ;
        RECT 319.000 50.180 319.320 50.240 ;
        RECT 325.440 50.180 325.760 50.240 ;
        RECT 325.900 50.380 326.220 50.440 ;
        RECT 328.200 50.380 328.520 50.440 ;
        RECT 329.595 50.380 329.885 50.425 ;
        RECT 325.900 50.240 327.970 50.380 ;
        RECT 325.900 50.180 326.220 50.240 ;
        RECT 299.220 49.900 300.905 50.040 ;
        RECT 303.165 49.900 303.680 50.040 ;
        RECT 299.220 49.840 299.540 49.900 ;
        RECT 300.615 49.855 300.905 49.900 ;
        RECT 303.360 49.840 303.680 49.900 ;
        RECT 315.795 49.855 316.085 50.085 ;
        RECT 317.175 49.855 317.465 50.085 ;
        RECT 324.075 50.040 324.365 50.085 ;
        RECT 326.820 50.040 327.140 50.100 ;
        RECT 327.830 50.085 327.970 50.240 ;
        RECT 328.200 50.240 329.885 50.380 ;
        RECT 328.200 50.180 328.520 50.240 ;
        RECT 329.595 50.195 329.885 50.240 ;
        RECT 324.075 49.900 327.335 50.040 ;
        RECT 324.075 49.855 324.365 49.900 ;
        RECT 227.000 49.700 227.320 49.760 ;
        RECT 234.820 49.700 235.140 49.760 ;
        RECT 227.000 49.560 235.140 49.700 ;
        RECT 227.000 49.500 227.320 49.560 ;
        RECT 234.820 49.500 235.140 49.560 ;
        RECT 238.055 49.515 238.345 49.745 ;
        RECT 239.900 49.700 240.190 49.745 ;
        RECT 242.680 49.700 242.970 49.745 ;
        RECT 239.900 49.560 242.970 49.700 ;
        RECT 239.900 49.515 240.190 49.560 ;
        RECT 242.680 49.515 242.970 49.560 ;
        RECT 256.000 49.700 256.290 49.745 ;
        RECT 258.780 49.700 259.070 49.745 ;
        RECT 256.000 49.560 259.070 49.700 ;
        RECT 256.000 49.515 256.290 49.560 ;
        RECT 258.780 49.515 259.070 49.560 ;
        RECT 259.660 49.700 259.980 49.760 ;
        RECT 270.240 49.700 270.560 49.760 ;
        RECT 259.660 49.560 266.330 49.700 ;
        RECT 270.045 49.560 270.560 49.700 ;
        RECT 235.740 49.360 236.060 49.420 ;
        RECT 225.250 49.220 236.060 49.360 ;
        RECT 238.130 49.360 238.270 49.515 ;
        RECT 259.660 49.500 259.980 49.560 ;
        RECT 246.320 49.360 246.640 49.420 ;
        RECT 265.655 49.360 265.945 49.405 ;
        RECT 238.130 49.220 244.710 49.360 ;
        RECT 202.620 49.160 202.940 49.220 ;
        RECT 223.320 49.160 223.640 49.220 ;
        RECT 235.740 49.160 236.060 49.220 ;
        RECT 197.100 49.020 197.420 49.080 ;
        RECT 194.430 48.880 197.420 49.020 ;
        RECT 185.140 48.820 185.460 48.880 ;
        RECT 188.820 48.820 189.140 48.880 ;
        RECT 197.100 48.820 197.420 48.880 ;
        RECT 197.560 49.020 197.880 49.080 ;
        RECT 202.160 49.020 202.480 49.080 ;
        RECT 197.560 48.880 202.480 49.020 ;
        RECT 197.560 48.820 197.880 48.880 ;
        RECT 202.160 48.820 202.480 48.880 ;
        RECT 203.080 49.020 203.400 49.080 ;
        RECT 204.475 49.020 204.765 49.065 ;
        RECT 203.080 48.880 204.765 49.020 ;
        RECT 203.080 48.820 203.400 48.880 ;
        RECT 204.475 48.835 204.765 48.880 ;
        RECT 205.380 49.020 205.700 49.080 ;
        RECT 215.975 49.020 216.265 49.065 ;
        RECT 205.380 48.880 216.265 49.020 ;
        RECT 205.380 48.820 205.700 48.880 ;
        RECT 215.975 48.835 216.265 48.880 ;
        RECT 217.800 49.020 218.120 49.080 ;
        RECT 228.380 49.020 228.700 49.080 ;
        RECT 217.800 48.880 228.700 49.020 ;
        RECT 217.800 48.820 218.120 48.880 ;
        RECT 228.380 48.820 228.700 48.880 ;
        RECT 232.075 49.020 232.365 49.065 ;
        RECT 241.720 49.020 242.040 49.080 ;
        RECT 232.075 48.880 242.040 49.020 ;
        RECT 232.075 48.835 232.365 48.880 ;
        RECT 241.720 48.820 242.040 48.880 ;
        RECT 243.100 49.020 243.420 49.080 ;
        RECT 243.575 49.020 243.865 49.065 ;
        RECT 243.100 48.880 243.865 49.020 ;
        RECT 244.570 49.020 244.710 49.220 ;
        RECT 246.320 49.220 265.945 49.360 ;
        RECT 266.190 49.360 266.330 49.560 ;
        RECT 270.240 49.500 270.560 49.560 ;
        RECT 272.560 49.700 272.850 49.745 ;
        RECT 275.340 49.700 275.630 49.745 ;
        RECT 272.560 49.560 275.630 49.700 ;
        RECT 272.560 49.515 272.850 49.560 ;
        RECT 275.340 49.515 275.630 49.560 ;
        RECT 276.220 49.700 276.540 49.760 ;
        RECT 284.515 49.700 284.805 49.745 ;
        RECT 276.220 49.560 284.805 49.700 ;
        RECT 276.220 49.500 276.540 49.560 ;
        RECT 284.515 49.515 284.805 49.560 ;
        RECT 290.035 49.515 290.325 49.745 ;
        RECT 291.880 49.700 292.170 49.745 ;
        RECT 294.660 49.700 294.950 49.745 ;
        RECT 291.880 49.560 294.950 49.700 ;
        RECT 291.880 49.515 292.170 49.560 ;
        RECT 294.660 49.515 294.950 49.560 ;
        RECT 296.460 49.700 296.780 49.760 ;
        RECT 302.915 49.700 303.205 49.745 ;
        RECT 296.460 49.560 303.205 49.700 ;
        RECT 287.720 49.360 288.040 49.420 ;
        RECT 266.190 49.220 288.040 49.360 ;
        RECT 290.110 49.360 290.250 49.515 ;
        RECT 296.460 49.500 296.780 49.560 ;
        RECT 302.915 49.515 303.205 49.560 ;
        RECT 304.280 49.700 304.600 49.760 ;
        RECT 310.720 49.700 311.040 49.760 ;
        RECT 304.280 49.560 311.040 49.700 ;
        RECT 304.280 49.500 304.600 49.560 ;
        RECT 310.720 49.500 311.040 49.560 ;
        RECT 295.080 49.360 295.400 49.420 ;
        RECT 290.110 49.220 295.400 49.360 ;
        RECT 246.320 49.160 246.640 49.220 ;
        RECT 265.655 49.175 265.945 49.220 ;
        RECT 287.720 49.160 288.040 49.220 ;
        RECT 295.080 49.160 295.400 49.220 ;
        RECT 259.660 49.020 259.980 49.080 ;
        RECT 244.570 48.880 259.980 49.020 ;
        RECT 243.100 48.820 243.420 48.880 ;
        RECT 243.575 48.835 243.865 48.880 ;
        RECT 259.660 48.820 259.980 48.880 ;
        RECT 270.240 49.020 270.560 49.080 ;
        RECT 274.380 49.020 274.700 49.080 ;
        RECT 270.240 48.880 274.700 49.020 ;
        RECT 270.240 48.820 270.560 48.880 ;
        RECT 274.380 48.820 274.700 48.880 ;
        RECT 276.220 49.020 276.540 49.080 ;
        RECT 283.120 49.020 283.440 49.080 ;
        RECT 290.480 49.020 290.800 49.080 ;
        RECT 276.220 48.880 276.735 49.020 ;
        RECT 283.120 48.880 290.800 49.020 ;
        RECT 276.220 48.820 276.540 48.880 ;
        RECT 283.120 48.820 283.440 48.880 ;
        RECT 290.480 48.820 290.800 48.880 ;
        RECT 292.320 49.020 292.640 49.080 ;
        RECT 314.860 49.020 315.180 49.080 ;
        RECT 292.320 48.880 315.180 49.020 ;
        RECT 315.870 49.020 316.010 49.855 ;
        RECT 326.820 49.840 327.140 49.900 ;
        RECT 327.755 49.855 328.045 50.085 ;
        RECT 331.420 50.040 331.740 50.100 ;
        RECT 336.020 50.040 336.340 50.100 ;
        RECT 331.420 49.900 336.340 50.040 ;
        RECT 331.420 49.840 331.740 49.900 ;
        RECT 336.020 49.840 336.340 49.900 ;
        RECT 337.400 50.040 337.720 50.100 ;
        RECT 344.390 50.085 344.530 50.580 ;
        RECT 345.220 50.380 345.540 50.440 ;
        RECT 345.220 50.240 346.830 50.380 ;
        RECT 345.220 50.180 345.540 50.240 ;
        RECT 346.690 50.085 346.830 50.240 ;
        RECT 347.150 50.085 347.290 50.580 ;
        RECT 347.980 50.580 349.665 50.720 ;
        RECT 354.685 50.580 355.200 50.720 ;
        RECT 347.980 50.520 348.300 50.580 ;
        RECT 349.375 50.535 349.665 50.580 ;
        RECT 354.880 50.520 355.200 50.580 ;
        RECT 367.390 50.580 374.980 50.720 ;
        RECT 347.520 50.380 347.840 50.440 ;
        RECT 359.020 50.380 359.340 50.440 ;
        RECT 367.390 50.380 367.530 50.580 ;
        RECT 374.660 50.520 374.980 50.580 ;
        RECT 375.135 50.720 375.425 50.765 ;
        RECT 376.040 50.720 376.360 50.780 ;
        RECT 375.135 50.580 376.360 50.720 ;
        RECT 375.135 50.535 375.425 50.580 ;
        RECT 376.040 50.520 376.360 50.580 ;
        RECT 382.020 50.720 382.340 50.780 ;
        RECT 394.900 50.720 395.220 50.780 ;
        RECT 382.020 50.580 395.220 50.720 ;
        RECT 382.020 50.520 382.340 50.580 ;
        RECT 394.900 50.520 395.220 50.580 ;
        RECT 382.480 50.380 382.800 50.440 ;
        RECT 347.520 50.240 356.950 50.380 ;
        RECT 347.520 50.180 347.840 50.240 ;
        RECT 337.875 50.040 338.165 50.085 ;
        RECT 337.400 49.900 338.165 50.040 ;
        RECT 337.400 49.840 337.720 49.900 ;
        RECT 337.875 49.855 338.165 49.900 ;
        RECT 344.315 49.855 344.605 50.085 ;
        RECT 346.645 49.855 346.935 50.085 ;
        RECT 347.075 50.040 347.365 50.085 ;
        RECT 353.040 50.040 353.360 50.100 ;
        RECT 356.810 50.085 356.950 50.240 ;
        RECT 359.020 50.240 367.530 50.380 ;
        RECT 367.850 50.240 382.800 50.380 ;
        RECT 359.020 50.180 359.340 50.240 ;
        RECT 347.075 49.900 353.730 50.040 ;
        RECT 347.075 49.855 347.365 49.900 ;
        RECT 353.040 49.840 353.360 49.900 ;
        RECT 323.615 49.515 323.905 49.745 ;
        RECT 325.460 49.700 325.750 49.745 ;
        RECT 328.240 49.700 328.530 49.745 ;
        RECT 325.460 49.560 328.530 49.700 ;
        RECT 325.460 49.515 325.750 49.560 ;
        RECT 328.240 49.515 328.530 49.560 ;
        RECT 343.380 49.700 343.700 49.760 ;
        RECT 345.700 49.700 345.990 49.745 ;
        RECT 348.480 49.700 348.770 49.745 ;
        RECT 343.380 49.560 343.895 49.700 ;
        RECT 345.700 49.560 348.770 49.700 ;
        RECT 323.690 49.360 323.830 49.515 ;
        RECT 343.380 49.500 343.700 49.560 ;
        RECT 345.700 49.515 345.990 49.560 ;
        RECT 348.480 49.515 348.770 49.560 ;
        RECT 344.300 49.360 344.620 49.420 ;
        RECT 353.040 49.360 353.360 49.420 ;
        RECT 323.690 49.220 339.470 49.360 ;
        RECT 327.280 49.020 327.600 49.080 ;
        RECT 315.870 48.880 327.600 49.020 ;
        RECT 339.330 49.020 339.470 49.220 ;
        RECT 344.300 49.220 353.360 49.360 ;
        RECT 353.590 49.360 353.730 49.900 ;
        RECT 355.815 49.855 356.105 50.085 ;
        RECT 356.735 49.855 357.025 50.085 ;
        RECT 367.315 50.040 367.605 50.085 ;
        RECT 367.850 50.040 367.990 50.240 ;
        RECT 382.480 50.180 382.800 50.240 ;
        RECT 382.940 50.380 383.260 50.440 ;
        RECT 391.220 50.380 391.540 50.440 ;
        RECT 382.940 50.240 391.540 50.380 ;
        RECT 382.940 50.180 383.260 50.240 ;
        RECT 391.220 50.180 391.540 50.240 ;
        RECT 367.315 49.900 367.990 50.040 ;
        RECT 368.680 50.085 369.000 50.100 ;
        RECT 367.315 49.855 367.605 49.900 ;
        RECT 368.680 49.855 369.215 50.085 ;
        RECT 374.675 49.855 374.965 50.085 ;
        RECT 375.120 50.040 375.440 50.100 ;
        RECT 376.055 50.040 376.345 50.085 ;
        RECT 400.880 50.040 401.200 50.100 ;
        RECT 375.120 49.900 376.345 50.040 ;
        RECT 355.890 49.700 356.030 49.855 ;
        RECT 368.680 49.840 369.000 49.855 ;
        RECT 360.400 49.700 360.720 49.760 ;
        RECT 368.235 49.700 368.525 49.745 ;
        RECT 355.890 49.560 360.720 49.700 ;
        RECT 360.400 49.500 360.720 49.560 ;
        RECT 360.950 49.560 368.525 49.700 ;
        RECT 374.750 49.700 374.890 49.855 ;
        RECT 375.120 49.840 375.440 49.900 ;
        RECT 376.055 49.855 376.345 49.900 ;
        RECT 377.050 49.900 401.200 50.040 ;
        RECT 377.050 49.700 377.190 49.900 ;
        RECT 400.880 49.840 401.200 49.900 ;
        RECT 374.750 49.560 377.190 49.700 ;
        RECT 360.950 49.360 361.090 49.560 ;
        RECT 368.235 49.515 368.525 49.560 ;
        RECT 353.590 49.220 361.090 49.360 ;
        RECT 366.840 49.360 367.160 49.420 ;
        RECT 387.555 49.360 387.845 49.405 ;
        RECT 366.840 49.220 387.845 49.360 ;
        RECT 344.300 49.160 344.620 49.220 ;
        RECT 353.040 49.160 353.360 49.220 ;
        RECT 366.840 49.160 367.160 49.220 ;
        RECT 387.555 49.175 387.845 49.220 ;
        RECT 342.920 49.020 343.240 49.080 ;
        RECT 339.330 48.880 343.240 49.020 ;
        RECT 292.320 48.820 292.640 48.880 ;
        RECT 314.860 48.820 315.180 48.880 ;
        RECT 327.280 48.820 327.600 48.880 ;
        RECT 342.920 48.820 343.240 48.880 ;
        RECT 350.280 49.020 350.600 49.080 ;
        RECT 357.640 49.020 357.960 49.080 ;
        RECT 350.280 48.880 357.960 49.020 ;
        RECT 350.280 48.820 350.600 48.880 ;
        RECT 357.640 48.820 357.960 48.880 ;
        RECT 359.480 49.020 359.800 49.080 ;
        RECT 382.495 49.020 382.785 49.065 ;
        RECT 359.480 48.880 382.785 49.020 ;
        RECT 359.480 48.820 359.800 48.880 ;
        RECT 382.495 48.835 382.785 48.880 ;
        RECT 392.140 49.020 392.460 49.080 ;
        RECT 394.915 49.020 395.205 49.065 ;
        RECT 392.140 48.880 395.205 49.020 ;
        RECT 392.140 48.820 392.460 48.880 ;
        RECT 394.915 48.835 395.205 48.880 ;
        RECT 395.820 49.020 396.140 49.080 ;
        RECT 399.975 49.020 400.265 49.065 ;
        RECT 395.820 48.880 400.265 49.020 ;
        RECT 395.820 48.820 396.140 48.880 ;
        RECT 399.975 48.835 400.265 48.880 ;
        RECT 403.180 49.020 403.500 49.080 ;
        RECT 405.035 49.020 405.325 49.065 ;
        RECT 414.220 49.020 414.540 49.080 ;
        RECT 428.940 49.020 429.260 49.080 ;
        RECT 436.300 49.020 436.620 49.080 ;
        RECT 403.180 48.880 405.325 49.020 ;
        RECT 414.025 48.880 414.540 49.020 ;
        RECT 428.745 48.880 429.260 49.020 ;
        RECT 436.105 48.880 436.620 49.020 ;
        RECT 403.180 48.820 403.500 48.880 ;
        RECT 405.035 48.835 405.325 48.880 ;
        RECT 414.220 48.820 414.540 48.880 ;
        RECT 428.940 48.820 429.260 48.880 ;
        RECT 436.300 48.820 436.620 48.880 ;
        RECT 447.340 49.020 447.660 49.080 ;
        RECT 451.035 49.020 451.325 49.065 ;
        RECT 458.380 49.020 458.700 49.080 ;
        RECT 469.420 49.020 469.740 49.080 ;
        RECT 480.460 49.020 480.780 49.080 ;
        RECT 487.820 49.020 488.140 49.080 ;
        RECT 513.580 49.020 513.900 49.080 ;
        RECT 520.940 49.020 521.260 49.080 ;
        RECT 535.660 49.020 535.980 49.080 ;
        RECT 543.020 49.020 543.340 49.080 ;
        RECT 554.060 49.020 554.380 49.080 ;
        RECT 564.640 49.020 564.960 49.080 ;
        RECT 572.000 49.020 572.320 49.080 ;
        RECT 597.760 49.020 598.080 49.080 ;
        RECT 619.840 49.020 620.160 49.080 ;
        RECT 447.340 48.880 451.325 49.020 ;
        RECT 458.185 48.880 458.700 49.020 ;
        RECT 469.225 48.880 469.740 49.020 ;
        RECT 480.265 48.880 480.780 49.020 ;
        RECT 487.625 48.880 488.140 49.020 ;
        RECT 513.385 48.880 513.900 49.020 ;
        RECT 520.745 48.880 521.260 49.020 ;
        RECT 535.465 48.880 535.980 49.020 ;
        RECT 542.825 48.880 543.340 49.020 ;
        RECT 553.865 48.880 554.380 49.020 ;
        RECT 564.445 48.880 564.960 49.020 ;
        RECT 571.805 48.880 572.320 49.020 ;
        RECT 597.565 48.880 598.080 49.020 ;
        RECT 619.645 48.880 620.160 49.020 ;
        RECT 447.340 48.820 447.660 48.880 ;
        RECT 451.035 48.835 451.325 48.880 ;
        RECT 458.380 48.820 458.700 48.880 ;
        RECT 469.420 48.820 469.740 48.880 ;
        RECT 480.460 48.820 480.780 48.880 ;
        RECT 487.820 48.820 488.140 48.880 ;
        RECT 513.580 48.820 513.900 48.880 ;
        RECT 520.940 48.820 521.260 48.880 ;
        RECT 535.660 48.820 535.980 48.880 ;
        RECT 543.020 48.820 543.340 48.880 ;
        RECT 554.060 48.820 554.380 48.880 ;
        RECT 564.640 48.820 564.960 48.880 ;
        RECT 572.000 48.820 572.320 48.880 ;
        RECT 597.760 48.820 598.080 48.880 ;
        RECT 619.840 48.820 620.160 48.880 ;
        RECT 624.915 49.020 625.205 49.065 ;
        RECT 627.200 49.020 627.520 49.080 ;
        RECT 624.915 48.880 627.520 49.020 ;
        RECT 624.915 48.835 625.205 48.880 ;
        RECT 627.200 48.820 627.520 48.880 ;
        RECT 42.470 48.200 631.270 48.680 ;
        RECT 83.940 48.000 84.260 48.060 ;
        RECT 99.120 48.000 99.440 48.060 ;
        RECT 83.940 47.860 99.440 48.000 ;
        RECT 83.940 47.800 84.260 47.860 ;
        RECT 99.120 47.800 99.440 47.860 ;
        RECT 106.940 48.000 107.260 48.060 ;
        RECT 146.500 48.000 146.820 48.060 ;
        RECT 149.720 48.000 150.040 48.060 ;
        RECT 106.940 47.860 146.820 48.000 ;
        RECT 149.525 47.860 150.040 48.000 ;
        RECT 106.940 47.800 107.260 47.860 ;
        RECT 146.500 47.800 146.820 47.860 ;
        RECT 149.720 47.800 150.040 47.860 ;
        RECT 153.400 48.000 153.720 48.060 ;
        RECT 176.860 48.000 177.180 48.060 ;
        RECT 153.400 47.860 177.180 48.000 ;
        RECT 153.400 47.800 153.720 47.860 ;
        RECT 176.860 47.800 177.180 47.860 ;
        RECT 184.680 48.000 185.000 48.060 ;
        RECT 212.755 48.000 213.045 48.045 ;
        RECT 213.660 48.000 213.980 48.060 ;
        RECT 184.680 47.860 213.980 48.000 ;
        RECT 184.680 47.800 185.000 47.860 ;
        RECT 212.755 47.815 213.045 47.860 ;
        RECT 213.660 47.800 213.980 47.860 ;
        RECT 219.640 48.000 219.960 48.060 ;
        RECT 223.780 48.000 224.100 48.060 ;
        RECT 219.640 47.860 224.100 48.000 ;
        RECT 219.640 47.800 219.960 47.860 ;
        RECT 223.780 47.800 224.100 47.860 ;
        RECT 224.700 48.000 225.020 48.060 ;
        RECT 230.680 48.000 231.000 48.060 ;
        RECT 224.700 47.860 231.000 48.000 ;
        RECT 224.700 47.800 225.020 47.860 ;
        RECT 230.680 47.800 231.000 47.860 ;
        RECT 232.075 48.000 232.365 48.045 ;
        RECT 233.900 48.000 234.220 48.060 ;
        RECT 232.075 47.860 234.220 48.000 ;
        RECT 232.075 47.815 232.365 47.860 ;
        RECT 233.900 47.800 234.220 47.860 ;
        RECT 234.360 48.000 234.680 48.060 ;
        RECT 240.340 48.000 240.660 48.060 ;
        RECT 246.780 48.000 247.100 48.060 ;
        RECT 234.360 47.860 240.660 48.000 ;
        RECT 234.360 47.800 234.680 47.860 ;
        RECT 240.340 47.800 240.660 47.860 ;
        RECT 242.270 47.860 247.100 48.000 ;
        RECT 55.420 47.660 55.740 47.720 ;
        RECT 91.760 47.660 92.080 47.720 ;
        RECT 105.560 47.660 105.880 47.720 ;
        RECT 119.360 47.660 119.680 47.720 ;
        RECT 120.280 47.660 120.600 47.720 ;
        RECT 55.420 47.520 91.070 47.660 ;
        RECT 55.420 47.460 55.740 47.520 ;
        RECT 42.080 47.320 42.400 47.380 ;
        RECT 77.515 47.320 77.805 47.365 ;
        RECT 42.080 47.180 77.805 47.320 ;
        RECT 42.080 47.120 42.400 47.180 ;
        RECT 77.515 47.135 77.805 47.180 ;
        RECT 78.420 47.320 78.740 47.380 ;
        RECT 89.000 47.320 89.320 47.380 ;
        RECT 78.420 47.180 89.320 47.320 ;
        RECT 78.420 47.120 78.740 47.180 ;
        RECT 89.000 47.120 89.320 47.180 ;
        RECT 43.460 46.980 43.780 47.040 ;
        RECT 72.455 46.980 72.745 47.025 ;
        RECT 43.460 46.840 72.745 46.980 ;
        RECT 43.460 46.780 43.780 46.840 ;
        RECT 72.455 46.795 72.745 46.840 ;
        RECT 77.975 46.795 78.265 47.025 ;
        RECT 85.335 46.980 85.625 47.025 ;
        RECT 90.380 46.980 90.700 47.040 ;
        RECT 90.930 47.025 91.070 47.520 ;
        RECT 91.760 47.520 105.880 47.660 ;
        RECT 91.760 47.460 92.080 47.520 ;
        RECT 105.560 47.460 105.880 47.520 ;
        RECT 113.930 47.520 119.680 47.660 ;
        RECT 120.085 47.520 120.600 47.660 ;
        RECT 91.300 47.320 91.620 47.380 ;
        RECT 94.535 47.320 94.825 47.365 ;
        RECT 113.930 47.320 114.070 47.520 ;
        RECT 119.360 47.460 119.680 47.520 ;
        RECT 120.280 47.460 120.600 47.520 ;
        RECT 125.800 47.660 126.120 47.720 ;
        RECT 128.120 47.660 128.410 47.705 ;
        RECT 130.440 47.660 130.730 47.705 ;
        RECT 131.820 47.660 132.110 47.705 ;
        RECT 134.540 47.660 134.860 47.720 ;
        RECT 147.420 47.660 147.740 47.720 ;
        RECT 125.800 47.520 127.870 47.660 ;
        RECT 125.800 47.460 126.120 47.520 ;
        RECT 114.760 47.320 115.080 47.380 ;
        RECT 117.980 47.320 118.300 47.380 ;
        RECT 91.300 47.180 93.830 47.320 ;
        RECT 91.300 47.120 91.620 47.180 ;
        RECT 85.335 46.840 90.700 46.980 ;
        RECT 85.335 46.795 85.625 46.840 ;
        RECT 48.060 46.640 48.380 46.700 ;
        RECT 63.700 46.640 64.020 46.700 ;
        RECT 78.050 46.640 78.190 46.795 ;
        RECT 90.380 46.780 90.700 46.840 ;
        RECT 90.855 46.795 91.145 47.025 ;
        RECT 93.140 46.980 93.460 47.040 ;
        RECT 92.945 46.840 93.460 46.980 ;
        RECT 93.690 46.980 93.830 47.180 ;
        RECT 94.535 47.180 114.070 47.320 ;
        RECT 114.565 47.180 115.080 47.320 ;
        RECT 94.535 47.135 94.825 47.180 ;
        RECT 114.760 47.120 115.080 47.180 ;
        RECT 115.770 47.180 118.300 47.320 ;
        RECT 103.275 46.980 103.565 47.025 ;
        RECT 106.020 46.980 106.340 47.040 ;
        RECT 93.690 46.840 103.565 46.980 ;
        RECT 105.825 46.840 106.340 46.980 ;
        RECT 93.140 46.780 93.460 46.840 ;
        RECT 103.275 46.795 103.565 46.840 ;
        RECT 106.020 46.780 106.340 46.840 ;
        RECT 111.555 46.795 111.845 47.025 ;
        RECT 112.460 46.980 112.780 47.040 ;
        RECT 113.855 46.980 114.145 47.025 ;
        RECT 115.770 46.980 115.910 47.180 ;
        RECT 117.980 47.120 118.300 47.180 ;
        RECT 118.440 47.320 118.760 47.380 ;
        RECT 127.730 47.365 127.870 47.520 ;
        RECT 128.120 47.520 132.110 47.660 ;
        RECT 134.345 47.520 134.860 47.660 ;
        RECT 128.120 47.475 128.410 47.520 ;
        RECT 130.440 47.475 130.730 47.520 ;
        RECT 131.820 47.475 132.110 47.520 ;
        RECT 134.540 47.460 134.860 47.520 ;
        RECT 144.750 47.520 147.740 47.660 ;
        RECT 120.755 47.320 121.045 47.365 ;
        RECT 118.440 47.180 121.045 47.320 ;
        RECT 118.440 47.120 118.760 47.180 ;
        RECT 120.755 47.135 121.045 47.180 ;
        RECT 127.690 47.135 127.980 47.365 ;
        RECT 128.560 47.320 128.880 47.380 ;
        RECT 129.035 47.320 129.325 47.365 ;
        RECT 136.840 47.320 137.160 47.380 ;
        RECT 128.560 47.180 129.325 47.320 ;
        RECT 128.560 47.120 128.880 47.180 ;
        RECT 129.035 47.135 129.325 47.180 ;
        RECT 129.570 47.180 137.160 47.320 ;
        RECT 112.460 46.840 115.910 46.980 ;
        RECT 119.360 47.025 119.680 47.040 ;
        RECT 48.060 46.500 64.020 46.640 ;
        RECT 48.060 46.440 48.380 46.500 ;
        RECT 63.700 46.440 64.020 46.500 ;
        RECT 64.250 46.500 78.190 46.640 ;
        RECT 80.275 46.640 80.565 46.685 ;
        RECT 84.860 46.640 85.180 46.700 ;
        RECT 80.275 46.500 85.180 46.640 ;
        RECT 40.700 46.300 41.020 46.360 ;
        RECT 64.250 46.300 64.390 46.500 ;
        RECT 80.275 46.455 80.565 46.500 ;
        RECT 84.860 46.440 85.180 46.500 ;
        RECT 102.340 46.640 102.660 46.700 ;
        RECT 111.630 46.640 111.770 46.795 ;
        RECT 112.460 46.780 112.780 46.840 ;
        RECT 113.855 46.795 114.145 46.840 ;
        RECT 119.360 46.795 119.940 47.025 ;
        RECT 122.595 46.980 122.885 47.025 ;
        RECT 129.570 46.980 129.710 47.180 ;
        RECT 136.840 47.120 137.160 47.180 ;
        RECT 122.595 46.840 129.710 46.980 ;
        RECT 143.740 46.980 144.060 47.040 ;
        RECT 144.750 47.025 144.890 47.520 ;
        RECT 147.420 47.460 147.740 47.520 ;
        RECT 155.720 47.660 156.010 47.705 ;
        RECT 158.040 47.660 158.330 47.705 ;
        RECT 159.420 47.660 159.710 47.705 ;
        RECT 155.720 47.520 159.710 47.660 ;
        RECT 155.720 47.475 156.010 47.520 ;
        RECT 158.040 47.475 158.330 47.520 ;
        RECT 159.420 47.475 159.710 47.520 ;
        RECT 167.200 47.660 167.520 47.720 ;
        RECT 169.520 47.660 169.810 47.705 ;
        RECT 171.840 47.660 172.130 47.705 ;
        RECT 173.220 47.660 173.510 47.705 ;
        RECT 167.200 47.520 169.270 47.660 ;
        RECT 167.200 47.460 167.520 47.520 ;
        RECT 146.060 47.320 146.350 47.365 ;
        RECT 148.840 47.320 149.130 47.365 ;
        RECT 146.060 47.180 149.130 47.320 ;
        RECT 146.060 47.135 146.350 47.180 ;
        RECT 148.840 47.135 149.130 47.180 ;
        RECT 153.860 47.320 154.180 47.380 ;
        RECT 155.255 47.320 155.545 47.365 ;
        RECT 153.860 47.180 155.545 47.320 ;
        RECT 169.130 47.320 169.270 47.520 ;
        RECT 169.520 47.520 173.510 47.660 ;
        RECT 169.520 47.475 169.810 47.520 ;
        RECT 171.840 47.475 172.130 47.520 ;
        RECT 173.220 47.475 173.510 47.520 ;
        RECT 185.160 47.660 185.450 47.705 ;
        RECT 187.480 47.660 187.770 47.705 ;
        RECT 188.860 47.660 189.150 47.705 ;
        RECT 185.160 47.520 189.150 47.660 ;
        RECT 185.160 47.475 185.450 47.520 ;
        RECT 187.480 47.475 187.770 47.520 ;
        RECT 188.860 47.475 189.150 47.520 ;
        RECT 189.740 47.660 190.060 47.720 ;
        RECT 191.595 47.660 191.885 47.705 ;
        RECT 189.740 47.520 191.885 47.660 ;
        RECT 189.740 47.460 190.060 47.520 ;
        RECT 191.595 47.475 191.885 47.520 ;
        RECT 197.580 47.660 197.870 47.705 ;
        RECT 199.900 47.660 200.190 47.705 ;
        RECT 201.280 47.660 201.570 47.705 ;
        RECT 197.580 47.520 201.570 47.660 ;
        RECT 197.580 47.475 197.870 47.520 ;
        RECT 199.900 47.475 200.190 47.520 ;
        RECT 201.280 47.475 201.570 47.520 ;
        RECT 214.595 47.660 214.885 47.705 ;
        RECT 217.800 47.660 218.120 47.720 ;
        RECT 219.180 47.660 219.500 47.720 ;
        RECT 226.540 47.660 226.860 47.720 ;
        RECT 214.595 47.520 218.120 47.660 ;
        RECT 218.745 47.520 226.860 47.660 ;
        RECT 214.595 47.475 214.885 47.520 ;
        RECT 217.800 47.460 218.120 47.520 ;
        RECT 219.180 47.460 219.500 47.520 ;
        RECT 226.540 47.460 226.860 47.520 ;
        RECT 228.380 47.660 228.700 47.720 ;
        RECT 238.960 47.660 239.280 47.720 ;
        RECT 242.270 47.660 242.410 47.860 ;
        RECT 246.780 47.800 247.100 47.860 ;
        RECT 247.240 48.000 247.560 48.060 ;
        RECT 252.775 48.000 253.065 48.045 ;
        RECT 268.400 48.000 268.720 48.060 ;
        RECT 276.220 48.000 276.540 48.060 ;
        RECT 247.240 47.860 253.065 48.000 ;
        RECT 268.205 47.860 268.720 48.000 ;
        RECT 247.240 47.800 247.560 47.860 ;
        RECT 252.775 47.815 253.065 47.860 ;
        RECT 268.400 47.800 268.720 47.860 ;
        RECT 271.250 47.860 276.540 48.000 ;
        RECT 228.380 47.520 239.280 47.660 ;
        RECT 228.380 47.460 228.700 47.520 ;
        RECT 238.960 47.460 239.280 47.520 ;
        RECT 239.510 47.520 242.410 47.660 ;
        RECT 242.640 47.660 242.960 47.720 ;
        RECT 251.165 47.660 251.455 47.705 ;
        RECT 242.640 47.520 251.455 47.660 ;
        RECT 170.405 47.320 170.695 47.365 ;
        RECT 169.130 47.180 170.695 47.320 ;
        RECT 153.860 47.120 154.180 47.180 ;
        RECT 155.255 47.135 155.545 47.180 ;
        RECT 170.405 47.135 170.695 47.180 ;
        RECT 170.880 47.320 171.200 47.380 ;
        RECT 186.075 47.320 186.365 47.365 ;
        RECT 205.380 47.320 205.700 47.380 ;
        RECT 218.260 47.320 218.580 47.380 ;
        RECT 170.880 47.180 185.370 47.320 ;
        RECT 170.880 47.120 171.200 47.180 ;
        RECT 144.675 46.980 144.965 47.025 ;
        RECT 143.740 46.840 144.965 46.980 ;
        RECT 122.595 46.795 122.885 46.840 ;
        RECT 119.360 46.780 119.680 46.795 ;
        RECT 143.740 46.780 144.060 46.840 ;
        RECT 144.675 46.795 144.965 46.840 ;
        RECT 145.120 46.980 145.440 47.040 ;
        RECT 145.120 46.840 145.635 46.980 ;
        RECT 145.120 46.780 145.440 46.840 ;
        RECT 146.975 46.795 147.265 47.025 ;
        RECT 147.420 46.980 147.740 47.040 ;
        RECT 156.635 46.980 156.925 47.025 ;
        RECT 160.300 46.980 160.620 47.040 ;
        RECT 147.420 46.840 147.935 46.980 ;
        RECT 156.635 46.840 160.620 46.980 ;
        RECT 102.340 46.500 111.770 46.640 ;
        RECT 112.920 46.640 113.240 46.700 ;
        RECT 115.680 46.640 116.000 46.700 ;
        RECT 118.900 46.640 119.220 46.700 ;
        RECT 112.920 46.500 116.000 46.640 ;
        RECT 118.705 46.500 119.220 46.640 ;
        RECT 102.340 46.440 102.660 46.500 ;
        RECT 112.920 46.440 113.240 46.500 ;
        RECT 115.680 46.440 116.000 46.500 ;
        RECT 118.900 46.440 119.220 46.500 ;
        RECT 120.740 46.640 121.060 46.700 ;
        RECT 128.580 46.640 128.870 46.685 ;
        RECT 129.980 46.640 130.270 46.685 ;
        RECT 131.820 46.640 132.110 46.685 ;
        RECT 120.740 46.500 122.810 46.640 ;
        RECT 120.740 46.440 121.060 46.500 ;
        RECT 40.700 46.160 64.390 46.300 ;
        RECT 72.915 46.300 73.205 46.345 ;
        RECT 85.320 46.300 85.640 46.360 ;
        RECT 86.240 46.300 86.560 46.360 ;
        RECT 72.915 46.160 85.640 46.300 ;
        RECT 86.045 46.160 86.560 46.300 ;
        RECT 40.700 46.100 41.020 46.160 ;
        RECT 72.915 46.115 73.205 46.160 ;
        RECT 85.320 46.100 85.640 46.160 ;
        RECT 86.240 46.100 86.560 46.160 ;
        RECT 92.680 46.300 93.000 46.360 ;
        RECT 98.200 46.300 98.520 46.360 ;
        RECT 104.640 46.300 104.960 46.360 ;
        RECT 92.680 46.160 98.520 46.300 ;
        RECT 104.445 46.160 104.960 46.300 ;
        RECT 122.670 46.300 122.810 46.500 ;
        RECT 128.580 46.500 132.110 46.640 ;
        RECT 128.580 46.455 128.870 46.500 ;
        RECT 129.980 46.455 130.270 46.500 ;
        RECT 131.820 46.455 132.110 46.500 ;
        RECT 137.760 46.640 138.080 46.700 ;
        RECT 147.050 46.640 147.190 46.795 ;
        RECT 147.420 46.780 147.740 46.840 ;
        RECT 156.635 46.795 156.925 46.840 ;
        RECT 160.300 46.780 160.620 46.840 ;
        RECT 169.055 46.980 169.345 47.025 ;
        RECT 177.780 46.980 178.100 47.040 ;
        RECT 184.680 46.980 185.000 47.040 ;
        RECT 169.055 46.840 185.000 46.980 ;
        RECT 185.230 46.980 185.370 47.180 ;
        RECT 186.075 47.180 205.700 47.320 ;
        RECT 186.075 47.135 186.365 47.180 ;
        RECT 205.380 47.120 205.700 47.180 ;
        RECT 209.150 47.180 218.580 47.320 ;
        RECT 194.800 46.980 195.120 47.040 ;
        RECT 197.100 46.980 197.420 47.040 ;
        RECT 185.230 46.840 195.120 46.980 ;
        RECT 196.905 46.840 197.420 46.980 ;
        RECT 169.055 46.795 169.345 46.840 ;
        RECT 177.780 46.780 178.100 46.840 ;
        RECT 184.680 46.780 185.000 46.840 ;
        RECT 194.800 46.780 195.120 46.840 ;
        RECT 197.100 46.780 197.420 46.840 ;
        RECT 198.495 46.980 198.785 47.025 ;
        RECT 209.150 46.980 209.290 47.180 ;
        RECT 218.260 47.120 218.580 47.180 ;
        RECT 222.875 47.320 223.165 47.365 ;
        RECT 230.220 47.320 230.540 47.380 ;
        RECT 222.875 47.180 230.540 47.320 ;
        RECT 222.875 47.135 223.165 47.180 ;
        RECT 230.220 47.120 230.540 47.180 ;
        RECT 230.680 47.120 231.000 47.380 ;
        RECT 231.600 47.365 231.920 47.380 ;
        RECT 231.430 47.135 231.920 47.365 ;
        RECT 232.535 47.320 232.825 47.365 ;
        RECT 232.980 47.320 233.300 47.380 ;
        RECT 232.535 47.180 233.300 47.320 ;
        RECT 232.535 47.135 232.825 47.180 ;
        RECT 231.600 47.120 231.920 47.135 ;
        RECT 232.980 47.120 233.300 47.180 ;
        RECT 234.375 47.320 234.665 47.365 ;
        RECT 234.820 47.320 235.140 47.380 ;
        RECT 239.510 47.365 239.650 47.520 ;
        RECT 242.640 47.460 242.960 47.520 ;
        RECT 251.165 47.475 251.455 47.520 ;
        RECT 251.855 47.660 252.145 47.705 ;
        RECT 253.680 47.660 254.000 47.720 ;
        RECT 251.855 47.520 254.000 47.660 ;
        RECT 251.855 47.475 252.145 47.520 ;
        RECT 253.680 47.460 254.000 47.520 ;
        RECT 264.260 47.660 264.580 47.720 ;
        RECT 271.250 47.660 271.390 47.860 ;
        RECT 276.220 47.800 276.540 47.860 ;
        RECT 283.580 48.000 283.900 48.060 ;
        RECT 311.640 48.000 311.960 48.060 ;
        RECT 317.620 48.000 317.940 48.060 ;
        RECT 283.580 47.860 311.410 48.000 ;
        RECT 283.580 47.800 283.900 47.860 ;
        RECT 264.260 47.520 271.390 47.660 ;
        RECT 274.380 47.660 274.700 47.720 ;
        RECT 309.800 47.660 310.120 47.720 ;
        RECT 274.380 47.520 310.120 47.660 ;
        RECT 311.270 47.660 311.410 47.860 ;
        RECT 311.640 47.860 317.940 48.000 ;
        RECT 311.640 47.800 311.960 47.860 ;
        RECT 317.620 47.800 317.940 47.860 ;
        RECT 325.900 48.000 326.220 48.060 ;
        RECT 333.720 48.000 334.040 48.060 ;
        RECT 325.900 47.860 334.040 48.000 ;
        RECT 325.900 47.800 326.220 47.860 ;
        RECT 333.720 47.800 334.040 47.860 ;
        RECT 334.180 48.000 334.500 48.060 ;
        RECT 342.920 48.000 343.240 48.060 ;
        RECT 361.780 48.000 362.100 48.060 ;
        RECT 334.180 47.860 339.010 48.000 ;
        RECT 334.180 47.800 334.500 47.860 ;
        RECT 332.340 47.660 332.660 47.720 ;
        RECT 311.270 47.520 332.660 47.660 ;
        RECT 264.260 47.460 264.580 47.520 ;
        RECT 274.380 47.460 274.700 47.520 ;
        RECT 309.800 47.460 310.120 47.520 ;
        RECT 332.340 47.460 332.660 47.520 ;
        RECT 234.375 47.180 235.140 47.320 ;
        RECT 234.375 47.135 234.665 47.180 ;
        RECT 234.820 47.120 235.140 47.180 ;
        RECT 239.435 47.135 239.725 47.365 ;
        RECT 241.740 47.320 242.030 47.365 ;
        RECT 244.520 47.320 244.810 47.365 ;
        RECT 245.400 47.320 245.720 47.380 ;
        RECT 252.300 47.320 252.620 47.380 ;
        RECT 292.320 47.320 292.640 47.380 ;
        RECT 239.970 47.180 241.490 47.320 ;
        RECT 198.495 46.840 209.290 46.980 ;
        RECT 198.495 46.795 198.785 46.840 ;
        RECT 212.110 46.795 212.400 47.025 ;
        RECT 213.070 46.980 213.360 47.025 ;
        RECT 214.120 46.980 214.440 47.040 ;
        RECT 220.100 46.980 220.420 47.040 ;
        RECT 213.070 46.840 214.440 46.980 ;
        RECT 219.905 46.840 220.420 46.980 ;
        RECT 213.070 46.795 213.360 46.840 ;
        RECT 137.760 46.500 147.190 46.640 ;
        RECT 156.180 46.640 156.470 46.685 ;
        RECT 157.580 46.640 157.870 46.685 ;
        RECT 159.420 46.640 159.710 46.685 ;
        RECT 156.180 46.500 159.710 46.640 ;
        RECT 137.760 46.440 138.080 46.500 ;
        RECT 156.180 46.455 156.470 46.500 ;
        RECT 157.580 46.455 157.870 46.500 ;
        RECT 159.420 46.455 159.710 46.500 ;
        RECT 169.980 46.640 170.270 46.685 ;
        RECT 171.380 46.640 171.670 46.685 ;
        RECT 173.220 46.640 173.510 46.685 ;
        RECT 185.620 46.640 185.910 46.685 ;
        RECT 187.020 46.640 187.310 46.685 ;
        RECT 188.860 46.640 189.150 46.685 ;
        RECT 196.640 46.640 196.960 46.700 ;
        RECT 169.980 46.500 173.510 46.640 ;
        RECT 169.980 46.455 170.270 46.500 ;
        RECT 171.380 46.455 171.670 46.500 ;
        RECT 173.220 46.455 173.510 46.500 ;
        RECT 173.730 46.500 176.630 46.640 ;
        RECT 140.980 46.300 141.300 46.360 ;
        RECT 122.670 46.160 141.300 46.300 ;
        RECT 92.680 46.100 93.000 46.160 ;
        RECT 98.200 46.100 98.520 46.160 ;
        RECT 104.640 46.100 104.960 46.160 ;
        RECT 140.980 46.100 141.300 46.160 ;
        RECT 142.360 46.300 142.680 46.360 ;
        RECT 156.620 46.300 156.940 46.360 ;
        RECT 142.360 46.160 156.940 46.300 ;
        RECT 142.360 46.100 142.680 46.160 ;
        RECT 156.620 46.100 156.940 46.160 ;
        RECT 160.300 46.300 160.620 46.360 ;
        RECT 162.155 46.300 162.445 46.345 ;
        RECT 160.300 46.160 162.445 46.300 ;
        RECT 160.300 46.100 160.620 46.160 ;
        RECT 162.155 46.115 162.445 46.160 ;
        RECT 165.820 46.300 166.140 46.360 ;
        RECT 173.730 46.300 173.870 46.500 ;
        RECT 165.820 46.160 173.870 46.300 ;
        RECT 176.490 46.300 176.630 46.500 ;
        RECT 185.620 46.500 189.150 46.640 ;
        RECT 185.620 46.455 185.910 46.500 ;
        RECT 187.020 46.455 187.310 46.500 ;
        RECT 188.860 46.455 189.150 46.500 ;
        RECT 189.370 46.500 196.960 46.640 ;
        RECT 189.370 46.300 189.510 46.500 ;
        RECT 196.640 46.440 196.960 46.500 ;
        RECT 198.040 46.640 198.330 46.685 ;
        RECT 199.440 46.640 199.730 46.685 ;
        RECT 201.280 46.640 201.570 46.685 ;
        RECT 198.040 46.500 201.570 46.640 ;
        RECT 198.040 46.455 198.330 46.500 ;
        RECT 199.440 46.455 199.730 46.500 ;
        RECT 201.280 46.455 201.570 46.500 ;
        RECT 202.160 46.640 202.480 46.700 ;
        RECT 205.395 46.640 205.685 46.685 ;
        RECT 202.160 46.500 205.685 46.640 ;
        RECT 202.160 46.440 202.480 46.500 ;
        RECT 205.395 46.455 205.685 46.500 ;
        RECT 211.375 46.455 211.665 46.685 ;
        RECT 212.185 46.640 212.325 46.795 ;
        RECT 214.120 46.780 214.440 46.840 ;
        RECT 220.100 46.780 220.420 46.840 ;
        RECT 220.575 46.980 220.865 47.025 ;
        RECT 228.380 46.980 228.700 47.040 ;
        RECT 220.575 46.840 228.700 46.980 ;
        RECT 230.770 46.980 230.910 47.120 ;
        RECT 239.970 46.980 240.110 47.180 ;
        RECT 230.770 46.840 240.110 46.980 ;
        RECT 240.340 46.980 240.660 47.040 ;
        RECT 240.340 46.840 240.855 46.980 ;
        RECT 220.575 46.795 220.865 46.840 ;
        RECT 228.380 46.780 228.700 46.840 ;
        RECT 240.340 46.780 240.660 46.840 ;
        RECT 227.460 46.640 227.780 46.700 ;
        RECT 212.185 46.500 227.780 46.640 ;
        RECT 176.490 46.160 189.510 46.300 ;
        RECT 211.450 46.300 211.590 46.455 ;
        RECT 227.460 46.440 227.780 46.500 ;
        RECT 230.695 46.640 230.985 46.685 ;
        RECT 231.140 46.640 231.460 46.700 ;
        RECT 230.695 46.500 231.460 46.640 ;
        RECT 230.695 46.455 230.985 46.500 ;
        RECT 231.140 46.440 231.460 46.500 ;
        RECT 231.600 46.640 231.920 46.700 ;
        RECT 233.440 46.640 233.760 46.700 ;
        RECT 231.600 46.500 233.760 46.640 ;
        RECT 231.600 46.440 231.920 46.500 ;
        RECT 233.440 46.440 233.760 46.500 ;
        RECT 233.900 46.640 234.220 46.700 ;
        RECT 238.040 46.640 238.360 46.700 ;
        RECT 238.960 46.640 239.280 46.700 ;
        RECT 233.900 46.500 239.280 46.640 ;
        RECT 241.350 46.640 241.490 47.180 ;
        RECT 241.740 47.180 244.810 47.320 ;
        RECT 245.205 47.180 245.720 47.320 ;
        RECT 252.105 47.180 252.620 47.320 ;
        RECT 241.740 47.135 242.030 47.180 ;
        RECT 244.520 47.135 244.810 47.180 ;
        RECT 245.400 47.120 245.720 47.180 ;
        RECT 252.300 47.120 252.620 47.180 ;
        RECT 254.230 47.180 287.950 47.320 ;
        RECT 242.685 46.795 242.975 47.025 ;
        RECT 243.115 46.980 243.405 47.025 ;
        RECT 243.560 46.980 243.880 47.040 ;
        RECT 243.115 46.840 243.880 46.980 ;
        RECT 243.115 46.795 243.405 46.840 ;
        RECT 242.730 46.640 242.870 46.795 ;
        RECT 243.560 46.780 243.880 46.840 ;
        RECT 244.020 46.980 244.340 47.040 ;
        RECT 250.475 46.980 250.765 47.025 ;
        RECT 251.840 46.980 252.160 47.040 ;
        RECT 244.020 46.840 246.550 46.980 ;
        RECT 244.020 46.780 244.340 46.840 ;
        RECT 241.350 46.500 242.870 46.640 ;
        RECT 246.410 46.640 246.550 46.840 ;
        RECT 250.475 46.840 252.160 46.980 ;
        RECT 250.475 46.795 250.765 46.840 ;
        RECT 251.840 46.780 252.160 46.840 ;
        RECT 253.220 46.980 253.540 47.040 ;
        RECT 254.230 46.980 254.370 47.180 ;
        RECT 253.220 46.840 254.370 46.980 ;
        RECT 255.980 46.980 256.300 47.040 ;
        RECT 259.215 46.980 259.505 47.025 ;
        RECT 261.040 46.980 261.360 47.040 ;
        RECT 255.980 46.840 259.505 46.980 ;
        RECT 260.845 46.840 261.360 46.980 ;
        RECT 253.220 46.780 253.540 46.840 ;
        RECT 255.980 46.780 256.300 46.840 ;
        RECT 259.215 46.795 259.505 46.840 ;
        RECT 261.040 46.780 261.360 46.840 ;
        RECT 267.495 46.980 267.785 47.025 ;
        RECT 270.700 46.980 271.020 47.040 ;
        RECT 267.495 46.840 271.020 46.980 ;
        RECT 267.495 46.795 267.785 46.840 ;
        RECT 270.700 46.780 271.020 46.840 ;
        RECT 274.395 46.795 274.685 47.025 ;
        RECT 275.760 46.980 276.080 47.040 ;
        RECT 284.040 46.980 284.360 47.040 ;
        RECT 287.275 46.980 287.565 47.025 ;
        RECT 275.565 46.840 276.080 46.980 ;
        RECT 283.845 46.840 287.565 46.980 ;
        RECT 254.600 46.640 254.920 46.700 ;
        RECT 246.410 46.500 254.920 46.640 ;
        RECT 233.900 46.440 234.220 46.500 ;
        RECT 238.040 46.440 238.360 46.500 ;
        RECT 238.960 46.440 239.280 46.500 ;
        RECT 254.600 46.440 254.920 46.500 ;
        RECT 256.440 46.640 256.760 46.700 ;
        RECT 258.295 46.640 258.585 46.685 ;
        RECT 274.470 46.640 274.610 46.795 ;
        RECT 275.760 46.780 276.080 46.840 ;
        RECT 284.040 46.780 284.360 46.840 ;
        RECT 287.275 46.795 287.565 46.840 ;
        RECT 286.800 46.640 287.120 46.700 ;
        RECT 256.440 46.500 258.585 46.640 ;
        RECT 256.440 46.440 256.760 46.500 ;
        RECT 258.295 46.455 258.585 46.500 ;
        RECT 262.050 46.500 274.150 46.640 ;
        RECT 274.470 46.500 287.120 46.640 ;
        RECT 214.580 46.300 214.900 46.360 ;
        RECT 211.450 46.160 214.900 46.300 ;
        RECT 165.820 46.100 166.140 46.160 ;
        RECT 214.580 46.100 214.900 46.160 ;
        RECT 228.380 46.300 228.700 46.360 ;
        RECT 246.320 46.300 246.640 46.360 ;
        RECT 228.380 46.160 246.640 46.300 ;
        RECT 228.380 46.100 228.700 46.160 ;
        RECT 246.320 46.100 246.640 46.160 ;
        RECT 246.780 46.300 247.100 46.360 ;
        RECT 262.050 46.300 262.190 46.500 ;
        RECT 246.780 46.160 262.190 46.300 ;
        RECT 262.420 46.300 262.740 46.360 ;
        RECT 273.475 46.300 273.765 46.345 ;
        RECT 262.420 46.160 273.765 46.300 ;
        RECT 274.010 46.300 274.150 46.500 ;
        RECT 286.800 46.440 287.120 46.500 ;
        RECT 284.500 46.300 284.820 46.360 ;
        RECT 285.420 46.300 285.740 46.360 ;
        RECT 274.010 46.160 284.820 46.300 ;
        RECT 285.225 46.160 285.740 46.300 ;
        RECT 287.810 46.300 287.950 47.180 ;
        RECT 288.270 47.180 292.640 47.320 ;
        RECT 288.270 47.025 288.410 47.180 ;
        RECT 292.320 47.120 292.640 47.180 ;
        RECT 293.240 47.320 293.560 47.380 ;
        RECT 297.855 47.320 298.145 47.365 ;
        RECT 316.240 47.320 316.560 47.380 ;
        RECT 338.320 47.320 338.640 47.380 ;
        RECT 293.240 47.180 298.145 47.320 ;
        RECT 293.240 47.120 293.560 47.180 ;
        RECT 297.855 47.135 298.145 47.180 ;
        RECT 304.830 47.180 316.560 47.320 ;
        RECT 288.195 46.795 288.485 47.025 ;
        RECT 289.100 46.980 289.420 47.040 ;
        RECT 290.035 46.980 290.325 47.025 ;
        RECT 290.940 46.980 291.260 47.040 ;
        RECT 298.300 46.980 298.620 47.040 ;
        RECT 289.100 46.840 290.325 46.980 ;
        RECT 290.745 46.840 291.260 46.980 ;
        RECT 298.105 46.840 298.620 46.980 ;
        RECT 289.100 46.780 289.420 46.840 ;
        RECT 290.035 46.795 290.325 46.840 ;
        RECT 290.940 46.780 291.260 46.840 ;
        RECT 298.300 46.780 298.620 46.840 ;
        RECT 299.680 46.980 300.000 47.040 ;
        RECT 304.830 47.025 304.970 47.180 ;
        RECT 316.240 47.120 316.560 47.180 ;
        RECT 316.790 47.180 338.640 47.320 ;
        RECT 338.870 47.320 339.010 47.860 ;
        RECT 342.920 47.860 362.100 48.000 ;
        RECT 342.920 47.800 343.240 47.860 ;
        RECT 361.780 47.800 362.100 47.860 ;
        RECT 362.240 48.000 362.560 48.060 ;
        RECT 380.180 48.000 380.500 48.060 ;
        RECT 362.240 47.860 380.500 48.000 ;
        RECT 362.240 47.800 362.560 47.860 ;
        RECT 380.180 47.800 380.500 47.860 ;
        RECT 390.775 47.660 391.065 47.705 ;
        RECT 381.650 47.520 391.065 47.660 ;
        RECT 350.740 47.320 351.060 47.380 ;
        RECT 370.520 47.320 370.840 47.380 ;
        RECT 373.740 47.320 374.060 47.380 ;
        RECT 381.650 47.320 381.790 47.520 ;
        RECT 390.775 47.475 391.065 47.520 ;
        RECT 338.870 47.180 351.060 47.320 ;
        RECT 299.680 46.840 304.050 46.980 ;
        RECT 299.680 46.780 300.000 46.840 ;
        RECT 295.630 46.500 296.690 46.640 ;
        RECT 295.630 46.300 295.770 46.500 ;
        RECT 287.810 46.160 295.770 46.300 ;
        RECT 296.550 46.300 296.690 46.500 ;
        RECT 302.900 46.300 303.220 46.360 ;
        RECT 303.910 46.345 304.050 46.840 ;
        RECT 304.755 46.795 305.045 47.025 ;
        RECT 306.120 46.980 306.440 47.040 ;
        RECT 305.925 46.840 306.440 46.980 ;
        RECT 306.120 46.780 306.440 46.840 ;
        RECT 311.195 46.795 311.485 47.025 ;
        RECT 313.955 46.980 314.245 47.025 ;
        RECT 314.400 46.980 314.720 47.040 ;
        RECT 313.955 46.840 314.720 46.980 ;
        RECT 313.955 46.795 314.245 46.840 ;
        RECT 311.270 46.360 311.410 46.795 ;
        RECT 314.400 46.780 314.720 46.840 ;
        RECT 314.860 46.980 315.180 47.040 ;
        RECT 316.790 46.980 316.930 47.180 ;
        RECT 338.320 47.120 338.640 47.180 ;
        RECT 350.740 47.120 351.060 47.180 ;
        RECT 354.050 47.180 362.010 47.320 ;
        RECT 314.860 46.840 316.930 46.980 ;
        RECT 314.860 46.780 315.180 46.840 ;
        RECT 324.995 46.795 325.285 47.025 ;
        RECT 326.360 46.980 326.680 47.040 ;
        RECT 332.800 46.980 333.120 47.040 ;
        RECT 326.165 46.840 326.680 46.980 ;
        RECT 332.605 46.840 333.120 46.980 ;
        RECT 325.070 46.640 325.210 46.795 ;
        RECT 326.360 46.780 326.680 46.840 ;
        RECT 332.800 46.780 333.120 46.840 ;
        RECT 333.260 46.980 333.580 47.040 ;
        RECT 333.735 46.980 334.025 47.025 ;
        RECT 340.160 46.980 340.480 47.040 ;
        RECT 333.260 46.840 340.480 46.980 ;
        RECT 333.260 46.780 333.580 46.840 ;
        RECT 333.735 46.795 334.025 46.840 ;
        RECT 340.160 46.780 340.480 46.840 ;
        RECT 340.635 46.980 340.925 47.025 ;
        RECT 341.540 46.980 341.860 47.040 ;
        RECT 342.015 46.980 342.305 47.025 ;
        RECT 347.520 46.980 347.840 47.040 ;
        RECT 340.635 46.840 341.235 46.980 ;
        RECT 340.635 46.795 340.925 46.840 ;
        RECT 330.960 46.640 331.280 46.700 ;
        RECT 325.070 46.500 331.280 46.640 ;
        RECT 330.960 46.440 331.280 46.500 ;
        RECT 334.180 46.640 334.500 46.700 ;
        RECT 335.115 46.640 335.405 46.685 ;
        RECT 334.180 46.500 335.405 46.640 ;
        RECT 334.180 46.440 334.500 46.500 ;
        RECT 335.115 46.455 335.405 46.500 ;
        RECT 296.550 46.160 303.220 46.300 ;
        RECT 246.780 46.100 247.100 46.160 ;
        RECT 262.420 46.100 262.740 46.160 ;
        RECT 273.475 46.115 273.765 46.160 ;
        RECT 284.500 46.100 284.820 46.160 ;
        RECT 285.420 46.100 285.740 46.160 ;
        RECT 302.900 46.100 303.220 46.160 ;
        RECT 303.835 46.115 304.125 46.345 ;
        RECT 311.180 46.100 311.500 46.360 ;
        RECT 312.560 46.300 312.880 46.360 ;
        RECT 324.060 46.300 324.380 46.360 ;
        RECT 312.365 46.160 312.880 46.300 ;
        RECT 323.865 46.160 324.380 46.300 ;
        RECT 312.560 46.100 312.880 46.160 ;
        RECT 324.060 46.100 324.380 46.160 ;
        RECT 325.440 46.300 325.760 46.360 ;
        RECT 338.780 46.300 339.100 46.360 ;
        RECT 339.700 46.300 340.020 46.360 ;
        RECT 325.440 46.160 339.100 46.300 ;
        RECT 339.505 46.160 340.020 46.300 ;
        RECT 341.095 46.300 341.235 46.840 ;
        RECT 341.540 46.840 347.840 46.980 ;
        RECT 341.540 46.780 341.860 46.840 ;
        RECT 342.015 46.795 342.305 46.840 ;
        RECT 347.520 46.780 347.840 46.840 ;
        RECT 353.055 46.795 353.345 47.025 ;
        RECT 353.500 46.980 353.820 47.040 ;
        RECT 354.050 47.025 354.190 47.180 ;
        RECT 361.870 47.025 362.010 47.180 ;
        RECT 368.310 47.180 370.290 47.320 ;
        RECT 353.975 46.980 354.265 47.025 ;
        RECT 353.500 46.840 354.265 46.980 ;
        RECT 342.460 46.640 342.780 46.700 ;
        RECT 353.130 46.640 353.270 46.795 ;
        RECT 353.500 46.780 353.820 46.840 ;
        RECT 353.975 46.795 354.265 46.840 ;
        RECT 360.875 46.795 361.165 47.025 ;
        RECT 361.795 46.795 362.085 47.025 ;
        RECT 356.720 46.640 357.040 46.700 ;
        RECT 360.950 46.640 361.090 46.795 ;
        RECT 367.760 46.640 368.080 46.700 ;
        RECT 342.460 46.500 352.350 46.640 ;
        RECT 353.130 46.500 357.040 46.640 ;
        RECT 342.460 46.440 342.780 46.500 ;
        RECT 345.680 46.300 346.000 46.360 ;
        RECT 352.210 46.345 352.350 46.500 ;
        RECT 356.720 46.440 357.040 46.500 ;
        RECT 357.270 46.500 360.630 46.640 ;
        RECT 360.950 46.500 368.080 46.640 ;
        RECT 341.095 46.160 346.000 46.300 ;
        RECT 325.440 46.100 325.760 46.160 ;
        RECT 338.780 46.100 339.100 46.160 ;
        RECT 339.700 46.100 340.020 46.160 ;
        RECT 345.680 46.100 346.000 46.160 ;
        RECT 352.135 46.115 352.425 46.345 ;
        RECT 352.580 46.300 352.900 46.360 ;
        RECT 357.270 46.300 357.410 46.500 ;
        RECT 352.580 46.160 357.410 46.300 ;
        RECT 357.640 46.300 357.960 46.360 ;
        RECT 359.955 46.300 360.245 46.345 ;
        RECT 357.640 46.160 360.245 46.300 ;
        RECT 360.490 46.300 360.630 46.500 ;
        RECT 367.760 46.440 368.080 46.500 ;
        RECT 368.310 46.300 368.450 47.180 ;
        RECT 368.695 46.795 368.985 47.025 ;
        RECT 369.140 46.980 369.460 47.040 ;
        RECT 369.615 46.980 369.905 47.025 ;
        RECT 369.140 46.840 369.905 46.980 ;
        RECT 370.150 46.980 370.290 47.180 ;
        RECT 370.520 47.180 371.035 47.320 ;
        RECT 373.740 47.180 381.790 47.320 ;
        RECT 370.520 47.120 370.840 47.180 ;
        RECT 373.740 47.120 374.060 47.180 ;
        RECT 385.715 46.980 386.005 47.025 ;
        RECT 370.150 46.840 386.005 46.980 ;
        RECT 368.770 46.640 368.910 46.795 ;
        RECT 369.140 46.780 369.460 46.840 ;
        RECT 369.615 46.795 369.905 46.840 ;
        RECT 385.715 46.795 386.005 46.840 ;
        RECT 399.500 46.980 399.820 47.040 ;
        RECT 400.895 46.980 401.185 47.025 ;
        RECT 399.500 46.840 401.185 46.980 ;
        RECT 399.500 46.780 399.820 46.840 ;
        RECT 400.895 46.795 401.185 46.840 ;
        RECT 406.860 46.980 407.180 47.040 ;
        RECT 408.715 46.980 409.005 47.025 ;
        RECT 406.860 46.840 409.005 46.980 ;
        RECT 406.860 46.780 407.180 46.840 ;
        RECT 408.715 46.795 409.005 46.840 ;
        RECT 410.540 46.980 410.860 47.040 ;
        RECT 413.775 46.980 414.065 47.025 ;
        RECT 410.540 46.840 414.065 46.980 ;
        RECT 410.540 46.780 410.860 46.840 ;
        RECT 413.775 46.795 414.065 46.840 ;
        RECT 417.900 46.980 418.220 47.040 ;
        RECT 418.835 46.980 419.125 47.025 ;
        RECT 417.900 46.840 419.125 46.980 ;
        RECT 417.900 46.780 418.220 46.840 ;
        RECT 418.835 46.795 419.125 46.840 ;
        RECT 421.580 46.980 421.900 47.040 ;
        RECT 423.895 46.980 424.185 47.025 ;
        RECT 421.580 46.840 424.185 46.980 ;
        RECT 421.580 46.780 421.900 46.840 ;
        RECT 423.895 46.795 424.185 46.840 ;
        RECT 425.260 46.980 425.580 47.040 ;
        RECT 428.955 46.980 429.245 47.025 ;
        RECT 425.260 46.840 429.245 46.980 ;
        RECT 425.260 46.780 425.580 46.840 ;
        RECT 428.955 46.795 429.245 46.840 ;
        RECT 439.980 46.980 440.300 47.040 ;
        RECT 441.835 46.980 442.125 47.025 ;
        RECT 439.980 46.840 442.125 46.980 ;
        RECT 439.980 46.780 440.300 46.840 ;
        RECT 441.835 46.795 442.125 46.840 ;
        RECT 443.660 46.980 443.980 47.040 ;
        RECT 446.895 46.980 447.185 47.025 ;
        RECT 443.660 46.840 447.185 46.980 ;
        RECT 443.660 46.780 443.980 46.840 ;
        RECT 446.895 46.795 447.185 46.840 ;
        RECT 451.020 46.980 451.340 47.040 ;
        RECT 451.955 46.980 452.245 47.025 ;
        RECT 451.020 46.840 452.245 46.980 ;
        RECT 451.020 46.780 451.340 46.840 ;
        RECT 451.955 46.795 452.245 46.840 ;
        RECT 454.700 46.980 455.020 47.040 ;
        RECT 457.015 46.980 457.305 47.025 ;
        RECT 454.700 46.840 457.305 46.980 ;
        RECT 454.700 46.780 455.020 46.840 ;
        RECT 457.015 46.795 457.305 46.840 ;
        RECT 465.740 46.980 466.060 47.040 ;
        RECT 469.895 46.980 470.185 47.025 ;
        RECT 465.740 46.840 470.185 46.980 ;
        RECT 465.740 46.780 466.060 46.840 ;
        RECT 469.895 46.795 470.185 46.840 ;
        RECT 473.100 46.980 473.420 47.040 ;
        RECT 474.955 46.980 475.245 47.025 ;
        RECT 473.100 46.840 475.245 46.980 ;
        RECT 473.100 46.780 473.420 46.840 ;
        RECT 474.955 46.795 475.245 46.840 ;
        RECT 476.780 46.980 477.100 47.040 ;
        RECT 480.015 46.980 480.305 47.025 ;
        RECT 476.780 46.840 480.305 46.980 ;
        RECT 476.780 46.780 477.100 46.840 ;
        RECT 480.015 46.795 480.305 46.840 ;
        RECT 484.140 46.980 484.460 47.040 ;
        RECT 485.075 46.980 485.365 47.025 ;
        RECT 484.140 46.840 485.365 46.980 ;
        RECT 484.140 46.780 484.460 46.840 ;
        RECT 485.075 46.795 485.365 46.840 ;
        RECT 491.500 46.980 491.820 47.040 ;
        RECT 492.895 46.980 493.185 47.025 ;
        RECT 491.500 46.840 493.185 46.980 ;
        RECT 491.500 46.780 491.820 46.840 ;
        RECT 492.895 46.795 493.185 46.840 ;
        RECT 495.180 46.980 495.500 47.040 ;
        RECT 497.955 46.980 498.245 47.025 ;
        RECT 495.180 46.840 498.245 46.980 ;
        RECT 495.180 46.780 495.500 46.840 ;
        RECT 497.955 46.795 498.245 46.840 ;
        RECT 498.860 46.980 499.180 47.040 ;
        RECT 503.015 46.980 503.305 47.025 ;
        RECT 498.860 46.840 503.305 46.980 ;
        RECT 498.860 46.780 499.180 46.840 ;
        RECT 503.015 46.795 503.305 46.840 ;
        RECT 506.220 46.980 506.540 47.040 ;
        RECT 508.075 46.980 508.365 47.025 ;
        RECT 506.220 46.840 508.365 46.980 ;
        RECT 506.220 46.780 506.540 46.840 ;
        RECT 508.075 46.795 508.365 46.840 ;
        RECT 517.260 46.980 517.580 47.040 ;
        RECT 520.955 46.980 521.245 47.025 ;
        RECT 517.260 46.840 521.245 46.980 ;
        RECT 517.260 46.780 517.580 46.840 ;
        RECT 520.955 46.795 521.245 46.840 ;
        RECT 524.620 46.980 524.940 47.040 ;
        RECT 526.015 46.980 526.305 47.025 ;
        RECT 524.620 46.840 526.305 46.980 ;
        RECT 524.620 46.780 524.940 46.840 ;
        RECT 526.015 46.795 526.305 46.840 ;
        RECT 528.300 46.980 528.620 47.040 ;
        RECT 531.075 46.980 531.365 47.025 ;
        RECT 528.300 46.840 531.365 46.980 ;
        RECT 528.300 46.780 528.620 46.840 ;
        RECT 531.075 46.795 531.365 46.840 ;
        RECT 531.980 46.980 532.300 47.040 ;
        RECT 536.135 46.980 536.425 47.025 ;
        RECT 531.980 46.840 536.425 46.980 ;
        RECT 531.980 46.780 532.300 46.840 ;
        RECT 536.135 46.795 536.425 46.840 ;
        RECT 539.340 46.980 539.660 47.040 ;
        RECT 541.195 46.980 541.485 47.025 ;
        RECT 539.340 46.840 541.485 46.980 ;
        RECT 539.340 46.780 539.660 46.840 ;
        RECT 541.195 46.795 541.485 46.840 ;
        RECT 546.700 46.980 547.020 47.040 ;
        RECT 549.015 46.980 549.305 47.025 ;
        RECT 546.700 46.840 549.305 46.980 ;
        RECT 546.700 46.780 547.020 46.840 ;
        RECT 549.015 46.795 549.305 46.840 ;
        RECT 550.380 46.980 550.700 47.040 ;
        RECT 554.075 46.980 554.365 47.025 ;
        RECT 550.380 46.840 554.365 46.980 ;
        RECT 550.380 46.780 550.700 46.840 ;
        RECT 554.075 46.795 554.365 46.840 ;
        RECT 557.740 46.980 558.060 47.040 ;
        RECT 559.135 46.980 559.425 47.025 ;
        RECT 557.740 46.840 559.425 46.980 ;
        RECT 557.740 46.780 558.060 46.840 ;
        RECT 559.135 46.795 559.425 46.840 ;
        RECT 561.420 46.980 561.740 47.040 ;
        RECT 564.195 46.980 564.485 47.025 ;
        RECT 561.420 46.840 564.485 46.980 ;
        RECT 561.420 46.780 561.740 46.840 ;
        RECT 564.195 46.795 564.485 46.840 ;
        RECT 568.320 46.980 568.640 47.040 ;
        RECT 569.255 46.980 569.545 47.025 ;
        RECT 568.320 46.840 569.545 46.980 ;
        RECT 568.320 46.780 568.640 46.840 ;
        RECT 569.255 46.795 569.545 46.840 ;
        RECT 575.680 46.980 576.000 47.040 ;
        RECT 577.075 46.980 577.365 47.025 ;
        RECT 575.680 46.840 577.365 46.980 ;
        RECT 575.680 46.780 576.000 46.840 ;
        RECT 577.075 46.795 577.365 46.840 ;
        RECT 579.360 46.980 579.680 47.040 ;
        RECT 582.135 46.980 582.425 47.025 ;
        RECT 579.360 46.840 582.425 46.980 ;
        RECT 579.360 46.780 579.680 46.840 ;
        RECT 582.135 46.795 582.425 46.840 ;
        RECT 583.040 46.980 583.360 47.040 ;
        RECT 587.195 46.980 587.485 47.025 ;
        RECT 583.040 46.840 587.485 46.980 ;
        RECT 583.040 46.780 583.360 46.840 ;
        RECT 587.195 46.795 587.485 46.840 ;
        RECT 590.400 46.980 590.720 47.040 ;
        RECT 592.255 46.980 592.545 47.025 ;
        RECT 590.400 46.840 592.545 46.980 ;
        RECT 590.400 46.780 590.720 46.840 ;
        RECT 592.255 46.795 592.545 46.840 ;
        RECT 594.080 46.980 594.400 47.040 ;
        RECT 597.315 46.980 597.605 47.025 ;
        RECT 594.080 46.840 597.605 46.980 ;
        RECT 594.080 46.780 594.400 46.840 ;
        RECT 597.315 46.795 597.605 46.840 ;
        RECT 601.440 46.980 601.760 47.040 ;
        RECT 605.135 46.980 605.425 47.025 ;
        RECT 601.440 46.840 605.425 46.980 ;
        RECT 601.440 46.780 601.760 46.840 ;
        RECT 605.135 46.795 605.425 46.840 ;
        RECT 608.800 46.980 609.120 47.040 ;
        RECT 610.195 46.980 610.485 47.025 ;
        RECT 608.800 46.840 610.485 46.980 ;
        RECT 608.800 46.780 609.120 46.840 ;
        RECT 610.195 46.795 610.485 46.840 ;
        RECT 612.480 46.980 612.800 47.040 ;
        RECT 615.255 46.980 615.545 47.025 ;
        RECT 612.480 46.840 615.545 46.980 ;
        RECT 612.480 46.780 612.800 46.840 ;
        RECT 615.255 46.795 615.545 46.840 ;
        RECT 616.160 46.980 616.480 47.040 ;
        RECT 620.315 46.980 620.605 47.025 ;
        RECT 616.160 46.840 620.605 46.980 ;
        RECT 616.160 46.780 616.480 46.840 ;
        RECT 620.315 46.795 620.605 46.840 ;
        RECT 623.520 46.980 623.840 47.040 ;
        RECT 625.375 46.980 625.665 47.025 ;
        RECT 623.520 46.840 625.665 46.980 ;
        RECT 623.520 46.780 623.840 46.840 ;
        RECT 625.375 46.795 625.665 46.840 ;
        RECT 375.120 46.640 375.440 46.700 ;
        RECT 368.770 46.500 375.440 46.640 ;
        RECT 375.120 46.440 375.440 46.500 ;
        RECT 381.100 46.640 381.420 46.700 ;
        RECT 389.840 46.640 390.160 46.700 ;
        RECT 381.100 46.500 390.160 46.640 ;
        RECT 381.100 46.440 381.420 46.500 ;
        RECT 389.840 46.440 390.160 46.500 ;
        RECT 360.490 46.160 368.450 46.300 ;
        RECT 370.060 46.300 370.380 46.360 ;
        RECT 386.160 46.300 386.480 46.360 ;
        RECT 370.060 46.160 386.480 46.300 ;
        RECT 352.580 46.100 352.900 46.160 ;
        RECT 357.640 46.100 357.960 46.160 ;
        RECT 359.955 46.115 360.245 46.160 ;
        RECT 370.060 46.100 370.380 46.160 ;
        RECT 386.160 46.100 386.480 46.160 ;
        RECT 386.620 46.300 386.940 46.360 ;
        RECT 398.580 46.300 398.900 46.360 ;
        RECT 386.620 46.160 398.900 46.300 ;
        RECT 386.620 46.100 386.940 46.160 ;
        RECT 398.580 46.100 398.900 46.160 ;
        RECT 42.470 45.480 631.270 45.960 ;
        RECT 101.435 45.280 101.725 45.325 ;
        RECT 118.455 45.280 118.745 45.325 ;
        RECT 128.100 45.280 128.420 45.340 ;
        RECT 64.710 45.140 101.190 45.280 ;
        RECT 39.780 44.260 40.100 44.320 ;
        RECT 64.710 44.260 64.850 45.140 ;
        RECT 78.420 44.940 78.740 45.000 ;
        RECT 78.225 44.800 78.740 44.940 ;
        RECT 78.420 44.740 78.740 44.800 ;
        RECT 81.195 44.940 81.485 44.985 ;
        RECT 89.460 44.940 89.780 45.000 ;
        RECT 81.195 44.800 89.780 44.940 ;
        RECT 81.195 44.755 81.485 44.800 ;
        RECT 89.460 44.740 89.780 44.800 ;
        RECT 95.455 44.940 95.745 44.985 ;
        RECT 97.280 44.940 97.600 45.000 ;
        RECT 95.455 44.800 97.600 44.940 ;
        RECT 95.455 44.755 95.745 44.800 ;
        RECT 97.280 44.740 97.600 44.800 ;
        RECT 65.540 44.600 65.860 44.660 ;
        RECT 79.355 44.600 79.645 44.645 ;
        RECT 86.675 44.600 86.965 44.645 ;
        RECT 65.540 44.460 79.645 44.600 ;
        RECT 65.540 44.400 65.860 44.460 ;
        RECT 79.355 44.415 79.645 44.460 ;
        RECT 79.890 44.460 86.965 44.600 ;
        RECT 79.890 44.260 80.030 44.460 ;
        RECT 86.675 44.415 86.965 44.460 ;
        RECT 87.175 44.600 87.465 44.645 ;
        RECT 90.840 44.600 91.160 44.660 ;
        RECT 94.060 44.600 94.380 44.660 ;
        RECT 100.500 44.600 100.820 44.660 ;
        RECT 87.175 44.460 91.160 44.600 ;
        RECT 93.865 44.460 94.380 44.600 ;
        RECT 100.305 44.460 100.820 44.600 ;
        RECT 101.050 44.600 101.190 45.140 ;
        RECT 101.435 45.140 117.750 45.280 ;
        RECT 101.435 45.095 101.725 45.140 ;
        RECT 101.880 44.940 102.200 45.000 ;
        RECT 106.035 44.940 106.325 44.985 ;
        RECT 101.880 44.800 106.325 44.940 ;
        RECT 101.880 44.740 102.200 44.800 ;
        RECT 106.035 44.755 106.325 44.800 ;
        RECT 109.715 44.940 110.005 44.985 ;
        RECT 110.160 44.940 110.480 45.000 ;
        RECT 109.715 44.800 110.480 44.940 ;
        RECT 117.610 44.940 117.750 45.140 ;
        RECT 118.455 45.140 128.420 45.280 ;
        RECT 118.455 45.095 118.745 45.140 ;
        RECT 128.100 45.080 128.420 45.140 ;
        RECT 140.980 45.280 141.300 45.340 ;
        RECT 150.195 45.280 150.485 45.325 ;
        RECT 186.060 45.280 186.380 45.340 ;
        RECT 140.980 45.140 149.030 45.280 ;
        RECT 140.980 45.080 141.300 45.140 ;
        RECT 123.500 44.940 123.820 45.000 ;
        RECT 117.610 44.800 119.130 44.940 ;
        RECT 109.715 44.755 110.005 44.800 ;
        RECT 110.160 44.740 110.480 44.800 ;
        RECT 115.220 44.600 115.540 44.660 ;
        RECT 101.050 44.460 108.090 44.600 ;
        RECT 115.025 44.460 115.540 44.600 ;
        RECT 87.175 44.415 87.465 44.460 ;
        RECT 90.840 44.400 91.160 44.460 ;
        RECT 94.060 44.400 94.380 44.460 ;
        RECT 100.500 44.400 100.820 44.460 ;
        RECT 107.950 44.305 108.090 44.460 ;
        RECT 115.220 44.400 115.540 44.460 ;
        RECT 39.780 44.120 64.850 44.260 ;
        RECT 65.170 44.120 80.030 44.260 ;
        RECT 107.875 44.260 108.165 44.305 ;
        RECT 117.075 44.260 117.365 44.305 ;
        RECT 118.440 44.260 118.760 44.320 ;
        RECT 107.875 44.120 118.760 44.260 ;
        RECT 118.990 44.260 119.130 44.800 ;
        RECT 123.130 44.800 123.820 44.940 ;
        RECT 123.130 44.645 123.270 44.800 ;
        RECT 123.500 44.740 123.820 44.800 ;
        RECT 127.640 44.940 127.960 45.000 ;
        RECT 128.575 44.940 128.865 44.985 ;
        RECT 127.640 44.800 128.865 44.940 ;
        RECT 127.640 44.740 127.960 44.800 ;
        RECT 128.575 44.755 128.865 44.800 ;
        RECT 123.055 44.415 123.345 44.645 ;
        RECT 135.920 44.600 136.240 44.660 ;
        RECT 136.840 44.600 137.160 44.660 ;
        RECT 123.590 44.460 136.240 44.600 ;
        RECT 136.645 44.460 137.160 44.600 ;
        RECT 123.590 44.260 123.730 44.460 ;
        RECT 135.920 44.400 136.240 44.460 ;
        RECT 136.840 44.400 137.160 44.460 ;
        RECT 137.300 44.600 137.620 44.660 ;
        RECT 148.890 44.645 149.030 45.140 ;
        RECT 150.195 45.140 186.380 45.280 ;
        RECT 150.195 45.095 150.485 45.140 ;
        RECT 186.060 45.080 186.380 45.140 ;
        RECT 191.120 45.280 191.440 45.340 ;
        RECT 192.975 45.280 193.265 45.325 ;
        RECT 191.120 45.140 193.265 45.280 ;
        RECT 191.120 45.080 191.440 45.140 ;
        RECT 192.975 45.095 193.265 45.140 ;
        RECT 216.420 45.280 216.740 45.340 ;
        RECT 222.875 45.280 223.165 45.325 ;
        RECT 216.420 45.140 223.165 45.280 ;
        RECT 216.420 45.080 216.740 45.140 ;
        RECT 222.875 45.095 223.165 45.140 ;
        RECT 226.080 45.280 226.400 45.340 ;
        RECT 232.060 45.280 232.380 45.340 ;
        RECT 237.135 45.280 237.425 45.325 ;
        RECT 258.295 45.280 258.585 45.325 ;
        RECT 226.080 45.140 229.530 45.280 ;
        RECT 226.080 45.080 226.400 45.140 ;
        RECT 158.020 44.940 158.310 44.985 ;
        RECT 159.420 44.940 159.710 44.985 ;
        RECT 161.260 44.940 161.550 44.985 ;
        RECT 158.020 44.800 161.550 44.940 ;
        RECT 158.020 44.755 158.310 44.800 ;
        RECT 159.420 44.755 159.710 44.800 ;
        RECT 161.260 44.755 161.550 44.800 ;
        RECT 162.600 44.940 162.920 45.000 ;
        RECT 172.260 44.940 172.580 45.000 ;
        RECT 185.140 44.940 185.460 45.000 ;
        RECT 162.600 44.800 185.460 44.940 ;
        RECT 162.600 44.740 162.920 44.800 ;
        RECT 172.260 44.740 172.580 44.800 ;
        RECT 185.140 44.740 185.460 44.800 ;
        RECT 187.000 44.940 187.290 44.985 ;
        RECT 188.400 44.940 188.690 44.985 ;
        RECT 190.240 44.940 190.530 44.985 ;
        RECT 209.980 44.940 210.300 45.000 ;
        RECT 219.180 44.940 219.500 45.000 ;
        RECT 187.000 44.800 190.530 44.940 ;
        RECT 187.000 44.755 187.290 44.800 ;
        RECT 188.400 44.755 188.690 44.800 ;
        RECT 190.240 44.755 190.530 44.800 ;
        RECT 206.390 44.800 210.300 44.940 ;
        RECT 143.295 44.600 143.585 44.645 ;
        RECT 137.300 44.460 143.585 44.600 ;
        RECT 137.300 44.400 137.620 44.460 ;
        RECT 143.295 44.415 143.585 44.460 ;
        RECT 148.815 44.415 149.105 44.645 ;
        RECT 151.115 44.415 151.405 44.645 ;
        RECT 153.860 44.600 154.180 44.660 ;
        RECT 157.095 44.600 157.385 44.645 ;
        RECT 174.560 44.600 174.880 44.660 ;
        RECT 177.335 44.600 177.625 44.645 ;
        RECT 178.240 44.600 178.560 44.660 ;
        RECT 153.860 44.460 157.385 44.600 ;
        RECT 174.365 44.460 177.625 44.600 ;
        RECT 178.045 44.460 178.560 44.600 ;
        RECT 118.990 44.120 123.730 44.260 ;
        RECT 129.020 44.305 129.340 44.320 ;
        RECT 39.780 44.060 40.100 44.120 ;
        RECT 62.780 43.920 63.100 43.980 ;
        RECT 65.170 43.920 65.310 44.120 ;
        RECT 107.875 44.075 108.165 44.120 ;
        RECT 117.075 44.075 117.365 44.120 ;
        RECT 118.440 44.060 118.760 44.120 ;
        RECT 129.020 44.075 129.600 44.305 ;
        RECT 130.415 44.260 130.705 44.305 ;
        RECT 151.190 44.260 151.330 44.415 ;
        RECT 153.860 44.400 154.180 44.460 ;
        RECT 157.095 44.415 157.385 44.460 ;
        RECT 174.560 44.400 174.880 44.460 ;
        RECT 177.335 44.415 177.625 44.460 ;
        RECT 178.240 44.400 178.560 44.460 ;
        RECT 184.680 44.600 185.000 44.660 ;
        RECT 186.075 44.600 186.365 44.645 ;
        RECT 184.680 44.460 186.365 44.600 ;
        RECT 184.680 44.400 185.000 44.460 ;
        RECT 186.075 44.415 186.365 44.460 ;
        RECT 187.455 44.600 187.745 44.645 ;
        RECT 205.840 44.600 206.160 44.660 ;
        RECT 206.390 44.645 206.530 44.800 ;
        RECT 209.980 44.740 210.300 44.800 ;
        RECT 214.670 44.800 219.500 44.940 ;
        RECT 229.390 44.940 229.530 45.140 ;
        RECT 232.060 45.140 237.425 45.280 ;
        RECT 232.060 45.080 232.380 45.140 ;
        RECT 237.135 45.095 237.425 45.140 ;
        RECT 238.590 45.140 258.585 45.280 ;
        RECT 238.590 44.940 238.730 45.140 ;
        RECT 258.295 45.095 258.585 45.140 ;
        RECT 259.200 45.280 259.520 45.340 ;
        RECT 277.155 45.280 277.445 45.325 ;
        RECT 293.700 45.280 294.020 45.340 ;
        RECT 259.200 45.140 277.445 45.280 ;
        RECT 259.200 45.080 259.520 45.140 ;
        RECT 277.155 45.095 277.445 45.140 ;
        RECT 278.150 45.140 294.020 45.280 ;
        RECT 229.390 44.800 238.730 44.940 ;
        RECT 240.800 44.940 241.120 45.000 ;
        RECT 247.240 44.940 247.560 45.000 ;
        RECT 249.555 44.940 249.845 44.985 ;
        RECT 256.915 44.940 257.205 44.985 ;
        RECT 240.800 44.800 244.250 44.940 ;
        RECT 187.455 44.460 206.160 44.600 ;
        RECT 187.455 44.415 187.745 44.460 ;
        RECT 205.840 44.400 206.160 44.460 ;
        RECT 206.315 44.415 206.605 44.645 ;
        RECT 208.140 44.600 208.460 44.660 ;
        RECT 214.670 44.645 214.810 44.800 ;
        RECT 219.180 44.740 219.500 44.800 ;
        RECT 240.800 44.740 241.120 44.800 ;
        RECT 207.945 44.460 208.460 44.600 ;
        RECT 208.140 44.400 208.460 44.460 ;
        RECT 214.595 44.415 214.885 44.645 ;
        RECT 215.040 44.600 215.360 44.660 ;
        RECT 215.720 44.600 216.010 44.645 ;
        RECT 216.420 44.600 216.740 44.660 ;
        RECT 215.040 44.460 215.555 44.600 ;
        RECT 215.720 44.460 216.740 44.600 ;
        RECT 215.040 44.400 215.360 44.460 ;
        RECT 215.720 44.415 216.010 44.460 ;
        RECT 216.420 44.400 216.740 44.460 ;
        RECT 217.815 44.600 218.105 44.645 ;
        RECT 221.020 44.600 221.340 44.660 ;
        RECT 217.815 44.460 221.340 44.600 ;
        RECT 217.815 44.415 218.105 44.460 ;
        RECT 221.020 44.400 221.340 44.460 ;
        RECT 221.480 44.600 221.800 44.660 ;
        RECT 221.985 44.600 222.275 44.645 ;
        RECT 228.380 44.600 228.700 44.660 ;
        RECT 229.760 44.600 230.080 44.660 ;
        RECT 221.480 44.460 222.275 44.600 ;
        RECT 228.185 44.460 228.700 44.600 ;
        RECT 229.565 44.460 230.080 44.600 ;
        RECT 221.480 44.400 221.800 44.460 ;
        RECT 221.985 44.415 222.275 44.460 ;
        RECT 228.380 44.400 228.700 44.460 ;
        RECT 229.760 44.400 230.080 44.460 ;
        RECT 235.740 44.600 236.060 44.660 ;
        RECT 236.215 44.600 236.505 44.645 ;
        RECT 235.740 44.460 236.505 44.600 ;
        RECT 235.740 44.400 236.060 44.460 ;
        RECT 236.215 44.415 236.505 44.460 ;
        RECT 238.960 44.600 239.280 44.660 ;
        RECT 242.655 44.600 242.945 44.645 ;
        RECT 243.560 44.600 243.880 44.660 ;
        RECT 238.960 44.460 242.945 44.600 ;
        RECT 243.365 44.460 243.880 44.600 ;
        RECT 244.110 44.600 244.250 44.800 ;
        RECT 247.240 44.800 249.845 44.940 ;
        RECT 247.240 44.740 247.560 44.800 ;
        RECT 249.555 44.755 249.845 44.800 ;
        RECT 250.090 44.800 257.205 44.940 ;
        RECT 250.090 44.600 250.230 44.800 ;
        RECT 256.915 44.755 257.205 44.800 ;
        RECT 244.110 44.460 250.230 44.600 ;
        RECT 238.960 44.400 239.280 44.460 ;
        RECT 242.655 44.415 242.945 44.460 ;
        RECT 243.560 44.400 243.880 44.460 ;
        RECT 250.475 44.415 250.765 44.645 ;
        RECT 257.820 44.600 258.140 44.660 ;
        RECT 257.625 44.460 258.140 44.600 ;
        RECT 156.160 44.260 156.480 44.320 ;
        RECT 130.415 44.120 137.070 44.260 ;
        RECT 130.415 44.075 130.705 44.120 ;
        RECT 129.020 44.060 129.340 44.075 ;
        RECT 136.930 43.980 137.070 44.120 ;
        RECT 137.850 44.120 156.480 44.260 ;
        RECT 115.925 43.920 116.215 43.965 ;
        RECT 119.360 43.920 119.680 43.980 ;
        RECT 129.955 43.920 130.245 43.965 ;
        RECT 62.780 43.780 65.310 43.920 ;
        RECT 106.800 43.780 119.680 43.920 ;
        RECT 62.780 43.720 63.100 43.780 ;
        RECT 85.320 43.580 85.640 43.640 ;
        RECT 106.800 43.625 106.940 43.780 ;
        RECT 115.925 43.735 116.215 43.780 ;
        RECT 119.360 43.720 119.680 43.780 ;
        RECT 120.370 43.780 132.440 43.920 ;
        RECT 120.370 43.640 120.510 43.780 ;
        RECT 129.955 43.735 130.245 43.780 ;
        RECT 106.725 43.580 107.015 43.625 ;
        RECT 85.320 43.440 107.015 43.580 ;
        RECT 85.320 43.380 85.640 43.440 ;
        RECT 106.725 43.395 107.015 43.440 ;
        RECT 107.415 43.580 107.705 43.625 ;
        RECT 116.615 43.580 116.905 43.625 ;
        RECT 120.280 43.580 120.600 43.640 ;
        RECT 123.500 43.580 123.820 43.640 ;
        RECT 131.780 43.580 132.100 43.640 ;
        RECT 107.415 43.440 120.600 43.580 ;
        RECT 123.305 43.440 123.820 43.580 ;
        RECT 131.585 43.440 132.100 43.580 ;
        RECT 132.300 43.580 132.440 43.780 ;
        RECT 136.840 43.720 137.160 43.980 ;
        RECT 137.850 43.965 137.990 44.120 ;
        RECT 156.160 44.060 156.480 44.120 ;
        RECT 158.475 44.260 158.765 44.305 ;
        RECT 174.100 44.260 174.420 44.320 ;
        RECT 158.475 44.120 169.270 44.260 ;
        RECT 173.905 44.120 174.420 44.260 ;
        RECT 158.475 44.075 158.765 44.120 ;
        RECT 137.775 43.735 138.065 43.965 ;
        RECT 156.620 43.920 156.940 43.980 ;
        RECT 138.310 43.780 156.940 43.920 ;
        RECT 138.310 43.580 138.450 43.780 ;
        RECT 156.620 43.720 156.940 43.780 ;
        RECT 157.560 43.920 157.850 43.965 ;
        RECT 159.880 43.920 160.170 43.965 ;
        RECT 161.260 43.920 161.550 43.965 ;
        RECT 157.560 43.780 161.550 43.920 ;
        RECT 169.130 43.920 169.270 44.120 ;
        RECT 174.100 44.060 174.420 44.120 ;
        RECT 175.960 44.260 176.250 44.305 ;
        RECT 178.740 44.260 179.030 44.305 ;
        RECT 175.960 44.120 179.030 44.260 ;
        RECT 175.960 44.075 176.250 44.120 ;
        RECT 178.740 44.075 179.030 44.120 ;
        RECT 179.620 44.260 179.940 44.320 ;
        RECT 204.015 44.260 204.305 44.305 ;
        RECT 179.620 44.120 204.305 44.260 ;
        RECT 179.620 44.060 179.940 44.120 ;
        RECT 204.015 44.075 204.305 44.120 ;
        RECT 207.680 44.260 208.000 44.320 ;
        RECT 208.615 44.260 208.905 44.305 ;
        RECT 230.680 44.260 231.000 44.320 ;
        RECT 207.680 44.120 208.905 44.260 ;
        RECT 230.485 44.120 231.000 44.260 ;
        RECT 207.680 44.060 208.000 44.120 ;
        RECT 208.615 44.075 208.905 44.120 ;
        RECT 230.680 44.060 231.000 44.120 ;
        RECT 232.980 44.260 233.300 44.320 ;
        RECT 243.650 44.260 243.790 44.400 ;
        RECT 232.980 44.120 243.790 44.260 ;
        RECT 232.980 44.060 233.300 44.120 ;
        RECT 245.415 44.075 245.705 44.305 ;
        RECT 250.550 44.260 250.690 44.415 ;
        RECT 257.820 44.400 258.140 44.460 ;
        RECT 258.740 44.600 259.060 44.660 ;
        RECT 263.815 44.600 264.105 44.645 ;
        RECT 258.740 44.460 264.105 44.600 ;
        RECT 258.740 44.400 259.060 44.460 ;
        RECT 263.815 44.415 264.105 44.460 ;
        RECT 270.700 44.600 271.020 44.660 ;
        RECT 278.150 44.645 278.290 45.140 ;
        RECT 293.700 45.080 294.020 45.140 ;
        RECT 294.175 45.280 294.465 45.325 ;
        RECT 297.840 45.280 298.160 45.340 ;
        RECT 294.175 45.140 298.160 45.280 ;
        RECT 294.175 45.095 294.465 45.140 ;
        RECT 292.320 44.940 292.640 45.000 ;
        RECT 286.890 44.800 292.640 44.940 ;
        RECT 271.175 44.600 271.465 44.645 ;
        RECT 270.700 44.460 271.465 44.600 ;
        RECT 270.700 44.400 271.020 44.460 ;
        RECT 271.175 44.415 271.465 44.460 ;
        RECT 278.075 44.415 278.365 44.645 ;
        RECT 278.995 44.415 279.285 44.645 ;
        RECT 279.440 44.600 279.760 44.660 ;
        RECT 286.890 44.645 287.030 44.800 ;
        RECT 292.320 44.740 292.640 44.800 ;
        RECT 292.780 44.940 293.100 45.000 ;
        RECT 294.250 44.940 294.390 45.095 ;
        RECT 297.840 45.080 298.160 45.140 ;
        RECT 299.220 45.280 299.540 45.340 ;
        RECT 305.200 45.280 305.520 45.340 ;
        RECT 299.220 45.140 305.520 45.280 ;
        RECT 299.220 45.080 299.540 45.140 ;
        RECT 305.200 45.080 305.520 45.140 ;
        RECT 305.660 45.280 305.980 45.340 ;
        RECT 328.675 45.280 328.965 45.325 ;
        RECT 357.180 45.280 357.500 45.340 ;
        RECT 305.660 45.140 328.965 45.280 ;
        RECT 356.985 45.140 357.500 45.280 ;
        RECT 305.660 45.080 305.980 45.140 ;
        RECT 328.675 45.095 328.965 45.140 ;
        RECT 357.180 45.080 357.500 45.140 ;
        RECT 358.100 45.280 358.420 45.340 ;
        RECT 371.455 45.280 371.745 45.325 ;
        RECT 358.100 45.140 371.745 45.280 ;
        RECT 358.100 45.080 358.420 45.140 ;
        RECT 371.455 45.095 371.745 45.140 ;
        RECT 312.560 44.940 312.880 45.000 ;
        RECT 326.360 44.940 326.680 45.000 ;
        RECT 292.780 44.800 294.390 44.940 ;
        RECT 301.150 44.800 312.880 44.940 ;
        RECT 292.780 44.740 293.100 44.800 ;
        RECT 288.640 44.645 288.960 44.660 ;
        RECT 279.440 44.460 284.730 44.600 ;
        RECT 267.940 44.260 268.260 44.320 ;
        RECT 275.760 44.260 276.080 44.320 ;
        RECT 279.070 44.260 279.210 44.415 ;
        RECT 279.440 44.400 279.760 44.460 ;
        RECT 250.550 44.120 268.260 44.260 ;
        RECT 179.175 43.920 179.465 43.965 ;
        RECT 169.130 43.780 179.465 43.920 ;
        RECT 157.560 43.735 157.850 43.780 ;
        RECT 159.880 43.735 160.170 43.780 ;
        RECT 161.260 43.735 161.550 43.780 ;
        RECT 179.175 43.735 179.465 43.780 ;
        RECT 186.540 43.920 186.830 43.965 ;
        RECT 188.860 43.920 189.150 43.965 ;
        RECT 190.240 43.920 190.530 43.965 ;
        RECT 186.540 43.780 190.530 43.920 ;
        RECT 186.540 43.735 186.830 43.780 ;
        RECT 188.860 43.735 189.150 43.780 ;
        RECT 190.240 43.735 190.530 43.780 ;
        RECT 213.660 43.920 213.980 43.980 ;
        RECT 228.855 43.920 229.145 43.965 ;
        RECT 232.520 43.920 232.840 43.980 ;
        RECT 213.660 43.780 232.840 43.920 ;
        RECT 213.660 43.720 213.980 43.780 ;
        RECT 228.855 43.735 229.145 43.780 ;
        RECT 232.520 43.720 232.840 43.780 ;
        RECT 237.580 43.920 237.900 43.980 ;
        RECT 244.940 43.920 245.260 43.980 ;
        RECT 237.580 43.780 245.260 43.920 ;
        RECT 245.490 43.920 245.630 44.075 ;
        RECT 267.940 44.060 268.260 44.120 ;
        RECT 272.170 44.120 279.210 44.260 ;
        RECT 284.590 44.260 284.730 44.460 ;
        RECT 286.815 44.415 287.105 44.645 ;
        RECT 288.425 44.415 288.960 44.645 ;
        RECT 293.255 44.600 293.545 44.645 ;
        RECT 298.760 44.600 299.080 44.660 ;
        RECT 301.150 44.645 301.290 44.800 ;
        RECT 312.560 44.740 312.880 44.800 ;
        RECT 313.110 44.800 321.990 44.940 ;
        RECT 288.640 44.400 288.960 44.415 ;
        RECT 292.870 44.460 299.080 44.600 ;
        RECT 292.870 44.320 293.010 44.460 ;
        RECT 293.255 44.415 293.545 44.460 ;
        RECT 298.760 44.400 299.080 44.460 ;
        RECT 301.075 44.415 301.365 44.645 ;
        RECT 302.455 44.600 302.745 44.645 ;
        RECT 306.120 44.600 306.440 44.660 ;
        RECT 302.455 44.460 306.440 44.600 ;
        RECT 302.455 44.415 302.745 44.460 ;
        RECT 306.120 44.400 306.440 44.460 ;
        RECT 307.515 44.600 307.805 44.645 ;
        RECT 313.110 44.600 313.250 44.800 ;
        RECT 321.850 44.645 321.990 44.800 ;
        RECT 326.360 44.800 373.510 44.940 ;
        RECT 326.360 44.740 326.680 44.800 ;
        RECT 330.590 44.645 330.730 44.800 ;
        RECT 307.515 44.460 313.250 44.600 ;
        RECT 307.515 44.415 307.805 44.460 ;
        RECT 315.335 44.415 315.625 44.645 ;
        RECT 316.715 44.415 317.005 44.645 ;
        RECT 321.775 44.415 322.065 44.645 ;
        RECT 329.595 44.415 329.885 44.645 ;
        RECT 330.515 44.415 330.805 44.645 ;
        RECT 336.035 44.600 336.325 44.645 ;
        RECT 336.480 44.600 336.800 44.660 ;
        RECT 345.220 44.600 345.540 44.660 ;
        RECT 347.995 44.600 348.285 44.645 ;
        RECT 336.035 44.460 336.800 44.600 ;
        RECT 344.785 44.460 348.285 44.600 ;
        RECT 336.035 44.415 336.325 44.460 ;
        RECT 287.735 44.260 288.025 44.305 ;
        RECT 284.590 44.120 288.025 44.260 ;
        RECT 258.280 43.920 258.600 43.980 ;
        RECT 272.170 43.965 272.310 44.120 ;
        RECT 275.760 44.060 276.080 44.120 ;
        RECT 245.490 43.780 258.600 43.920 ;
        RECT 237.580 43.720 237.900 43.780 ;
        RECT 244.940 43.720 245.260 43.780 ;
        RECT 258.280 43.720 258.600 43.780 ;
        RECT 272.095 43.735 272.385 43.965 ;
        RECT 279.070 43.920 279.210 44.120 ;
        RECT 287.735 44.075 288.025 44.120 ;
        RECT 292.780 44.060 293.100 44.320 ;
        RECT 298.300 44.260 298.620 44.320 ;
        RECT 301.980 44.260 302.300 44.320 ;
        RECT 298.300 44.120 300.370 44.260 ;
        RECT 301.785 44.120 302.300 44.260 ;
        RECT 298.300 44.060 298.620 44.120 ;
        RECT 300.230 43.920 300.370 44.120 ;
        RECT 301.980 44.060 302.300 44.120 ;
        RECT 307.590 43.920 307.730 44.415 ;
        RECT 313.480 43.920 313.800 43.980 ;
        RECT 279.070 43.780 293.010 43.920 ;
        RECT 300.230 43.780 307.730 43.920 ;
        RECT 308.510 43.780 313.800 43.920 ;
        RECT 315.410 43.920 315.550 44.415 ;
        RECT 315.780 44.260 316.100 44.320 ;
        RECT 316.255 44.260 316.545 44.305 ;
        RECT 315.780 44.120 316.545 44.260 ;
        RECT 316.790 44.260 316.930 44.415 ;
        RECT 316.790 44.120 322.910 44.260 ;
        RECT 315.780 44.060 316.100 44.120 ;
        RECT 316.255 44.075 316.545 44.120 ;
        RECT 319.920 43.920 320.240 43.980 ;
        RECT 315.410 43.780 320.240 43.920 ;
        RECT 132.300 43.440 138.450 43.580 ;
        RECT 144.215 43.580 144.505 43.625 ;
        RECT 163.060 43.580 163.380 43.640 ;
        RECT 163.980 43.580 164.300 43.640 ;
        RECT 144.215 43.440 163.380 43.580 ;
        RECT 163.785 43.440 164.300 43.580 ;
        RECT 107.415 43.395 107.705 43.440 ;
        RECT 116.615 43.395 116.905 43.440 ;
        RECT 120.280 43.380 120.600 43.440 ;
        RECT 123.500 43.380 123.820 43.440 ;
        RECT 131.780 43.380 132.100 43.440 ;
        RECT 144.215 43.395 144.505 43.440 ;
        RECT 163.060 43.380 163.380 43.440 ;
        RECT 163.980 43.380 164.300 43.440 ;
        RECT 216.420 43.580 216.740 43.640 ;
        RECT 221.940 43.580 222.260 43.640 ;
        RECT 216.420 43.440 222.260 43.580 ;
        RECT 216.420 43.380 216.740 43.440 ;
        RECT 221.940 43.380 222.260 43.440 ;
        RECT 236.660 43.580 236.980 43.640 ;
        RECT 250.935 43.580 251.225 43.625 ;
        RECT 264.720 43.580 265.040 43.640 ;
        RECT 236.660 43.440 251.225 43.580 ;
        RECT 264.525 43.440 265.040 43.580 ;
        RECT 292.870 43.580 293.010 43.780 ;
        RECT 308.510 43.640 308.650 43.780 ;
        RECT 313.480 43.720 313.800 43.780 ;
        RECT 319.920 43.720 320.240 43.780 ;
        RECT 298.300 43.580 298.620 43.640 ;
        RECT 308.420 43.580 308.740 43.640 ;
        RECT 292.870 43.440 298.620 43.580 ;
        RECT 308.225 43.440 308.740 43.580 ;
        RECT 236.660 43.380 236.980 43.440 ;
        RECT 250.935 43.395 251.225 43.440 ;
        RECT 264.720 43.380 265.040 43.440 ;
        RECT 298.300 43.380 298.620 43.440 ;
        RECT 308.420 43.380 308.740 43.440 ;
        RECT 309.800 43.580 310.120 43.640 ;
        RECT 317.620 43.580 317.940 43.640 ;
        RECT 322.770 43.625 322.910 44.120 ;
        RECT 329.670 43.920 329.810 44.415 ;
        RECT 336.480 44.400 336.800 44.460 ;
        RECT 345.220 44.400 345.540 44.460 ;
        RECT 347.995 44.415 348.285 44.460 ;
        RECT 348.915 44.415 349.205 44.645 ;
        RECT 350.755 44.415 351.045 44.645 ;
        RECT 351.675 44.600 351.965 44.645 ;
        RECT 352.120 44.600 352.440 44.660 ;
        RECT 358.100 44.600 358.420 44.660 ;
        RECT 351.675 44.460 352.440 44.600 ;
        RECT 357.905 44.460 358.420 44.600 ;
        RECT 351.675 44.415 351.965 44.460 ;
        RECT 342.920 44.260 343.240 44.320 ;
        RECT 345.695 44.260 345.985 44.305 ;
        RECT 342.920 44.120 345.985 44.260 ;
        RECT 342.920 44.060 343.240 44.120 ;
        RECT 345.695 44.075 345.985 44.120 ;
        RECT 338.320 43.920 338.640 43.980 ;
        RECT 329.670 43.780 338.640 43.920 ;
        RECT 348.990 43.920 349.130 44.415 ;
        RECT 350.830 44.260 350.970 44.415 ;
        RECT 352.120 44.400 352.440 44.460 ;
        RECT 358.100 44.400 358.420 44.460 ;
        RECT 358.560 44.600 358.880 44.660 ;
        RECT 373.370 44.645 373.510 44.800 ;
        RECT 359.035 44.600 359.325 44.645 ;
        RECT 358.560 44.460 359.325 44.600 ;
        RECT 358.560 44.400 358.880 44.460 ;
        RECT 359.035 44.415 359.325 44.460 ;
        RECT 364.555 44.600 364.845 44.645 ;
        RECT 364.555 44.460 365.690 44.600 ;
        RECT 364.555 44.415 364.845 44.460 ;
        RECT 365.550 44.260 365.690 44.460 ;
        RECT 372.375 44.415 372.665 44.645 ;
        RECT 373.295 44.415 373.585 44.645 ;
        RECT 381.100 44.600 381.420 44.660 ;
        RECT 386.160 44.600 386.480 44.660 ;
        RECT 373.830 44.460 381.420 44.600 ;
        RECT 385.965 44.460 386.480 44.600 ;
        RECT 350.830 44.120 365.690 44.260 ;
        RECT 372.450 44.260 372.590 44.415 ;
        RECT 373.830 44.260 373.970 44.460 ;
        RECT 381.100 44.400 381.420 44.460 ;
        RECT 386.160 44.400 386.480 44.460 ;
        RECT 372.450 44.120 373.970 44.260 ;
        RECT 365.015 43.920 365.305 43.965 ;
        RECT 348.990 43.780 365.305 43.920 ;
        RECT 365.550 43.920 365.690 44.120 ;
        RECT 381.100 43.920 381.420 43.980 ;
        RECT 391.235 43.920 391.525 43.965 ;
        RECT 365.550 43.780 380.410 43.920 ;
        RECT 338.320 43.720 338.640 43.780 ;
        RECT 365.015 43.735 365.305 43.780 ;
        RECT 309.800 43.440 317.940 43.580 ;
        RECT 309.800 43.380 310.120 43.440 ;
        RECT 317.620 43.380 317.940 43.440 ;
        RECT 322.695 43.580 322.985 43.625 ;
        RECT 333.260 43.580 333.580 43.640 ;
        RECT 336.940 43.580 337.260 43.640 ;
        RECT 322.695 43.440 333.580 43.580 ;
        RECT 336.745 43.440 337.260 43.580 ;
        RECT 322.695 43.395 322.985 43.440 ;
        RECT 333.260 43.380 333.580 43.440 ;
        RECT 336.940 43.380 337.260 43.440 ;
        RECT 358.100 43.580 358.420 43.640 ;
        RECT 371.440 43.580 371.760 43.640 ;
        RECT 379.720 43.580 380.040 43.640 ;
        RECT 358.100 43.440 371.760 43.580 ;
        RECT 379.525 43.440 380.040 43.580 ;
        RECT 380.270 43.580 380.410 43.780 ;
        RECT 381.100 43.780 391.525 43.920 ;
        RECT 381.100 43.720 381.420 43.780 ;
        RECT 391.235 43.735 391.525 43.780 ;
        RECT 404.560 43.580 404.880 43.640 ;
        RECT 502.540 43.580 502.860 43.640 ;
        RECT 586.720 43.580 587.040 43.640 ;
        RECT 380.270 43.440 404.880 43.580 ;
        RECT 502.345 43.440 502.860 43.580 ;
        RECT 586.525 43.440 587.040 43.580 ;
        RECT 358.100 43.380 358.420 43.440 ;
        RECT 371.440 43.380 371.760 43.440 ;
        RECT 379.720 43.380 380.040 43.440 ;
        RECT 404.560 43.380 404.880 43.440 ;
        RECT 502.540 43.380 502.860 43.440 ;
        RECT 586.720 43.380 587.040 43.440 ;
        RECT 42.470 42.760 631.270 43.240 ;
        RECT 77.500 42.560 77.820 42.620 ;
        RECT 115.220 42.560 115.540 42.620 ;
        RECT 77.500 42.420 115.540 42.560 ;
        RECT 77.500 42.360 77.820 42.420 ;
        RECT 115.220 42.360 115.540 42.420 ;
        RECT 117.520 42.560 117.840 42.620 ;
        RECT 156.620 42.560 156.940 42.620 ;
        RECT 213.660 42.560 213.980 42.620 ;
        RECT 215.040 42.560 215.360 42.620 ;
        RECT 221.480 42.560 221.800 42.620 ;
        RECT 117.520 42.420 156.390 42.560 ;
        RECT 117.520 42.360 117.840 42.420 ;
        RECT 84.860 42.220 85.180 42.280 ;
        RECT 137.300 42.220 137.620 42.280 ;
        RECT 84.860 42.080 137.620 42.220 ;
        RECT 84.860 42.020 85.180 42.080 ;
        RECT 137.300 42.020 137.620 42.080 ;
        RECT 137.760 42.220 138.080 42.280 ;
        RECT 155.715 42.220 156.005 42.265 ;
        RECT 137.760 42.080 156.005 42.220 ;
        RECT 156.250 42.220 156.390 42.420 ;
        RECT 156.620 42.420 213.980 42.560 ;
        RECT 214.845 42.420 215.360 42.560 ;
        RECT 221.285 42.420 221.800 42.560 ;
        RECT 156.620 42.360 156.940 42.420 ;
        RECT 213.660 42.360 213.980 42.420 ;
        RECT 215.040 42.360 215.360 42.420 ;
        RECT 221.480 42.360 221.800 42.420 ;
        RECT 221.940 42.560 222.260 42.620 ;
        RECT 237.120 42.560 237.440 42.620 ;
        RECT 221.940 42.420 237.440 42.560 ;
        RECT 221.940 42.360 222.260 42.420 ;
        RECT 237.120 42.360 237.440 42.420 ;
        RECT 243.560 42.560 243.880 42.620 ;
        RECT 282.200 42.560 282.520 42.620 ;
        RECT 336.940 42.560 337.260 42.620 ;
        RECT 357.180 42.560 357.500 42.620 ;
        RECT 243.560 42.420 281.970 42.560 ;
        RECT 243.560 42.360 243.880 42.420 ;
        RECT 178.240 42.220 178.560 42.280 ;
        RECT 156.250 42.080 178.560 42.220 ;
        RECT 137.760 42.020 138.080 42.080 ;
        RECT 155.715 42.035 156.005 42.080 ;
        RECT 178.240 42.020 178.560 42.080 ;
        RECT 224.715 42.220 225.005 42.265 ;
        RECT 232.980 42.220 233.300 42.280 ;
        RECT 224.715 42.080 233.300 42.220 ;
        RECT 281.830 42.220 281.970 42.420 ;
        RECT 282.200 42.420 337.260 42.560 ;
        RECT 282.200 42.360 282.520 42.420 ;
        RECT 336.940 42.360 337.260 42.420 ;
        RECT 337.490 42.420 357.500 42.560 ;
        RECT 287.260 42.220 287.580 42.280 ;
        RECT 281.830 42.080 287.580 42.220 ;
        RECT 224.715 42.035 225.005 42.080 ;
        RECT 232.980 42.020 233.300 42.080 ;
        RECT 287.260 42.020 287.580 42.080 ;
        RECT 289.560 42.220 289.880 42.280 ;
        RECT 301.060 42.220 301.380 42.280 ;
        RECT 289.560 42.080 301.380 42.220 ;
        RECT 289.560 42.020 289.880 42.080 ;
        RECT 301.060 42.020 301.380 42.080 ;
        RECT 329.580 42.220 329.900 42.280 ;
        RECT 337.490 42.220 337.630 42.420 ;
        RECT 357.180 42.360 357.500 42.420 ;
        RECT 329.580 42.080 337.630 42.220 ;
        RECT 352.120 42.220 352.440 42.280 ;
        RECT 402.260 42.220 402.580 42.280 ;
        RECT 352.120 42.080 402.580 42.220 ;
        RECT 329.580 42.020 329.900 42.080 ;
        RECT 352.120 42.020 352.440 42.080 ;
        RECT 402.260 42.020 402.580 42.080 ;
        RECT 86.240 41.880 86.560 41.940 ;
        RECT 163.075 41.880 163.365 41.925 ;
        RECT 86.240 41.740 163.365 41.880 ;
        RECT 86.240 41.680 86.560 41.740 ;
        RECT 163.075 41.695 163.365 41.740 ;
        RECT 164.440 41.880 164.760 41.940 ;
        RECT 175.035 41.880 175.325 41.925 ;
        RECT 164.440 41.740 175.325 41.880 ;
        RECT 164.440 41.680 164.760 41.740 ;
        RECT 175.035 41.695 175.325 41.740 ;
        RECT 201.240 41.880 201.560 41.940 ;
        RECT 223.795 41.880 224.085 41.925 ;
        RECT 201.240 41.740 224.085 41.880 ;
        RECT 201.240 41.680 201.560 41.740 ;
        RECT 223.795 41.695 224.085 41.740 ;
        RECT 224.255 41.880 224.545 41.925 ;
        RECT 264.720 41.880 265.040 41.940 ;
        RECT 224.255 41.740 265.040 41.880 ;
        RECT 224.255 41.695 224.545 41.740 ;
        RECT 264.720 41.680 265.040 41.740 ;
        RECT 273.920 41.880 274.240 41.940 ;
        RECT 301.980 41.880 302.300 41.940 ;
        RECT 273.920 41.740 302.300 41.880 ;
        RECT 273.920 41.680 274.240 41.740 ;
        RECT 301.980 41.680 302.300 41.740 ;
        RECT 344.300 41.880 344.620 41.940 ;
        RECT 379.720 41.880 380.040 41.940 ;
        RECT 344.300 41.740 380.040 41.880 ;
        RECT 344.300 41.680 344.620 41.740 ;
        RECT 379.720 41.680 380.040 41.740 ;
        RECT 37.480 41.540 37.800 41.600 ;
        RECT 345.220 41.540 345.540 41.600 ;
        RECT 37.480 41.400 345.540 41.540 ;
        RECT 37.480 41.340 37.800 41.400 ;
        RECT 345.220 41.340 345.540 41.400 ;
        RECT 87.160 41.200 87.480 41.260 ;
        RECT 175.480 41.200 175.800 41.260 ;
        RECT 87.160 41.060 175.800 41.200 ;
        RECT 87.160 41.000 87.480 41.060 ;
        RECT 175.480 41.000 175.800 41.060 ;
        RECT 208.140 41.200 208.460 41.260 ;
        RECT 223.335 41.200 223.625 41.245 ;
        RECT 208.140 41.060 223.625 41.200 ;
        RECT 208.140 41.000 208.460 41.060 ;
        RECT 223.335 41.015 223.625 41.060 ;
        RECT 239.880 41.200 240.200 41.260 ;
        RECT 342.920 41.200 343.240 41.260 ;
        RECT 239.880 41.060 343.240 41.200 ;
        RECT 239.880 41.000 240.200 41.060 ;
        RECT 342.920 41.000 343.240 41.060 ;
        RECT 118.440 40.860 118.760 40.920 ;
        RECT 136.840 40.860 137.160 40.920 ;
        RECT 118.440 40.720 137.160 40.860 ;
        RECT 118.440 40.660 118.760 40.720 ;
        RECT 136.840 40.660 137.160 40.720 ;
        RECT 143.740 40.860 144.060 40.920 ;
        RECT 154.780 40.860 155.100 40.920 ;
        RECT 143.740 40.720 155.100 40.860 ;
        RECT 143.740 40.660 144.060 40.720 ;
        RECT 154.780 40.660 155.100 40.720 ;
        RECT 155.715 40.860 156.005 40.905 ;
        RECT 162.600 40.860 162.920 40.920 ;
        RECT 155.715 40.720 162.920 40.860 ;
        RECT 155.715 40.675 156.005 40.720 ;
        RECT 162.600 40.660 162.920 40.720 ;
        RECT 163.060 40.860 163.380 40.920 ;
        RECT 258.295 40.860 258.585 40.905 ;
        RECT 163.060 40.720 258.585 40.860 ;
        RECT 163.060 40.660 163.380 40.720 ;
        RECT 258.295 40.675 258.585 40.720 ;
        RECT 280.360 40.860 280.680 40.920 ;
        RECT 315.780 40.860 316.100 40.920 ;
        RECT 280.360 40.720 316.100 40.860 ;
        RECT 280.360 40.660 280.680 40.720 ;
        RECT 315.780 40.660 316.100 40.720 ;
        RECT 336.480 40.860 336.800 40.920 ;
        RECT 358.100 40.860 358.420 40.920 ;
        RECT 336.480 40.720 358.420 40.860 ;
        RECT 336.480 40.660 336.800 40.720 ;
        RECT 358.100 40.660 358.420 40.720 ;
        RECT 111.540 40.520 111.860 40.580 ;
        RECT 230.680 40.520 231.000 40.580 ;
        RECT 111.540 40.380 231.000 40.520 ;
        RECT 111.540 40.320 111.860 40.380 ;
        RECT 230.680 40.320 231.000 40.380 ;
        RECT 244.940 40.520 245.260 40.580 ;
        RECT 308.420 40.520 308.740 40.580 ;
        RECT 244.940 40.380 308.740 40.520 ;
        RECT 244.940 40.320 245.260 40.380 ;
        RECT 308.420 40.320 308.740 40.380 ;
        RECT 311.180 40.520 311.500 40.580 ;
        RECT 323.600 40.520 323.920 40.580 ;
        RECT 311.180 40.380 323.920 40.520 ;
        RECT 311.180 40.320 311.500 40.380 ;
        RECT 323.600 40.320 323.920 40.380 ;
        RECT 329.120 40.520 329.440 40.580 ;
        RECT 369.140 40.520 369.460 40.580 ;
        RECT 329.120 40.380 369.460 40.520 ;
        RECT 329.120 40.320 329.440 40.380 ;
        RECT 369.140 40.320 369.460 40.380 ;
        RECT 123.500 40.180 123.820 40.240 ;
        RECT 169.040 40.180 169.360 40.240 ;
        RECT 123.500 40.040 169.360 40.180 ;
        RECT 123.500 39.980 123.820 40.040 ;
        RECT 169.040 39.980 169.360 40.040 ;
        RECT 174.100 40.180 174.420 40.240 ;
        RECT 220.560 40.180 220.880 40.240 ;
        RECT 174.100 40.040 220.880 40.180 ;
        RECT 174.100 39.980 174.420 40.040 ;
        RECT 220.560 39.980 220.880 40.040 ;
        RECT 228.380 40.180 228.700 40.240 ;
        RECT 285.420 40.180 285.740 40.240 ;
        RECT 228.380 40.040 285.740 40.180 ;
        RECT 228.380 39.980 228.700 40.040 ;
        RECT 285.420 39.980 285.740 40.040 ;
        RECT 341.080 40.180 341.400 40.240 ;
        RECT 372.820 40.180 373.140 40.240 ;
        RECT 341.080 40.040 373.140 40.180 ;
        RECT 341.080 39.980 341.400 40.040 ;
        RECT 372.820 39.980 373.140 40.040 ;
        RECT 88.540 39.840 88.860 39.900 ;
        RECT 130.400 39.840 130.720 39.900 ;
        RECT 88.540 39.700 130.720 39.840 ;
        RECT 88.540 39.640 88.860 39.700 ;
        RECT 130.400 39.640 130.720 39.700 ;
        RECT 131.780 39.840 132.100 39.900 ;
        RECT 155.700 39.840 156.020 39.900 ;
        RECT 131.780 39.700 156.020 39.840 ;
        RECT 131.780 39.640 132.100 39.700 ;
        RECT 155.700 39.640 156.020 39.700 ;
        RECT 163.075 39.840 163.365 39.885 ;
        RECT 179.160 39.840 179.480 39.900 ;
        RECT 163.075 39.700 179.480 39.840 ;
        RECT 163.075 39.655 163.365 39.700 ;
        RECT 179.160 39.640 179.480 39.700 ;
        RECT 230.680 39.840 231.000 39.900 ;
        RECT 255.060 39.840 255.380 39.900 ;
        RECT 230.680 39.700 255.380 39.840 ;
        RECT 230.680 39.640 231.000 39.700 ;
        RECT 255.060 39.640 255.380 39.700 ;
        RECT 258.295 39.840 258.585 39.885 ;
        RECT 270.700 39.840 271.020 39.900 ;
        RECT 292.780 39.840 293.100 39.900 ;
        RECT 258.295 39.700 293.100 39.840 ;
        RECT 258.295 39.655 258.585 39.700 ;
        RECT 270.700 39.640 271.020 39.700 ;
        RECT 292.780 39.640 293.100 39.700 ;
        RECT 293.240 39.840 293.560 39.900 ;
        RECT 303.820 39.840 304.140 39.900 ;
        RECT 293.240 39.700 304.140 39.840 ;
        RECT 293.240 39.640 293.560 39.700 ;
        RECT 303.820 39.640 304.140 39.700 ;
        RECT 332.800 39.840 333.120 39.900 ;
        RECT 342.000 39.840 342.320 39.900 ;
        RECT 332.800 39.700 342.320 39.840 ;
        RECT 332.800 39.640 333.120 39.700 ;
        RECT 342.000 39.640 342.320 39.700 ;
        RECT 117.060 39.500 117.380 39.560 ;
        RECT 117.980 39.500 118.300 39.560 ;
        RECT 163.980 39.500 164.300 39.560 ;
        RECT 117.060 39.360 164.300 39.500 ;
        RECT 117.060 39.300 117.380 39.360 ;
        RECT 117.980 39.300 118.300 39.360 ;
        RECT 163.980 39.300 164.300 39.360 ;
        RECT 165.360 39.500 165.680 39.560 ;
        RECT 221.495 39.500 221.785 39.545 ;
        RECT 165.360 39.360 221.785 39.500 ;
        RECT 165.360 39.300 165.680 39.360 ;
        RECT 221.495 39.315 221.785 39.360 ;
        RECT 238.040 39.500 238.360 39.560 ;
        RECT 245.860 39.500 246.180 39.560 ;
        RECT 238.040 39.360 246.180 39.500 ;
        RECT 238.040 39.300 238.360 39.360 ;
        RECT 245.860 39.300 246.180 39.360 ;
        RECT 256.440 39.500 256.760 39.560 ;
        RECT 276.680 39.500 277.000 39.560 ;
        RECT 256.440 39.360 277.000 39.500 ;
        RECT 256.440 39.300 256.760 39.360 ;
        RECT 276.680 39.300 277.000 39.360 ;
        RECT 281.740 39.500 282.060 39.560 ;
        RECT 299.220 39.500 299.540 39.560 ;
        RECT 281.740 39.360 299.540 39.500 ;
        RECT 281.740 39.300 282.060 39.360 ;
        RECT 299.220 39.300 299.540 39.360 ;
        RECT 106.020 39.160 106.340 39.220 ;
        RECT 126.720 39.160 127.040 39.220 ;
        RECT 106.020 39.020 127.040 39.160 ;
        RECT 106.020 38.960 106.340 39.020 ;
        RECT 126.720 38.960 127.040 39.020 ;
        RECT 158.460 39.160 158.780 39.220 ;
        RECT 170.880 39.160 171.200 39.220 ;
        RECT 158.460 39.020 171.200 39.160 ;
        RECT 158.460 38.960 158.780 39.020 ;
        RECT 170.880 38.960 171.200 39.020 ;
        RECT 172.720 39.160 173.040 39.220 ;
        RECT 215.055 39.160 215.345 39.205 ;
        RECT 172.720 39.020 215.345 39.160 ;
        RECT 172.720 38.960 173.040 39.020 ;
        RECT 215.055 38.975 215.345 39.020 ;
        RECT 245.400 39.160 245.720 39.220 ;
        RECT 250.460 39.160 250.780 39.220 ;
        RECT 245.400 39.020 250.780 39.160 ;
        RECT 245.400 38.960 245.720 39.020 ;
        RECT 250.460 38.960 250.780 39.020 ;
        RECT 286.340 39.160 286.660 39.220 ;
        RECT 291.860 39.160 292.180 39.220 ;
        RECT 286.340 39.020 292.180 39.160 ;
        RECT 286.340 38.960 286.660 39.020 ;
        RECT 291.860 38.960 292.180 39.020 ;
        RECT 292.320 39.160 292.640 39.220 ;
        RECT 297.840 39.160 298.160 39.220 ;
        RECT 292.320 39.020 298.160 39.160 ;
        RECT 292.320 38.960 292.640 39.020 ;
        RECT 297.840 38.960 298.160 39.020 ;
        RECT 135.920 38.820 136.240 38.880 ;
        RECT 171.800 38.820 172.120 38.880 ;
        RECT 135.920 38.680 172.120 38.820 ;
        RECT 135.920 38.620 136.240 38.680 ;
        RECT 171.800 38.620 172.120 38.680 ;
        RECT 175.035 38.820 175.325 38.865 ;
        RECT 222.860 38.820 223.180 38.880 ;
        RECT 175.035 38.680 223.180 38.820 ;
        RECT 175.035 38.635 175.325 38.680 ;
        RECT 222.860 38.620 223.180 38.680 ;
        RECT 127.640 38.480 127.960 38.540 ;
        RECT 129.940 38.480 130.260 38.540 ;
        RECT 127.640 38.340 130.260 38.480 ;
        RECT 127.640 38.280 127.960 38.340 ;
        RECT 129.940 38.280 130.260 38.340 ;
        RECT 147.420 38.480 147.740 38.540 ;
        RECT 175.940 38.480 176.260 38.540 ;
        RECT 147.420 38.340 176.260 38.480 ;
        RECT 147.420 38.280 147.740 38.340 ;
        RECT 175.940 38.280 176.260 38.340 ;
        RECT 282.660 38.480 282.980 38.540 ;
        RECT 324.980 38.480 325.300 38.540 ;
        RECT 282.660 38.340 325.300 38.480 ;
        RECT 282.660 38.280 282.980 38.340 ;
        RECT 324.980 38.280 325.300 38.340 ;
        RECT 154.780 38.140 155.100 38.200 ;
        RECT 175.020 38.140 175.340 38.200 ;
        RECT 154.780 38.000 175.340 38.140 ;
        RECT 154.780 37.940 155.100 38.000 ;
        RECT 175.020 37.940 175.340 38.000 ;
        RECT 347.980 37.800 348.300 37.860 ;
        RECT 359.480 37.800 359.800 37.860 ;
        RECT 347.980 37.660 359.800 37.800 ;
        RECT 347.980 37.600 348.300 37.660 ;
        RECT 359.480 37.600 359.800 37.660 ;
        RECT 149.720 37.460 150.040 37.520 ;
        RECT 178.700 37.460 179.020 37.520 ;
        RECT 149.720 37.320 179.020 37.460 ;
        RECT 149.720 37.260 150.040 37.320 ;
        RECT 178.700 37.260 179.020 37.320 ;
      LAYER via ;
        RECT 58.180 53.750 58.440 54.010 ;
        RECT 58.500 53.750 58.760 54.010 ;
        RECT 58.820 53.750 59.080 54.010 ;
        RECT 59.140 53.750 59.400 54.010 ;
        RECT 211.780 53.750 212.040 54.010 ;
        RECT 212.100 53.750 212.360 54.010 ;
        RECT 212.420 53.750 212.680 54.010 ;
        RECT 212.740 53.750 213.000 54.010 ;
        RECT 365.380 53.750 365.640 54.010 ;
        RECT 365.700 53.750 365.960 54.010 ;
        RECT 366.020 53.750 366.280 54.010 ;
        RECT 366.340 53.750 366.600 54.010 ;
        RECT 518.980 53.750 519.240 54.010 ;
        RECT 519.300 53.750 519.560 54.010 ;
        RECT 519.620 53.750 519.880 54.010 ;
        RECT 519.940 53.750 520.200 54.010 ;
        RECT 50.850 52.560 51.110 52.820 ;
        RECT 65.110 52.560 65.370 52.820 ;
        RECT 72.930 52.560 73.190 52.820 ;
        RECT 92.710 53.240 92.970 53.500 ;
        RECT 88.110 52.900 88.370 53.160 ;
        RECT 138.710 53.240 138.970 53.500 ;
        RECT 53.150 52.220 53.410 52.480 ;
        RECT 85.350 52.220 85.610 52.480 ;
        RECT 91.790 52.560 92.050 52.820 ;
        RECT 99.150 52.900 99.410 53.160 ;
        RECT 133.190 52.900 133.450 53.160 ;
        RECT 139.170 52.900 139.430 53.160 ;
        RECT 145.150 53.240 145.410 53.500 ;
        RECT 152.050 53.240 152.310 53.500 ;
        RECT 152.510 53.240 152.770 53.500 ;
        RECT 163.550 53.240 163.810 53.500 ;
        RECT 184.250 53.240 184.510 53.500 ;
        RECT 186.550 53.240 186.810 53.500 ;
        RECT 188.390 53.240 188.650 53.500 ;
        RECT 148.370 52.900 148.630 53.160 ;
        RECT 210.930 53.240 211.190 53.500 ;
        RECT 219.210 53.240 219.470 53.500 ;
        RECT 248.190 53.240 248.450 53.500 ;
        RECT 249.110 53.240 249.370 53.500 ;
        RECT 260.150 53.240 260.410 53.500 ;
        RECT 98.690 52.560 98.950 52.820 ;
        RECT 100.070 52.560 100.330 52.820 ;
        RECT 107.430 52.560 107.690 52.820 ;
        RECT 121.690 52.560 121.950 52.820 ;
        RECT 113.410 52.220 113.670 52.480 ;
        RECT 114.330 52.220 114.590 52.480 ;
        RECT 141.930 52.560 142.190 52.820 ;
        RECT 153.890 52.560 154.150 52.820 ;
        RECT 125.830 52.220 126.090 52.480 ;
        RECT 128.590 52.220 128.850 52.480 ;
        RECT 132.270 52.220 132.530 52.480 ;
        RECT 139.630 52.220 139.890 52.480 ;
        RECT 149.750 52.220 150.010 52.480 ;
        RECT 156.650 52.560 156.910 52.820 ;
        RECT 158.950 52.560 159.210 52.820 ;
        RECT 170.450 52.220 170.710 52.480 ;
        RECT 171.830 52.560 172.090 52.820 ;
        RECT 178.730 52.560 178.990 52.820 ;
        RECT 181.950 52.220 182.210 52.480 ;
        RECT 183.790 52.220 184.050 52.480 ;
        RECT 190.690 52.560 190.950 52.820 ;
        RECT 212.310 52.560 212.570 52.820 ;
        RECT 197.590 52.220 197.850 52.480 ;
        RECT 202.650 52.220 202.910 52.480 ;
        RECT 47.170 51.540 47.430 51.800 ;
        RECT 81.670 51.880 81.930 52.140 ;
        RECT 125.370 51.880 125.630 52.140 ;
        RECT 127.670 51.880 127.930 52.140 ;
        RECT 136.870 51.880 137.130 52.140 ;
        RECT 140.090 51.880 140.350 52.140 ;
        RECT 77.530 51.540 77.790 51.800 ;
        RECT 89.950 51.540 90.210 51.800 ;
        RECT 108.350 51.540 108.610 51.800 ;
        RECT 119.390 51.540 119.650 51.800 ;
        RECT 133.190 51.540 133.450 51.800 ;
        RECT 138.710 51.540 138.970 51.800 ;
        RECT 154.810 51.880 155.070 52.140 ;
        RECT 178.270 51.880 178.530 52.140 ;
        RECT 190.690 51.880 190.950 52.140 ;
        RECT 191.610 51.540 191.870 51.800 ;
        RECT 197.130 51.540 197.390 51.800 ;
        RECT 213.230 52.220 213.490 52.480 ;
        RECT 220.130 52.220 220.390 52.480 ;
        RECT 228.870 52.900 229.130 53.160 ;
        RECT 238.070 52.900 238.330 53.160 ;
        RECT 238.990 52.900 239.250 53.160 ;
        RECT 252.790 52.900 253.050 53.160 ;
        RECT 204.030 51.540 204.290 51.800 ;
        RECT 205.410 51.540 205.670 51.800 ;
        RECT 225.190 51.540 225.450 51.800 ;
        RECT 226.570 52.220 226.830 52.480 ;
        RECT 228.870 52.220 229.130 52.480 ;
        RECT 243.130 52.560 243.390 52.820 ;
        RECT 256.470 52.560 256.730 52.820 ;
        RECT 235.310 52.220 235.570 52.480 ;
        RECT 238.070 52.220 238.330 52.480 ;
        RECT 230.250 51.880 230.510 52.140 ;
        RECT 235.770 51.880 236.030 52.140 ;
        RECT 249.110 52.220 249.370 52.480 ;
        RECT 249.570 52.220 249.830 52.480 ;
        RECT 258.770 52.220 259.030 52.480 ;
        RECT 261.990 53.240 262.250 53.500 ;
        RECT 279.470 53.240 279.730 53.500 ;
        RECT 279.930 53.240 280.190 53.500 ;
        RECT 290.510 53.240 290.770 53.500 ;
        RECT 328.690 53.240 328.950 53.500 ;
        RECT 350.310 53.240 350.570 53.500 ;
        RECT 268.430 52.900 268.690 53.160 ;
        RECT 302.930 52.900 303.190 53.160 ;
        RECT 261.990 52.560 262.250 52.820 ;
        RECT 273.030 52.560 273.290 52.820 ;
        RECT 277.170 52.560 277.430 52.820 ;
        RECT 277.630 52.560 277.890 52.820 ;
        RECT 284.070 52.560 284.330 52.820 ;
        RECT 288.210 52.560 288.470 52.820 ;
        RECT 327.770 52.900 328.030 53.160 ;
        RECT 270.270 52.220 270.530 52.480 ;
        RECT 272.570 52.220 272.830 52.480 ;
        RECT 274.410 52.220 274.670 52.480 ;
        RECT 275.330 52.220 275.590 52.480 ;
        RECT 282.690 52.220 282.950 52.480 ;
        RECT 227.030 51.540 227.290 51.800 ;
        RECT 241.750 51.540 242.010 51.800 ;
        RECT 244.970 51.540 245.230 51.800 ;
        RECT 251.410 51.540 251.670 51.800 ;
        RECT 251.870 51.540 252.130 51.800 ;
        RECT 253.710 51.540 253.970 51.800 ;
        RECT 256.470 51.540 256.730 51.800 ;
        RECT 281.770 51.880 282.030 52.140 ;
        RECT 283.610 52.220 283.870 52.480 ;
        RECT 285.450 52.220 285.710 52.480 ;
        RECT 295.570 52.220 295.830 52.480 ;
        RECT 286.370 51.880 286.630 52.140 ;
        RECT 274.870 51.540 275.130 51.800 ;
        RECT 280.390 51.540 280.650 51.800 ;
        RECT 287.750 51.540 288.010 51.800 ;
        RECT 298.330 52.220 298.590 52.480 ;
        RECT 315.350 52.560 315.610 52.820 ;
        RECT 320.870 52.560 321.130 52.820 ;
        RECT 308.910 52.220 309.170 52.480 ;
        RECT 309.830 52.220 310.090 52.480 ;
        RECT 311.670 52.220 311.930 52.480 ;
        RECT 317.190 52.220 317.450 52.480 ;
        RECT 318.110 52.220 318.370 52.480 ;
        RECT 323.630 52.220 323.890 52.480 ;
        RECT 326.850 52.560 327.110 52.820 ;
        RECT 329.610 52.560 329.870 52.820 ;
        RECT 335.130 52.560 335.390 52.820 ;
        RECT 342.950 52.900 343.210 53.160 ;
        RECT 346.170 52.560 346.430 52.820 ;
        RECT 352.610 52.900 352.870 53.160 ;
        RECT 371.930 53.240 372.190 53.500 ;
        RECT 382.050 53.240 382.310 53.500 ;
        RECT 357.670 52.560 357.930 52.820 ;
        RECT 358.590 52.560 358.850 52.820 ;
        RECT 327.770 52.220 328.030 52.480 ;
        RECT 329.150 52.220 329.410 52.480 ;
        RECT 330.070 52.220 330.330 52.480 ;
        RECT 332.370 52.220 332.630 52.480 ;
        RECT 332.830 52.220 333.090 52.480 ;
        RECT 334.210 51.880 334.470 52.140 ;
        RECT 343.410 52.220 343.670 52.480 ;
        RECT 351.690 52.220 351.950 52.480 ;
        RECT 353.530 52.220 353.790 52.480 ;
        RECT 358.130 52.220 358.390 52.480 ;
        RECT 359.510 51.880 359.770 52.140 ;
        RECT 368.710 52.220 368.970 52.480 ;
        RECT 372.850 52.220 373.110 52.480 ;
        RECT 377.450 52.900 377.710 53.160 ;
        RECT 375.150 52.560 375.410 52.820 ;
        RECT 387.570 52.220 387.830 52.480 ;
        RECT 388.490 52.220 388.750 52.480 ;
        RECT 630.910 52.220 631.170 52.480 ;
        RECT 308.910 51.540 309.170 51.800 ;
        RECT 312.130 51.540 312.390 51.800 ;
        RECT 318.110 51.540 318.370 51.800 ;
        RECT 318.570 51.540 318.830 51.800 ;
        RECT 327.310 51.540 327.570 51.800 ;
        RECT 328.230 51.540 328.490 51.800 ;
        RECT 330.070 51.540 330.330 51.800 ;
        RECT 332.830 51.540 333.090 51.800 ;
        RECT 336.050 51.540 336.310 51.800 ;
        RECT 354.910 51.540 355.170 51.800 ;
        RECT 393.550 51.880 393.810 52.140 ;
        RECT 385.730 51.540 385.990 51.800 ;
        RECT 134.980 51.030 135.240 51.290 ;
        RECT 135.300 51.030 135.560 51.290 ;
        RECT 135.620 51.030 135.880 51.290 ;
        RECT 135.940 51.030 136.200 51.290 ;
        RECT 288.580 51.030 288.840 51.290 ;
        RECT 288.900 51.030 289.160 51.290 ;
        RECT 289.220 51.030 289.480 51.290 ;
        RECT 289.540 51.030 289.800 51.290 ;
        RECT 442.180 51.030 442.440 51.290 ;
        RECT 442.500 51.030 442.760 51.290 ;
        RECT 442.820 51.030 443.080 51.290 ;
        RECT 443.140 51.030 443.400 51.290 ;
        RECT 595.780 51.030 596.040 51.290 ;
        RECT 596.100 51.030 596.360 51.290 ;
        RECT 596.420 51.030 596.680 51.290 ;
        RECT 596.740 51.030 597.000 51.290 ;
        RECT 56.830 50.520 57.090 50.780 ;
        RECT 72.470 50.520 72.730 50.780 ;
        RECT 98.690 50.520 98.950 50.780 ;
        RECT 100.530 50.520 100.790 50.780 ;
        RECT 60.050 50.180 60.310 50.440 ;
        RECT 86.730 50.180 86.990 50.440 ;
        RECT 61.890 49.500 62.150 49.760 ;
        RECT 77.990 49.840 78.250 50.100 ;
        RECT 78.910 49.840 79.170 50.100 ;
        RECT 80.750 49.840 81.010 50.100 ;
        RECT 91.790 49.840 92.050 50.100 ;
        RECT 106.050 50.180 106.310 50.440 ;
        RECT 99.610 49.840 99.870 50.100 ;
        RECT 89.950 49.500 90.210 49.760 ;
        RECT 91.330 49.500 91.590 49.760 ;
        RECT 106.050 49.500 106.310 49.760 ;
        RECT 112.030 49.840 112.290 50.100 ;
        RECT 133.190 50.520 133.450 50.780 ;
        RECT 157.110 50.520 157.370 50.780 ;
        RECT 162.630 50.520 162.890 50.780 ;
        RECT 130.890 50.180 131.150 50.440 ;
        RECT 141.930 50.180 142.190 50.440 ;
        RECT 112.490 49.500 112.750 49.760 ;
        RECT 120.310 49.840 120.570 50.100 ;
        RECT 126.290 49.840 126.550 50.100 ;
        RECT 133.650 49.840 133.910 50.100 ;
        RECT 139.630 49.840 139.890 50.100 ;
        RECT 148.830 50.180 149.090 50.440 ;
        RECT 162.170 50.180 162.430 50.440 ;
        RECT 194.830 50.520 195.090 50.780 ;
        RECT 191.610 50.180 191.870 50.440 ;
        RECT 213.690 50.520 213.950 50.780 ;
        RECT 249.570 50.520 249.830 50.780 ;
        RECT 250.030 50.520 250.290 50.780 ;
        RECT 256.930 50.520 257.190 50.780 ;
        RECT 259.690 50.520 259.950 50.780 ;
        RECT 272.570 50.520 272.830 50.780 ;
        RECT 282.690 50.520 282.950 50.780 ;
        RECT 147.910 49.840 148.170 50.100 ;
        RECT 125.830 49.500 126.090 49.760 ;
        RECT 130.430 49.500 130.690 49.760 ;
        RECT 134.570 49.500 134.830 49.760 ;
        RECT 153.890 49.500 154.150 49.760 ;
        RECT 155.270 49.840 155.530 50.100 ;
        RECT 163.090 49.840 163.350 50.100 ;
        RECT 170.910 49.840 171.170 50.100 ;
        RECT 181.950 49.840 182.210 50.100 ;
        RECT 192.070 49.840 192.330 50.100 ;
        RECT 194.370 49.840 194.630 50.100 ;
        RECT 205.410 49.840 205.670 50.100 ;
        RECT 213.230 49.840 213.490 50.100 ;
        RECT 214.610 49.840 214.870 50.100 ;
        RECT 219.670 49.840 219.930 50.100 ;
        RECT 224.730 49.840 224.990 50.100 ;
        RECT 66.490 49.160 66.750 49.420 ;
        RECT 90.870 49.160 91.130 49.420 ;
        RECT 70.170 48.820 70.430 49.080 ;
        RECT 86.270 48.820 86.530 49.080 ;
        RECT 87.190 48.820 87.450 49.080 ;
        RECT 96.850 48.820 97.110 49.080 ;
        RECT 108.810 48.820 109.070 49.080 ;
        RECT 150.670 48.820 150.930 49.080 ;
        RECT 175.970 49.500 176.230 49.760 ;
        RECT 191.150 49.500 191.410 49.760 ;
        RECT 185.170 48.820 185.430 49.080 ;
        RECT 193.450 49.160 193.710 49.420 ;
        RECT 188.850 48.820 189.110 49.080 ;
        RECT 197.590 49.500 197.850 49.760 ;
        RECT 210.470 49.500 210.730 49.760 ;
        RECT 202.650 49.160 202.910 49.420 ;
        RECT 223.350 49.160 223.610 49.420 ;
        RECT 230.710 50.180 230.970 50.440 ;
        RECT 228.870 49.840 229.130 50.100 ;
        RECT 238.990 50.180 239.250 50.440 ;
        RECT 241.290 49.840 241.550 50.100 ;
        RECT 242.210 49.840 242.470 50.100 ;
        RECT 252.790 49.840 253.050 50.100 ;
        RECT 256.930 49.840 257.190 50.100 ;
        RECT 257.850 50.180 258.110 50.440 ;
        RECT 258.770 50.180 259.030 50.440 ;
        RECT 260.610 49.840 260.870 50.100 ;
        RECT 265.670 49.840 265.930 50.100 ;
        RECT 272.110 49.840 272.370 50.100 ;
        RECT 275.790 50.180 276.050 50.440 ;
        RECT 291.890 50.520 292.150 50.780 ;
        RECT 292.350 50.520 292.610 50.780 ;
        RECT 280.390 49.840 280.650 50.100 ;
        RECT 282.230 49.840 282.490 50.100 ;
        RECT 283.150 49.840 283.410 50.100 ;
        RECT 295.110 50.180 295.370 50.440 ;
        RECT 284.990 49.840 285.250 50.100 ;
        RECT 287.750 49.840 288.010 50.100 ;
        RECT 292.810 49.840 293.070 50.100 ;
        RECT 294.190 49.840 294.450 50.100 ;
        RECT 299.250 49.840 299.510 50.100 ;
        RECT 303.390 49.840 303.650 50.100 ;
        RECT 318.110 50.520 318.370 50.780 ;
        RECT 331.910 50.520 332.170 50.780 ;
        RECT 319.030 50.180 319.290 50.440 ;
        RECT 325.470 50.180 325.730 50.440 ;
        RECT 325.930 50.180 326.190 50.440 ;
        RECT 227.030 49.500 227.290 49.760 ;
        RECT 234.850 49.500 235.110 49.760 ;
        RECT 235.770 49.160 236.030 49.420 ;
        RECT 259.690 49.500 259.950 49.760 ;
        RECT 197.130 48.820 197.390 49.080 ;
        RECT 197.590 48.820 197.850 49.080 ;
        RECT 202.190 48.820 202.450 49.080 ;
        RECT 203.110 48.820 203.370 49.080 ;
        RECT 205.410 48.820 205.670 49.080 ;
        RECT 217.830 48.820 218.090 49.080 ;
        RECT 228.410 48.820 228.670 49.080 ;
        RECT 241.750 48.820 242.010 49.080 ;
        RECT 243.130 48.820 243.390 49.080 ;
        RECT 246.350 49.160 246.610 49.420 ;
        RECT 270.270 49.500 270.530 49.760 ;
        RECT 276.250 49.500 276.510 49.760 ;
        RECT 287.750 49.160 288.010 49.420 ;
        RECT 296.490 49.500 296.750 49.760 ;
        RECT 304.310 49.500 304.570 49.760 ;
        RECT 310.750 49.500 311.010 49.760 ;
        RECT 295.110 49.160 295.370 49.420 ;
        RECT 259.690 48.820 259.950 49.080 ;
        RECT 270.270 48.820 270.530 49.080 ;
        RECT 274.410 48.820 274.670 49.080 ;
        RECT 276.250 48.820 276.510 49.080 ;
        RECT 283.150 48.820 283.410 49.080 ;
        RECT 290.510 48.820 290.770 49.080 ;
        RECT 292.350 48.820 292.610 49.080 ;
        RECT 314.890 48.820 315.150 49.080 ;
        RECT 326.850 49.840 327.110 50.100 ;
        RECT 328.230 50.180 328.490 50.440 ;
        RECT 331.450 49.840 331.710 50.100 ;
        RECT 336.050 49.840 336.310 50.100 ;
        RECT 337.430 49.840 337.690 50.100 ;
        RECT 345.250 50.180 345.510 50.440 ;
        RECT 348.010 50.520 348.270 50.780 ;
        RECT 354.910 50.520 355.170 50.780 ;
        RECT 347.550 50.180 347.810 50.440 ;
        RECT 353.070 49.840 353.330 50.100 ;
        RECT 359.050 50.180 359.310 50.440 ;
        RECT 374.690 50.520 374.950 50.780 ;
        RECT 376.070 50.520 376.330 50.780 ;
        RECT 382.050 50.520 382.310 50.780 ;
        RECT 394.930 50.520 395.190 50.780 ;
        RECT 343.410 49.500 343.670 49.760 ;
        RECT 327.310 48.820 327.570 49.080 ;
        RECT 344.330 49.160 344.590 49.420 ;
        RECT 353.070 49.160 353.330 49.420 ;
        RECT 382.510 50.180 382.770 50.440 ;
        RECT 382.970 50.180 383.230 50.440 ;
        RECT 391.250 50.180 391.510 50.440 ;
        RECT 368.710 49.840 368.970 50.100 ;
        RECT 360.430 49.500 360.690 49.760 ;
        RECT 375.150 49.840 375.410 50.100 ;
        RECT 400.910 49.840 401.170 50.100 ;
        RECT 366.870 49.160 367.130 49.420 ;
        RECT 342.950 48.820 343.210 49.080 ;
        RECT 350.310 48.820 350.570 49.080 ;
        RECT 357.670 48.820 357.930 49.080 ;
        RECT 359.510 48.820 359.770 49.080 ;
        RECT 392.170 48.820 392.430 49.080 ;
        RECT 395.850 48.820 396.110 49.080 ;
        RECT 403.210 48.820 403.470 49.080 ;
        RECT 414.250 48.820 414.510 49.080 ;
        RECT 428.970 48.820 429.230 49.080 ;
        RECT 436.330 48.820 436.590 49.080 ;
        RECT 447.370 48.820 447.630 49.080 ;
        RECT 458.410 48.820 458.670 49.080 ;
        RECT 469.450 48.820 469.710 49.080 ;
        RECT 480.490 48.820 480.750 49.080 ;
        RECT 487.850 48.820 488.110 49.080 ;
        RECT 513.610 48.820 513.870 49.080 ;
        RECT 520.970 48.820 521.230 49.080 ;
        RECT 535.690 48.820 535.950 49.080 ;
        RECT 543.050 48.820 543.310 49.080 ;
        RECT 554.090 48.820 554.350 49.080 ;
        RECT 564.670 48.820 564.930 49.080 ;
        RECT 572.030 48.820 572.290 49.080 ;
        RECT 597.790 48.820 598.050 49.080 ;
        RECT 619.870 48.820 620.130 49.080 ;
        RECT 627.230 48.820 627.490 49.080 ;
        RECT 58.180 48.310 58.440 48.570 ;
        RECT 58.500 48.310 58.760 48.570 ;
        RECT 58.820 48.310 59.080 48.570 ;
        RECT 59.140 48.310 59.400 48.570 ;
        RECT 211.780 48.310 212.040 48.570 ;
        RECT 212.100 48.310 212.360 48.570 ;
        RECT 212.420 48.310 212.680 48.570 ;
        RECT 212.740 48.310 213.000 48.570 ;
        RECT 365.380 48.310 365.640 48.570 ;
        RECT 365.700 48.310 365.960 48.570 ;
        RECT 366.020 48.310 366.280 48.570 ;
        RECT 366.340 48.310 366.600 48.570 ;
        RECT 518.980 48.310 519.240 48.570 ;
        RECT 519.300 48.310 519.560 48.570 ;
        RECT 519.620 48.310 519.880 48.570 ;
        RECT 519.940 48.310 520.200 48.570 ;
        RECT 83.970 47.800 84.230 48.060 ;
        RECT 99.150 47.800 99.410 48.060 ;
        RECT 106.970 47.800 107.230 48.060 ;
        RECT 146.530 47.800 146.790 48.060 ;
        RECT 149.750 47.800 150.010 48.060 ;
        RECT 153.430 47.800 153.690 48.060 ;
        RECT 176.890 47.800 177.150 48.060 ;
        RECT 184.710 47.800 184.970 48.060 ;
        RECT 213.690 47.800 213.950 48.060 ;
        RECT 219.670 47.800 219.930 48.060 ;
        RECT 223.810 47.800 224.070 48.060 ;
        RECT 224.730 47.800 224.990 48.060 ;
        RECT 230.710 47.800 230.970 48.060 ;
        RECT 233.930 47.800 234.190 48.060 ;
        RECT 234.390 47.800 234.650 48.060 ;
        RECT 240.370 47.800 240.630 48.060 ;
        RECT 55.450 47.460 55.710 47.720 ;
        RECT 42.110 47.120 42.370 47.380 ;
        RECT 78.450 47.120 78.710 47.380 ;
        RECT 89.030 47.120 89.290 47.380 ;
        RECT 43.490 46.780 43.750 47.040 ;
        RECT 48.090 46.440 48.350 46.700 ;
        RECT 63.730 46.440 63.990 46.700 ;
        RECT 90.410 46.780 90.670 47.040 ;
        RECT 91.790 47.460 92.050 47.720 ;
        RECT 105.590 47.460 105.850 47.720 ;
        RECT 91.330 47.120 91.590 47.380 ;
        RECT 119.390 47.460 119.650 47.720 ;
        RECT 120.310 47.460 120.570 47.720 ;
        RECT 125.830 47.460 126.090 47.720 ;
        RECT 93.170 46.780 93.430 47.040 ;
        RECT 114.790 47.120 115.050 47.380 ;
        RECT 106.050 46.780 106.310 47.040 ;
        RECT 40.730 46.100 40.990 46.360 ;
        RECT 84.890 46.440 85.150 46.700 ;
        RECT 102.370 46.440 102.630 46.700 ;
        RECT 112.490 46.780 112.750 47.040 ;
        RECT 118.010 47.120 118.270 47.380 ;
        RECT 118.470 47.120 118.730 47.380 ;
        RECT 134.570 47.460 134.830 47.720 ;
        RECT 128.590 47.120 128.850 47.380 ;
        RECT 119.390 46.780 119.650 47.040 ;
        RECT 136.870 47.120 137.130 47.380 ;
        RECT 143.770 46.780 144.030 47.040 ;
        RECT 147.450 47.460 147.710 47.720 ;
        RECT 167.230 47.460 167.490 47.720 ;
        RECT 153.890 47.120 154.150 47.380 ;
        RECT 189.770 47.460 190.030 47.720 ;
        RECT 217.830 47.460 218.090 47.720 ;
        RECT 219.210 47.460 219.470 47.720 ;
        RECT 226.570 47.460 226.830 47.720 ;
        RECT 228.410 47.460 228.670 47.720 ;
        RECT 238.990 47.460 239.250 47.720 ;
        RECT 246.810 47.800 247.070 48.060 ;
        RECT 247.270 47.800 247.530 48.060 ;
        RECT 268.430 47.800 268.690 48.060 ;
        RECT 170.910 47.120 171.170 47.380 ;
        RECT 145.150 46.780 145.410 47.040 ;
        RECT 112.950 46.440 113.210 46.700 ;
        RECT 115.710 46.440 115.970 46.700 ;
        RECT 118.930 46.440 119.190 46.700 ;
        RECT 120.770 46.440 121.030 46.700 ;
        RECT 85.350 46.100 85.610 46.360 ;
        RECT 86.270 46.100 86.530 46.360 ;
        RECT 92.710 46.100 92.970 46.360 ;
        RECT 98.230 46.100 98.490 46.360 ;
        RECT 104.670 46.100 104.930 46.360 ;
        RECT 137.790 46.440 138.050 46.700 ;
        RECT 147.450 46.780 147.710 47.040 ;
        RECT 160.330 46.780 160.590 47.040 ;
        RECT 177.810 46.780 178.070 47.040 ;
        RECT 184.710 46.780 184.970 47.040 ;
        RECT 205.410 47.120 205.670 47.380 ;
        RECT 194.830 46.780 195.090 47.040 ;
        RECT 197.130 46.780 197.390 47.040 ;
        RECT 218.290 47.120 218.550 47.380 ;
        RECT 230.250 47.120 230.510 47.380 ;
        RECT 230.710 47.120 230.970 47.380 ;
        RECT 231.630 47.120 231.890 47.380 ;
        RECT 233.010 47.120 233.270 47.380 ;
        RECT 234.850 47.120 235.110 47.380 ;
        RECT 242.670 47.460 242.930 47.720 ;
        RECT 253.710 47.460 253.970 47.720 ;
        RECT 264.290 47.460 264.550 47.720 ;
        RECT 276.250 47.800 276.510 48.060 ;
        RECT 283.610 47.800 283.870 48.060 ;
        RECT 274.410 47.460 274.670 47.720 ;
        RECT 309.830 47.460 310.090 47.720 ;
        RECT 311.670 47.800 311.930 48.060 ;
        RECT 317.650 47.800 317.910 48.060 ;
        RECT 325.930 47.800 326.190 48.060 ;
        RECT 333.750 47.800 334.010 48.060 ;
        RECT 334.210 47.800 334.470 48.060 ;
        RECT 332.370 47.460 332.630 47.720 ;
        RECT 141.010 46.100 141.270 46.360 ;
        RECT 142.390 46.100 142.650 46.360 ;
        RECT 156.650 46.100 156.910 46.360 ;
        RECT 160.330 46.100 160.590 46.360 ;
        RECT 165.850 46.100 166.110 46.360 ;
        RECT 196.670 46.440 196.930 46.700 ;
        RECT 202.190 46.440 202.450 46.700 ;
        RECT 214.150 46.780 214.410 47.040 ;
        RECT 220.130 46.780 220.390 47.040 ;
        RECT 228.410 46.780 228.670 47.040 ;
        RECT 240.370 46.780 240.630 47.040 ;
        RECT 227.490 46.440 227.750 46.700 ;
        RECT 231.170 46.440 231.430 46.700 ;
        RECT 231.630 46.440 231.890 46.700 ;
        RECT 233.470 46.440 233.730 46.700 ;
        RECT 233.930 46.440 234.190 46.700 ;
        RECT 238.070 46.440 238.330 46.700 ;
        RECT 238.990 46.440 239.250 46.700 ;
        RECT 245.430 47.120 245.690 47.380 ;
        RECT 252.330 47.120 252.590 47.380 ;
        RECT 243.590 46.780 243.850 47.040 ;
        RECT 244.050 46.780 244.310 47.040 ;
        RECT 251.870 46.780 252.130 47.040 ;
        RECT 253.250 46.780 253.510 47.040 ;
        RECT 256.010 46.780 256.270 47.040 ;
        RECT 261.070 46.780 261.330 47.040 ;
        RECT 270.730 46.780 270.990 47.040 ;
        RECT 254.630 46.440 254.890 46.700 ;
        RECT 256.470 46.440 256.730 46.700 ;
        RECT 275.790 46.780 276.050 47.040 ;
        RECT 284.070 46.780 284.330 47.040 ;
        RECT 214.610 46.100 214.870 46.360 ;
        RECT 228.410 46.100 228.670 46.360 ;
        RECT 246.350 46.100 246.610 46.360 ;
        RECT 246.810 46.100 247.070 46.360 ;
        RECT 262.450 46.100 262.710 46.360 ;
        RECT 286.830 46.440 287.090 46.700 ;
        RECT 284.530 46.100 284.790 46.360 ;
        RECT 285.450 46.100 285.710 46.360 ;
        RECT 292.350 47.120 292.610 47.380 ;
        RECT 293.270 47.120 293.530 47.380 ;
        RECT 289.130 46.780 289.390 47.040 ;
        RECT 290.970 46.780 291.230 47.040 ;
        RECT 298.330 46.780 298.590 47.040 ;
        RECT 299.710 46.780 299.970 47.040 ;
        RECT 316.270 47.120 316.530 47.380 ;
        RECT 302.930 46.100 303.190 46.360 ;
        RECT 306.150 46.780 306.410 47.040 ;
        RECT 314.430 46.780 314.690 47.040 ;
        RECT 314.890 46.780 315.150 47.040 ;
        RECT 338.350 47.120 338.610 47.380 ;
        RECT 342.950 47.800 343.210 48.060 ;
        RECT 361.810 47.800 362.070 48.060 ;
        RECT 362.270 47.800 362.530 48.060 ;
        RECT 380.210 47.800 380.470 48.060 ;
        RECT 350.770 47.120 351.030 47.380 ;
        RECT 326.390 46.780 326.650 47.040 ;
        RECT 332.830 46.780 333.090 47.040 ;
        RECT 333.290 46.780 333.550 47.040 ;
        RECT 340.190 46.780 340.450 47.040 ;
        RECT 330.990 46.440 331.250 46.700 ;
        RECT 334.210 46.440 334.470 46.700 ;
        RECT 311.210 46.100 311.470 46.360 ;
        RECT 312.590 46.100 312.850 46.360 ;
        RECT 324.090 46.100 324.350 46.360 ;
        RECT 325.470 46.100 325.730 46.360 ;
        RECT 338.810 46.100 339.070 46.360 ;
        RECT 339.730 46.100 339.990 46.360 ;
        RECT 341.570 46.780 341.830 47.040 ;
        RECT 347.550 46.780 347.810 47.040 ;
        RECT 342.490 46.440 342.750 46.700 ;
        RECT 353.530 46.780 353.790 47.040 ;
        RECT 345.710 46.100 345.970 46.360 ;
        RECT 356.750 46.440 357.010 46.700 ;
        RECT 352.610 46.100 352.870 46.360 ;
        RECT 357.670 46.100 357.930 46.360 ;
        RECT 367.790 46.440 368.050 46.700 ;
        RECT 369.170 46.780 369.430 47.040 ;
        RECT 370.550 47.120 370.810 47.380 ;
        RECT 373.770 47.120 374.030 47.380 ;
        RECT 399.530 46.780 399.790 47.040 ;
        RECT 406.890 46.780 407.150 47.040 ;
        RECT 410.570 46.780 410.830 47.040 ;
        RECT 417.930 46.780 418.190 47.040 ;
        RECT 421.610 46.780 421.870 47.040 ;
        RECT 425.290 46.780 425.550 47.040 ;
        RECT 440.010 46.780 440.270 47.040 ;
        RECT 443.690 46.780 443.950 47.040 ;
        RECT 451.050 46.780 451.310 47.040 ;
        RECT 454.730 46.780 454.990 47.040 ;
        RECT 465.770 46.780 466.030 47.040 ;
        RECT 473.130 46.780 473.390 47.040 ;
        RECT 476.810 46.780 477.070 47.040 ;
        RECT 484.170 46.780 484.430 47.040 ;
        RECT 491.530 46.780 491.790 47.040 ;
        RECT 495.210 46.780 495.470 47.040 ;
        RECT 498.890 46.780 499.150 47.040 ;
        RECT 506.250 46.780 506.510 47.040 ;
        RECT 517.290 46.780 517.550 47.040 ;
        RECT 524.650 46.780 524.910 47.040 ;
        RECT 528.330 46.780 528.590 47.040 ;
        RECT 532.010 46.780 532.270 47.040 ;
        RECT 539.370 46.780 539.630 47.040 ;
        RECT 546.730 46.780 546.990 47.040 ;
        RECT 550.410 46.780 550.670 47.040 ;
        RECT 557.770 46.780 558.030 47.040 ;
        RECT 561.450 46.780 561.710 47.040 ;
        RECT 568.350 46.780 568.610 47.040 ;
        RECT 575.710 46.780 575.970 47.040 ;
        RECT 579.390 46.780 579.650 47.040 ;
        RECT 583.070 46.780 583.330 47.040 ;
        RECT 590.430 46.780 590.690 47.040 ;
        RECT 594.110 46.780 594.370 47.040 ;
        RECT 601.470 46.780 601.730 47.040 ;
        RECT 608.830 46.780 609.090 47.040 ;
        RECT 612.510 46.780 612.770 47.040 ;
        RECT 616.190 46.780 616.450 47.040 ;
        RECT 623.550 46.780 623.810 47.040 ;
        RECT 375.150 46.440 375.410 46.700 ;
        RECT 381.130 46.440 381.390 46.700 ;
        RECT 389.870 46.440 390.130 46.700 ;
        RECT 370.090 46.100 370.350 46.360 ;
        RECT 386.190 46.100 386.450 46.360 ;
        RECT 386.650 46.100 386.910 46.360 ;
        RECT 398.610 46.100 398.870 46.360 ;
        RECT 134.980 45.590 135.240 45.850 ;
        RECT 135.300 45.590 135.560 45.850 ;
        RECT 135.620 45.590 135.880 45.850 ;
        RECT 135.940 45.590 136.200 45.850 ;
        RECT 288.580 45.590 288.840 45.850 ;
        RECT 288.900 45.590 289.160 45.850 ;
        RECT 289.220 45.590 289.480 45.850 ;
        RECT 289.540 45.590 289.800 45.850 ;
        RECT 442.180 45.590 442.440 45.850 ;
        RECT 442.500 45.590 442.760 45.850 ;
        RECT 442.820 45.590 443.080 45.850 ;
        RECT 443.140 45.590 443.400 45.850 ;
        RECT 595.780 45.590 596.040 45.850 ;
        RECT 596.100 45.590 596.360 45.850 ;
        RECT 596.420 45.590 596.680 45.850 ;
        RECT 596.740 45.590 597.000 45.850 ;
        RECT 39.810 44.060 40.070 44.320 ;
        RECT 78.450 44.740 78.710 45.000 ;
        RECT 89.490 44.740 89.750 45.000 ;
        RECT 97.310 44.740 97.570 45.000 ;
        RECT 65.570 44.400 65.830 44.660 ;
        RECT 90.870 44.400 91.130 44.660 ;
        RECT 94.090 44.400 94.350 44.660 ;
        RECT 100.530 44.400 100.790 44.660 ;
        RECT 101.910 44.740 102.170 45.000 ;
        RECT 110.190 44.740 110.450 45.000 ;
        RECT 128.130 45.080 128.390 45.340 ;
        RECT 141.010 45.080 141.270 45.340 ;
        RECT 115.250 44.400 115.510 44.660 ;
        RECT 62.810 43.720 63.070 43.980 ;
        RECT 118.470 44.060 118.730 44.320 ;
        RECT 123.530 44.740 123.790 45.000 ;
        RECT 127.670 44.740 127.930 45.000 ;
        RECT 135.950 44.400 136.210 44.660 ;
        RECT 136.870 44.400 137.130 44.660 ;
        RECT 137.330 44.400 137.590 44.660 ;
        RECT 186.090 45.080 186.350 45.340 ;
        RECT 191.150 45.080 191.410 45.340 ;
        RECT 216.450 45.080 216.710 45.340 ;
        RECT 226.110 45.080 226.370 45.340 ;
        RECT 162.630 44.740 162.890 45.000 ;
        RECT 172.290 44.740 172.550 45.000 ;
        RECT 185.170 44.740 185.430 45.000 ;
        RECT 129.050 44.060 129.310 44.320 ;
        RECT 153.890 44.400 154.150 44.660 ;
        RECT 174.590 44.400 174.850 44.660 ;
        RECT 178.270 44.400 178.530 44.660 ;
        RECT 184.710 44.400 184.970 44.660 ;
        RECT 205.870 44.400 206.130 44.660 ;
        RECT 210.010 44.740 210.270 45.000 ;
        RECT 208.170 44.400 208.430 44.660 ;
        RECT 219.210 44.740 219.470 45.000 ;
        RECT 232.090 45.080 232.350 45.340 ;
        RECT 259.230 45.080 259.490 45.340 ;
        RECT 240.830 44.740 241.090 45.000 ;
        RECT 215.070 44.400 215.330 44.660 ;
        RECT 216.450 44.400 216.710 44.660 ;
        RECT 221.050 44.400 221.310 44.660 ;
        RECT 221.510 44.400 221.770 44.660 ;
        RECT 228.410 44.400 228.670 44.660 ;
        RECT 229.790 44.400 230.050 44.660 ;
        RECT 235.770 44.400 236.030 44.660 ;
        RECT 238.990 44.400 239.250 44.660 ;
        RECT 243.590 44.400 243.850 44.660 ;
        RECT 247.270 44.740 247.530 45.000 ;
        RECT 85.350 43.380 85.610 43.640 ;
        RECT 119.390 43.720 119.650 43.980 ;
        RECT 120.310 43.380 120.570 43.640 ;
        RECT 123.530 43.380 123.790 43.640 ;
        RECT 131.810 43.380 132.070 43.640 ;
        RECT 136.870 43.720 137.130 43.980 ;
        RECT 156.190 44.060 156.450 44.320 ;
        RECT 156.650 43.720 156.910 43.980 ;
        RECT 174.130 44.060 174.390 44.320 ;
        RECT 179.650 44.060 179.910 44.320 ;
        RECT 207.710 44.060 207.970 44.320 ;
        RECT 230.710 44.060 230.970 44.320 ;
        RECT 233.010 44.060 233.270 44.320 ;
        RECT 257.850 44.400 258.110 44.660 ;
        RECT 258.770 44.400 259.030 44.660 ;
        RECT 270.730 44.400 270.990 44.660 ;
        RECT 293.730 45.080 293.990 45.340 ;
        RECT 213.690 43.720 213.950 43.980 ;
        RECT 232.550 43.720 232.810 43.980 ;
        RECT 237.610 43.720 237.870 43.980 ;
        RECT 244.970 43.720 245.230 43.980 ;
        RECT 267.970 44.060 268.230 44.320 ;
        RECT 258.310 43.720 258.570 43.980 ;
        RECT 275.790 44.060 276.050 44.320 ;
        RECT 279.470 44.400 279.730 44.660 ;
        RECT 292.350 44.740 292.610 45.000 ;
        RECT 292.810 44.740 293.070 45.000 ;
        RECT 297.870 45.080 298.130 45.340 ;
        RECT 299.250 45.080 299.510 45.340 ;
        RECT 305.230 45.080 305.490 45.340 ;
        RECT 305.690 45.080 305.950 45.340 ;
        RECT 357.210 45.080 357.470 45.340 ;
        RECT 358.130 45.080 358.390 45.340 ;
        RECT 288.670 44.400 288.930 44.660 ;
        RECT 298.790 44.400 299.050 44.660 ;
        RECT 312.590 44.740 312.850 45.000 ;
        RECT 306.150 44.400 306.410 44.660 ;
        RECT 326.390 44.740 326.650 45.000 ;
        RECT 292.810 44.060 293.070 44.320 ;
        RECT 298.330 44.060 298.590 44.320 ;
        RECT 302.010 44.060 302.270 44.320 ;
        RECT 163.090 43.380 163.350 43.640 ;
        RECT 164.010 43.380 164.270 43.640 ;
        RECT 216.450 43.380 216.710 43.640 ;
        RECT 221.970 43.380 222.230 43.640 ;
        RECT 236.690 43.380 236.950 43.640 ;
        RECT 264.750 43.380 265.010 43.640 ;
        RECT 313.510 43.720 313.770 43.980 ;
        RECT 315.810 44.060 316.070 44.320 ;
        RECT 319.950 43.720 320.210 43.980 ;
        RECT 298.330 43.380 298.590 43.640 ;
        RECT 308.450 43.380 308.710 43.640 ;
        RECT 309.830 43.380 310.090 43.640 ;
        RECT 317.650 43.380 317.910 43.640 ;
        RECT 336.510 44.400 336.770 44.660 ;
        RECT 345.250 44.400 345.510 44.660 ;
        RECT 342.950 44.060 343.210 44.320 ;
        RECT 338.350 43.720 338.610 43.980 ;
        RECT 352.150 44.400 352.410 44.660 ;
        RECT 358.130 44.400 358.390 44.660 ;
        RECT 358.590 44.400 358.850 44.660 ;
        RECT 381.130 44.400 381.390 44.660 ;
        RECT 386.190 44.400 386.450 44.660 ;
        RECT 333.290 43.380 333.550 43.640 ;
        RECT 336.970 43.380 337.230 43.640 ;
        RECT 358.130 43.380 358.390 43.640 ;
        RECT 371.470 43.380 371.730 43.640 ;
        RECT 379.750 43.380 380.010 43.640 ;
        RECT 381.130 43.720 381.390 43.980 ;
        RECT 404.590 43.380 404.850 43.640 ;
        RECT 502.570 43.380 502.830 43.640 ;
        RECT 586.750 43.380 587.010 43.640 ;
        RECT 58.180 42.870 58.440 43.130 ;
        RECT 58.500 42.870 58.760 43.130 ;
        RECT 58.820 42.870 59.080 43.130 ;
        RECT 59.140 42.870 59.400 43.130 ;
        RECT 211.780 42.870 212.040 43.130 ;
        RECT 212.100 42.870 212.360 43.130 ;
        RECT 212.420 42.870 212.680 43.130 ;
        RECT 212.740 42.870 213.000 43.130 ;
        RECT 365.380 42.870 365.640 43.130 ;
        RECT 365.700 42.870 365.960 43.130 ;
        RECT 366.020 42.870 366.280 43.130 ;
        RECT 366.340 42.870 366.600 43.130 ;
        RECT 518.980 42.870 519.240 43.130 ;
        RECT 519.300 42.870 519.560 43.130 ;
        RECT 519.620 42.870 519.880 43.130 ;
        RECT 519.940 42.870 520.200 43.130 ;
        RECT 77.530 42.360 77.790 42.620 ;
        RECT 115.250 42.360 115.510 42.620 ;
        RECT 117.550 42.360 117.810 42.620 ;
        RECT 84.890 42.020 85.150 42.280 ;
        RECT 137.330 42.020 137.590 42.280 ;
        RECT 137.790 42.020 138.050 42.280 ;
        RECT 156.650 42.360 156.910 42.620 ;
        RECT 213.690 42.360 213.950 42.620 ;
        RECT 215.070 42.360 215.330 42.620 ;
        RECT 221.510 42.360 221.770 42.620 ;
        RECT 221.970 42.360 222.230 42.620 ;
        RECT 237.150 42.360 237.410 42.620 ;
        RECT 243.590 42.360 243.850 42.620 ;
        RECT 178.270 42.020 178.530 42.280 ;
        RECT 233.010 42.020 233.270 42.280 ;
        RECT 282.230 42.360 282.490 42.620 ;
        RECT 336.970 42.360 337.230 42.620 ;
        RECT 287.290 42.020 287.550 42.280 ;
        RECT 289.590 42.020 289.850 42.280 ;
        RECT 301.090 42.020 301.350 42.280 ;
        RECT 329.610 42.020 329.870 42.280 ;
        RECT 357.210 42.360 357.470 42.620 ;
        RECT 352.150 42.020 352.410 42.280 ;
        RECT 402.290 42.020 402.550 42.280 ;
        RECT 86.270 41.680 86.530 41.940 ;
        RECT 164.470 41.680 164.730 41.940 ;
        RECT 201.270 41.680 201.530 41.940 ;
        RECT 264.750 41.680 265.010 41.940 ;
        RECT 273.950 41.680 274.210 41.940 ;
        RECT 302.010 41.680 302.270 41.940 ;
        RECT 344.330 41.680 344.590 41.940 ;
        RECT 379.750 41.680 380.010 41.940 ;
        RECT 37.510 41.340 37.770 41.600 ;
        RECT 345.250 41.340 345.510 41.600 ;
        RECT 87.190 41.000 87.450 41.260 ;
        RECT 175.510 41.000 175.770 41.260 ;
        RECT 208.170 41.000 208.430 41.260 ;
        RECT 239.910 41.000 240.170 41.260 ;
        RECT 342.950 41.000 343.210 41.260 ;
        RECT 118.470 40.660 118.730 40.920 ;
        RECT 136.870 40.660 137.130 40.920 ;
        RECT 143.770 40.660 144.030 40.920 ;
        RECT 154.810 40.660 155.070 40.920 ;
        RECT 162.630 40.660 162.890 40.920 ;
        RECT 163.090 40.660 163.350 40.920 ;
        RECT 280.390 40.660 280.650 40.920 ;
        RECT 315.810 40.660 316.070 40.920 ;
        RECT 336.510 40.660 336.770 40.920 ;
        RECT 358.130 40.660 358.390 40.920 ;
        RECT 111.570 40.320 111.830 40.580 ;
        RECT 230.710 40.320 230.970 40.580 ;
        RECT 244.970 40.320 245.230 40.580 ;
        RECT 308.450 40.320 308.710 40.580 ;
        RECT 311.210 40.320 311.470 40.580 ;
        RECT 323.630 40.320 323.890 40.580 ;
        RECT 329.150 40.320 329.410 40.580 ;
        RECT 369.170 40.320 369.430 40.580 ;
        RECT 123.530 39.980 123.790 40.240 ;
        RECT 169.070 39.980 169.330 40.240 ;
        RECT 174.130 39.980 174.390 40.240 ;
        RECT 220.590 39.980 220.850 40.240 ;
        RECT 228.410 39.980 228.670 40.240 ;
        RECT 285.450 39.980 285.710 40.240 ;
        RECT 341.110 39.980 341.370 40.240 ;
        RECT 372.850 39.980 373.110 40.240 ;
        RECT 88.570 39.640 88.830 39.900 ;
        RECT 130.430 39.640 130.690 39.900 ;
        RECT 131.810 39.640 132.070 39.900 ;
        RECT 155.730 39.640 155.990 39.900 ;
        RECT 179.190 39.640 179.450 39.900 ;
        RECT 230.710 39.640 230.970 39.900 ;
        RECT 255.090 39.640 255.350 39.900 ;
        RECT 270.730 39.640 270.990 39.900 ;
        RECT 292.810 39.640 293.070 39.900 ;
        RECT 293.270 39.640 293.530 39.900 ;
        RECT 303.850 39.640 304.110 39.900 ;
        RECT 332.830 39.640 333.090 39.900 ;
        RECT 342.030 39.640 342.290 39.900 ;
        RECT 117.090 39.300 117.350 39.560 ;
        RECT 118.010 39.300 118.270 39.560 ;
        RECT 164.010 39.300 164.270 39.560 ;
        RECT 165.390 39.300 165.650 39.560 ;
        RECT 238.070 39.300 238.330 39.560 ;
        RECT 245.890 39.300 246.150 39.560 ;
        RECT 256.470 39.300 256.730 39.560 ;
        RECT 276.710 39.300 276.970 39.560 ;
        RECT 281.770 39.300 282.030 39.560 ;
        RECT 299.250 39.300 299.510 39.560 ;
        RECT 106.050 38.960 106.310 39.220 ;
        RECT 126.750 38.960 127.010 39.220 ;
        RECT 158.490 38.960 158.750 39.220 ;
        RECT 170.910 38.960 171.170 39.220 ;
        RECT 172.750 38.960 173.010 39.220 ;
        RECT 245.430 38.960 245.690 39.220 ;
        RECT 250.490 38.960 250.750 39.220 ;
        RECT 286.370 38.960 286.630 39.220 ;
        RECT 291.890 38.960 292.150 39.220 ;
        RECT 292.350 38.960 292.610 39.220 ;
        RECT 297.870 38.960 298.130 39.220 ;
        RECT 135.950 38.620 136.210 38.880 ;
        RECT 171.830 38.620 172.090 38.880 ;
        RECT 222.890 38.620 223.150 38.880 ;
        RECT 127.670 38.280 127.930 38.540 ;
        RECT 129.970 38.280 130.230 38.540 ;
        RECT 147.450 38.280 147.710 38.540 ;
        RECT 175.970 38.280 176.230 38.540 ;
        RECT 282.690 38.280 282.950 38.540 ;
        RECT 325.010 38.280 325.270 38.540 ;
        RECT 154.810 37.940 155.070 38.200 ;
        RECT 175.050 37.940 175.310 38.200 ;
        RECT 348.010 37.600 348.270 37.860 ;
        RECT 359.510 37.600 359.770 37.860 ;
        RECT 149.750 37.260 150.010 37.520 ;
        RECT 178.730 37.260 178.990 37.520 ;
        RECT 44.410 610.840 44.670 611.100 ;
        RECT 49.470 609.140 49.730 609.400 ;
      LAYER met2 ;
        RECT 39.340 629.720 39.620 632.120 ;
        RECT 44.400 629.720 44.680 632.120 ;
        RECT 49.460 629.720 49.740 632.120 ;
        RECT 44.470 611.130 44.610 629.720 ;
        RECT 44.410 610.810 44.670 611.130 ;
        RECT 49.530 609.430 49.670 629.720 ;
        RECT 49.470 609.110 49.730 609.430 ;
        RECT 54.000 54.000 636.240 632.120 ;
        RECT 58.050 53.640 59.530 54.000 ;
        RECT 50.850 52.530 51.110 52.850 ;
        RECT 47.170 51.510 47.430 51.830 ;
        RECT 42.110 47.090 42.370 47.410 ;
        RECT 38.420 46.555 38.700 46.925 ;
        RECT 37.510 41.310 37.770 41.630 ;
        RECT 37.570 34.520 37.710 41.310 ;
        RECT 38.490 34.520 38.630 46.555 ;
        RECT 40.730 46.070 40.990 46.390 ;
        RECT 39.810 44.030 40.070 44.350 ;
        RECT 39.870 34.520 40.010 44.030 ;
        RECT 40.790 34.520 40.930 46.070 ;
        RECT 42.170 34.520 42.310 47.090 ;
        RECT 43.490 46.750 43.750 47.070 ;
        RECT 43.550 34.520 43.690 46.750 ;
        RECT 47.230 34.520 47.370 51.510 ;
        RECT 48.090 46.410 48.350 46.730 ;
        RECT 48.150 34.520 48.290 46.410 ;
        RECT 50.910 34.520 51.050 52.530 ;
        RECT 53.150 52.190 53.410 52.510 ;
        RECT 53.210 34.520 53.350 52.190 ;
        RECT 56.830 50.490 57.090 50.810 ;
        RECT 55.450 47.430 55.710 47.750 ;
        RECT 55.510 34.520 55.650 47.430 ;
        RECT 56.890 34.520 57.030 50.490 ;
        RECT 60.050 50.150 60.310 50.470 ;
        RECT 58.050 48.200 59.530 48.680 ;
        RECT 58.050 42.760 59.530 43.240 ;
        RECT 60.110 39.330 60.250 50.150 ;
        RECT 58.270 39.190 60.250 39.330 ;
        RECT 58.270 34.520 58.410 39.190 ;
        RECT 60.570 34.520 60.710 54.000 ;
        RECT 61.890 49.470 62.150 49.790 ;
        RECT 61.950 34.520 62.090 49.470 ;
        RECT 64.710 46.810 64.850 54.000 ;
        RECT 65.170 52.850 65.310 54.000 ;
        RECT 65.110 52.530 65.370 52.850 ;
        RECT 72.930 52.530 73.190 52.850 ;
        RECT 72.470 50.490 72.730 50.810 ;
        RECT 72.530 50.325 72.670 50.490 ;
        RECT 72.460 49.955 72.740 50.325 ;
        RECT 66.490 49.130 66.750 49.450 ;
        RECT 69.240 49.275 69.520 49.645 ;
        RECT 63.790 46.730 64.850 46.810 ;
        RECT 63.730 46.670 64.850 46.730 ;
        RECT 63.730 46.410 63.990 46.670 ;
        RECT 65.570 44.370 65.830 44.690 ;
        RECT 62.810 43.690 63.070 44.010 ;
        RECT 62.870 34.520 63.010 43.690 ;
        RECT 65.630 34.520 65.770 44.370 ;
        RECT 66.550 34.520 66.690 49.130 ;
        RECT 69.310 34.520 69.450 49.275 ;
        RECT 70.170 48.790 70.430 49.110 ;
        RECT 70.230 34.520 70.370 48.790 ;
        RECT 72.990 34.520 73.130 52.530 ;
        RECT 73.910 34.520 74.050 54.000 ;
        RECT 76.670 34.520 76.810 54.000 ;
        RECT 77.530 51.510 77.790 51.830 ;
        RECT 77.060 50.635 77.340 51.005 ;
        RECT 77.130 37.290 77.270 50.635 ;
        RECT 77.590 42.650 77.730 51.510 ;
        RECT 77.990 49.810 78.250 50.130 ;
        RECT 78.910 49.810 79.170 50.130 ;
        RECT 78.050 49.530 78.190 49.810 ;
        RECT 78.970 49.645 79.110 49.810 ;
        RECT 78.050 49.390 78.650 49.530 ;
        RECT 78.510 47.410 78.650 49.390 ;
        RECT 78.900 49.275 79.180 49.645 ;
        RECT 78.450 47.090 78.710 47.410 ;
        RECT 78.510 45.030 78.650 47.090 ;
        RECT 78.450 44.710 78.710 45.030 ;
        RECT 77.530 42.330 77.790 42.650 ;
        RECT 77.130 37.150 77.730 37.290 ;
        RECT 77.590 34.520 77.730 37.150 ;
        RECT 80.350 34.520 80.490 54.000 ;
        RECT 80.810 50.130 80.950 54.000 ;
        RECT 81.730 52.170 81.870 54.000 ;
        RECT 85.410 52.510 85.550 54.000 ;
        RECT 85.350 52.190 85.610 52.510 ;
        RECT 81.670 51.850 81.930 52.170 ;
        RECT 86.790 50.470 86.930 54.000 ;
        RECT 86.730 50.150 86.990 50.470 ;
        RECT 80.750 49.810 81.010 50.130 ;
        RECT 87.250 49.700 87.390 54.000 ;
        RECT 88.170 53.190 88.310 54.000 ;
        RECT 88.110 52.870 88.370 53.190 ;
        RECT 84.420 49.275 84.700 49.645 ;
        RECT 86.330 49.560 87.390 49.700 ;
        RECT 81.200 48.595 81.480 48.965 ;
        RECT 81.270 34.520 81.410 48.595 ;
        RECT 83.970 47.770 84.230 48.090 ;
        RECT 84.030 34.520 84.170 47.770 ;
        RECT 84.490 37.290 84.630 49.275 ;
        RECT 86.330 49.110 86.470 49.560 ;
        RECT 86.270 48.790 86.530 49.110 ;
        RECT 87.190 48.790 87.450 49.110 ;
        RECT 84.890 46.410 85.150 46.730 ;
        RECT 84.950 42.310 85.090 46.410 ;
        RECT 85.350 46.070 85.610 46.390 ;
        RECT 86.270 46.070 86.530 46.390 ;
        RECT 85.410 43.670 85.550 46.070 ;
        RECT 85.350 43.350 85.610 43.670 ;
        RECT 84.890 41.990 85.150 42.310 ;
        RECT 86.330 41.970 86.470 46.070 ;
        RECT 86.270 41.650 86.530 41.970 ;
        RECT 87.250 41.290 87.390 48.790 ;
        RECT 89.090 47.410 89.230 54.000 ;
        RECT 89.030 47.090 89.290 47.410 ;
        RECT 89.550 45.030 89.690 54.000 ;
        RECT 89.950 51.510 90.210 51.830 ;
        RECT 90.010 49.790 90.150 51.510 ;
        RECT 89.950 49.470 90.210 49.790 ;
        RECT 90.470 47.070 90.610 54.000 ;
        RECT 91.390 49.790 91.530 54.000 ;
        RECT 92.770 53.530 92.910 54.000 ;
        RECT 92.710 53.210 92.970 53.530 ;
        RECT 91.790 52.530 92.050 52.850 ;
        RECT 91.850 50.130 91.990 52.530 ;
        RECT 91.790 49.810 92.050 50.130 ;
        RECT 91.330 49.470 91.590 49.790 ;
        RECT 90.870 49.130 91.130 49.450 ;
        RECT 90.930 48.170 91.070 49.130 ;
        RECT 90.930 48.030 91.990 48.170 ;
        RECT 91.850 47.750 91.990 48.030 ;
        RECT 91.790 47.430 92.050 47.750 ;
        RECT 91.330 47.090 91.590 47.410 ;
        RECT 90.410 46.750 90.670 47.070 ;
        RECT 89.490 44.710 89.750 45.030 ;
        RECT 90.860 44.515 91.140 44.885 ;
        RECT 90.870 44.370 91.130 44.515 ;
        RECT 87.190 40.970 87.450 41.290 ;
        RECT 88.570 39.610 88.830 39.930 ;
        RECT 84.490 37.150 85.090 37.290 ;
        RECT 84.950 34.520 85.090 37.150 ;
        RECT 88.630 34.520 88.770 39.610 ;
        RECT 91.390 34.520 91.530 47.090 ;
        RECT 93.230 47.070 93.370 54.000 ;
        RECT 93.690 50.325 93.830 54.000 ;
        RECT 93.620 49.955 93.900 50.325 ;
        RECT 93.170 46.810 93.430 47.070 ;
        RECT 93.170 46.750 94.290 46.810 ;
        RECT 93.230 46.670 94.290 46.750 ;
        RECT 92.710 46.070 92.970 46.390 ;
        RECT 92.770 37.290 92.910 46.070 ;
        RECT 94.150 44.690 94.290 46.670 ;
        RECT 94.090 44.370 94.350 44.690 ;
        RECT 92.310 37.150 92.910 37.290 ;
        RECT 92.310 34.520 92.450 37.150 ;
        RECT 95.070 34.520 95.210 54.000 ;
        RECT 95.990 34.520 96.130 54.000 ;
        RECT 96.840 49.955 97.120 50.325 ;
        RECT 96.910 49.110 97.050 49.955 ;
        RECT 96.850 48.790 97.110 49.110 ;
        RECT 97.370 45.030 97.510 54.000 ;
        RECT 97.310 44.710 97.570 45.030 ;
        RECT 97.830 39.330 97.970 54.000 ;
        RECT 99.140 53.355 99.420 53.725 ;
        RECT 99.210 53.190 99.350 53.355 ;
        RECT 99.150 52.870 99.410 53.190 ;
        RECT 100.130 52.850 100.270 54.000 ;
        RECT 98.690 52.530 98.950 52.850 ;
        RECT 100.070 52.530 100.330 52.850 ;
        RECT 98.750 50.810 98.890 52.530 ;
        RECT 100.590 50.810 100.730 54.000 ;
        RECT 98.690 50.490 98.950 50.810 ;
        RECT 100.530 50.490 100.790 50.810 ;
        RECT 99.610 50.040 99.870 50.130 ;
        RECT 99.210 49.900 99.870 50.040 ;
        RECT 99.210 48.090 99.350 49.900 ;
        RECT 99.610 49.810 99.870 49.900 ;
        RECT 99.150 47.770 99.410 48.090 ;
        RECT 98.220 47.235 98.500 47.605 ;
        RECT 98.290 46.390 98.430 47.235 ;
        RECT 98.230 46.070 98.490 46.390 ;
        RECT 100.530 44.600 100.790 44.690 ;
        RECT 101.050 44.600 101.190 54.000 ;
        RECT 101.970 45.030 102.110 54.000 ;
        RECT 103.350 53.725 103.490 54.000 ;
        RECT 103.280 53.355 103.560 53.725 ;
        RECT 103.280 52.675 103.560 53.045 ;
        RECT 102.370 46.410 102.630 46.730 ;
        RECT 101.910 44.710 102.170 45.030 ;
        RECT 100.530 44.460 101.190 44.600 ;
        RECT 100.530 44.370 100.790 44.460 ;
        RECT 97.830 39.190 98.890 39.330 ;
        RECT 98.750 34.520 98.890 39.190 ;
        RECT 102.430 34.520 102.570 46.410 ;
        RECT 103.350 34.520 103.490 52.675 ;
        RECT 104.730 46.390 104.870 54.000 ;
        RECT 105.650 47.750 105.790 54.000 ;
        RECT 106.110 50.470 106.250 54.000 ;
        RECT 107.490 52.850 107.630 54.000 ;
        RECT 107.430 52.530 107.690 52.850 ;
        RECT 108.410 51.830 108.550 54.000 ;
        RECT 108.350 51.510 108.610 51.830 ;
        RECT 108.870 51.005 109.010 54.000 ;
        RECT 108.800 50.635 109.080 51.005 ;
        RECT 106.050 50.150 106.310 50.470 ;
        RECT 106.050 49.470 106.310 49.790 ;
        RECT 105.590 47.430 105.850 47.750 ;
        RECT 106.110 47.070 106.250 49.470 ;
        RECT 108.870 49.110 109.010 50.635 ;
        RECT 108.810 48.790 109.070 49.110 ;
        RECT 109.330 48.170 109.470 54.000 ;
        RECT 109.790 51.685 109.930 54.000 ;
        RECT 109.720 51.315 110.000 51.685 ;
        RECT 109.790 48.965 109.930 51.315 ;
        RECT 109.720 48.595 110.000 48.965 ;
        RECT 106.970 47.770 107.230 48.090 ;
        RECT 109.330 48.030 109.930 48.170 ;
        RECT 106.050 46.750 106.310 47.070 ;
        RECT 104.670 46.070 104.930 46.390 ;
        RECT 106.050 38.930 106.310 39.250 ;
        RECT 106.110 34.520 106.250 38.930 ;
        RECT 107.030 34.520 107.170 47.770 ;
        RECT 109.790 34.520 109.930 48.030 ;
        RECT 110.250 45.030 110.390 54.000 ;
        RECT 110.640 51.995 110.920 52.365 ;
        RECT 110.190 44.710 110.450 45.030 ;
        RECT 110.710 34.520 110.850 51.995 ;
        RECT 111.630 40.610 111.770 54.000 ;
        RECT 112.090 50.130 112.230 54.000 ;
        RECT 113.470 52.510 113.610 54.000 ;
        RECT 113.410 52.190 113.670 52.510 ;
        RECT 114.330 52.190 114.590 52.510 ;
        RECT 114.390 51.685 114.530 52.190 ;
        RECT 114.320 51.315 114.600 51.685 ;
        RECT 112.030 49.810 112.290 50.130 ;
        RECT 114.780 49.955 115.060 50.325 ;
        RECT 112.490 49.470 112.750 49.790 ;
        RECT 112.550 47.070 112.690 49.470 ;
        RECT 114.320 49.275 114.600 49.645 ;
        RECT 112.490 46.750 112.750 47.070 ;
        RECT 112.950 46.410 113.210 46.730 ;
        RECT 111.570 40.290 111.830 40.610 ;
        RECT 113.010 34.520 113.150 46.410 ;
        RECT 114.390 34.520 114.530 49.275 ;
        RECT 114.850 47.410 114.990 49.955 ;
        RECT 114.790 47.090 115.050 47.410 ;
        RECT 115.770 46.730 115.910 54.000 ;
        RECT 116.230 48.965 116.370 54.000 ;
        RECT 116.160 48.595 116.440 48.965 ;
        RECT 115.710 46.410 115.970 46.730 ;
        RECT 115.250 44.370 115.510 44.690 ;
        RECT 115.310 42.650 115.450 44.370 ;
        RECT 115.250 42.330 115.510 42.650 ;
        RECT 116.690 34.520 116.830 54.000 ;
        RECT 117.150 39.590 117.290 54.000 ;
        RECT 117.610 42.650 117.750 54.000 ;
        RECT 118.070 47.410 118.210 54.000 ;
        RECT 118.010 47.090 118.270 47.410 ;
        RECT 118.470 47.090 118.730 47.410 ;
        RECT 118.530 44.350 118.670 47.090 ;
        RECT 118.990 46.730 119.130 54.000 ;
        RECT 119.390 51.510 119.650 51.830 ;
        RECT 119.450 48.965 119.590 51.510 ;
        RECT 119.380 48.595 119.660 48.965 ;
        RECT 119.390 47.660 119.650 47.750 ;
        RECT 119.910 47.660 120.050 54.000 ;
        RECT 120.370 50.130 120.510 54.000 ;
        RECT 121.750 52.850 121.890 54.000 ;
        RECT 121.690 52.530 121.950 52.850 ;
        RECT 120.310 49.810 120.570 50.130 ;
        RECT 119.390 47.520 120.050 47.660 ;
        RECT 119.390 47.430 119.650 47.520 ;
        RECT 120.310 47.430 120.570 47.750 ;
        RECT 119.390 46.750 119.650 47.070 ;
        RECT 118.930 46.410 119.190 46.730 ;
        RECT 118.470 44.030 118.730 44.350 ;
        RECT 119.450 44.205 119.590 46.750 ;
        RECT 117.550 42.330 117.810 42.650 ;
        RECT 118.530 40.950 118.670 44.030 ;
        RECT 119.380 43.835 119.660 44.205 ;
        RECT 119.390 43.690 119.650 43.835 ;
        RECT 119.450 43.535 119.590 43.690 ;
        RECT 120.370 43.670 120.510 47.430 ;
        RECT 120.770 46.410 121.030 46.730 ;
        RECT 120.310 43.350 120.570 43.670 ;
        RECT 118.470 40.630 118.730 40.950 ;
        RECT 117.090 39.270 117.350 39.590 ;
        RECT 118.010 39.270 118.270 39.590 ;
        RECT 120.830 39.330 120.970 46.410 ;
        RECT 123.130 46.300 123.270 54.000 ;
        RECT 118.070 34.520 118.210 39.270 ;
        RECT 120.370 39.190 120.970 39.330 ;
        RECT 121.750 46.160 123.270 46.300 ;
        RECT 120.370 34.520 120.510 39.190 ;
        RECT 121.750 34.520 121.890 46.160 ;
        RECT 123.590 45.030 123.730 54.000 ;
        RECT 123.530 44.710 123.790 45.030 ;
        RECT 123.530 43.350 123.790 43.670 ;
        RECT 123.590 40.270 123.730 43.350 ;
        RECT 123.530 39.950 123.790 40.270 ;
        RECT 124.050 34.520 124.190 54.000 ;
        RECT 125.830 52.190 126.090 52.510 ;
        RECT 125.370 51.850 125.630 52.170 ;
        RECT 125.430 34.520 125.570 51.850 ;
        RECT 125.890 51.685 126.030 52.190 ;
        RECT 125.820 51.315 126.100 51.685 ;
        RECT 125.890 49.790 126.030 51.315 ;
        RECT 126.350 50.130 126.490 54.000 ;
        RECT 126.290 49.810 126.550 50.130 ;
        RECT 125.830 49.470 126.090 49.790 ;
        RECT 125.890 47.750 126.030 49.470 ;
        RECT 125.830 47.430 126.090 47.750 ;
        RECT 126.810 39.250 126.950 54.000 ;
        RECT 127.730 53.045 127.870 54.000 ;
        RECT 127.660 52.675 127.940 53.045 ;
        RECT 127.730 52.170 127.870 52.675 ;
        RECT 127.670 51.850 127.930 52.170 ;
        RECT 128.190 45.370 128.330 54.000 ;
        RECT 128.650 52.510 128.790 54.000 ;
        RECT 128.590 52.190 128.850 52.510 ;
        RECT 128.590 47.320 128.850 47.410 ;
        RECT 129.110 47.320 129.250 54.000 ;
        RECT 128.590 47.180 129.250 47.320 ;
        RECT 128.590 47.090 128.850 47.180 ;
        RECT 128.130 45.050 128.390 45.370 ;
        RECT 127.670 44.885 127.930 45.030 ;
        RECT 127.660 44.515 127.940 44.885 ;
        RECT 129.050 44.205 129.310 44.350 ;
        RECT 129.040 43.835 129.320 44.205 ;
        RECT 126.750 38.930 127.010 39.250 ;
        RECT 130.030 38.570 130.170 54.000 ;
        RECT 130.950 50.470 131.090 54.000 ;
        RECT 130.890 50.150 131.150 50.470 ;
        RECT 130.430 49.470 130.690 49.790 ;
        RECT 130.490 39.930 130.630 49.470 ;
        RECT 130.950 47.605 131.090 50.150 ;
        RECT 130.880 47.235 131.160 47.605 ;
        RECT 130.430 39.610 130.690 39.930 ;
        RECT 127.670 38.250 127.930 38.570 ;
        RECT 129.970 38.250 130.230 38.570 ;
        RECT 127.730 34.520 127.870 38.250 ;
        RECT 131.410 34.520 131.550 54.000 ;
        RECT 132.270 52.190 132.530 52.510 ;
        RECT 132.330 51.685 132.470 52.190 ;
        RECT 132.260 51.315 132.540 51.685 ;
        RECT 131.810 43.350 132.070 43.670 ;
        RECT 131.870 39.930 132.010 43.350 ;
        RECT 131.810 39.610 132.070 39.930 ;
        RECT 132.790 34.520 132.930 54.000 ;
        RECT 133.250 53.190 133.390 54.000 ;
        RECT 133.190 52.870 133.450 53.190 ;
        RECT 133.190 51.510 133.450 51.830 ;
        RECT 133.250 50.810 133.390 51.510 ;
        RECT 133.190 50.490 133.450 50.810 ;
        RECT 133.710 50.130 133.850 54.000 ;
        RECT 136.870 51.850 137.130 52.170 ;
        RECT 134.850 50.920 136.330 51.400 ;
        RECT 133.650 49.810 133.910 50.130 ;
        RECT 134.570 49.470 134.830 49.790 ;
        RECT 134.630 47.750 134.770 49.470 ;
        RECT 136.400 48.595 136.680 48.965 ;
        RECT 134.570 47.430 134.830 47.750 ;
        RECT 134.850 45.480 136.330 45.960 ;
        RECT 135.950 44.370 136.210 44.690 ;
        RECT 136.010 38.910 136.150 44.370 ;
        RECT 135.950 38.590 136.210 38.910 ;
        RECT 136.470 34.520 136.610 48.595 ;
        RECT 136.930 47.410 137.070 51.850 ;
        RECT 136.870 47.090 137.130 47.410 ;
        RECT 136.930 44.690 137.070 47.090 ;
        RECT 137.850 46.730 137.990 54.000 ;
        RECT 138.770 53.530 138.910 54.000 ;
        RECT 138.710 53.210 138.970 53.530 ;
        RECT 139.230 53.190 139.370 54.000 ;
        RECT 139.170 52.870 139.430 53.190 ;
        RECT 139.690 52.510 139.830 54.000 ;
        RECT 139.630 52.190 139.890 52.510 ;
        RECT 138.710 51.510 138.970 51.830 ;
        RECT 137.790 46.410 138.050 46.730 ;
        RECT 136.870 44.370 137.130 44.690 ;
        RECT 137.330 44.370 137.590 44.690 ;
        RECT 136.870 43.690 137.130 44.010 ;
        RECT 136.930 41.370 137.070 43.690 ;
        RECT 137.390 42.310 137.530 44.370 ;
        RECT 137.330 41.990 137.590 42.310 ;
        RECT 137.790 41.990 138.050 42.310 ;
        RECT 137.850 41.370 137.990 41.990 ;
        RECT 136.930 41.230 137.990 41.370 ;
        RECT 136.930 40.950 137.070 41.230 ;
        RECT 136.870 40.630 137.130 40.950 ;
        RECT 138.770 34.520 138.910 51.510 ;
        RECT 139.690 50.130 139.830 52.190 ;
        RECT 140.150 52.170 140.290 54.000 ;
        RECT 141.930 52.530 142.190 52.850 ;
        RECT 140.090 51.850 140.350 52.170 ;
        RECT 141.990 50.470 142.130 52.530 ;
        RECT 141.930 50.150 142.190 50.470 ;
        RECT 139.630 49.810 139.890 50.130 ;
        RECT 140.080 47.235 140.360 47.605 ;
        RECT 140.150 34.520 140.290 47.235 ;
        RECT 143.830 47.070 143.970 54.000 ;
        RECT 145.670 53.725 145.810 54.000 ;
        RECT 145.150 53.210 145.410 53.530 ;
        RECT 145.600 53.355 145.880 53.725 ;
        RECT 145.210 47.070 145.350 53.210 ;
        RECT 143.770 46.750 144.030 47.070 ;
        RECT 145.150 46.750 145.410 47.070 ;
        RECT 141.010 46.070 141.270 46.390 ;
        RECT 142.390 46.070 142.650 46.390 ;
        RECT 141.070 45.370 141.210 46.070 ;
        RECT 141.010 45.050 141.270 45.370 ;
        RECT 142.450 34.520 142.590 46.070 ;
        RECT 143.770 40.630 144.030 40.950 ;
        RECT 143.830 34.520 143.970 40.630 ;
        RECT 146.130 34.520 146.270 54.000 ;
        RECT 146.520 51.995 146.800 52.365 ;
        RECT 146.590 48.090 146.730 51.995 ;
        RECT 147.970 50.130 148.110 54.000 ;
        RECT 148.430 53.190 148.570 54.000 ;
        RECT 148.370 52.870 148.630 53.190 ;
        RECT 148.890 50.470 149.030 54.000 ;
        RECT 149.750 52.190 150.010 52.510 ;
        RECT 150.730 52.365 150.870 54.000 ;
        RECT 152.110 53.530 152.250 54.000 ;
        RECT 152.570 53.530 152.710 54.000 ;
        RECT 152.050 53.210 152.310 53.530 ;
        RECT 152.510 53.210 152.770 53.530 ;
        RECT 148.830 50.150 149.090 50.470 ;
        RECT 147.910 49.810 148.170 50.130 ;
        RECT 149.810 48.090 149.950 52.190 ;
        RECT 150.660 51.995 150.940 52.365 ;
        RECT 150.730 49.110 150.870 51.995 ;
        RECT 152.570 51.685 152.710 53.210 ;
        RECT 152.500 51.315 152.780 51.685 ;
        RECT 150.670 48.790 150.930 49.110 ;
        RECT 153.030 49.020 153.170 54.000 ;
        RECT 153.950 52.850 154.090 54.000 ;
        RECT 153.890 52.530 154.150 52.850 ;
        RECT 154.870 52.170 155.010 54.000 ;
        RECT 154.810 51.850 155.070 52.170 ;
        RECT 154.800 51.315 155.080 51.685 ;
        RECT 153.890 49.470 154.150 49.790 ;
        RECT 153.950 49.020 154.090 49.470 ;
        RECT 151.120 48.595 151.400 48.965 ;
        RECT 153.030 48.880 154.090 49.020 ;
        RECT 146.530 47.770 146.790 48.090 ;
        RECT 149.750 47.770 150.010 48.090 ;
        RECT 147.450 47.430 147.710 47.750 ;
        RECT 147.510 47.070 147.650 47.430 ;
        RECT 147.450 46.750 147.710 47.070 ;
        RECT 147.450 38.250 147.710 38.570 ;
        RECT 147.510 34.520 147.650 38.250 ;
        RECT 149.750 37.230 150.010 37.550 ;
        RECT 149.810 34.520 149.950 37.230 ;
        RECT 151.190 34.520 151.330 48.595 ;
        RECT 153.430 47.770 153.690 48.090 ;
        RECT 153.490 34.520 153.630 47.770 ;
        RECT 153.950 47.410 154.090 48.880 ;
        RECT 153.890 47.090 154.150 47.410 ;
        RECT 153.950 44.690 154.090 47.090 ;
        RECT 153.890 44.370 154.150 44.690 ;
        RECT 154.870 40.950 155.010 51.315 ;
        RECT 155.330 50.130 155.470 54.000 ;
        RECT 155.270 49.810 155.530 50.130 ;
        RECT 154.810 40.630 155.070 40.950 ;
        RECT 155.790 39.930 155.930 54.000 ;
        RECT 156.710 52.850 156.850 54.000 ;
        RECT 156.650 52.530 156.910 52.850 ;
        RECT 157.630 52.250 157.770 54.000 ;
        RECT 156.250 52.110 157.770 52.250 ;
        RECT 156.250 44.350 156.390 52.110 ;
        RECT 158.020 51.995 158.300 52.365 ;
        RECT 157.110 50.490 157.370 50.810 ;
        RECT 156.640 49.275 156.920 49.645 ;
        RECT 156.710 46.390 156.850 49.275 ;
        RECT 156.650 46.070 156.910 46.390 ;
        RECT 156.190 44.030 156.450 44.350 ;
        RECT 156.650 43.690 156.910 44.010 ;
        RECT 156.710 42.650 156.850 43.690 ;
        RECT 156.650 42.330 156.910 42.650 ;
        RECT 155.730 39.610 155.990 39.930 ;
        RECT 154.810 37.910 155.070 38.230 ;
        RECT 154.870 34.520 155.010 37.910 ;
        RECT 157.170 34.520 157.310 50.490 ;
        RECT 158.090 47.605 158.230 51.995 ;
        RECT 158.550 48.000 158.690 54.000 ;
        RECT 158.940 52.675 159.220 53.045 ;
        RECT 158.950 52.530 159.210 52.675 ;
        RECT 159.470 50.325 159.610 54.000 ;
        RECT 159.400 49.955 159.680 50.325 ;
        RECT 158.550 47.860 159.150 48.000 ;
        RECT 159.010 47.605 159.150 47.860 ;
        RECT 158.020 47.235 158.300 47.605 ;
        RECT 158.940 47.235 159.220 47.605 ;
        RECT 159.470 46.130 159.610 49.955 ;
        RECT 160.390 47.070 160.530 54.000 ;
        RECT 160.330 46.750 160.590 47.070 ;
        RECT 160.330 46.130 160.590 46.390 ;
        RECT 159.470 46.070 160.590 46.130 ;
        RECT 159.470 45.990 160.530 46.070 ;
        RECT 158.490 38.930 158.750 39.250 ;
        RECT 158.550 34.520 158.690 38.930 ;
        RECT 160.850 34.520 160.990 54.000 ;
        RECT 162.230 51.005 162.370 54.000 ;
        RECT 162.160 50.635 162.440 51.005 ;
        RECT 162.690 50.810 162.830 54.000 ;
        RECT 162.630 50.490 162.890 50.810 ;
        RECT 162.170 50.150 162.430 50.470 ;
        RECT 162.230 34.520 162.370 50.150 ;
        RECT 163.150 50.130 163.290 54.000 ;
        RECT 163.610 53.530 163.750 54.000 ;
        RECT 163.550 53.210 163.810 53.530 ;
        RECT 164.990 50.325 165.130 54.000 ;
        RECT 163.090 49.810 163.350 50.130 ;
        RECT 164.920 49.955 165.200 50.325 ;
        RECT 162.630 44.710 162.890 45.030 ;
        RECT 162.690 40.950 162.830 44.710 ;
        RECT 163.090 43.350 163.350 43.670 ;
        RECT 164.010 43.350 164.270 43.670 ;
        RECT 163.150 40.950 163.290 43.350 ;
        RECT 162.630 40.630 162.890 40.950 ;
        RECT 163.090 40.630 163.350 40.950 ;
        RECT 164.070 39.590 164.210 43.350 ;
        RECT 164.470 41.650 164.730 41.970 ;
        RECT 164.010 39.270 164.270 39.590 ;
        RECT 164.530 34.520 164.670 41.650 ;
        RECT 165.450 39.590 165.590 54.000 ;
        RECT 167.290 47.750 167.430 54.000 ;
        RECT 167.230 47.430 167.490 47.750 ;
        RECT 165.850 46.070 166.110 46.390 ;
        RECT 165.390 39.270 165.650 39.590 ;
        RECT 165.910 34.520 166.050 46.070 ;
        RECT 168.210 34.520 168.350 54.000 ;
        RECT 169.130 40.270 169.270 54.000 ;
        RECT 170.440 52.675 170.720 53.045 ;
        RECT 170.510 52.510 170.650 52.675 ;
        RECT 170.450 52.190 170.710 52.510 ;
        RECT 170.970 50.130 171.110 54.000 ;
        RECT 171.890 52.850 172.030 54.000 ;
        RECT 171.830 52.530 172.090 52.850 ;
        RECT 170.910 49.810 171.170 50.130 ;
        RECT 170.910 47.090 171.170 47.410 ;
        RECT 169.070 39.950 169.330 40.270 ;
        RECT 170.970 39.250 171.110 47.090 ;
        RECT 172.350 45.030 172.490 54.000 ;
        RECT 172.290 44.710 172.550 45.030 ;
        RECT 172.810 39.250 172.950 54.000 ;
        RECT 174.650 44.690 174.790 54.000 ;
        RECT 174.590 44.370 174.850 44.690 ;
        RECT 174.130 44.030 174.390 44.350 ;
        RECT 174.190 40.270 174.330 44.030 ;
        RECT 174.130 39.950 174.390 40.270 ;
        RECT 170.910 38.930 171.170 39.250 ;
        RECT 172.750 38.930 173.010 39.250 ;
        RECT 171.830 38.590 172.090 38.910 ;
        RECT 171.890 34.520 172.030 38.590 ;
        RECT 175.110 38.230 175.250 54.000 ;
        RECT 175.970 49.470 176.230 49.790 ;
        RECT 176.490 49.645 176.630 54.000 ;
        RECT 175.510 40.970 175.770 41.290 ;
        RECT 175.050 37.910 175.310 38.230 ;
        RECT 175.570 34.520 175.710 40.970 ;
        RECT 176.030 38.570 176.170 49.470 ;
        RECT 176.420 49.275 176.700 49.645 ;
        RECT 176.950 48.090 177.090 54.000 ;
        RECT 177.870 53.045 178.010 54.000 ;
        RECT 177.800 52.675 178.080 53.045 ;
        RECT 176.890 47.770 177.150 48.090 ;
        RECT 177.870 47.070 178.010 52.675 ;
        RECT 178.330 52.170 178.470 54.000 ;
        RECT 178.730 52.530 178.990 52.850 ;
        RECT 178.270 51.850 178.530 52.170 ;
        RECT 177.810 46.750 178.070 47.070 ;
        RECT 178.270 44.370 178.530 44.690 ;
        RECT 178.330 42.310 178.470 44.370 ;
        RECT 178.270 41.990 178.530 42.310 ;
        RECT 175.970 38.250 176.230 38.570 ;
        RECT 178.790 37.550 178.930 52.530 ;
        RECT 179.710 44.350 179.850 54.000 ;
        RECT 183.850 52.510 183.990 54.000 ;
        RECT 184.310 53.530 184.450 54.000 ;
        RECT 184.250 53.210 184.510 53.530 ;
        RECT 181.950 52.190 182.210 52.510 ;
        RECT 183.790 52.190 184.050 52.510 ;
        RECT 182.010 50.130 182.150 52.190 ;
        RECT 181.950 49.810 182.210 50.130 ;
        RECT 184.770 48.090 184.910 54.000 ;
        RECT 185.230 52.365 185.370 54.000 ;
        RECT 185.160 51.995 185.440 52.365 ;
        RECT 185.170 48.790 185.430 49.110 ;
        RECT 184.710 47.770 184.970 48.090 ;
        RECT 184.710 46.980 184.970 47.070 ;
        RECT 185.230 46.980 185.370 48.790 ;
        RECT 184.710 46.840 185.370 46.980 ;
        RECT 184.710 46.750 184.970 46.840 ;
        RECT 184.770 44.690 184.910 46.750 ;
        RECT 186.150 45.370 186.290 54.000 ;
        RECT 186.610 53.530 186.750 54.000 ;
        RECT 186.550 53.210 186.810 53.530 ;
        RECT 187.070 50.040 187.210 54.000 ;
        RECT 188.450 53.530 188.590 54.000 ;
        RECT 188.390 53.210 188.650 53.530 ;
        RECT 188.910 51.685 189.050 54.000 ;
        RECT 188.840 51.315 189.120 51.685 ;
        RECT 189.760 51.315 190.040 51.685 ;
        RECT 186.610 49.900 187.210 50.040 ;
        RECT 186.090 45.050 186.350 45.370 ;
        RECT 185.170 44.885 185.430 45.030 ;
        RECT 184.710 44.370 184.970 44.690 ;
        RECT 185.160 44.515 185.440 44.885 ;
        RECT 179.650 44.030 179.910 44.350 ;
        RECT 179.190 39.610 179.450 39.930 ;
        RECT 178.730 37.230 178.990 37.550 ;
        RECT 179.250 34.520 179.390 39.610 ;
        RECT 186.610 34.520 186.750 49.900 ;
        RECT 188.850 48.790 189.110 49.110 ;
        RECT 188.910 48.285 189.050 48.790 ;
        RECT 188.840 47.915 189.120 48.285 ;
        RECT 189.830 47.750 189.970 51.315 ;
        RECT 189.770 47.430 190.030 47.750 ;
        RECT 190.290 34.520 190.430 54.000 ;
        RECT 190.750 52.850 190.890 54.000 ;
        RECT 190.690 52.530 190.950 52.850 ;
        RECT 190.680 51.995 190.960 52.365 ;
        RECT 190.690 51.850 190.950 51.995 ;
        RECT 191.210 49.790 191.350 54.000 ;
        RECT 191.610 51.510 191.870 51.830 ;
        RECT 191.670 50.470 191.810 51.510 ;
        RECT 191.610 50.150 191.870 50.470 ;
        RECT 192.130 50.130 192.270 54.000 ;
        RECT 192.070 49.810 192.330 50.130 ;
        RECT 191.150 49.470 191.410 49.790 ;
        RECT 191.210 45.370 191.350 49.470 ;
        RECT 193.510 49.450 193.650 54.000 ;
        RECT 194.430 50.130 194.570 54.000 ;
        RECT 194.820 51.995 195.100 52.365 ;
        RECT 194.890 50.810 195.030 51.995 ;
        RECT 194.830 50.490 195.090 50.810 ;
        RECT 194.370 49.810 194.630 50.130 ;
        RECT 195.350 49.645 195.490 54.000 ;
        RECT 196.270 52.365 196.410 54.000 ;
        RECT 196.200 51.995 196.480 52.365 ;
        RECT 193.450 49.130 193.710 49.450 ;
        RECT 195.280 49.275 195.560 49.645 ;
        RECT 194.830 46.750 195.090 47.070 ;
        RECT 194.890 46.245 195.030 46.750 ;
        RECT 196.730 46.730 196.870 54.000 ;
        RECT 197.190 51.830 197.330 54.000 ;
        RECT 197.590 52.190 197.850 52.510 ;
        RECT 197.130 51.510 197.390 51.830 ;
        RECT 197.650 49.790 197.790 52.190 ;
        RECT 199.490 51.685 199.630 54.000 ;
        RECT 201.260 51.995 201.540 52.365 ;
        RECT 199.420 51.315 199.700 51.685 ;
        RECT 197.590 49.470 197.850 49.790 ;
        RECT 197.130 48.790 197.390 49.110 ;
        RECT 197.590 48.790 197.850 49.110 ;
        RECT 197.190 47.070 197.330 48.790 ;
        RECT 197.130 46.750 197.390 47.070 ;
        RECT 196.670 46.410 196.930 46.730 ;
        RECT 194.820 45.875 195.100 46.245 ;
        RECT 191.150 45.050 191.410 45.370 ;
        RECT 193.900 45.195 194.180 45.565 ;
        RECT 193.970 34.520 194.110 45.195 ;
        RECT 197.650 34.520 197.790 48.790 ;
        RECT 199.490 46.245 199.630 51.315 ;
        RECT 201.330 47.490 201.470 51.995 ;
        RECT 201.790 48.965 201.930 54.000 ;
        RECT 202.250 49.110 202.390 54.000 ;
        RECT 202.650 52.190 202.910 52.510 ;
        RECT 202.710 49.450 202.850 52.190 ;
        RECT 202.650 49.130 202.910 49.450 ;
        RECT 201.720 48.595 202.000 48.965 ;
        RECT 202.190 48.790 202.450 49.110 ;
        RECT 203.110 48.790 203.370 49.110 ;
        RECT 201.790 48.170 201.930 48.595 ;
        RECT 203.170 48.170 203.310 48.790 ;
        RECT 201.790 48.030 203.310 48.170 ;
        RECT 203.630 48.170 203.770 54.000 ;
        RECT 204.030 51.685 204.290 51.830 ;
        RECT 204.020 51.315 204.300 51.685 ;
        RECT 205.410 51.510 205.670 51.830 ;
        RECT 205.470 50.130 205.610 51.510 ;
        RECT 205.410 49.810 205.670 50.130 ;
        RECT 205.410 48.790 205.670 49.110 ;
        RECT 203.630 48.030 205.150 48.170 ;
        RECT 201.330 47.350 202.390 47.490 ;
        RECT 202.250 46.730 202.390 47.350 ;
        RECT 202.190 46.410 202.450 46.730 ;
        RECT 199.420 45.875 199.700 46.245 ;
        RECT 201.270 41.650 201.530 41.970 ;
        RECT 201.330 34.520 201.470 41.650 ;
        RECT 205.010 34.520 205.150 48.030 ;
        RECT 205.470 47.410 205.610 48.790 ;
        RECT 205.410 47.090 205.670 47.410 ;
        RECT 205.930 44.690 206.070 54.000 ;
        RECT 205.870 44.370 206.130 44.690 ;
        RECT 207.770 44.350 207.910 54.000 ;
        RECT 208.620 51.995 208.900 52.365 ;
        RECT 208.170 44.370 208.430 44.690 ;
        RECT 207.710 44.030 207.970 44.350 ;
        RECT 208.230 41.290 208.370 44.370 ;
        RECT 208.170 40.970 208.430 41.290 ;
        RECT 208.690 34.520 208.830 51.995 ;
        RECT 210.070 45.030 210.210 54.000 ;
        RECT 210.990 53.530 211.130 54.000 ;
        RECT 211.650 53.640 213.130 54.000 ;
        RECT 210.930 53.210 211.190 53.530 ;
        RECT 212.310 52.530 212.570 52.850 ;
        RECT 212.370 51.685 212.510 52.530 ;
        RECT 213.290 52.510 213.430 54.000 ;
        RECT 214.140 52.675 214.420 53.045 ;
        RECT 213.230 52.190 213.490 52.510 ;
        RECT 212.300 51.315 212.580 51.685 ;
        RECT 210.460 50.635 210.740 51.005 ;
        RECT 210.530 49.790 210.670 50.635 ;
        RECT 213.290 50.130 213.430 52.190 ;
        RECT 214.210 51.005 214.350 52.675 ;
        RECT 213.690 50.490 213.950 50.810 ;
        RECT 214.140 50.635 214.420 51.005 ;
        RECT 213.230 49.810 213.490 50.130 ;
        RECT 210.470 49.470 210.730 49.790 ;
        RECT 211.650 48.200 213.130 48.680 ;
        RECT 213.750 48.090 213.890 50.490 ;
        RECT 213.690 47.770 213.950 48.090 ;
        RECT 214.210 47.070 214.350 50.635 ;
        RECT 214.610 49.810 214.870 50.130 ;
        RECT 214.670 49.645 214.810 49.810 ;
        RECT 214.600 49.275 214.880 49.645 ;
        RECT 214.150 46.750 214.410 47.070 ;
        RECT 214.610 46.300 214.870 46.390 ;
        RECT 215.130 46.300 215.270 54.000 ;
        RECT 215.590 49.020 215.730 54.000 ;
        RECT 216.050 51.685 216.190 54.000 ;
        RECT 215.980 51.315 216.260 51.685 ;
        RECT 215.590 48.880 216.190 49.020 ;
        RECT 214.610 46.160 215.270 46.300 ;
        RECT 214.610 46.070 214.870 46.160 ;
        RECT 210.010 44.710 210.270 45.030 ;
        RECT 215.070 44.370 215.330 44.690 ;
        RECT 213.690 43.690 213.950 44.010 ;
        RECT 211.650 42.760 213.130 43.240 ;
        RECT 213.750 42.650 213.890 43.690 ;
        RECT 215.130 42.650 215.270 44.370 ;
        RECT 213.690 42.330 213.950 42.650 ;
        RECT 215.070 42.330 215.330 42.650 ;
        RECT 216.050 34.520 216.190 48.880 ;
        RECT 216.510 45.370 216.650 54.000 ;
        RECT 217.830 48.790 218.090 49.110 ;
        RECT 217.890 47.750 218.030 48.790 ;
        RECT 217.830 47.430 218.090 47.750 ;
        RECT 218.350 47.410 218.490 54.000 ;
        RECT 219.270 53.530 219.410 54.000 ;
        RECT 219.210 53.210 219.470 53.530 ;
        RECT 219.730 50.130 219.870 54.000 ;
        RECT 220.190 52.510 220.330 54.000 ;
        RECT 220.130 52.190 220.390 52.510 ;
        RECT 219.670 49.810 219.930 50.130 ;
        RECT 219.670 47.770 219.930 48.090 ;
        RECT 219.210 47.430 219.470 47.750 ;
        RECT 218.290 47.090 218.550 47.410 ;
        RECT 216.450 45.050 216.710 45.370 ;
        RECT 219.270 45.030 219.410 47.430 ;
        RECT 219.210 44.710 219.470 45.030 ;
        RECT 216.450 44.370 216.710 44.690 ;
        RECT 216.510 43.670 216.650 44.370 ;
        RECT 216.450 43.350 216.710 43.670 ;
        RECT 219.730 34.520 219.870 47.770 ;
        RECT 220.120 47.235 220.400 47.605 ;
        RECT 220.190 47.070 220.330 47.235 ;
        RECT 220.130 46.750 220.390 47.070 ;
        RECT 220.650 40.270 220.790 54.000 ;
        RECT 221.570 45.280 221.710 54.000 ;
        RECT 223.410 49.450 223.550 54.000 ;
        RECT 223.350 49.130 223.610 49.450 ;
        RECT 223.870 48.090 224.010 54.000 ;
        RECT 223.810 47.770 224.070 48.090 ;
        RECT 221.110 45.140 221.710 45.280 ;
        RECT 221.110 44.690 221.250 45.140 ;
        RECT 221.050 44.370 221.310 44.690 ;
        RECT 221.510 44.370 221.770 44.690 ;
        RECT 221.570 42.650 221.710 44.370 ;
        RECT 221.970 43.350 222.230 43.670 ;
        RECT 222.030 42.650 222.170 43.350 ;
        RECT 221.510 42.330 221.770 42.650 ;
        RECT 221.970 42.330 222.230 42.650 ;
        RECT 222.950 42.165 224.010 42.220 ;
        RECT 222.950 42.080 224.080 42.165 ;
        RECT 220.590 39.950 220.850 40.270 ;
        RECT 222.950 38.910 223.090 42.080 ;
        RECT 223.800 41.795 224.080 42.080 ;
        RECT 224.330 41.370 224.470 54.000 ;
        RECT 225.180 52.675 225.460 53.045 ;
        RECT 225.250 51.830 225.390 52.675 ;
        RECT 225.190 51.510 225.450 51.830 ;
        RECT 224.730 49.810 224.990 50.130 ;
        RECT 224.790 48.090 224.930 49.810 ;
        RECT 225.710 49.645 225.850 54.000 ;
        RECT 225.640 49.275 225.920 49.645 ;
        RECT 224.730 47.770 224.990 48.090 ;
        RECT 226.170 45.370 226.310 54.000 ;
        RECT 226.630 52.510 226.770 54.000 ;
        RECT 226.570 52.190 226.830 52.510 ;
        RECT 226.630 47.750 226.770 52.190 ;
        RECT 227.090 51.830 227.230 54.000 ;
        RECT 227.030 51.510 227.290 51.830 ;
        RECT 227.030 49.470 227.290 49.790 ;
        RECT 226.570 47.430 226.830 47.750 ;
        RECT 226.110 45.050 226.370 45.370 ;
        RECT 223.410 41.230 224.470 41.370 ;
        RECT 222.890 38.590 223.150 38.910 ;
        RECT 223.410 34.520 223.550 41.230 ;
        RECT 227.090 34.520 227.230 49.470 ;
        RECT 227.550 46.730 227.690 54.000 ;
        RECT 227.490 46.410 227.750 46.730 ;
        RECT 228.010 44.770 228.150 54.000 ;
        RECT 228.470 49.110 228.610 54.000 ;
        RECT 228.870 53.045 229.130 53.190 ;
        RECT 228.860 52.675 229.140 53.045 ;
        RECT 228.870 52.190 229.130 52.510 ;
        RECT 228.930 50.130 229.070 52.190 ;
        RECT 230.250 51.850 230.510 52.170 ;
        RECT 228.870 49.810 229.130 50.130 ;
        RECT 228.410 48.790 228.670 49.110 ;
        RECT 228.410 47.430 228.670 47.750 ;
        RECT 228.470 47.070 228.610 47.430 ;
        RECT 230.310 47.410 230.450 51.850 ;
        RECT 230.710 50.325 230.970 50.470 ;
        RECT 230.700 49.955 230.980 50.325 ;
        RECT 230.710 47.770 230.970 48.090 ;
        RECT 231.160 47.915 231.440 48.285 ;
        RECT 230.770 47.410 230.910 47.770 ;
        RECT 230.250 47.090 230.510 47.410 ;
        RECT 230.710 47.090 230.970 47.410 ;
        RECT 228.410 46.750 228.670 47.070 ;
        RECT 231.230 46.730 231.370 47.915 ;
        RECT 231.630 47.090 231.890 47.410 ;
        RECT 231.690 46.730 231.830 47.090 ;
        RECT 231.170 46.410 231.430 46.730 ;
        RECT 231.630 46.410 231.890 46.730 ;
        RECT 228.410 46.070 228.670 46.390 ;
        RECT 228.470 45.565 228.610 46.070 ;
        RECT 228.400 45.195 228.680 45.565 ;
        RECT 232.150 45.370 232.290 54.000 ;
        RECT 232.090 45.050 232.350 45.370 ;
        RECT 228.010 44.690 228.610 44.770 ;
        RECT 228.010 44.630 228.670 44.690 ;
        RECT 228.410 44.370 228.670 44.630 ;
        RECT 229.780 44.515 230.060 44.885 ;
        RECT 229.790 44.370 230.050 44.515 ;
        RECT 228.470 40.270 228.610 44.370 ;
        RECT 230.710 44.030 230.970 44.350 ;
        RECT 230.770 40.610 230.910 44.030 ;
        RECT 232.610 44.010 232.750 54.000 ;
        RECT 233.070 47.410 233.210 54.000 ;
        RECT 233.010 47.090 233.270 47.410 ;
        RECT 233.070 44.350 233.210 47.090 ;
        RECT 233.530 46.730 233.670 54.000 ;
        RECT 234.450 48.850 234.590 54.000 ;
        RECT 234.910 49.790 235.050 54.000 ;
        RECT 235.370 52.510 235.510 54.000 ;
        RECT 235.310 52.190 235.570 52.510 ;
        RECT 235.830 52.170 235.970 54.000 ;
        RECT 235.770 51.850 236.030 52.170 ;
        RECT 236.220 51.995 236.500 52.365 ;
        RECT 236.290 50.720 236.430 51.995 ;
        RECT 235.830 50.580 236.430 50.720 ;
        RECT 234.850 49.470 235.110 49.790 ;
        RECT 235.830 49.450 235.970 50.580 ;
        RECT 235.770 49.130 236.030 49.450 ;
        RECT 233.990 48.710 234.590 48.850 ;
        RECT 233.990 48.090 234.130 48.710 ;
        RECT 233.930 47.770 234.190 48.090 ;
        RECT 234.390 47.770 234.650 48.090 ;
        RECT 234.840 47.915 235.120 48.285 ;
        RECT 233.990 46.730 234.130 47.770 ;
        RECT 233.470 46.410 233.730 46.730 ;
        RECT 233.930 46.410 234.190 46.730 ;
        RECT 233.010 44.030 233.270 44.350 ;
        RECT 232.550 43.690 232.810 44.010 ;
        RECT 233.070 42.310 233.210 44.030 ;
        RECT 233.010 41.990 233.270 42.310 ;
        RECT 230.710 40.290 230.970 40.610 ;
        RECT 228.410 39.950 228.670 40.270 ;
        RECT 230.710 39.610 230.970 39.930 ;
        RECT 230.770 34.520 230.910 39.610 ;
        RECT 234.450 34.520 234.590 47.770 ;
        RECT 234.910 47.410 235.050 47.915 ;
        RECT 234.850 47.090 235.110 47.410 ;
        RECT 235.830 44.690 235.970 49.130 ;
        RECT 235.770 44.370 236.030 44.690 ;
        RECT 236.750 43.670 236.890 54.000 ;
        RECT 236.690 43.350 236.950 43.670 ;
        RECT 237.210 42.650 237.350 54.000 ;
        RECT 237.670 44.010 237.810 54.000 ;
        RECT 238.130 53.190 238.270 54.000 ;
        RECT 238.070 52.870 238.330 53.190 ;
        RECT 238.990 52.870 239.250 53.190 ;
        RECT 238.070 52.365 238.330 52.510 ;
        RECT 238.060 51.995 238.340 52.365 ;
        RECT 238.060 51.315 238.340 51.685 ;
        RECT 238.130 46.730 238.270 51.315 ;
        RECT 239.050 50.470 239.190 52.870 ;
        RECT 238.990 50.150 239.250 50.470 ;
        RECT 238.990 47.660 239.250 47.750 ;
        RECT 239.510 47.660 239.650 54.000 ;
        RECT 238.990 47.520 239.650 47.660 ;
        RECT 238.990 47.430 239.250 47.520 ;
        RECT 238.070 46.410 238.330 46.730 ;
        RECT 238.990 46.410 239.250 46.730 ;
        RECT 239.050 44.690 239.190 46.410 ;
        RECT 238.990 44.370 239.250 44.690 ;
        RECT 237.610 43.690 237.870 44.010 ;
        RECT 237.150 42.330 237.410 42.650 ;
        RECT 239.970 41.290 240.110 54.000 ;
        RECT 240.430 48.090 240.570 54.000 ;
        RECT 240.370 47.770 240.630 48.090 ;
        RECT 240.360 47.235 240.640 47.605 ;
        RECT 240.430 47.070 240.570 47.235 ;
        RECT 240.370 46.750 240.630 47.070 ;
        RECT 240.890 45.030 241.030 54.000 ;
        RECT 241.750 51.510 242.010 51.830 ;
        RECT 241.280 49.955 241.560 50.325 ;
        RECT 241.290 49.810 241.550 49.955 ;
        RECT 241.810 49.110 241.950 51.510 ;
        RECT 242.270 50.130 242.410 54.000 ;
        RECT 242.210 49.810 242.470 50.130 ;
        RECT 241.750 48.790 242.010 49.110 ;
        RECT 242.730 47.750 242.870 54.000 ;
        RECT 243.120 52.675 243.400 53.045 ;
        RECT 243.130 52.530 243.390 52.675 ;
        RECT 245.030 51.830 245.170 54.000 ;
        RECT 244.970 51.510 245.230 51.830 ;
        RECT 243.120 49.275 243.400 49.645 ;
        RECT 243.190 49.110 243.330 49.275 ;
        RECT 243.130 48.790 243.390 49.110 ;
        RECT 244.500 48.170 244.780 48.285 ;
        RECT 243.650 48.030 244.780 48.170 ;
        RECT 242.670 47.430 242.930 47.750 ;
        RECT 243.650 47.605 243.790 48.030 ;
        RECT 244.500 47.915 244.780 48.030 ;
        RECT 243.580 47.235 243.860 47.605 ;
        RECT 245.490 47.410 245.630 54.000 ;
        RECT 243.650 47.070 243.790 47.235 ;
        RECT 245.430 47.090 245.690 47.410 ;
        RECT 243.590 46.750 243.850 47.070 ;
        RECT 244.050 46.750 244.310 47.070 ;
        RECT 244.110 46.130 244.250 46.750 ;
        RECT 241.810 45.990 244.250 46.130 ;
        RECT 240.830 44.710 241.090 45.030 ;
        RECT 239.910 40.970 240.170 41.290 ;
        RECT 238.070 39.270 238.330 39.590 ;
        RECT 238.130 34.520 238.270 39.270 ;
        RECT 241.810 34.520 241.950 45.990 ;
        RECT 243.590 44.370 243.850 44.690 ;
        RECT 243.650 42.650 243.790 44.370 ;
        RECT 244.970 43.690 245.230 44.010 ;
        RECT 243.590 42.330 243.850 42.650 ;
        RECT 245.030 40.610 245.170 43.690 ;
        RECT 244.970 40.290 245.230 40.610 ;
        RECT 245.950 39.590 246.090 54.000 ;
        RECT 246.350 49.130 246.610 49.450 ;
        RECT 246.410 46.390 246.550 49.130 ;
        RECT 247.330 48.090 247.470 54.000 ;
        RECT 248.250 53.530 248.390 54.000 ;
        RECT 248.190 53.210 248.450 53.530 ;
        RECT 246.810 47.770 247.070 48.090 ;
        RECT 247.270 47.770 247.530 48.090 ;
        RECT 246.870 46.390 247.010 47.770 ;
        RECT 246.350 46.070 246.610 46.390 ;
        RECT 246.810 46.070 247.070 46.390 ;
        RECT 247.330 45.030 247.470 47.770 ;
        RECT 247.270 44.710 247.530 45.030 ;
        RECT 248.710 44.940 248.850 54.000 ;
        RECT 249.110 53.210 249.370 53.530 ;
        RECT 249.170 52.510 249.310 53.210 ;
        RECT 249.110 52.190 249.370 52.510 ;
        RECT 249.570 52.190 249.830 52.510 ;
        RECT 249.630 50.810 249.770 52.190 ;
        RECT 250.090 51.570 250.230 54.000 ;
        RECT 250.090 51.430 250.690 51.570 ;
        RECT 249.570 50.490 249.830 50.810 ;
        RECT 250.020 50.635 250.300 51.005 ;
        RECT 250.030 50.490 250.290 50.635 ;
        RECT 248.710 44.800 249.310 44.940 ;
        RECT 245.890 39.270 246.150 39.590 ;
        RECT 245.430 38.930 245.690 39.250 ;
        RECT 245.490 34.520 245.630 38.930 ;
        RECT 249.170 34.520 249.310 44.800 ;
        RECT 250.550 39.250 250.690 51.430 ;
        RECT 251.010 51.005 251.150 54.000 ;
        RECT 251.470 51.830 251.610 54.000 ;
        RECT 251.930 53.045 252.070 54.000 ;
        RECT 251.860 52.675 252.140 53.045 ;
        RECT 251.410 51.510 251.670 51.830 ;
        RECT 251.870 51.510 252.130 51.830 ;
        RECT 250.940 50.635 251.220 51.005 ;
        RECT 251.930 47.070 252.070 51.510 ;
        RECT 252.390 48.965 252.530 54.000 ;
        RECT 252.850 53.190 252.990 54.000 ;
        RECT 252.790 52.870 253.050 53.190 ;
        RECT 253.770 51.830 253.910 54.000 ;
        RECT 254.230 53.045 254.370 54.000 ;
        RECT 254.160 52.675 254.440 53.045 ;
        RECT 253.710 51.510 253.970 51.830 ;
        RECT 252.790 49.810 253.050 50.130 ;
        RECT 252.320 48.595 252.600 48.965 ;
        RECT 252.320 47.235 252.600 47.605 ;
        RECT 252.330 47.090 252.590 47.235 ;
        RECT 251.870 46.750 252.130 47.070 ;
        RECT 252.850 46.980 252.990 49.810 ;
        RECT 254.230 48.850 254.370 52.675 ;
        RECT 253.770 48.710 254.370 48.850 ;
        RECT 253.770 47.750 253.910 48.710 ;
        RECT 253.710 47.430 253.970 47.750 ;
        RECT 253.250 46.980 253.510 47.070 ;
        RECT 252.850 46.840 253.510 46.980 ;
        RECT 253.250 46.750 253.510 46.840 ;
        RECT 254.690 46.730 254.830 54.000 ;
        RECT 254.630 46.410 254.890 46.730 ;
        RECT 252.780 45.875 253.060 46.245 ;
        RECT 250.490 38.930 250.750 39.250 ;
        RECT 252.850 34.520 252.990 45.875 ;
        RECT 255.150 39.930 255.290 54.000 ;
        RECT 256.070 47.070 256.210 54.000 ;
        RECT 256.470 52.530 256.730 52.850 ;
        RECT 256.530 52.365 256.670 52.530 ;
        RECT 256.460 51.995 256.740 52.365 ;
        RECT 256.470 51.510 256.730 51.830 ;
        RECT 256.990 51.570 257.130 54.000 ;
        RECT 256.010 46.750 256.270 47.070 ;
        RECT 256.530 46.730 256.670 51.510 ;
        RECT 256.990 51.430 258.050 51.570 ;
        RECT 256.930 50.490 257.190 50.810 ;
        RECT 256.990 50.130 257.130 50.490 ;
        RECT 257.910 50.470 258.050 51.430 ;
        RECT 257.850 50.150 258.110 50.470 ;
        RECT 256.930 49.810 257.190 50.130 ;
        RECT 256.470 46.410 256.730 46.730 ;
        RECT 257.850 44.370 258.110 44.690 ;
        RECT 257.910 42.165 258.050 44.370 ;
        RECT 258.370 44.010 258.510 54.000 ;
        RECT 258.830 52.510 258.970 54.000 ;
        RECT 258.770 52.190 259.030 52.510 ;
        RECT 258.770 50.150 259.030 50.470 ;
        RECT 258.830 44.690 258.970 50.150 ;
        RECT 259.290 45.370 259.430 54.000 ;
        RECT 259.750 50.810 259.890 54.000 ;
        RECT 260.210 53.530 260.350 54.000 ;
        RECT 260.150 53.210 260.410 53.530 ;
        RECT 259.690 50.490 259.950 50.810 ;
        RECT 260.670 50.130 260.810 54.000 ;
        RECT 260.610 49.810 260.870 50.130 ;
        RECT 259.690 49.470 259.950 49.790 ;
        RECT 259.750 49.110 259.890 49.470 ;
        RECT 259.690 48.790 259.950 49.110 ;
        RECT 261.130 47.070 261.270 54.000 ;
        RECT 261.520 53.355 261.800 53.725 ;
        RECT 262.050 53.530 262.190 54.000 ;
        RECT 261.590 52.760 261.730 53.355 ;
        RECT 261.990 53.210 262.250 53.530 ;
        RECT 261.990 52.760 262.250 52.850 ;
        RECT 261.590 52.620 262.250 52.760 ;
        RECT 261.990 52.530 262.250 52.620 ;
        RECT 262.510 48.285 262.650 54.000 ;
        RECT 262.970 53.725 263.110 54.000 ;
        RECT 262.900 53.355 263.180 53.725 ;
        RECT 262.970 50.325 263.110 53.355 ;
        RECT 262.900 49.955 263.180 50.325 ;
        RECT 262.440 47.915 262.720 48.285 ;
        RECT 261.070 46.750 261.330 47.070 ;
        RECT 262.510 46.390 262.650 47.915 ;
        RECT 262.450 46.070 262.710 46.390 ;
        RECT 259.230 45.050 259.490 45.370 ;
        RECT 258.770 44.370 259.030 44.690 ;
        RECT 258.310 43.690 258.570 44.010 ;
        RECT 257.840 41.795 258.120 42.165 ;
        RECT 255.090 39.610 255.350 39.930 ;
        RECT 256.470 39.270 256.730 39.590 ;
        RECT 256.530 34.520 256.670 39.270 ;
        RECT 263.890 34.520 264.030 54.000 ;
        RECT 264.350 47.750 264.490 54.000 ;
        RECT 265.730 50.130 265.870 54.000 ;
        RECT 266.190 53.045 266.330 54.000 ;
        RECT 266.120 52.675 266.400 53.045 ;
        RECT 265.670 49.810 265.930 50.130 ;
        RECT 264.290 47.430 264.550 47.750 ;
        RECT 266.650 47.605 266.790 54.000 ;
        RECT 266.580 47.235 266.860 47.605 ;
        RECT 264.750 43.350 265.010 43.670 ;
        RECT 264.810 41.970 264.950 43.350 ;
        RECT 264.750 41.650 265.010 41.970 ;
        RECT 267.570 34.520 267.710 54.000 ;
        RECT 268.030 47.605 268.170 54.000 ;
        RECT 268.490 53.190 268.630 54.000 ;
        RECT 268.430 52.870 268.690 53.190 ;
        RECT 270.260 52.675 270.540 53.045 ;
        RECT 270.330 52.510 270.470 52.675 ;
        RECT 270.270 52.190 270.530 52.510 ;
        RECT 270.790 50.325 270.930 54.000 ;
        RECT 270.720 49.955 271.000 50.325 ;
        RECT 270.270 49.470 270.530 49.790 ;
        RECT 270.330 49.110 270.470 49.470 ;
        RECT 270.270 48.790 270.530 49.110 ;
        RECT 268.420 47.915 268.700 48.285 ;
        RECT 268.430 47.770 268.690 47.915 ;
        RECT 267.960 47.235 268.240 47.605 ;
        RECT 268.030 44.350 268.170 47.235 ;
        RECT 270.730 46.750 270.990 47.070 ;
        RECT 270.790 44.690 270.930 46.750 ;
        RECT 270.730 44.370 270.990 44.690 ;
        RECT 267.970 44.030 268.230 44.350 ;
        RECT 270.790 39.930 270.930 44.370 ;
        RECT 270.730 39.610 270.990 39.930 ;
        RECT 271.250 34.520 271.390 54.000 ;
        RECT 272.170 50.130 272.310 54.000 ;
        RECT 273.030 52.760 273.290 52.850 ;
        RECT 274.010 52.760 274.150 54.000 ;
        RECT 273.030 52.620 274.150 52.760 ;
        RECT 273.030 52.530 273.290 52.620 ;
        RECT 272.570 52.190 272.830 52.510 ;
        RECT 272.630 50.810 272.770 52.190 ;
        RECT 272.570 50.490 272.830 50.810 ;
        RECT 272.110 49.810 272.370 50.130 ;
        RECT 274.010 41.970 274.150 52.620 ;
        RECT 274.470 52.510 274.610 54.000 ;
        RECT 276.240 53.355 276.520 53.725 ;
        RECT 275.320 52.675 275.600 53.045 ;
        RECT 275.390 52.510 275.530 52.675 ;
        RECT 274.410 52.190 274.670 52.510 ;
        RECT 275.330 52.190 275.590 52.510 ;
        RECT 274.870 51.510 275.130 51.830 ;
        RECT 274.410 48.790 274.670 49.110 ;
        RECT 274.470 47.750 274.610 48.790 ;
        RECT 274.410 47.430 274.670 47.750 ;
        RECT 273.950 41.650 274.210 41.970 ;
        RECT 274.930 34.520 275.070 51.510 ;
        RECT 275.790 50.150 276.050 50.470 ;
        RECT 275.850 48.285 275.990 50.150 ;
        RECT 276.310 49.790 276.450 53.355 ;
        RECT 276.250 49.470 276.510 49.790 ;
        RECT 276.250 48.790 276.510 49.110 ;
        RECT 275.780 47.915 276.060 48.285 ;
        RECT 276.310 48.090 276.450 48.790 ;
        RECT 276.250 47.770 276.510 48.090 ;
        RECT 275.790 46.750 276.050 47.070 ;
        RECT 275.850 44.350 275.990 46.750 ;
        RECT 275.790 44.030 276.050 44.350 ;
        RECT 276.770 39.590 276.910 54.000 ;
        RECT 277.230 52.850 277.370 54.000 ;
        RECT 277.690 52.850 277.830 54.000 ;
        RECT 277.170 52.530 277.430 52.850 ;
        RECT 277.630 52.530 277.890 52.850 ;
        RECT 276.710 39.270 276.970 39.590 ;
        RECT 278.610 34.520 278.750 54.000 ;
        RECT 279.990 53.530 280.130 54.000 ;
        RECT 279.470 53.210 279.730 53.530 ;
        RECT 279.930 53.210 280.190 53.530 ;
        RECT 279.530 44.690 279.670 53.210 ;
        RECT 280.450 51.830 280.590 54.000 ;
        RECT 281.770 51.850 282.030 52.170 ;
        RECT 280.390 51.510 280.650 51.830 ;
        RECT 280.390 49.810 280.650 50.130 ;
        RECT 279.470 44.370 279.730 44.690 ;
        RECT 280.450 40.950 280.590 49.810 ;
        RECT 280.390 40.630 280.650 40.950 ;
        RECT 281.830 39.590 281.970 51.850 ;
        RECT 282.290 50.130 282.430 54.000 ;
        RECT 282.750 53.045 282.890 54.000 ;
        RECT 282.680 52.675 282.960 53.045 ;
        RECT 284.070 52.760 284.330 52.850 ;
        RECT 282.750 52.510 282.890 52.675 ;
        RECT 284.070 52.620 285.190 52.760 ;
        RECT 284.070 52.530 284.330 52.620 ;
        RECT 282.690 52.190 282.950 52.510 ;
        RECT 283.610 52.190 283.870 52.510 ;
        RECT 282.690 50.490 282.950 50.810 ;
        RECT 282.230 49.810 282.490 50.130 ;
        RECT 282.230 42.330 282.490 42.650 ;
        RECT 281.770 39.270 282.030 39.590 ;
        RECT 282.290 34.520 282.430 42.330 ;
        RECT 282.750 38.570 282.890 50.490 ;
        RECT 283.150 49.810 283.410 50.130 ;
        RECT 283.210 49.110 283.350 49.810 ;
        RECT 283.150 48.790 283.410 49.110 ;
        RECT 283.670 48.090 283.810 52.190 ;
        RECT 285.050 50.130 285.190 52.620 ;
        RECT 285.450 52.190 285.710 52.510 ;
        RECT 285.510 51.685 285.650 52.190 ;
        RECT 286.430 52.170 286.570 54.000 ;
        RECT 286.370 51.850 286.630 52.170 ;
        RECT 285.440 51.315 285.720 51.685 ;
        RECT 286.890 51.570 287.030 54.000 ;
        RECT 287.810 52.760 287.950 54.000 ;
        RECT 288.210 52.760 288.470 52.850 ;
        RECT 287.810 52.620 288.470 52.760 ;
        RECT 288.210 52.530 288.470 52.620 ;
        RECT 288.730 52.250 288.870 54.000 ;
        RECT 290.570 53.530 290.710 54.000 ;
        RECT 290.510 53.210 290.770 53.530 ;
        RECT 285.970 51.430 287.030 51.570 ;
        RECT 287.350 52.110 288.870 52.250 ;
        RECT 284.990 49.810 285.250 50.130 ;
        RECT 283.610 47.770 283.870 48.090 ;
        RECT 284.070 46.925 284.330 47.070 ;
        RECT 284.060 46.555 284.340 46.925 ;
        RECT 284.530 46.070 284.790 46.390 ;
        RECT 285.450 46.070 285.710 46.390 ;
        RECT 282.690 38.250 282.950 38.570 ;
        RECT 284.590 34.520 284.730 46.070 ;
        RECT 285.510 40.270 285.650 46.070 ;
        RECT 285.450 39.950 285.710 40.270 ;
        RECT 285.970 34.520 286.110 51.430 ;
        RECT 286.360 50.635 286.640 51.005 ;
        RECT 286.430 39.250 286.570 50.635 ;
        RECT 286.830 46.410 287.090 46.730 ;
        RECT 286.370 38.930 286.630 39.250 ;
        RECT 286.890 34.520 287.030 46.410 ;
        RECT 287.350 42.310 287.490 52.110 ;
        RECT 287.750 51.510 288.010 51.830 ;
        RECT 287.810 50.130 287.950 51.510 ;
        RECT 288.450 50.920 289.930 51.400 ;
        RECT 290.500 50.890 290.780 51.005 ;
        RECT 290.110 50.750 290.780 50.890 ;
        RECT 291.950 50.810 292.090 54.000 ;
        RECT 292.340 52.675 292.620 53.045 ;
        RECT 292.410 50.810 292.550 52.675 ;
        RECT 287.750 49.810 288.010 50.130 ;
        RECT 287.750 49.130 288.010 49.450 ;
        RECT 287.290 41.990 287.550 42.310 ;
        RECT 287.810 38.650 287.950 49.130 ;
        RECT 289.120 47.915 289.400 48.285 ;
        RECT 289.190 47.070 289.330 47.915 ;
        RECT 290.110 47.605 290.250 50.750 ;
        RECT 290.500 50.635 290.780 50.750 ;
        RECT 291.890 50.490 292.150 50.810 ;
        RECT 292.350 50.490 292.610 50.810 ;
        RECT 292.810 49.810 293.070 50.130 ;
        RECT 290.510 48.790 290.770 49.110 ;
        RECT 292.350 48.790 292.610 49.110 ;
        RECT 290.040 47.235 290.320 47.605 ;
        RECT 289.130 46.750 289.390 47.070 ;
        RECT 288.450 45.480 289.930 45.960 ;
        RECT 288.660 44.515 288.940 44.885 ;
        RECT 288.670 44.370 288.930 44.515 ;
        RECT 289.590 41.990 289.850 42.310 ;
        RECT 287.810 38.510 288.410 38.650 ;
        RECT 288.270 34.520 288.410 38.510 ;
        RECT 289.650 34.520 289.790 41.990 ;
        RECT 290.570 34.520 290.710 48.790 ;
        RECT 290.960 47.235 291.240 47.605 ;
        RECT 292.410 47.410 292.550 48.790 ;
        RECT 291.030 47.070 291.170 47.235 ;
        RECT 292.350 47.090 292.610 47.410 ;
        RECT 290.970 46.750 291.230 47.070 ;
        RECT 292.870 46.245 293.010 49.810 ;
        RECT 293.330 47.410 293.470 54.000 ;
        RECT 294.250 50.130 294.390 54.000 ;
        RECT 295.170 50.470 295.310 54.000 ;
        RECT 295.630 52.510 295.770 54.000 ;
        RECT 295.570 52.190 295.830 52.510 ;
        RECT 295.110 50.150 295.370 50.470 ;
        RECT 294.190 49.810 294.450 50.130 ;
        RECT 295.110 49.130 295.370 49.450 ;
        RECT 293.270 47.090 293.530 47.410 ;
        RECT 292.800 45.875 293.080 46.245 ;
        RECT 293.730 45.050 293.990 45.370 ;
        RECT 292.350 44.710 292.610 45.030 ;
        RECT 292.810 44.885 293.070 45.030 ;
        RECT 292.410 39.250 292.550 44.710 ;
        RECT 292.800 44.515 293.080 44.885 ;
        RECT 293.790 44.770 293.930 45.050 ;
        RECT 295.170 44.885 295.310 49.130 ;
        RECT 296.090 46.245 296.230 54.000 ;
        RECT 296.550 49.790 296.690 54.000 ;
        RECT 296.490 49.470 296.750 49.790 ;
        RECT 296.020 45.875 296.300 46.245 ;
        RECT 293.790 44.630 294.390 44.770 ;
        RECT 292.810 44.030 293.070 44.350 ;
        RECT 292.870 39.930 293.010 44.030 ;
        RECT 292.810 39.610 293.070 39.930 ;
        RECT 293.270 39.610 293.530 39.930 ;
        RECT 291.890 38.930 292.150 39.250 ;
        RECT 292.350 38.930 292.610 39.250 ;
        RECT 291.950 34.520 292.090 38.930 ;
        RECT 293.330 34.520 293.470 39.610 ;
        RECT 294.250 34.520 294.390 44.630 ;
        RECT 295.100 44.515 295.380 44.885 ;
        RECT 297.010 34.520 297.150 54.000 ;
        RECT 298.390 53.725 298.530 54.000 ;
        RECT 298.320 53.355 298.600 53.725 ;
        RECT 298.390 52.930 298.530 53.355 ;
        RECT 298.390 52.790 298.990 52.930 ;
        RECT 298.330 52.365 298.590 52.510 ;
        RECT 298.320 52.250 298.600 52.365 ;
        RECT 297.930 52.110 298.600 52.250 ;
        RECT 297.930 45.370 298.070 52.110 ;
        RECT 298.320 51.995 298.600 52.110 ;
        RECT 298.330 46.750 298.590 47.070 ;
        RECT 297.870 45.050 298.130 45.370 ;
        RECT 298.390 44.350 298.530 46.750 ;
        RECT 298.850 44.690 298.990 52.790 ;
        RECT 299.250 49.810 299.510 50.130 ;
        RECT 299.310 45.370 299.450 49.810 ;
        RECT 299.770 47.070 299.910 54.000 ;
        RECT 299.710 46.750 299.970 47.070 ;
        RECT 299.250 45.050 299.510 45.370 ;
        RECT 298.790 44.370 299.050 44.690 ;
        RECT 298.330 44.030 298.590 44.350 ;
        RECT 298.390 43.670 298.530 44.030 ;
        RECT 298.330 43.350 298.590 43.670 ;
        RECT 299.250 39.270 299.510 39.590 ;
        RECT 297.870 38.930 298.130 39.250 ;
        RECT 297.930 34.520 298.070 38.930 ;
        RECT 299.310 34.520 299.450 39.270 ;
        RECT 300.690 34.520 300.830 54.000 ;
        RECT 301.150 42.310 301.290 54.000 ;
        RECT 302.990 53.190 303.130 54.000 ;
        RECT 302.930 52.870 303.190 53.190 ;
        RECT 303.450 53.045 303.590 54.000 ;
        RECT 303.380 52.675 303.660 53.045 ;
        RECT 303.450 50.130 303.590 52.675 ;
        RECT 303.390 49.810 303.650 50.130 ;
        RECT 302.930 46.070 303.190 46.390 ;
        RECT 302.010 44.030 302.270 44.350 ;
        RECT 301.090 41.990 301.350 42.310 ;
        RECT 302.070 41.970 302.210 44.030 ;
        RECT 302.010 41.650 302.270 41.970 ;
        RECT 302.990 34.520 303.130 46.070 ;
        RECT 303.910 39.930 304.050 54.000 ;
        RECT 304.310 49.470 304.570 49.790 ;
        RECT 303.850 39.610 304.110 39.930 ;
        RECT 304.370 34.520 304.510 49.470 ;
        RECT 304.830 46.640 304.970 54.000 ;
        RECT 305.290 46.980 305.430 54.000 ;
        RECT 306.600 48.595 306.880 48.965 ;
        RECT 306.150 46.980 306.410 47.070 ;
        RECT 305.290 46.840 306.410 46.980 ;
        RECT 306.150 46.750 306.410 46.840 ;
        RECT 304.830 46.500 305.890 46.640 ;
        RECT 305.750 45.370 305.890 46.500 ;
        RECT 306.210 45.565 306.350 46.750 ;
        RECT 305.230 45.050 305.490 45.370 ;
        RECT 305.690 45.050 305.950 45.370 ;
        RECT 306.140 45.195 306.420 45.565 ;
        RECT 305.290 34.520 305.430 45.050 ;
        RECT 306.210 44.690 306.350 45.195 ;
        RECT 306.150 44.370 306.410 44.690 ;
        RECT 306.670 34.520 306.810 48.595 ;
        RECT 308.050 34.520 308.190 54.000 ;
        RECT 309.890 52.510 310.030 54.000 ;
        RECT 308.910 52.420 309.170 52.510 ;
        RECT 309.830 52.420 310.090 52.510 ;
        RECT 308.910 52.280 310.090 52.420 ;
        RECT 308.910 52.190 309.170 52.280 ;
        RECT 309.830 52.190 310.090 52.280 ;
        RECT 308.910 51.510 309.170 51.830 ;
        RECT 308.450 43.350 308.710 43.670 ;
        RECT 308.510 40.610 308.650 43.350 ;
        RECT 308.450 40.290 308.710 40.610 ;
        RECT 308.970 34.520 309.110 51.510 ;
        RECT 310.280 51.315 310.560 51.685 ;
        RECT 309.830 47.430 310.090 47.750 ;
        RECT 309.890 43.670 310.030 47.430 ;
        RECT 309.830 43.350 310.090 43.670 ;
        RECT 310.350 34.520 310.490 51.315 ;
        RECT 310.810 49.790 310.950 54.000 ;
        RECT 311.670 52.190 311.930 52.510 ;
        RECT 311.730 51.005 311.870 52.190 ;
        RECT 312.190 51.830 312.330 54.000 ;
        RECT 312.130 51.510 312.390 51.830 ;
        RECT 311.660 50.635 311.940 51.005 ;
        RECT 310.750 49.470 311.010 49.790 ;
        RECT 311.670 47.770 311.930 48.090 ;
        RECT 311.210 46.070 311.470 46.390 ;
        RECT 311.270 40.610 311.410 46.070 ;
        RECT 311.210 40.290 311.470 40.610 ;
        RECT 311.730 34.520 311.870 47.770 ;
        RECT 312.650 46.390 312.790 54.000 ;
        RECT 312.590 46.070 312.850 46.390 ;
        RECT 312.590 44.710 312.850 45.030 ;
        RECT 312.650 34.520 312.790 44.710 ;
        RECT 313.570 44.010 313.710 54.000 ;
        RECT 313.510 43.690 313.770 44.010 ;
        RECT 314.030 34.520 314.170 54.000 ;
        RECT 317.180 53.355 317.460 53.725 ;
        RECT 315.350 52.530 315.610 52.850 ;
        RECT 314.890 48.790 315.150 49.110 ;
        RECT 314.950 47.070 315.090 48.790 ;
        RECT 314.430 46.750 314.690 47.070 ;
        RECT 314.890 46.750 315.150 47.070 ;
        RECT 314.490 45.565 314.630 46.750 ;
        RECT 314.420 45.195 314.700 45.565 ;
        RECT 315.410 34.520 315.550 52.530 ;
        RECT 317.250 52.510 317.390 53.355 ;
        RECT 317.190 52.190 317.450 52.510 ;
        RECT 317.710 48.090 317.850 54.000 ;
        RECT 318.170 52.510 318.310 54.000 ;
        RECT 320.930 52.850 321.070 54.000 ;
        RECT 320.870 52.530 321.130 52.850 ;
        RECT 318.110 52.190 318.370 52.510 ;
        RECT 318.110 51.510 318.370 51.830 ;
        RECT 318.570 51.510 318.830 51.830 ;
        RECT 318.170 50.810 318.310 51.510 ;
        RECT 318.110 50.490 318.370 50.810 ;
        RECT 317.650 47.770 317.910 48.090 ;
        RECT 316.270 47.090 316.530 47.410 ;
        RECT 315.810 44.030 316.070 44.350 ;
        RECT 315.870 40.950 316.010 44.030 ;
        RECT 315.810 40.630 316.070 40.950 ;
        RECT 316.330 34.520 316.470 47.090 ;
        RECT 318.630 46.925 318.770 51.510 ;
        RECT 319.030 50.150 319.290 50.470 ;
        RECT 318.560 46.555 318.840 46.925 ;
        RECT 317.650 43.350 317.910 43.670 ;
        RECT 317.710 34.520 317.850 43.350 ;
        RECT 319.090 34.520 319.230 50.150 ;
        RECT 321.320 49.955 321.600 50.325 ;
        RECT 319.950 43.690 320.210 44.010 ;
        RECT 320.010 34.520 320.150 43.690 ;
        RECT 321.390 34.520 321.530 49.955 ;
        RECT 322.770 34.520 322.910 54.000 ;
        RECT 323.690 52.510 323.830 54.000 ;
        RECT 323.630 52.190 323.890 52.510 ;
        RECT 324.150 46.390 324.290 54.000 ;
        RECT 325.530 50.470 325.670 54.000 ;
        RECT 325.990 50.470 326.130 54.000 ;
        RECT 326.380 52.675 326.660 53.045 ;
        RECT 325.470 50.150 325.730 50.470 ;
        RECT 325.930 50.150 326.190 50.470 ;
        RECT 325.930 47.770 326.190 48.090 ;
        RECT 324.090 46.070 324.350 46.390 ;
        RECT 325.470 46.070 325.730 46.390 ;
        RECT 325.530 44.885 325.670 46.070 ;
        RECT 325.460 44.515 325.740 44.885 ;
        RECT 323.630 40.290 323.890 40.610 ;
        RECT 323.690 34.520 323.830 40.290 ;
        RECT 325.010 38.250 325.270 38.570 ;
        RECT 325.070 34.520 325.210 38.250 ;
        RECT 325.990 37.290 326.130 47.770 ;
        RECT 326.450 47.070 326.590 52.675 ;
        RECT 326.850 52.530 327.110 52.850 ;
        RECT 326.910 50.130 327.050 52.530 ;
        RECT 327.370 51.830 327.510 54.000 ;
        RECT 327.830 53.610 327.970 54.000 ;
        RECT 327.830 53.470 328.430 53.610 ;
        RECT 328.750 53.530 328.890 54.000 ;
        RECT 327.770 53.045 328.030 53.190 ;
        RECT 327.760 52.675 328.040 53.045 ;
        RECT 328.290 52.930 328.430 53.470 ;
        RECT 328.690 53.210 328.950 53.530 ;
        RECT 328.290 52.790 328.890 52.930 ;
        RECT 329.670 52.850 329.810 54.000 ;
        RECT 327.770 52.190 328.030 52.510 ;
        RECT 327.310 51.510 327.570 51.830 ;
        RECT 326.850 49.810 327.110 50.130 ;
        RECT 327.310 48.790 327.570 49.110 ;
        RECT 327.830 48.965 327.970 52.190 ;
        RECT 328.230 51.510 328.490 51.830 ;
        RECT 328.290 50.470 328.430 51.510 ;
        RECT 328.230 50.150 328.490 50.470 ;
        RECT 326.390 46.750 326.650 47.070 ;
        RECT 326.450 45.030 326.590 46.750 ;
        RECT 326.390 44.710 326.650 45.030 ;
        RECT 325.990 37.150 326.590 37.290 ;
        RECT 326.450 34.520 326.590 37.150 ;
        RECT 327.370 34.520 327.510 48.790 ;
        RECT 327.760 48.595 328.040 48.965 ;
        RECT 328.750 34.520 328.890 52.790 ;
        RECT 329.610 52.530 329.870 52.850 ;
        RECT 330.130 52.510 330.270 54.000 ;
        RECT 329.150 52.190 329.410 52.510 ;
        RECT 330.070 52.190 330.330 52.510 ;
        RECT 329.210 40.610 329.350 52.190 ;
        RECT 330.130 51.830 330.270 52.190 ;
        RECT 330.070 51.740 330.330 51.830 ;
        RECT 329.670 51.600 330.330 51.740 ;
        RECT 329.670 42.310 329.810 51.600 ;
        RECT 330.070 51.510 330.330 51.600 ;
        RECT 331.050 49.700 331.190 54.000 ;
        RECT 331.440 52.675 331.720 53.045 ;
        RECT 331.510 50.130 331.650 52.675 ;
        RECT 331.970 52.365 332.110 54.000 ;
        RECT 332.430 52.510 332.570 54.000 ;
        RECT 331.900 51.995 332.180 52.365 ;
        RECT 332.370 52.190 332.630 52.510 ;
        RECT 332.830 52.190 333.090 52.510 ;
        RECT 332.890 51.830 333.030 52.190 ;
        RECT 332.830 51.510 333.090 51.830 ;
        RECT 331.910 50.490 332.170 50.810 ;
        RECT 331.450 49.810 331.710 50.130 ;
        RECT 330.130 49.560 331.190 49.700 ;
        RECT 329.610 41.990 329.870 42.310 ;
        RECT 329.150 40.290 329.410 40.610 ;
        RECT 330.130 34.520 330.270 49.560 ;
        RECT 330.990 46.410 331.250 46.730 ;
        RECT 331.050 34.520 331.190 46.410 ;
        RECT 331.970 44.885 332.110 50.490 ;
        RECT 333.810 48.090 333.950 54.000 ;
        RECT 334.210 51.850 334.470 52.170 ;
        RECT 334.270 48.090 334.410 51.850 ;
        RECT 333.750 47.770 334.010 48.090 ;
        RECT 334.210 47.770 334.470 48.090 ;
        RECT 332.370 47.430 332.630 47.750 ;
        RECT 334.730 47.490 334.870 54.000 ;
        RECT 335.190 52.850 335.330 54.000 ;
        RECT 335.130 52.530 335.390 52.850 ;
        RECT 331.900 44.515 332.180 44.885 ;
        RECT 332.430 34.520 332.570 47.430 ;
        RECT 333.810 47.350 334.870 47.490 ;
        RECT 332.830 46.750 333.090 47.070 ;
        RECT 333.290 46.750 333.550 47.070 ;
        RECT 332.890 39.930 333.030 46.750 ;
        RECT 333.350 43.670 333.490 46.750 ;
        RECT 333.290 43.350 333.550 43.670 ;
        RECT 332.830 39.610 333.090 39.930 ;
        RECT 333.810 34.520 333.950 47.350 ;
        RECT 334.210 46.410 334.470 46.730 ;
        RECT 334.270 46.245 334.410 46.410 ;
        RECT 335.650 46.300 335.790 54.000 ;
        RECT 336.110 51.830 336.250 54.000 ;
        RECT 336.050 51.510 336.310 51.830 ;
        RECT 336.050 49.810 336.310 50.130 ;
        RECT 334.200 45.875 334.480 46.245 ;
        RECT 334.730 46.160 335.790 46.300 ;
        RECT 334.730 34.520 334.870 46.160 ;
        RECT 336.110 34.520 336.250 49.810 ;
        RECT 336.570 44.690 336.710 54.000 ;
        RECT 336.510 44.370 336.770 44.690 ;
        RECT 337.030 44.090 337.170 54.000 ;
        RECT 337.490 50.130 337.630 54.000 ;
        RECT 337.950 50.325 338.090 54.000 ;
        RECT 337.430 49.810 337.690 50.130 ;
        RECT 337.880 49.955 338.160 50.325 ;
        RECT 337.950 48.285 338.090 49.955 ;
        RECT 337.880 47.915 338.160 48.285 ;
        RECT 338.410 47.410 338.550 54.000 ;
        RECT 339.720 48.595 340.000 48.965 ;
        RECT 338.350 47.090 338.610 47.410 ;
        RECT 339.790 46.390 339.930 48.595 ;
        RECT 340.190 46.980 340.450 47.070 ;
        RECT 340.710 46.980 340.850 54.000 ;
        RECT 340.190 46.840 340.850 46.980 ;
        RECT 340.190 46.750 340.450 46.840 ;
        RECT 338.810 46.070 339.070 46.390 ;
        RECT 339.730 46.070 339.990 46.390 ;
        RECT 338.870 45.450 339.010 46.070 ;
        RECT 340.640 45.875 340.920 46.245 ;
        RECT 338.870 45.310 339.930 45.450 ;
        RECT 336.570 43.950 337.170 44.090 ;
        RECT 336.570 40.950 336.710 43.950 ;
        RECT 338.350 43.690 338.610 44.010 ;
        RECT 336.970 43.350 337.230 43.670 ;
        RECT 337.030 42.650 337.170 43.350 ;
        RECT 336.970 42.330 337.230 42.650 ;
        RECT 336.510 40.630 336.770 40.950 ;
        RECT 338.410 34.520 338.550 43.690 ;
        RECT 339.790 34.520 339.930 45.310 ;
        RECT 340.710 34.520 340.850 45.875 ;
        RECT 341.170 40.270 341.310 54.000 ;
        RECT 341.560 51.995 341.840 52.365 ;
        RECT 341.630 47.070 341.770 51.995 ;
        RECT 341.570 46.750 341.830 47.070 ;
        RECT 342.550 46.730 342.690 54.000 ;
        RECT 342.950 52.870 343.210 53.190 ;
        RECT 343.010 52.365 343.150 52.870 ;
        RECT 343.470 52.510 343.610 54.000 ;
        RECT 342.940 51.995 343.220 52.365 ;
        RECT 343.410 52.190 343.670 52.510 ;
        RECT 343.410 49.700 343.670 49.790 ;
        RECT 343.410 49.560 344.070 49.700 ;
        RECT 343.410 49.470 343.670 49.560 ;
        RECT 342.950 48.790 343.210 49.110 ;
        RECT 343.930 48.965 344.070 49.560 ;
        RECT 344.390 49.450 344.530 54.000 ;
        RECT 345.310 50.470 345.450 54.000 ;
        RECT 346.230 52.850 346.370 54.000 ;
        RECT 346.170 52.530 346.430 52.850 ;
        RECT 345.250 50.150 345.510 50.470 ;
        RECT 344.330 49.130 344.590 49.450 ;
        RECT 343.010 48.090 343.150 48.790 ;
        RECT 343.860 48.595 344.140 48.965 ;
        RECT 342.950 47.770 343.210 48.090 ;
        RECT 342.490 46.410 342.750 46.730 ;
        RECT 345.710 46.070 345.970 46.390 ;
        RECT 345.250 44.370 345.510 44.690 ;
        RECT 342.950 44.030 343.210 44.350 ;
        RECT 343.010 41.290 343.150 44.030 ;
        RECT 344.330 41.650 344.590 41.970 ;
        RECT 342.950 40.970 343.210 41.290 ;
        RECT 341.110 39.950 341.370 40.270 ;
        RECT 342.030 39.610 342.290 39.930 ;
        RECT 342.090 34.520 342.230 39.610 ;
        RECT 344.390 34.520 344.530 41.650 ;
        RECT 345.310 41.630 345.450 44.370 ;
        RECT 345.250 41.310 345.510 41.630 ;
        RECT 345.770 34.520 345.910 46.070 ;
        RECT 347.150 34.520 347.290 54.000 ;
        RECT 348.070 50.810 348.210 54.000 ;
        RECT 348.010 50.490 348.270 50.810 ;
        RECT 347.550 50.150 347.810 50.470 ;
        RECT 347.610 47.070 347.750 50.150 ;
        RECT 347.550 46.750 347.810 47.070 ;
        RECT 348.530 46.245 348.670 54.000 ;
        RECT 350.310 53.210 350.570 53.530 ;
        RECT 350.370 49.110 350.510 53.210 ;
        RECT 351.750 52.510 351.890 54.000 ;
        RECT 352.670 53.190 352.810 54.000 ;
        RECT 352.610 52.870 352.870 53.190 ;
        RECT 351.690 52.190 351.950 52.510 ;
        RECT 353.130 50.130 353.270 54.000 ;
        RECT 353.590 52.510 353.730 54.000 ;
        RECT 353.530 52.190 353.790 52.510 ;
        RECT 353.070 49.810 353.330 50.130 ;
        RECT 353.070 49.130 353.330 49.450 ;
        RECT 350.310 48.790 350.570 49.110 ;
        RECT 350.770 47.090 351.030 47.410 ;
        RECT 348.460 45.875 348.740 46.245 ;
        RECT 348.010 37.570 348.270 37.890 ;
        RECT 348.070 34.520 348.210 37.570 ;
        RECT 350.830 34.520 350.970 47.090 ;
        RECT 352.610 46.070 352.870 46.390 ;
        RECT 352.150 44.370 352.410 44.690 ;
        RECT 352.210 42.310 352.350 44.370 ;
        RECT 352.150 41.990 352.410 42.310 ;
        RECT 352.670 39.330 352.810 46.070 ;
        RECT 351.750 39.190 352.810 39.330 ;
        RECT 351.750 34.520 351.890 39.190 ;
        RECT 353.130 34.520 353.270 49.130 ;
        RECT 353.530 46.750 353.790 47.070 ;
        RECT 353.590 45.565 353.730 46.750 ;
        RECT 353.520 45.195 353.800 45.565 ;
        RECT 354.510 34.520 354.650 54.000 ;
        RECT 357.730 52.850 357.870 54.000 ;
        RECT 357.670 52.530 357.930 52.850 ;
        RECT 358.190 52.510 358.330 54.000 ;
        RECT 358.590 52.530 358.850 52.850 ;
        RECT 358.130 52.190 358.390 52.510 ;
        RECT 354.910 51.510 355.170 51.830 ;
        RECT 354.970 50.810 355.110 51.510 ;
        RECT 354.910 50.490 355.170 50.810 ;
        RECT 357.670 48.790 357.930 49.110 ;
        RECT 356.750 46.410 357.010 46.730 ;
        RECT 356.810 34.520 356.950 46.410 ;
        RECT 357.730 46.390 357.870 48.790 ;
        RECT 357.670 46.070 357.930 46.390 ;
        RECT 358.190 45.370 358.330 52.190 ;
        RECT 357.210 45.050 357.470 45.370 ;
        RECT 358.130 45.050 358.390 45.370 ;
        RECT 357.270 42.650 357.410 45.050 ;
        RECT 358.650 44.885 358.790 52.530 ;
        RECT 359.570 52.170 359.710 54.000 ;
        RECT 359.510 51.850 359.770 52.170 ;
        RECT 359.050 50.150 359.310 50.470 ;
        RECT 358.130 44.370 358.390 44.690 ;
        RECT 358.580 44.515 358.860 44.885 ;
        RECT 358.590 44.370 358.850 44.515 ;
        RECT 358.190 43.670 358.330 44.370 ;
        RECT 358.130 43.350 358.390 43.670 ;
        RECT 357.210 42.330 357.470 42.650 ;
        RECT 358.130 40.630 358.390 40.950 ;
        RECT 358.190 34.520 358.330 40.630 ;
        RECT 359.110 34.520 359.250 50.150 ;
        RECT 360.430 49.470 360.690 49.790 ;
        RECT 359.510 48.790 359.770 49.110 ;
        RECT 359.570 37.890 359.710 48.790 ;
        RECT 359.510 37.570 359.770 37.890 ;
        RECT 360.490 34.520 360.630 49.470 ;
        RECT 362.260 48.595 362.540 48.965 ;
        RECT 362.330 48.090 362.470 48.595 ;
        RECT 361.810 47.770 362.070 48.090 ;
        RECT 362.270 47.770 362.530 48.090 ;
        RECT 361.870 34.520 362.010 47.770 ;
        RECT 362.790 34.520 362.930 54.000 ;
        RECT 364.170 34.520 364.310 54.000 ;
        RECT 364.630 42.560 364.770 54.000 ;
        RECT 365.250 53.640 366.730 54.000 ;
        RECT 368.710 52.190 368.970 52.510 ;
        RECT 368.770 50.130 368.910 52.190 ;
        RECT 368.710 49.810 368.970 50.130 ;
        RECT 366.870 49.130 367.130 49.450 ;
        RECT 365.250 48.200 366.730 48.680 ;
        RECT 365.250 42.760 366.730 43.240 ;
        RECT 364.630 42.420 365.690 42.560 ;
        RECT 365.550 34.520 365.690 42.420 ;
        RECT 366.930 39.330 367.070 49.130 ;
        RECT 368.770 46.980 368.910 49.810 ;
        RECT 370.610 47.410 370.750 54.000 ;
        RECT 371.990 53.530 372.130 54.000 ;
        RECT 371.930 53.210 372.190 53.530 ;
        RECT 372.910 52.510 373.050 54.000 ;
        RECT 375.150 52.530 375.410 52.850 ;
        RECT 372.850 52.420 373.110 52.510 ;
        RECT 372.850 52.280 374.430 52.420 ;
        RECT 372.850 52.190 373.110 52.280 ;
        RECT 374.290 50.210 374.430 52.280 ;
        RECT 374.690 50.720 374.950 50.810 ;
        RECT 375.210 50.720 375.350 52.530 ;
        RECT 376.130 50.810 376.270 54.000 ;
        RECT 382.050 53.210 382.310 53.530 ;
        RECT 377.450 52.870 377.710 53.190 ;
        RECT 376.520 51.995 376.800 52.365 ;
        RECT 374.690 50.580 375.350 50.720 ;
        RECT 374.690 50.490 374.950 50.580 ;
        RECT 376.070 50.490 376.330 50.810 ;
        RECT 374.290 50.130 375.350 50.210 ;
        RECT 374.290 50.070 375.410 50.130 ;
        RECT 375.150 49.810 375.410 50.070 ;
        RECT 370.550 47.090 370.810 47.410 ;
        RECT 373.770 47.090 374.030 47.410 ;
        RECT 369.170 46.980 369.430 47.070 ;
        RECT 368.770 46.840 369.430 46.980 ;
        RECT 369.170 46.750 369.430 46.840 ;
        RECT 367.790 46.410 368.050 46.730 ;
        RECT 366.470 39.190 367.070 39.330 ;
        RECT 366.470 34.520 366.610 39.190 ;
        RECT 367.850 34.520 367.990 46.410 ;
        RECT 370.090 46.070 370.350 46.390 ;
        RECT 369.170 40.290 369.430 40.610 ;
        RECT 369.230 34.520 369.370 40.290 ;
        RECT 370.150 34.520 370.290 46.070 ;
        RECT 371.470 43.350 371.730 43.670 ;
        RECT 371.530 34.520 371.670 43.350 ;
        RECT 372.850 39.950 373.110 40.270 ;
        RECT 372.910 34.520 373.050 39.950 ;
        RECT 373.830 34.520 373.970 47.090 ;
        RECT 375.150 46.410 375.410 46.730 ;
        RECT 375.210 34.520 375.350 46.410 ;
        RECT 376.590 34.520 376.730 51.995 ;
        RECT 377.510 34.520 377.650 52.870 ;
        RECT 382.110 50.810 382.250 53.210 ;
        RECT 382.050 50.490 382.310 50.810 ;
        RECT 383.030 50.470 383.170 54.000 ;
        RECT 382.510 50.150 382.770 50.470 ;
        RECT 382.970 50.150 383.230 50.470 ;
        RECT 380.210 47.770 380.470 48.090 ;
        RECT 379.750 43.350 380.010 43.670 ;
        RECT 379.810 41.970 379.950 43.350 ;
        RECT 379.750 41.650 380.010 41.970 ;
        RECT 380.270 34.520 380.410 47.770 ;
        RECT 381.130 46.410 381.390 46.730 ;
        RECT 381.190 44.690 381.330 46.410 ;
        RECT 381.130 44.370 381.390 44.690 ;
        RECT 381.130 43.690 381.390 44.010 ;
        RECT 381.190 34.520 381.330 43.690 ;
        RECT 382.570 34.520 382.710 50.150 ;
        RECT 383.950 34.520 384.090 54.000 ;
        RECT 385.730 51.510 385.990 51.830 ;
        RECT 385.790 37.290 385.930 51.510 ;
        RECT 386.710 46.390 386.850 54.000 ;
        RECT 387.570 52.190 387.830 52.510 ;
        RECT 388.490 52.190 388.750 52.510 ;
        RECT 395.450 52.420 395.590 54.000 ;
        RECT 518.850 53.640 520.330 54.000 ;
        RECT 395.450 52.280 397.430 52.420 ;
        RECT 386.190 46.070 386.450 46.390 ;
        RECT 386.650 46.070 386.910 46.390 ;
        RECT 386.250 44.690 386.390 46.070 ;
        RECT 386.190 44.370 386.450 44.690 ;
        RECT 385.790 37.150 386.390 37.290 ;
        RECT 386.250 34.520 386.390 37.150 ;
        RECT 387.630 34.520 387.770 52.190 ;
        RECT 388.550 34.520 388.690 52.190 ;
        RECT 393.550 51.850 393.810 52.170 ;
        RECT 391.250 50.150 391.510 50.470 ;
        RECT 389.870 46.410 390.130 46.730 ;
        RECT 389.930 34.520 390.070 46.410 ;
        RECT 391.310 34.520 391.450 50.150 ;
        RECT 392.170 48.790 392.430 49.110 ;
        RECT 392.230 34.520 392.370 48.790 ;
        RECT 393.610 34.520 393.750 51.850 ;
        RECT 394.930 50.490 395.190 50.810 ;
        RECT 394.990 34.520 395.130 50.490 ;
        RECT 395.850 48.790 396.110 49.110 ;
        RECT 395.910 34.520 396.050 48.790 ;
        RECT 397.290 34.520 397.430 52.280 ;
        RECT 630.910 52.190 631.170 52.510 ;
        RECT 442.050 50.920 443.530 51.400 ;
        RECT 595.650 50.920 597.130 51.400 ;
        RECT 400.910 49.810 401.170 50.130 ;
        RECT 408.260 49.955 408.540 50.325 ;
        RECT 399.530 46.750 399.790 47.070 ;
        RECT 398.610 46.070 398.870 46.390 ;
        RECT 398.670 34.520 398.810 46.070 ;
        RECT 399.590 34.520 399.730 46.750 ;
        RECT 400.970 34.520 401.110 49.810 ;
        RECT 403.210 48.790 403.470 49.110 ;
        RECT 402.290 41.990 402.550 42.310 ;
        RECT 402.350 34.520 402.490 41.990 ;
        RECT 403.270 34.520 403.410 48.790 ;
        RECT 405.960 47.235 406.240 47.605 ;
        RECT 404.590 43.350 404.850 43.670 ;
        RECT 404.650 34.520 404.790 43.350 ;
        RECT 406.030 34.520 406.170 47.235 ;
        RECT 406.890 46.750 407.150 47.070 ;
        RECT 406.950 34.520 407.090 46.750 ;
        RECT 408.330 34.520 408.470 49.955 ;
        RECT 414.250 48.790 414.510 49.110 ;
        RECT 428.970 48.790 429.230 49.110 ;
        RECT 436.330 48.790 436.590 49.110 ;
        RECT 447.370 48.790 447.630 49.110 ;
        RECT 458.410 48.790 458.670 49.110 ;
        RECT 469.450 48.790 469.710 49.110 ;
        RECT 480.490 48.790 480.750 49.110 ;
        RECT 487.850 48.790 488.110 49.110 ;
        RECT 513.610 48.790 513.870 49.110 ;
        RECT 520.970 48.790 521.230 49.110 ;
        RECT 535.690 48.790 535.950 49.110 ;
        RECT 543.050 48.790 543.310 49.110 ;
        RECT 554.090 48.790 554.350 49.110 ;
        RECT 564.670 48.790 564.930 49.110 ;
        RECT 572.030 48.790 572.290 49.110 ;
        RECT 597.790 48.790 598.050 49.110 ;
        RECT 619.870 48.790 620.130 49.110 ;
        RECT 627.230 48.790 627.490 49.110 ;
        RECT 410.570 46.750 410.830 47.070 ;
        RECT 410.630 34.520 410.770 46.750 ;
        RECT 414.310 34.520 414.450 48.790 ;
        RECT 417.930 46.750 418.190 47.070 ;
        RECT 421.610 46.750 421.870 47.070 ;
        RECT 425.290 46.750 425.550 47.070 ;
        RECT 417.990 34.520 418.130 46.750 ;
        RECT 421.670 34.520 421.810 46.750 ;
        RECT 425.350 34.520 425.490 46.750 ;
        RECT 429.030 34.520 429.170 48.790 ;
        RECT 436.390 34.520 436.530 48.790 ;
        RECT 440.010 46.750 440.270 47.070 ;
        RECT 443.690 46.750 443.950 47.070 ;
        RECT 440.070 34.520 440.210 46.750 ;
        RECT 442.050 45.480 443.530 45.960 ;
        RECT 443.750 34.520 443.890 46.750 ;
        RECT 447.430 34.520 447.570 48.790 ;
        RECT 451.050 46.750 451.310 47.070 ;
        RECT 454.730 46.750 454.990 47.070 ;
        RECT 451.110 34.520 451.250 46.750 ;
        RECT 454.790 34.520 454.930 46.750 ;
        RECT 458.470 34.520 458.610 48.790 ;
        RECT 465.770 46.750 466.030 47.070 ;
        RECT 465.830 34.520 465.970 46.750 ;
        RECT 469.510 34.520 469.650 48.790 ;
        RECT 473.130 46.750 473.390 47.070 ;
        RECT 476.810 46.750 477.070 47.070 ;
        RECT 473.190 34.520 473.330 46.750 ;
        RECT 476.870 34.520 477.010 46.750 ;
        RECT 480.550 34.520 480.690 48.790 ;
        RECT 484.170 46.750 484.430 47.070 ;
        RECT 484.230 34.520 484.370 46.750 ;
        RECT 487.910 34.520 488.050 48.790 ;
        RECT 491.530 46.750 491.790 47.070 ;
        RECT 495.210 46.750 495.470 47.070 ;
        RECT 498.890 46.750 499.150 47.070 ;
        RECT 506.250 46.750 506.510 47.070 ;
        RECT 491.590 34.520 491.730 46.750 ;
        RECT 495.270 34.520 495.410 46.750 ;
        RECT 498.950 34.520 499.090 46.750 ;
        RECT 502.570 43.350 502.830 43.670 ;
        RECT 502.630 34.520 502.770 43.350 ;
        RECT 506.310 34.520 506.450 46.750 ;
        RECT 513.670 34.520 513.810 48.790 ;
        RECT 518.850 48.200 520.330 48.680 ;
        RECT 517.290 46.750 517.550 47.070 ;
        RECT 517.350 34.520 517.490 46.750 ;
        RECT 518.850 42.760 520.330 43.240 ;
        RECT 521.030 34.520 521.170 48.790 ;
        RECT 524.650 46.750 524.910 47.070 ;
        RECT 528.330 46.750 528.590 47.070 ;
        RECT 532.010 46.750 532.270 47.070 ;
        RECT 524.710 34.520 524.850 46.750 ;
        RECT 528.390 34.520 528.530 46.750 ;
        RECT 532.070 34.520 532.210 46.750 ;
        RECT 535.750 34.520 535.890 48.790 ;
        RECT 539.370 46.750 539.630 47.070 ;
        RECT 539.430 34.520 539.570 46.750 ;
        RECT 543.110 34.520 543.250 48.790 ;
        RECT 546.730 46.750 546.990 47.070 ;
        RECT 550.410 46.750 550.670 47.070 ;
        RECT 546.790 34.520 546.930 46.750 ;
        RECT 550.470 34.520 550.610 46.750 ;
        RECT 554.150 34.520 554.290 48.790 ;
        RECT 557.770 46.750 558.030 47.070 ;
        RECT 561.450 46.750 561.710 47.070 ;
        RECT 557.830 34.520 557.970 46.750 ;
        RECT 561.510 34.520 561.650 46.750 ;
        RECT 564.730 34.520 564.870 48.790 ;
        RECT 568.350 46.750 568.610 47.070 ;
        RECT 568.410 34.520 568.550 46.750 ;
        RECT 572.090 34.520 572.230 48.790 ;
        RECT 575.710 46.750 575.970 47.070 ;
        RECT 579.390 46.750 579.650 47.070 ;
        RECT 583.070 46.750 583.330 47.070 ;
        RECT 590.430 46.750 590.690 47.070 ;
        RECT 594.110 46.750 594.370 47.070 ;
        RECT 575.770 34.520 575.910 46.750 ;
        RECT 579.450 34.520 579.590 46.750 ;
        RECT 583.130 34.520 583.270 46.750 ;
        RECT 586.750 43.350 587.010 43.670 ;
        RECT 586.810 34.520 586.950 43.350 ;
        RECT 590.490 34.520 590.630 46.750 ;
        RECT 594.170 34.520 594.310 46.750 ;
        RECT 595.650 45.480 597.130 45.960 ;
        RECT 597.850 34.520 597.990 48.790 ;
        RECT 601.470 46.750 601.730 47.070 ;
        RECT 608.830 46.750 609.090 47.070 ;
        RECT 612.510 46.750 612.770 47.070 ;
        RECT 616.190 46.750 616.450 47.070 ;
        RECT 601.530 34.520 601.670 46.750 ;
        RECT 608.890 34.520 609.030 46.750 ;
        RECT 612.570 34.520 612.710 46.750 ;
        RECT 616.250 34.520 616.390 46.750 ;
        RECT 619.930 34.520 620.070 48.790 ;
        RECT 623.550 46.750 623.810 47.070 ;
        RECT 623.610 34.520 623.750 46.750 ;
        RECT 627.290 34.520 627.430 48.790 ;
        RECT 630.970 34.520 631.110 52.190 ;
        RECT 37.500 32.120 37.780 34.520 ;
        RECT 38.420 32.120 38.700 34.520 ;
        RECT 39.800 32.120 40.080 34.520 ;
        RECT 40.720 32.120 41.000 34.520 ;
        RECT 42.100 32.120 42.380 34.520 ;
        RECT 43.480 32.120 43.760 34.520 ;
        RECT 44.400 32.120 44.680 34.520 ;
        RECT 47.160 32.120 47.440 34.520 ;
        RECT 48.080 32.120 48.360 34.520 ;
        RECT 49.460 32.120 49.740 34.520 ;
        RECT 50.840 32.120 51.120 34.520 ;
        RECT 53.140 32.120 53.420 34.520 ;
        RECT 54.520 32.120 54.800 34.520 ;
        RECT 55.440 32.120 55.720 34.520 ;
        RECT 56.820 32.120 57.100 34.520 ;
        RECT 58.200 32.120 58.480 34.520 ;
        RECT 59.120 32.120 59.400 34.520 ;
        RECT 60.500 32.120 60.780 34.520 ;
        RECT 61.880 32.120 62.160 34.520 ;
        RECT 62.800 32.120 63.080 34.520 ;
        RECT 64.180 32.120 64.460 34.520 ;
        RECT 65.560 32.120 65.840 34.520 ;
        RECT 66.480 32.120 66.760 34.520 ;
        RECT 67.860 32.120 68.140 34.520 ;
        RECT 69.240 32.120 69.520 34.520 ;
        RECT 70.160 32.120 70.440 34.520 ;
        RECT 71.540 32.120 71.820 34.520 ;
        RECT 72.920 32.120 73.200 34.520 ;
        RECT 73.840 32.120 74.120 34.520 ;
        RECT 75.220 32.120 75.500 34.520 ;
        RECT 76.600 32.120 76.880 34.520 ;
        RECT 77.520 32.120 77.800 34.520 ;
        RECT 78.900 32.120 79.180 34.520 ;
        RECT 80.280 32.120 80.560 34.520 ;
        RECT 81.200 32.120 81.480 34.520 ;
        RECT 82.580 32.120 82.860 34.520 ;
        RECT 83.960 32.120 84.240 34.520 ;
        RECT 84.880 32.120 85.160 34.520 ;
        RECT 86.260 32.120 86.540 34.520 ;
        RECT 88.560 32.120 88.840 34.520 ;
        RECT 89.940 32.120 90.220 34.520 ;
        RECT 91.320 32.120 91.600 34.520 ;
        RECT 92.240 32.120 92.520 34.520 ;
        RECT 95.000 32.120 95.280 34.520 ;
        RECT 95.920 32.120 96.200 34.520 ;
        RECT 97.300 32.120 97.580 34.520 ;
        RECT 98.680 32.120 98.960 34.520 ;
        RECT 100.980 32.120 101.260 34.520 ;
        RECT 102.360 32.120 102.640 34.520 ;
        RECT 103.280 32.120 103.560 34.520 ;
        RECT 104.660 32.120 104.940 34.520 ;
        RECT 106.040 32.120 106.320 34.520 ;
        RECT 106.960 32.120 107.240 34.520 ;
        RECT 108.340 32.120 108.620 34.520 ;
        RECT 109.720 32.120 110.000 34.520 ;
        RECT 110.640 32.120 110.920 34.520 ;
        RECT 112.020 32.120 112.300 34.520 ;
        RECT 112.940 32.120 113.220 34.520 ;
        RECT 114.320 32.120 114.600 34.520 ;
        RECT 115.700 32.120 115.980 34.520 ;
        RECT 116.620 32.120 116.900 34.520 ;
        RECT 118.000 32.120 118.280 34.520 ;
        RECT 119.380 32.120 119.660 34.520 ;
        RECT 120.300 32.120 120.580 34.520 ;
        RECT 121.680 32.120 121.960 34.520 ;
        RECT 123.060 32.120 123.340 34.520 ;
        RECT 123.980 32.120 124.260 34.520 ;
        RECT 125.360 32.120 125.640 34.520 ;
        RECT 126.740 32.120 127.020 34.520 ;
        RECT 127.660 32.120 127.940 34.520 ;
        RECT 130.420 32.120 130.700 34.520 ;
        RECT 131.340 32.120 131.620 34.520 ;
        RECT 132.720 32.120 133.000 34.520 ;
        RECT 134.100 32.120 134.380 34.520 ;
        RECT 136.400 32.120 136.680 34.520 ;
        RECT 137.780 32.120 138.060 34.520 ;
        RECT 138.700 32.120 138.980 34.520 ;
        RECT 140.080 32.120 140.360 34.520 ;
        RECT 141.460 32.120 141.740 34.520 ;
        RECT 142.380 32.120 142.660 34.520 ;
        RECT 143.760 32.120 144.040 34.520 ;
        RECT 145.140 32.120 145.420 34.520 ;
        RECT 146.060 32.120 146.340 34.520 ;
        RECT 147.440 32.120 147.720 34.520 ;
        RECT 148.820 32.120 149.100 34.520 ;
        RECT 149.740 32.120 150.020 34.520 ;
        RECT 151.120 32.120 151.400 34.520 ;
        RECT 152.500 32.120 152.780 34.520 ;
        RECT 153.420 32.120 153.700 34.520 ;
        RECT 154.800 32.120 155.080 34.520 ;
        RECT 156.180 32.120 156.460 34.520 ;
        RECT 157.100 32.120 157.380 34.520 ;
        RECT 158.480 32.120 158.760 34.520 ;
        RECT 159.860 32.120 160.140 34.520 ;
        RECT 160.780 32.120 161.060 34.520 ;
        RECT 162.160 32.120 162.440 34.520 ;
        RECT 163.540 32.120 163.820 34.520 ;
        RECT 164.460 32.120 164.740 34.520 ;
        RECT 165.840 32.120 166.120 34.520 ;
        RECT 167.220 32.120 167.500 34.520 ;
        RECT 168.140 32.120 168.420 34.520 ;
        RECT 169.520 32.120 169.800 34.520 ;
        RECT 171.820 32.120 172.100 34.520 ;
        RECT 173.200 32.120 173.480 34.520 ;
        RECT 174.580 32.120 174.860 34.520 ;
        RECT 175.500 32.120 175.780 34.520 ;
        RECT 178.260 32.120 178.540 34.520 ;
        RECT 179.180 32.120 179.460 34.520 ;
        RECT 180.560 32.120 180.840 34.520 ;
        RECT 181.940 32.120 182.220 34.520 ;
        RECT 184.240 32.120 184.520 34.520 ;
        RECT 185.620 32.120 185.900 34.520 ;
        RECT 186.540 32.120 186.820 34.520 ;
        RECT 187.920 32.120 188.200 34.520 ;
        RECT 190.220 32.120 190.500 34.520 ;
        RECT 191.600 32.120 191.880 34.520 ;
        RECT 192.520 32.120 192.800 34.520 ;
        RECT 193.900 32.120 194.180 34.520 ;
        RECT 195.280 32.120 195.560 34.520 ;
        RECT 196.200 32.120 196.480 34.520 ;
        RECT 197.580 32.120 197.860 34.520 ;
        RECT 198.960 32.120 199.240 34.520 ;
        RECT 199.880 32.120 200.160 34.520 ;
        RECT 201.260 32.120 201.540 34.520 ;
        RECT 202.640 32.120 202.920 34.520 ;
        RECT 203.560 32.120 203.840 34.520 ;
        RECT 204.940 32.120 205.220 34.520 ;
        RECT 206.320 32.120 206.600 34.520 ;
        RECT 207.240 32.120 207.520 34.520 ;
        RECT 208.620 32.120 208.900 34.520 ;
        RECT 210.000 32.120 210.280 34.520 ;
        RECT 210.920 32.120 211.200 34.520 ;
        RECT 213.680 32.120 213.960 34.520 ;
        RECT 214.600 32.120 214.880 34.520 ;
        RECT 215.980 32.120 216.260 34.520 ;
        RECT 217.360 32.120 217.640 34.520 ;
        RECT 219.660 32.120 219.940 34.520 ;
        RECT 221.040 32.120 221.320 34.520 ;
        RECT 221.960 32.120 222.240 34.520 ;
        RECT 223.340 32.120 223.620 34.520 ;
        RECT 224.720 32.120 225.000 34.520 ;
        RECT 225.640 32.120 225.920 34.520 ;
        RECT 227.020 32.120 227.300 34.520 ;
        RECT 228.400 32.120 228.680 34.520 ;
        RECT 229.320 32.120 229.600 34.520 ;
        RECT 230.700 32.120 230.980 34.520 ;
        RECT 232.080 32.120 232.360 34.520 ;
        RECT 233.000 32.120 233.280 34.520 ;
        RECT 234.380 32.120 234.660 34.520 ;
        RECT 235.760 32.120 236.040 34.520 ;
        RECT 236.680 32.120 236.960 34.520 ;
        RECT 238.060 32.120 238.340 34.520 ;
        RECT 239.440 32.120 239.720 34.520 ;
        RECT 240.360 32.120 240.640 34.520 ;
        RECT 241.740 32.120 242.020 34.520 ;
        RECT 243.120 32.120 243.400 34.520 ;
        RECT 244.040 32.120 244.320 34.520 ;
        RECT 245.420 32.120 245.700 34.520 ;
        RECT 246.800 32.120 247.080 34.520 ;
        RECT 247.720 32.120 248.000 34.520 ;
        RECT 249.100 32.120 249.380 34.520 ;
        RECT 250.480 32.120 250.760 34.520 ;
        RECT 251.400 32.120 251.680 34.520 ;
        RECT 252.780 32.120 253.060 34.520 ;
        RECT 255.080 32.120 255.360 34.520 ;
        RECT 256.460 32.120 256.740 34.520 ;
        RECT 257.840 32.120 258.120 34.520 ;
        RECT 258.760 32.120 259.040 34.520 ;
        RECT 261.520 32.120 261.800 34.520 ;
        RECT 262.440 32.120 262.720 34.520 ;
        RECT 263.820 32.120 264.100 34.520 ;
        RECT 264.740 32.120 265.020 34.520 ;
        RECT 267.500 32.120 267.780 34.520 ;
        RECT 268.420 32.120 268.700 34.520 ;
        RECT 269.800 32.120 270.080 34.520 ;
        RECT 271.180 32.120 271.460 34.520 ;
        RECT 273.480 32.120 273.760 34.520 ;
        RECT 274.860 32.120 275.140 34.520 ;
        RECT 275.780 32.120 276.060 34.520 ;
        RECT 277.160 32.120 277.440 34.520 ;
        RECT 278.540 32.120 278.820 34.520 ;
        RECT 279.460 32.120 279.740 34.520 ;
        RECT 280.840 32.120 281.120 34.520 ;
        RECT 282.220 32.120 282.500 34.520 ;
        RECT 283.140 32.120 283.420 34.520 ;
        RECT 284.520 32.120 284.800 34.520 ;
        RECT 285.900 32.120 286.180 34.520 ;
        RECT 286.820 32.120 287.100 34.520 ;
        RECT 288.200 32.120 288.480 34.520 ;
        RECT 289.580 32.120 289.860 34.520 ;
        RECT 290.500 32.120 290.780 34.520 ;
        RECT 291.880 32.120 292.160 34.520 ;
        RECT 293.260 32.120 293.540 34.520 ;
        RECT 294.180 32.120 294.460 34.520 ;
        RECT 296.940 32.120 297.220 34.520 ;
        RECT 297.860 32.120 298.140 34.520 ;
        RECT 299.240 32.120 299.520 34.520 ;
        RECT 300.620 32.120 300.900 34.520 ;
        RECT 302.920 32.120 303.200 34.520 ;
        RECT 304.300 32.120 304.580 34.520 ;
        RECT 305.220 32.120 305.500 34.520 ;
        RECT 306.600 32.120 306.880 34.520 ;
        RECT 307.980 32.120 308.260 34.520 ;
        RECT 308.900 32.120 309.180 34.520 ;
        RECT 310.280 32.120 310.560 34.520 ;
        RECT 311.660 32.120 311.940 34.520 ;
        RECT 312.580 32.120 312.860 34.520 ;
        RECT 313.960 32.120 314.240 34.520 ;
        RECT 315.340 32.120 315.620 34.520 ;
        RECT 316.260 32.120 316.540 34.520 ;
        RECT 317.640 32.120 317.920 34.520 ;
        RECT 319.020 32.120 319.300 34.520 ;
        RECT 319.940 32.120 320.220 34.520 ;
        RECT 321.320 32.120 321.600 34.520 ;
        RECT 322.700 32.120 322.980 34.520 ;
        RECT 323.620 32.120 323.900 34.520 ;
        RECT 325.000 32.120 325.280 34.520 ;
        RECT 326.380 32.120 326.660 34.520 ;
        RECT 327.300 32.120 327.580 34.520 ;
        RECT 328.680 32.120 328.960 34.520 ;
        RECT 330.060 32.120 330.340 34.520 ;
        RECT 330.980 32.120 331.260 34.520 ;
        RECT 332.360 32.120 332.640 34.520 ;
        RECT 333.740 32.120 334.020 34.520 ;
        RECT 334.660 32.120 334.940 34.520 ;
        RECT 336.040 32.120 336.320 34.520 ;
        RECT 338.340 32.120 338.620 34.520 ;
        RECT 339.720 32.120 340.000 34.520 ;
        RECT 340.640 32.120 340.920 34.520 ;
        RECT 342.020 32.120 342.300 34.520 ;
        RECT 344.320 32.120 344.600 34.520 ;
        RECT 345.700 32.120 345.980 34.520 ;
        RECT 347.080 32.120 347.360 34.520 ;
        RECT 348.000 32.120 348.280 34.520 ;
        RECT 350.760 32.120 351.040 34.520 ;
        RECT 351.680 32.120 351.960 34.520 ;
        RECT 353.060 32.120 353.340 34.520 ;
        RECT 354.440 32.120 354.720 34.520 ;
        RECT 356.740 32.120 357.020 34.520 ;
        RECT 358.120 32.120 358.400 34.520 ;
        RECT 359.040 32.120 359.320 34.520 ;
        RECT 360.420 32.120 360.700 34.520 ;
        RECT 361.800 32.120 362.080 34.520 ;
        RECT 362.720 32.120 363.000 34.520 ;
        RECT 364.100 32.120 364.380 34.520 ;
        RECT 365.480 32.120 365.760 34.520 ;
        RECT 366.400 32.120 366.680 34.520 ;
        RECT 367.780 32.120 368.060 34.520 ;
        RECT 369.160 32.120 369.440 34.520 ;
        RECT 370.080 32.120 370.360 34.520 ;
        RECT 371.460 32.120 371.740 34.520 ;
        RECT 372.840 32.120 373.120 34.520 ;
        RECT 373.760 32.120 374.040 34.520 ;
        RECT 375.140 32.120 375.420 34.520 ;
        RECT 376.520 32.120 376.800 34.520 ;
        RECT 377.440 32.120 377.720 34.520 ;
        RECT 380.200 32.120 380.480 34.520 ;
        RECT 381.120 32.120 381.400 34.520 ;
        RECT 382.500 32.120 382.780 34.520 ;
        RECT 383.880 32.120 384.160 34.520 ;
        RECT 386.180 32.120 386.460 34.520 ;
        RECT 387.560 32.120 387.840 34.520 ;
        RECT 388.480 32.120 388.760 34.520 ;
        RECT 389.860 32.120 390.140 34.520 ;
        RECT 391.240 32.120 391.520 34.520 ;
        RECT 392.160 32.120 392.440 34.520 ;
        RECT 393.540 32.120 393.820 34.520 ;
        RECT 394.920 32.120 395.200 34.520 ;
        RECT 395.840 32.120 396.120 34.520 ;
        RECT 397.220 32.120 397.500 34.520 ;
        RECT 398.600 32.120 398.880 34.520 ;
        RECT 399.520 32.120 399.800 34.520 ;
        RECT 400.900 32.120 401.180 34.520 ;
        RECT 402.280 32.120 402.560 34.520 ;
        RECT 403.200 32.120 403.480 34.520 ;
        RECT 404.580 32.120 404.860 34.520 ;
        RECT 405.960 32.120 406.240 34.520 ;
        RECT 406.880 32.120 407.160 34.520 ;
        RECT 408.260 32.120 408.540 34.520 ;
        RECT 409.640 32.120 409.920 34.520 ;
        RECT 410.560 32.120 410.840 34.520 ;
        RECT 411.940 32.120 412.220 34.520 ;
        RECT 412.860 32.120 413.140 34.520 ;
        RECT 414.240 32.120 414.520 34.520 ;
        RECT 415.620 32.120 415.900 34.520 ;
        RECT 416.540 32.120 416.820 34.520 ;
        RECT 417.920 32.120 418.200 34.520 ;
        RECT 419.300 32.120 419.580 34.520 ;
        RECT 420.220 32.120 420.500 34.520 ;
        RECT 421.600 32.120 421.880 34.520 ;
        RECT 422.980 32.120 423.260 34.520 ;
        RECT 423.900 32.120 424.180 34.520 ;
        RECT 425.280 32.120 425.560 34.520 ;
        RECT 427.580 32.120 427.860 34.520 ;
        RECT 428.960 32.120 429.240 34.520 ;
        RECT 430.340 32.120 430.620 34.520 ;
        RECT 431.260 32.120 431.540 34.520 ;
        RECT 434.020 32.120 434.300 34.520 ;
        RECT 434.940 32.120 435.220 34.520 ;
        RECT 436.320 32.120 436.600 34.520 ;
        RECT 437.700 32.120 437.980 34.520 ;
        RECT 440.000 32.120 440.280 34.520 ;
        RECT 441.380 32.120 441.660 34.520 ;
        RECT 442.300 32.120 442.580 34.520 ;
        RECT 443.680 32.120 443.960 34.520 ;
        RECT 445.060 32.120 445.340 34.520 ;
        RECT 445.980 32.120 446.260 34.520 ;
        RECT 447.360 32.120 447.640 34.520 ;
        RECT 448.740 32.120 449.020 34.520 ;
        RECT 449.660 32.120 449.940 34.520 ;
        RECT 451.040 32.120 451.320 34.520 ;
        RECT 452.420 32.120 452.700 34.520 ;
        RECT 453.340 32.120 453.620 34.520 ;
        RECT 454.720 32.120 455.000 34.520 ;
        RECT 456.100 32.120 456.380 34.520 ;
        RECT 457.020 32.120 457.300 34.520 ;
        RECT 458.400 32.120 458.680 34.520 ;
        RECT 459.780 32.120 460.060 34.520 ;
        RECT 460.700 32.120 460.980 34.520 ;
        RECT 463.460 32.120 463.740 34.520 ;
        RECT 464.380 32.120 464.660 34.520 ;
        RECT 465.760 32.120 466.040 34.520 ;
        RECT 467.140 32.120 467.420 34.520 ;
        RECT 469.440 32.120 469.720 34.520 ;
        RECT 470.820 32.120 471.100 34.520 ;
        RECT 471.740 32.120 472.020 34.520 ;
        RECT 473.120 32.120 473.400 34.520 ;
        RECT 474.500 32.120 474.780 34.520 ;
        RECT 475.420 32.120 475.700 34.520 ;
        RECT 476.800 32.120 477.080 34.520 ;
        RECT 478.180 32.120 478.460 34.520 ;
        RECT 479.100 32.120 479.380 34.520 ;
        RECT 480.480 32.120 480.760 34.520 ;
        RECT 481.860 32.120 482.140 34.520 ;
        RECT 482.780 32.120 483.060 34.520 ;
        RECT 484.160 32.120 484.440 34.520 ;
        RECT 485.540 32.120 485.820 34.520 ;
        RECT 486.460 32.120 486.740 34.520 ;
        RECT 487.840 32.120 488.120 34.520 ;
        RECT 488.760 32.120 489.040 34.520 ;
        RECT 490.140 32.120 490.420 34.520 ;
        RECT 491.520 32.120 491.800 34.520 ;
        RECT 492.440 32.120 492.720 34.520 ;
        RECT 493.820 32.120 494.100 34.520 ;
        RECT 495.200 32.120 495.480 34.520 ;
        RECT 496.120 32.120 496.400 34.520 ;
        RECT 497.500 32.120 497.780 34.520 ;
        RECT 498.880 32.120 499.160 34.520 ;
        RECT 499.800 32.120 500.080 34.520 ;
        RECT 501.180 32.120 501.460 34.520 ;
        RECT 502.560 32.120 502.840 34.520 ;
        RECT 503.480 32.120 503.760 34.520 ;
        RECT 504.860 32.120 505.140 34.520 ;
        RECT 506.240 32.120 506.520 34.520 ;
        RECT 507.160 32.120 507.440 34.520 ;
        RECT 508.540 32.120 508.820 34.520 ;
        RECT 510.840 32.120 511.120 34.520 ;
        RECT 512.220 32.120 512.500 34.520 ;
        RECT 513.600 32.120 513.880 34.520 ;
        RECT 514.520 32.120 514.800 34.520 ;
        RECT 517.280 32.120 517.560 34.520 ;
        RECT 518.200 32.120 518.480 34.520 ;
        RECT 519.580 32.120 519.860 34.520 ;
        RECT 520.960 32.120 521.240 34.520 ;
        RECT 523.260 32.120 523.540 34.520 ;
        RECT 524.640 32.120 524.920 34.520 ;
        RECT 525.560 32.120 525.840 34.520 ;
        RECT 526.940 32.120 527.220 34.520 ;
        RECT 528.320 32.120 528.600 34.520 ;
        RECT 529.240 32.120 529.520 34.520 ;
        RECT 530.620 32.120 530.900 34.520 ;
        RECT 532.000 32.120 532.280 34.520 ;
        RECT 532.920 32.120 533.200 34.520 ;
        RECT 534.300 32.120 534.580 34.520 ;
        RECT 535.680 32.120 535.960 34.520 ;
        RECT 536.600 32.120 536.880 34.520 ;
        RECT 537.980 32.120 538.260 34.520 ;
        RECT 539.360 32.120 539.640 34.520 ;
        RECT 540.280 32.120 540.560 34.520 ;
        RECT 541.660 32.120 541.940 34.520 ;
        RECT 543.040 32.120 543.320 34.520 ;
        RECT 543.960 32.120 544.240 34.520 ;
        RECT 546.720 32.120 547.000 34.520 ;
        RECT 547.640 32.120 547.920 34.520 ;
        RECT 549.020 32.120 549.300 34.520 ;
        RECT 550.400 32.120 550.680 34.520 ;
        RECT 552.700 32.120 552.980 34.520 ;
        RECT 554.080 32.120 554.360 34.520 ;
        RECT 555.000 32.120 555.280 34.520 ;
        RECT 556.380 32.120 556.660 34.520 ;
        RECT 557.760 32.120 558.040 34.520 ;
        RECT 558.680 32.120 558.960 34.520 ;
        RECT 560.060 32.120 560.340 34.520 ;
        RECT 561.440 32.120 561.720 34.520 ;
        RECT 562.360 32.120 562.640 34.520 ;
        RECT 563.740 32.120 564.020 34.520 ;
        RECT 564.660 32.120 564.940 34.520 ;
        RECT 566.040 32.120 566.320 34.520 ;
        RECT 567.420 32.120 567.700 34.520 ;
        RECT 568.340 32.120 568.620 34.520 ;
        RECT 569.720 32.120 570.000 34.520 ;
        RECT 571.100 32.120 571.380 34.520 ;
        RECT 572.020 32.120 572.300 34.520 ;
        RECT 573.400 32.120 573.680 34.520 ;
        RECT 574.780 32.120 575.060 34.520 ;
        RECT 575.700 32.120 575.980 34.520 ;
        RECT 577.080 32.120 577.360 34.520 ;
        RECT 578.460 32.120 578.740 34.520 ;
        RECT 579.380 32.120 579.660 34.520 ;
        RECT 580.760 32.120 581.040 34.520 ;
        RECT 582.140 32.120 582.420 34.520 ;
        RECT 583.060 32.120 583.340 34.520 ;
        RECT 584.440 32.120 584.720 34.520 ;
        RECT 585.820 32.120 586.100 34.520 ;
        RECT 586.740 32.120 587.020 34.520 ;
        RECT 588.120 32.120 588.400 34.520 ;
        RECT 589.500 32.120 589.780 34.520 ;
        RECT 590.420 32.120 590.700 34.520 ;
        RECT 591.800 32.120 592.080 34.520 ;
        RECT 594.100 32.120 594.380 34.520 ;
        RECT 595.480 32.120 595.760 34.520 ;
        RECT 596.860 32.120 597.140 34.520 ;
        RECT 597.780 32.120 598.060 34.520 ;
        RECT 600.540 32.120 600.820 34.520 ;
        RECT 601.460 32.120 601.740 34.520 ;
        RECT 602.840 32.120 603.120 34.520 ;
        RECT 604.220 32.120 604.500 34.520 ;
        RECT 606.520 32.120 606.800 34.520 ;
        RECT 607.900 32.120 608.180 34.520 ;
        RECT 608.820 32.120 609.100 34.520 ;
        RECT 610.200 32.120 610.480 34.520 ;
        RECT 611.580 32.120 611.860 34.520 ;
        RECT 612.500 32.120 612.780 34.520 ;
        RECT 613.880 32.120 614.160 34.520 ;
        RECT 615.260 32.120 615.540 34.520 ;
        RECT 616.180 32.120 616.460 34.520 ;
        RECT 617.560 32.120 617.840 34.520 ;
        RECT 618.940 32.120 619.220 34.520 ;
        RECT 619.860 32.120 620.140 34.520 ;
        RECT 621.240 32.120 621.520 34.520 ;
        RECT 622.620 32.120 622.900 34.520 ;
        RECT 623.540 32.120 623.820 34.520 ;
        RECT 624.920 32.120 625.200 34.520 ;
        RECT 626.300 32.120 626.580 34.520 ;
        RECT 627.220 32.120 627.500 34.520 ;
        RECT 629.980 32.120 630.260 34.520 ;
        RECT 630.900 32.120 631.180 34.520 ;
        RECT 632.280 32.120 632.560 34.520 ;
        RECT 633.660 32.120 633.940 34.520 ;
        RECT 635.960 32.120 636.240 34.520 ;
      LAYER via2 ;
        RECT 58.050 53.740 58.330 54.010 ;
        RECT 58.450 53.740 58.730 54.010 ;
        RECT 58.850 53.740 59.130 54.010 ;
        RECT 59.250 53.740 59.530 54.010 ;
        RECT 38.420 46.600 38.700 46.880 ;
        RECT 58.050 48.300 58.330 48.580 ;
        RECT 58.450 48.300 58.730 48.580 ;
        RECT 58.850 48.300 59.130 48.580 ;
        RECT 59.250 48.300 59.530 48.580 ;
        RECT 58.050 42.860 58.330 43.140 ;
        RECT 58.450 42.860 58.730 43.140 ;
        RECT 58.850 42.860 59.130 43.140 ;
        RECT 59.250 42.860 59.530 43.140 ;
        RECT 72.460 50.000 72.740 50.280 ;
        RECT 69.240 49.320 69.520 49.600 ;
        RECT 77.060 50.680 77.340 50.960 ;
        RECT 78.900 49.320 79.180 49.600 ;
        RECT 84.420 49.320 84.700 49.600 ;
        RECT 81.200 48.640 81.480 48.920 ;
        RECT 90.860 44.560 91.140 44.840 ;
        RECT 93.620 50.000 93.900 50.280 ;
        RECT 96.840 50.000 97.120 50.280 ;
        RECT 99.140 53.400 99.420 53.680 ;
        RECT 98.220 47.280 98.500 47.560 ;
        RECT 103.280 53.400 103.560 53.680 ;
        RECT 103.280 52.720 103.560 53.000 ;
        RECT 108.800 50.680 109.080 50.960 ;
        RECT 109.720 51.360 110.000 51.640 ;
        RECT 109.720 48.640 110.000 48.920 ;
        RECT 110.640 52.040 110.920 52.320 ;
        RECT 114.320 51.360 114.600 51.640 ;
        RECT 114.780 50.000 115.060 50.280 ;
        RECT 114.320 49.320 114.600 49.600 ;
        RECT 116.160 48.640 116.440 48.920 ;
        RECT 119.380 48.640 119.660 48.920 ;
        RECT 119.380 43.880 119.660 44.160 ;
        RECT 125.820 51.360 126.100 51.640 ;
        RECT 127.660 52.720 127.940 53.000 ;
        RECT 127.660 44.560 127.940 44.840 ;
        RECT 129.040 43.880 129.320 44.160 ;
        RECT 130.880 47.280 131.160 47.560 ;
        RECT 132.260 51.360 132.540 51.640 ;
        RECT 134.850 51.020 135.130 51.300 ;
        RECT 135.250 51.020 135.530 51.300 ;
        RECT 135.650 51.020 135.930 51.300 ;
        RECT 136.050 51.020 136.330 51.300 ;
        RECT 136.400 48.640 136.680 48.920 ;
        RECT 134.850 45.580 135.130 45.860 ;
        RECT 135.250 45.580 135.530 45.860 ;
        RECT 135.650 45.580 135.930 45.860 ;
        RECT 136.050 45.580 136.330 45.860 ;
        RECT 140.080 47.280 140.360 47.560 ;
        RECT 145.600 53.400 145.880 53.680 ;
        RECT 146.520 52.040 146.800 52.320 ;
        RECT 150.660 52.040 150.940 52.320 ;
        RECT 152.500 51.360 152.780 51.640 ;
        RECT 154.800 51.360 155.080 51.640 ;
        RECT 151.120 48.640 151.400 48.920 ;
        RECT 158.020 52.040 158.300 52.320 ;
        RECT 156.640 49.320 156.920 49.600 ;
        RECT 158.940 52.720 159.220 53.000 ;
        RECT 159.400 50.000 159.680 50.280 ;
        RECT 158.020 47.280 158.300 47.560 ;
        RECT 158.940 47.280 159.220 47.560 ;
        RECT 162.160 50.680 162.440 50.960 ;
        RECT 164.920 50.000 165.200 50.280 ;
        RECT 170.440 52.720 170.720 53.000 ;
        RECT 176.420 49.320 176.700 49.600 ;
        RECT 177.800 52.720 178.080 53.000 ;
        RECT 185.160 52.040 185.440 52.320 ;
        RECT 188.840 51.360 189.120 51.640 ;
        RECT 189.760 51.360 190.040 51.640 ;
        RECT 185.160 44.560 185.440 44.840 ;
        RECT 188.840 47.960 189.120 48.240 ;
        RECT 190.680 52.040 190.960 52.320 ;
        RECT 194.820 52.040 195.100 52.320 ;
        RECT 196.200 52.040 196.480 52.320 ;
        RECT 195.280 49.320 195.560 49.600 ;
        RECT 201.260 52.040 201.540 52.320 ;
        RECT 199.420 51.360 199.700 51.640 ;
        RECT 194.820 45.920 195.100 46.200 ;
        RECT 193.900 45.240 194.180 45.520 ;
        RECT 201.720 48.640 202.000 48.920 ;
        RECT 204.020 51.360 204.300 51.640 ;
        RECT 199.420 45.920 199.700 46.200 ;
        RECT 208.620 52.040 208.900 52.320 ;
        RECT 211.650 53.740 211.930 54.010 ;
        RECT 212.050 53.740 212.330 54.010 ;
        RECT 212.450 53.740 212.730 54.010 ;
        RECT 212.850 53.740 213.130 54.010 ;
        RECT 214.140 52.720 214.420 53.000 ;
        RECT 212.300 51.360 212.580 51.640 ;
        RECT 210.460 50.680 210.740 50.960 ;
        RECT 214.140 50.680 214.420 50.960 ;
        RECT 211.650 48.300 211.930 48.580 ;
        RECT 212.050 48.300 212.330 48.580 ;
        RECT 212.450 48.300 212.730 48.580 ;
        RECT 212.850 48.300 213.130 48.580 ;
        RECT 214.600 49.320 214.880 49.600 ;
        RECT 215.980 51.360 216.260 51.640 ;
        RECT 211.650 42.860 211.930 43.140 ;
        RECT 212.050 42.860 212.330 43.140 ;
        RECT 212.450 42.860 212.730 43.140 ;
        RECT 212.850 42.860 213.130 43.140 ;
        RECT 220.120 47.280 220.400 47.560 ;
        RECT 223.800 41.840 224.080 42.120 ;
        RECT 225.180 52.720 225.460 53.000 ;
        RECT 225.640 49.320 225.920 49.600 ;
        RECT 228.860 52.720 229.140 53.000 ;
        RECT 230.700 50.000 230.980 50.280 ;
        RECT 231.160 47.960 231.440 48.240 ;
        RECT 228.400 45.240 228.680 45.520 ;
        RECT 229.780 44.560 230.060 44.840 ;
        RECT 236.220 52.040 236.500 52.320 ;
        RECT 234.840 47.960 235.120 48.240 ;
        RECT 238.060 52.040 238.340 52.320 ;
        RECT 238.060 51.360 238.340 51.640 ;
        RECT 240.360 47.280 240.640 47.560 ;
        RECT 241.280 50.000 241.560 50.280 ;
        RECT 243.120 52.720 243.400 53.000 ;
        RECT 243.120 49.320 243.400 49.600 ;
        RECT 244.500 47.960 244.780 48.240 ;
        RECT 243.580 47.280 243.860 47.560 ;
        RECT 250.020 50.680 250.300 50.960 ;
        RECT 251.860 52.720 252.140 53.000 ;
        RECT 250.940 50.680 251.220 50.960 ;
        RECT 254.160 52.720 254.440 53.000 ;
        RECT 252.320 48.640 252.600 48.920 ;
        RECT 252.320 47.280 252.600 47.560 ;
        RECT 252.780 45.920 253.060 46.200 ;
        RECT 256.460 52.040 256.740 52.320 ;
        RECT 261.520 53.400 261.800 53.680 ;
        RECT 262.900 53.400 263.180 53.680 ;
        RECT 262.900 50.000 263.180 50.280 ;
        RECT 262.440 47.960 262.720 48.240 ;
        RECT 257.840 41.840 258.120 42.120 ;
        RECT 266.120 52.720 266.400 53.000 ;
        RECT 266.580 47.280 266.860 47.560 ;
        RECT 270.260 52.720 270.540 53.000 ;
        RECT 270.720 50.000 271.000 50.280 ;
        RECT 268.420 47.960 268.700 48.240 ;
        RECT 267.960 47.280 268.240 47.560 ;
        RECT 276.240 53.400 276.520 53.680 ;
        RECT 275.320 52.720 275.600 53.000 ;
        RECT 275.780 47.960 276.060 48.240 ;
        RECT 282.680 52.720 282.960 53.000 ;
        RECT 285.440 51.360 285.720 51.640 ;
        RECT 284.060 46.600 284.340 46.880 ;
        RECT 286.360 50.680 286.640 50.960 ;
        RECT 288.450 51.020 288.730 51.300 ;
        RECT 288.850 51.020 289.130 51.300 ;
        RECT 289.250 51.020 289.530 51.300 ;
        RECT 289.650 51.020 289.930 51.300 ;
        RECT 289.120 47.960 289.400 48.240 ;
        RECT 290.500 50.680 290.780 50.960 ;
        RECT 292.340 52.720 292.620 53.000 ;
        RECT 290.040 47.280 290.320 47.560 ;
        RECT 288.450 45.580 288.730 45.860 ;
        RECT 288.850 45.580 289.130 45.860 ;
        RECT 289.250 45.580 289.530 45.860 ;
        RECT 289.650 45.580 289.930 45.860 ;
        RECT 288.660 44.560 288.940 44.840 ;
        RECT 290.960 47.280 291.240 47.560 ;
        RECT 292.800 45.920 293.080 46.200 ;
        RECT 292.800 44.560 293.080 44.840 ;
        RECT 296.020 45.920 296.300 46.200 ;
        RECT 295.100 44.560 295.380 44.840 ;
        RECT 298.320 53.400 298.600 53.680 ;
        RECT 298.320 52.040 298.600 52.320 ;
        RECT 303.380 52.720 303.660 53.000 ;
        RECT 306.600 48.640 306.880 48.920 ;
        RECT 306.140 45.240 306.420 45.520 ;
        RECT 310.280 51.360 310.560 51.640 ;
        RECT 311.660 50.680 311.940 50.960 ;
        RECT 317.180 53.400 317.460 53.680 ;
        RECT 314.420 45.240 314.700 45.520 ;
        RECT 318.560 46.600 318.840 46.880 ;
        RECT 321.320 50.000 321.600 50.280 ;
        RECT 326.380 52.720 326.660 53.000 ;
        RECT 325.460 44.560 325.740 44.840 ;
        RECT 327.760 52.720 328.040 53.000 ;
        RECT 327.760 48.640 328.040 48.920 ;
        RECT 331.440 52.720 331.720 53.000 ;
        RECT 331.900 52.040 332.180 52.320 ;
        RECT 331.900 44.560 332.180 44.840 ;
        RECT 334.200 45.920 334.480 46.200 ;
        RECT 337.880 50.000 338.160 50.280 ;
        RECT 337.880 47.960 338.160 48.240 ;
        RECT 339.720 48.640 340.000 48.920 ;
        RECT 340.640 45.920 340.920 46.200 ;
        RECT 341.560 52.040 341.840 52.320 ;
        RECT 342.940 52.040 343.220 52.320 ;
        RECT 343.860 48.640 344.140 48.920 ;
        RECT 348.460 45.920 348.740 46.200 ;
        RECT 353.520 45.240 353.800 45.520 ;
        RECT 358.580 44.560 358.860 44.840 ;
        RECT 362.260 48.640 362.540 48.920 ;
        RECT 365.250 53.740 365.530 54.010 ;
        RECT 365.650 53.740 365.930 54.010 ;
        RECT 366.050 53.740 366.330 54.010 ;
        RECT 366.450 53.740 366.730 54.010 ;
        RECT 365.250 48.300 365.530 48.580 ;
        RECT 365.650 48.300 365.930 48.580 ;
        RECT 366.050 48.300 366.330 48.580 ;
        RECT 366.450 48.300 366.730 48.580 ;
        RECT 365.250 42.860 365.530 43.140 ;
        RECT 365.650 42.860 365.930 43.140 ;
        RECT 366.050 42.860 366.330 43.140 ;
        RECT 366.450 42.860 366.730 43.140 ;
        RECT 376.520 52.040 376.800 52.320 ;
        RECT 518.850 53.740 519.130 54.010 ;
        RECT 519.250 53.740 519.530 54.010 ;
        RECT 519.650 53.740 519.930 54.010 ;
        RECT 520.050 53.740 520.330 54.010 ;
        RECT 442.050 51.020 442.330 51.300 ;
        RECT 442.450 51.020 442.730 51.300 ;
        RECT 442.850 51.020 443.130 51.300 ;
        RECT 443.250 51.020 443.530 51.300 ;
        RECT 595.650 51.020 595.930 51.300 ;
        RECT 596.050 51.020 596.330 51.300 ;
        RECT 596.450 51.020 596.730 51.300 ;
        RECT 596.850 51.020 597.130 51.300 ;
        RECT 408.260 50.000 408.540 50.280 ;
        RECT 405.960 47.280 406.240 47.560 ;
        RECT 442.050 45.580 442.330 45.860 ;
        RECT 442.450 45.580 442.730 45.860 ;
        RECT 442.850 45.580 443.130 45.860 ;
        RECT 443.250 45.580 443.530 45.860 ;
        RECT 518.850 48.300 519.130 48.580 ;
        RECT 519.250 48.300 519.530 48.580 ;
        RECT 519.650 48.300 519.930 48.580 ;
        RECT 520.050 48.300 520.330 48.580 ;
        RECT 518.850 42.860 519.130 43.140 ;
        RECT 519.250 42.860 519.530 43.140 ;
        RECT 519.650 42.860 519.930 43.140 ;
        RECT 520.050 42.860 520.330 43.140 ;
        RECT 595.650 45.580 595.930 45.860 ;
        RECT 596.050 45.580 596.330 45.860 ;
        RECT 596.450 45.580 596.730 45.860 ;
        RECT 596.850 45.580 597.130 45.860 ;
      LAYER met3 ;
        RECT 54.000 54.000 597.190 619.805 ;
        RECT 57.990 53.715 59.590 54.000 ;
        RECT 211.590 53.715 213.190 54.000 ;
        RECT 365.190 53.715 366.790 54.000 ;
        RECT 518.790 53.715 520.390 54.000 ;
        RECT 99.115 53.690 99.445 53.705 ;
        RECT 103.255 53.690 103.585 53.705 ;
        RECT 145.575 53.690 145.905 53.705 ;
        RECT 99.115 53.390 103.585 53.690 ;
        RECT 99.115 53.375 99.445 53.390 ;
        RECT 103.255 53.375 103.585 53.390 ;
        RECT 104.420 53.390 145.905 53.690 ;
        RECT 103.255 53.010 103.585 53.025 ;
        RECT 104.420 53.010 104.720 53.390 ;
        RECT 145.575 53.375 145.905 53.390 ;
        RECT 237.780 53.690 238.160 53.700 ;
        RECT 261.495 53.690 261.825 53.705 ;
        RECT 237.780 53.390 261.825 53.690 ;
        RECT 237.780 53.380 238.160 53.390 ;
        RECT 261.495 53.375 261.825 53.390 ;
        RECT 262.875 53.690 263.205 53.705 ;
        RECT 276.215 53.690 276.545 53.705 ;
        RECT 262.875 53.390 276.545 53.690 ;
        RECT 262.875 53.375 263.205 53.390 ;
        RECT 276.215 53.375 276.545 53.390 ;
        RECT 298.295 53.690 298.625 53.705 ;
        RECT 317.155 53.690 317.485 53.705 ;
        RECT 298.295 53.390 317.485 53.690 ;
        RECT 298.295 53.375 298.625 53.390 ;
        RECT 317.155 53.375 317.485 53.390 ;
        RECT 103.255 52.710 104.720 53.010 ;
        RECT 127.635 53.010 127.965 53.025 ;
        RECT 158.915 53.010 159.245 53.025 ;
        RECT 127.635 52.710 159.245 53.010 ;
        RECT 103.255 52.695 103.585 52.710 ;
        RECT 127.635 52.695 127.965 52.710 ;
        RECT 158.915 52.695 159.245 52.710 ;
        RECT 170.415 53.010 170.745 53.025 ;
        RECT 177.775 53.010 178.105 53.025 ;
        RECT 214.115 53.020 214.445 53.025 ;
        RECT 170.415 52.710 178.105 53.010 ;
        RECT 170.415 52.695 170.745 52.710 ;
        RECT 177.775 52.695 178.105 52.710 ;
        RECT 213.860 53.010 214.445 53.020 ;
        RECT 225.155 53.010 225.485 53.025 ;
        RECT 228.835 53.010 229.165 53.025 ;
        RECT 213.860 52.710 214.670 53.010 ;
        RECT 225.155 52.710 229.165 53.010 ;
        RECT 213.860 52.700 214.445 52.710 ;
        RECT 214.115 52.695 214.445 52.700 ;
        RECT 225.155 52.695 225.485 52.710 ;
        RECT 228.835 52.695 229.165 52.710 ;
        RECT 243.095 53.010 243.425 53.025 ;
        RECT 251.835 53.010 252.165 53.025 ;
        RECT 243.095 52.710 252.165 53.010 ;
        RECT 243.095 52.695 243.425 52.710 ;
        RECT 251.835 52.695 252.165 52.710 ;
        RECT 254.135 53.010 254.465 53.025 ;
        RECT 266.095 53.010 266.425 53.025 ;
        RECT 254.135 52.710 266.425 53.010 ;
        RECT 254.135 52.695 254.465 52.710 ;
        RECT 266.095 52.695 266.425 52.710 ;
        RECT 270.235 53.010 270.565 53.025 ;
        RECT 275.295 53.010 275.625 53.025 ;
        RECT 270.235 52.710 275.625 53.010 ;
        RECT 270.235 52.695 270.565 52.710 ;
        RECT 275.295 52.695 275.625 52.710 ;
        RECT 282.655 53.010 282.985 53.025 ;
        RECT 292.315 53.010 292.645 53.025 ;
        RECT 282.655 52.710 292.645 53.010 ;
        RECT 282.655 52.695 282.985 52.710 ;
        RECT 292.315 52.695 292.645 52.710 ;
        RECT 303.355 53.010 303.685 53.025 ;
        RECT 326.355 53.010 326.685 53.025 ;
        RECT 303.355 52.710 326.685 53.010 ;
        RECT 303.355 52.695 303.685 52.710 ;
        RECT 326.355 52.695 326.685 52.710 ;
        RECT 327.735 53.010 328.065 53.025 ;
        RECT 331.415 53.010 331.745 53.025 ;
        RECT 327.735 52.710 331.745 53.010 ;
        RECT 327.735 52.695 328.065 52.710 ;
        RECT 331.415 52.695 331.745 52.710 ;
        RECT 110.615 52.330 110.945 52.345 ;
        RECT 146.495 52.330 146.825 52.345 ;
        RECT 150.635 52.330 150.965 52.345 ;
        RECT 110.615 52.030 137.840 52.330 ;
        RECT 110.615 52.015 110.945 52.030 ;
        RECT 109.695 51.650 110.025 51.665 ;
        RECT 114.295 51.650 114.625 51.665 ;
        RECT 109.695 51.350 114.625 51.650 ;
        RECT 109.695 51.335 110.025 51.350 ;
        RECT 114.295 51.335 114.625 51.350 ;
        RECT 125.795 51.650 126.125 51.665 ;
        RECT 132.235 51.650 132.565 51.665 ;
        RECT 125.795 51.350 132.565 51.650 ;
        RECT 137.540 51.650 137.840 52.030 ;
        RECT 146.495 52.030 150.965 52.330 ;
        RECT 146.495 52.015 146.825 52.030 ;
        RECT 150.635 52.015 150.965 52.030 ;
        RECT 157.995 52.330 158.325 52.345 ;
        RECT 185.135 52.330 185.465 52.345 ;
        RECT 190.655 52.330 190.985 52.345 ;
        RECT 157.995 52.030 190.985 52.330 ;
        RECT 157.995 52.015 158.325 52.030 ;
        RECT 185.135 52.015 185.465 52.030 ;
        RECT 190.655 52.015 190.985 52.030 ;
        RECT 194.795 52.330 195.125 52.345 ;
        RECT 196.175 52.330 196.505 52.345 ;
        RECT 201.235 52.330 201.565 52.345 ;
        RECT 194.795 52.030 201.565 52.330 ;
        RECT 194.795 52.015 195.125 52.030 ;
        RECT 196.175 52.015 196.505 52.030 ;
        RECT 201.235 52.015 201.565 52.030 ;
        RECT 208.595 52.330 208.925 52.345 ;
        RECT 235.020 52.330 235.400 52.340 ;
        RECT 208.595 52.030 235.400 52.330 ;
        RECT 208.595 52.015 208.925 52.030 ;
        RECT 235.020 52.020 235.400 52.030 ;
        RECT 236.195 52.330 236.525 52.345 ;
        RECT 238.035 52.330 238.365 52.345 ;
        RECT 236.195 52.030 238.365 52.330 ;
        RECT 236.195 52.015 236.525 52.030 ;
        RECT 238.035 52.015 238.365 52.030 ;
        RECT 256.435 52.330 256.765 52.345 ;
        RECT 298.295 52.330 298.625 52.345 ;
        RECT 331.875 52.330 332.205 52.345 ;
        RECT 341.535 52.330 341.865 52.345 ;
        RECT 256.435 52.030 291.480 52.330 ;
        RECT 256.435 52.015 256.765 52.030 ;
        RECT 152.475 51.650 152.805 51.665 ;
        RECT 137.540 51.350 152.805 51.650 ;
        RECT 125.795 51.335 126.125 51.350 ;
        RECT 132.235 51.335 132.565 51.350 ;
        RECT 152.475 51.335 152.805 51.350 ;
        RECT 154.775 51.650 155.105 51.665 ;
        RECT 188.815 51.650 189.145 51.665 ;
        RECT 189.735 51.650 190.065 51.665 ;
        RECT 154.775 51.350 190.065 51.650 ;
        RECT 154.775 51.335 155.105 51.350 ;
        RECT 188.815 51.335 189.145 51.350 ;
        RECT 189.735 51.335 190.065 51.350 ;
        RECT 199.395 51.650 199.725 51.665 ;
        RECT 203.995 51.650 204.325 51.665 ;
        RECT 199.395 51.350 204.325 51.650 ;
        RECT 199.395 51.335 199.725 51.350 ;
        RECT 203.995 51.335 204.325 51.350 ;
        RECT 212.275 51.650 212.605 51.665 ;
        RECT 215.955 51.650 216.285 51.665 ;
        RECT 212.275 51.350 216.285 51.650 ;
        RECT 212.275 51.335 212.605 51.350 ;
        RECT 215.955 51.335 216.285 51.350 ;
        RECT 238.035 51.650 238.365 51.665 ;
        RECT 285.415 51.650 285.745 51.665 ;
        RECT 238.035 51.350 285.745 51.650 ;
        RECT 291.180 51.650 291.480 52.030 ;
        RECT 298.295 52.030 341.865 52.330 ;
        RECT 298.295 52.015 298.625 52.030 ;
        RECT 331.875 52.015 332.205 52.030 ;
        RECT 341.535 52.015 341.865 52.030 ;
        RECT 342.915 52.330 343.245 52.345 ;
        RECT 376.495 52.330 376.825 52.345 ;
        RECT 342.915 52.030 376.825 52.330 ;
        RECT 342.915 52.015 343.245 52.030 ;
        RECT 376.495 52.015 376.825 52.030 ;
        RECT 310.255 51.650 310.585 51.665 ;
        RECT 291.180 51.350 310.585 51.650 ;
        RECT 238.035 51.335 238.365 51.350 ;
        RECT 285.415 51.335 285.745 51.350 ;
        RECT 310.255 51.335 310.585 51.350 ;
        RECT 134.790 50.995 136.390 51.325 ;
        RECT 288.390 50.995 289.990 51.325 ;
        RECT 441.990 50.995 443.590 51.325 ;
        RECT 595.590 50.995 597.190 51.325 ;
        RECT 77.035 50.970 77.365 50.985 ;
        RECT 108.775 50.970 109.105 50.985 ;
        RECT 162.135 50.970 162.465 50.985 ;
        RECT 210.435 50.980 210.765 50.985 ;
        RECT 77.035 50.670 109.105 50.970 ;
        RECT 77.035 50.655 77.365 50.670 ;
        RECT 108.775 50.655 109.105 50.670 ;
        RECT 137.540 50.670 162.465 50.970 ;
        RECT 72.435 50.290 72.765 50.305 ;
        RECT 93.595 50.290 93.925 50.305 ;
        RECT 96.815 50.290 97.145 50.305 ;
        RECT 72.435 49.990 97.145 50.290 ;
        RECT 72.435 49.975 72.765 49.990 ;
        RECT 93.595 49.975 93.925 49.990 ;
        RECT 96.815 49.975 97.145 49.990 ;
        RECT 114.755 50.290 115.085 50.305 ;
        RECT 137.540 50.290 137.840 50.670 ;
        RECT 162.135 50.655 162.465 50.670 ;
        RECT 210.180 50.970 210.765 50.980 ;
        RECT 214.115 50.970 214.445 50.985 ;
        RECT 249.995 50.970 250.325 50.985 ;
        RECT 210.180 50.670 210.990 50.970 ;
        RECT 214.115 50.670 250.325 50.970 ;
        RECT 210.180 50.660 210.765 50.670 ;
        RECT 210.435 50.655 210.765 50.660 ;
        RECT 214.115 50.655 214.445 50.670 ;
        RECT 249.995 50.655 250.325 50.670 ;
        RECT 250.915 50.970 251.245 50.985 ;
        RECT 286.335 50.970 286.665 50.985 ;
        RECT 250.915 50.670 286.665 50.970 ;
        RECT 250.915 50.655 251.245 50.670 ;
        RECT 286.335 50.655 286.665 50.670 ;
        RECT 290.475 50.970 290.805 50.985 ;
        RECT 311.635 50.970 311.965 50.985 ;
        RECT 290.475 50.670 311.965 50.970 ;
        RECT 290.475 50.655 290.805 50.670 ;
        RECT 311.635 50.655 311.965 50.670 ;
        RECT 159.375 50.290 159.705 50.305 ;
        RECT 114.755 49.990 137.840 50.290 ;
        RECT 138.460 49.990 159.705 50.290 ;
        RECT 114.755 49.975 115.085 49.990 ;
        RECT 69.215 49.610 69.545 49.625 ;
        RECT 78.875 49.610 79.205 49.625 ;
        RECT 69.215 49.310 79.205 49.610 ;
        RECT 69.215 49.295 69.545 49.310 ;
        RECT 78.875 49.295 79.205 49.310 ;
        RECT 84.395 49.610 84.725 49.625 ;
        RECT 114.295 49.610 114.625 49.625 ;
        RECT 138.460 49.610 138.760 49.990 ;
        RECT 159.375 49.975 159.705 49.990 ;
        RECT 164.895 50.290 165.225 50.305 ;
        RECT 230.675 50.290 231.005 50.305 ;
        RECT 164.895 49.990 231.005 50.290 ;
        RECT 164.895 49.975 165.225 49.990 ;
        RECT 230.675 49.975 231.005 49.990 ;
        RECT 241.255 50.290 241.585 50.305 ;
        RECT 262.875 50.290 263.205 50.305 ;
        RECT 241.255 49.990 263.205 50.290 ;
        RECT 241.255 49.975 241.585 49.990 ;
        RECT 262.875 49.975 263.205 49.990 ;
        RECT 270.695 50.290 271.025 50.305 ;
        RECT 321.295 50.290 321.625 50.305 ;
        RECT 270.695 49.990 321.625 50.290 ;
        RECT 270.695 49.975 271.025 49.990 ;
        RECT 321.295 49.975 321.625 49.990 ;
        RECT 337.855 50.290 338.185 50.305 ;
        RECT 408.235 50.290 408.565 50.305 ;
        RECT 337.855 49.990 408.565 50.290 ;
        RECT 337.855 49.975 338.185 49.990 ;
        RECT 408.235 49.975 408.565 49.990 ;
        RECT 84.395 49.310 113.920 49.610 ;
        RECT 84.395 49.295 84.725 49.310 ;
        RECT 81.175 48.930 81.505 48.945 ;
        RECT 109.695 48.930 110.025 48.945 ;
        RECT 81.175 48.630 110.025 48.930 ;
        RECT 113.620 48.930 113.920 49.310 ;
        RECT 114.295 49.310 138.760 49.610 ;
        RECT 156.615 49.610 156.945 49.625 ;
        RECT 176.395 49.610 176.725 49.625 ;
        RECT 156.615 49.310 176.725 49.610 ;
        RECT 114.295 49.295 114.625 49.310 ;
        RECT 156.615 49.295 156.945 49.310 ;
        RECT 176.395 49.295 176.725 49.310 ;
        RECT 195.255 49.610 195.585 49.625 ;
        RECT 214.575 49.610 214.905 49.625 ;
        RECT 195.255 49.310 214.905 49.610 ;
        RECT 195.255 49.295 195.585 49.310 ;
        RECT 214.575 49.295 214.905 49.310 ;
        RECT 225.615 49.610 225.945 49.625 ;
        RECT 243.095 49.610 243.425 49.625 ;
        RECT 225.615 49.310 243.425 49.610 ;
        RECT 225.615 49.295 225.945 49.310 ;
        RECT 243.095 49.295 243.425 49.310 ;
        RECT 116.135 48.930 116.465 48.945 ;
        RECT 119.355 48.930 119.685 48.945 ;
        RECT 113.620 48.630 119.685 48.930 ;
        RECT 81.175 48.615 81.505 48.630 ;
        RECT 109.695 48.615 110.025 48.630 ;
        RECT 116.135 48.615 116.465 48.630 ;
        RECT 119.355 48.615 119.685 48.630 ;
        RECT 136.375 48.930 136.705 48.945 ;
        RECT 151.095 48.930 151.425 48.945 ;
        RECT 201.695 48.930 202.025 48.945 ;
        RECT 136.375 48.630 147.960 48.930 ;
        RECT 136.375 48.615 136.705 48.630 ;
        RECT 57.990 48.275 59.590 48.605 ;
        RECT 147.660 48.250 147.960 48.630 ;
        RECT 151.095 48.630 202.025 48.930 ;
        RECT 151.095 48.615 151.425 48.630 ;
        RECT 201.695 48.615 202.025 48.630 ;
        RECT 252.295 48.930 252.625 48.945 ;
        RECT 306.575 48.930 306.905 48.945 ;
        RECT 252.295 48.630 306.905 48.930 ;
        RECT 252.295 48.615 252.625 48.630 ;
        RECT 306.575 48.615 306.905 48.630 ;
        RECT 327.735 48.930 328.065 48.945 ;
        RECT 339.695 48.930 340.025 48.945 ;
        RECT 327.735 48.630 340.025 48.930 ;
        RECT 327.735 48.615 328.065 48.630 ;
        RECT 339.695 48.615 340.025 48.630 ;
        RECT 343.835 48.930 344.165 48.945 ;
        RECT 362.235 48.930 362.565 48.945 ;
        RECT 343.835 48.630 362.565 48.930 ;
        RECT 343.835 48.615 344.165 48.630 ;
        RECT 362.235 48.615 362.565 48.630 ;
        RECT 211.590 48.275 213.190 48.605 ;
        RECT 365.190 48.275 366.790 48.605 ;
        RECT 518.790 48.275 520.390 48.605 ;
        RECT 181.660 48.250 182.040 48.260 ;
        RECT 188.815 48.250 189.145 48.265 ;
        RECT 147.660 47.950 189.145 48.250 ;
        RECT 181.660 47.940 182.040 47.950 ;
        RECT 188.815 47.935 189.145 47.950 ;
        RECT 231.135 48.260 231.465 48.265 ;
        RECT 231.135 48.250 231.720 48.260 ;
        RECT 233.180 48.250 233.560 48.260 ;
        RECT 234.815 48.250 235.145 48.265 ;
        RECT 231.135 47.950 231.920 48.250 ;
        RECT 233.180 47.950 235.145 48.250 ;
        RECT 231.135 47.940 231.720 47.950 ;
        RECT 233.180 47.940 233.560 47.950 ;
        RECT 231.135 47.935 231.465 47.940 ;
        RECT 234.815 47.935 235.145 47.950 ;
        RECT 244.475 48.250 244.805 48.265 ;
        RECT 262.415 48.250 262.745 48.265 ;
        RECT 244.475 47.950 262.745 48.250 ;
        RECT 244.475 47.935 244.805 47.950 ;
        RECT 262.415 47.935 262.745 47.950 ;
        RECT 268.395 48.250 268.725 48.265 ;
        RECT 275.755 48.250 276.085 48.265 ;
        RECT 268.395 47.950 276.085 48.250 ;
        RECT 268.395 47.935 268.725 47.950 ;
        RECT 275.755 47.935 276.085 47.950 ;
        RECT 289.095 48.250 289.425 48.265 ;
        RECT 337.855 48.250 338.185 48.265 ;
        RECT 289.095 47.950 338.185 48.250 ;
        RECT 289.095 47.935 289.425 47.950 ;
        RECT 337.855 47.935 338.185 47.950 ;
        RECT 98.195 47.570 98.525 47.585 ;
        RECT 130.855 47.570 131.185 47.585 ;
        RECT 98.195 47.270 131.185 47.570 ;
        RECT 98.195 47.255 98.525 47.270 ;
        RECT 130.855 47.255 131.185 47.270 ;
        RECT 140.055 47.570 140.385 47.585 ;
        RECT 157.995 47.570 158.325 47.585 ;
        RECT 140.055 47.270 158.325 47.570 ;
        RECT 140.055 47.255 140.385 47.270 ;
        RECT 157.995 47.255 158.325 47.270 ;
        RECT 158.915 47.570 159.245 47.585 ;
        RECT 220.095 47.570 220.425 47.585 ;
        RECT 158.915 47.270 220.425 47.570 ;
        RECT 158.915 47.255 159.245 47.270 ;
        RECT 220.095 47.255 220.425 47.270 ;
        RECT 240.335 47.570 240.665 47.585 ;
        RECT 243.555 47.570 243.885 47.585 ;
        RECT 240.335 47.270 243.885 47.570 ;
        RECT 240.335 47.255 240.665 47.270 ;
        RECT 243.555 47.255 243.885 47.270 ;
        RECT 252.295 47.570 252.625 47.585 ;
        RECT 266.555 47.570 266.885 47.585 ;
        RECT 252.295 47.270 266.885 47.570 ;
        RECT 252.295 47.255 252.625 47.270 ;
        RECT 266.555 47.255 266.885 47.270 ;
        RECT 267.935 47.570 268.265 47.585 ;
        RECT 290.015 47.570 290.345 47.585 ;
        RECT 267.935 47.270 290.345 47.570 ;
        RECT 267.935 47.255 268.265 47.270 ;
        RECT 290.015 47.255 290.345 47.270 ;
        RECT 290.935 47.570 291.265 47.585 ;
        RECT 405.935 47.570 406.265 47.585 ;
        RECT 290.935 47.270 406.265 47.570 ;
        RECT 290.935 47.255 291.265 47.270 ;
        RECT 405.935 47.255 406.265 47.270 ;
        RECT 38.395 46.890 38.725 46.905 ;
        RECT 284.035 46.890 284.365 46.905 ;
        RECT 318.535 46.890 318.865 46.905 ;
        RECT 38.395 46.590 284.365 46.890 ;
        RECT 38.395 46.575 38.725 46.590 ;
        RECT 284.035 46.575 284.365 46.590 ;
        RECT 284.740 46.590 318.865 46.890 ;
        RECT 194.795 46.210 195.125 46.225 ;
        RECT 199.395 46.210 199.725 46.225 ;
        RECT 194.795 45.910 199.725 46.210 ;
        RECT 194.795 45.895 195.125 45.910 ;
        RECT 199.395 45.895 199.725 45.910 ;
        RECT 252.755 46.210 253.085 46.225 ;
        RECT 284.740 46.210 285.040 46.590 ;
        RECT 318.535 46.575 318.865 46.590 ;
        RECT 252.755 45.910 285.040 46.210 ;
        RECT 292.775 46.210 293.105 46.225 ;
        RECT 295.995 46.210 296.325 46.225 ;
        RECT 334.175 46.210 334.505 46.225 ;
        RECT 292.775 45.910 334.505 46.210 ;
        RECT 252.755 45.895 253.085 45.910 ;
        RECT 292.775 45.895 293.105 45.910 ;
        RECT 295.995 45.895 296.325 45.910 ;
        RECT 334.175 45.895 334.505 45.910 ;
        RECT 340.615 46.210 340.945 46.225 ;
        RECT 348.435 46.210 348.765 46.225 ;
        RECT 340.615 45.910 348.765 46.210 ;
        RECT 340.615 45.895 340.945 45.910 ;
        RECT 348.435 45.895 348.765 45.910 ;
        RECT 134.790 45.555 136.390 45.885 ;
        RECT 288.390 45.555 289.990 45.885 ;
        RECT 441.990 45.555 443.590 45.885 ;
        RECT 595.590 45.555 597.190 45.885 ;
        RECT 193.875 45.530 194.205 45.545 ;
        RECT 228.375 45.530 228.705 45.545 ;
        RECT 193.875 45.230 228.705 45.530 ;
        RECT 193.875 45.215 194.205 45.230 ;
        RECT 228.375 45.215 228.705 45.230 ;
        RECT 306.115 45.530 306.445 45.545 ;
        RECT 314.395 45.530 314.725 45.545 ;
        RECT 353.495 45.530 353.825 45.545 ;
        RECT 306.115 45.230 353.825 45.530 ;
        RECT 306.115 45.215 306.445 45.230 ;
        RECT 314.395 45.215 314.725 45.230 ;
        RECT 353.495 45.215 353.825 45.230 ;
        RECT 90.835 44.850 91.165 44.865 ;
        RECT 127.635 44.850 127.965 44.865 ;
        RECT 90.835 44.550 127.965 44.850 ;
        RECT 90.835 44.535 91.165 44.550 ;
        RECT 127.635 44.535 127.965 44.550 ;
        RECT 185.135 44.850 185.465 44.865 ;
        RECT 229.755 44.850 230.085 44.865 ;
        RECT 185.135 44.550 230.085 44.850 ;
        RECT 185.135 44.535 185.465 44.550 ;
        RECT 229.755 44.535 230.085 44.550 ;
        RECT 288.635 44.850 288.965 44.865 ;
        RECT 292.775 44.850 293.105 44.865 ;
        RECT 288.635 44.550 293.105 44.850 ;
        RECT 288.635 44.535 288.965 44.550 ;
        RECT 292.775 44.535 293.105 44.550 ;
        RECT 295.075 44.850 295.405 44.865 ;
        RECT 325.435 44.850 325.765 44.865 ;
        RECT 295.075 44.550 325.765 44.850 ;
        RECT 295.075 44.535 295.405 44.550 ;
        RECT 325.435 44.535 325.765 44.550 ;
        RECT 331.875 44.850 332.205 44.865 ;
        RECT 358.555 44.850 358.885 44.865 ;
        RECT 331.875 44.550 358.885 44.850 ;
        RECT 331.875 44.535 332.205 44.550 ;
        RECT 358.555 44.535 358.885 44.550 ;
        RECT 119.355 44.170 119.685 44.185 ;
        RECT 129.015 44.170 129.345 44.185 ;
        RECT 119.355 43.870 129.345 44.170 ;
        RECT 119.355 43.855 119.685 43.870 ;
        RECT 129.015 43.855 129.345 43.870 ;
        RECT 57.990 42.835 59.590 43.165 ;
        RECT 211.590 42.835 213.190 43.165 ;
        RECT 365.190 42.835 366.790 43.165 ;
        RECT 518.790 42.835 520.390 43.165 ;
        RECT 223.775 42.130 224.105 42.145 ;
        RECT 257.815 42.130 258.145 42.145 ;
        RECT 223.775 41.830 258.145 42.130 ;
        RECT 223.775 41.815 224.105 41.830 ;
        RECT 257.815 41.815 258.145 41.830 ;
      LAYER via3 ;
        RECT 58.030 53.720 58.350 54.020 ;
        RECT 58.430 53.720 58.750 54.020 ;
        RECT 58.830 53.720 59.150 54.020 ;
        RECT 59.230 53.720 59.550 54.020 ;
        RECT 211.630 53.720 211.950 54.020 ;
        RECT 212.030 53.720 212.350 54.020 ;
        RECT 212.430 53.720 212.750 54.020 ;
        RECT 212.830 53.720 213.150 54.020 ;
        RECT 365.230 53.720 365.550 54.020 ;
        RECT 365.630 53.720 365.950 54.020 ;
        RECT 366.030 53.720 366.350 54.020 ;
        RECT 366.430 53.720 366.750 54.020 ;
        RECT 518.830 53.720 519.150 54.020 ;
        RECT 519.230 53.720 519.550 54.020 ;
        RECT 519.630 53.720 519.950 54.020 ;
        RECT 520.030 53.720 520.350 54.020 ;
        RECT 237.810 53.380 238.130 53.700 ;
        RECT 213.890 52.700 214.210 53.020 ;
        RECT 235.050 52.020 235.370 52.340 ;
        RECT 134.830 51.000 135.150 51.320 ;
        RECT 135.230 51.000 135.550 51.320 ;
        RECT 135.630 51.000 135.950 51.320 ;
        RECT 136.030 51.000 136.350 51.320 ;
        RECT 288.430 51.000 288.750 51.320 ;
        RECT 288.830 51.000 289.150 51.320 ;
        RECT 289.230 51.000 289.550 51.320 ;
        RECT 289.630 51.000 289.950 51.320 ;
        RECT 442.030 51.000 442.350 51.320 ;
        RECT 442.430 51.000 442.750 51.320 ;
        RECT 442.830 51.000 443.150 51.320 ;
        RECT 443.230 51.000 443.550 51.320 ;
        RECT 595.630 51.000 595.950 51.320 ;
        RECT 596.030 51.000 596.350 51.320 ;
        RECT 596.430 51.000 596.750 51.320 ;
        RECT 596.830 51.000 597.150 51.320 ;
        RECT 210.210 50.660 210.530 50.980 ;
        RECT 58.030 48.280 58.350 48.600 ;
        RECT 58.430 48.280 58.750 48.600 ;
        RECT 58.830 48.280 59.150 48.600 ;
        RECT 59.230 48.280 59.550 48.600 ;
        RECT 211.630 48.280 211.950 48.600 ;
        RECT 212.030 48.280 212.350 48.600 ;
        RECT 212.430 48.280 212.750 48.600 ;
        RECT 212.830 48.280 213.150 48.600 ;
        RECT 365.230 48.280 365.550 48.600 ;
        RECT 365.630 48.280 365.950 48.600 ;
        RECT 366.030 48.280 366.350 48.600 ;
        RECT 366.430 48.280 366.750 48.600 ;
        RECT 518.830 48.280 519.150 48.600 ;
        RECT 519.230 48.280 519.550 48.600 ;
        RECT 519.630 48.280 519.950 48.600 ;
        RECT 520.030 48.280 520.350 48.600 ;
        RECT 181.690 47.940 182.010 48.260 ;
        RECT 231.370 47.940 231.690 48.260 ;
        RECT 233.210 47.940 233.530 48.260 ;
        RECT 134.830 45.560 135.150 45.880 ;
        RECT 135.230 45.560 135.550 45.880 ;
        RECT 135.630 45.560 135.950 45.880 ;
        RECT 136.030 45.560 136.350 45.880 ;
        RECT 288.430 45.560 288.750 45.880 ;
        RECT 288.830 45.560 289.150 45.880 ;
        RECT 289.230 45.560 289.550 45.880 ;
        RECT 289.630 45.560 289.950 45.880 ;
        RECT 442.030 45.560 442.350 45.880 ;
        RECT 442.430 45.560 442.750 45.880 ;
        RECT 442.830 45.560 443.150 45.880 ;
        RECT 443.230 45.560 443.550 45.880 ;
        RECT 595.630 45.560 595.950 45.880 ;
        RECT 596.030 45.560 596.350 45.880 ;
        RECT 596.430 45.560 596.750 45.880 ;
        RECT 596.830 45.560 597.150 45.880 ;
        RECT 58.030 42.840 58.350 43.160 ;
        RECT 58.430 42.840 58.750 43.160 ;
        RECT 58.830 42.840 59.150 43.160 ;
        RECT 59.230 42.840 59.550 43.160 ;
        RECT 211.630 42.840 211.950 43.160 ;
        RECT 212.030 42.840 212.350 43.160 ;
        RECT 212.430 42.840 212.750 43.160 ;
        RECT 212.830 42.840 213.150 43.160 ;
        RECT 365.230 42.840 365.550 43.160 ;
        RECT 365.630 42.840 365.950 43.160 ;
        RECT 366.030 42.840 366.350 43.160 ;
        RECT 366.430 42.840 366.750 43.160 ;
        RECT 518.830 42.840 519.150 43.160 ;
        RECT 519.230 42.840 519.550 43.160 ;
        RECT 519.630 42.840 519.950 43.160 ;
        RECT 520.030 42.840 520.350 43.160 ;
      LAYER met4 ;
        RECT 57.990 54.000 597.190 619.880 ;
        RECT 57.990 42.760 59.590 54.000 ;
        RECT 134.790 42.760 136.390 54.000 ;
        RECT 181.700 48.265 182.000 54.000 ;
        RECT 210.220 50.985 210.520 54.000 ;
        RECT 210.205 50.655 210.535 50.985 ;
        RECT 181.685 47.935 182.015 48.265 ;
        RECT 211.590 42.760 213.190 54.000 ;
        RECT 213.900 53.025 214.200 54.000 ;
        RECT 213.885 52.695 214.215 53.025 ;
        RECT 231.380 48.265 231.680 54.000 ;
        RECT 233.220 48.265 233.520 54.000 ;
        RECT 235.060 52.345 235.360 54.000 ;
        RECT 237.820 53.705 238.120 54.000 ;
        RECT 237.805 53.375 238.135 53.705 ;
        RECT 235.045 52.015 235.375 52.345 ;
        RECT 231.365 47.935 231.695 48.265 ;
        RECT 233.205 47.935 233.535 48.265 ;
        RECT 288.390 42.760 289.990 54.000 ;
        RECT 365.190 42.760 366.790 54.000 ;
        RECT 441.990 42.760 443.590 54.000 ;
        RECT 518.790 42.760 520.390 54.000 ;
        RECT 595.590 42.760 597.190 54.000 ;
  END
END user_project_wrapper
END LIBRARY

