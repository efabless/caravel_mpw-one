magic
tech sky130A
magscale 12 1
timestamp 1598787509
<< metal5 >>
rect 30 85 45 90
rect 25 80 45 85
rect 20 75 45 80
rect 15 70 40 75
rect 10 65 35 70
rect 5 60 30 65
rect 0 45 25 60
rect 5 40 30 45
rect 10 35 35 40
rect 15 30 40 35
rect 20 25 45 30
rect 25 20 45 25
rect 30 15 45 20
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
