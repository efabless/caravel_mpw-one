magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1288 -1260 1388 1527
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_0
timestamp 1623348570
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_1
timestamp 1623348570
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 5765212
string GDS_START 5764162
<< end >>
