VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io_alt
  CLASS BLOCK ;
  FOREIGN chip_io_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.900 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.900 95.440 ;
    END
  END flash_clk
  PIN flash_clk_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_clk_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.215 208.565 1787.495 210.965 ;
    END
  END flash_clk_ieb_core
  PIN flash_clk_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.475 208.565 1824.755 210.965 ;
    END
  END flash_clk_oeb_core
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.900 95.440 ;
    END
  END flash_csb
  PIN flash_csb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_csb_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.215 208.565 1513.495 210.965 ;
    END
  END flash_csb_ieb_core
  PIN flash_csb_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.475 208.565 1550.755 210.965 ;
    END
  END flash_csb_oeb_core
  PIN flash_io0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.900 95.440 ;
    END
  END flash_io0
  PIN flash_io0_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2046.610 209.000 2046.930 209.060 ;
        RECT 2061.790 209.000 2062.110 209.060 ;
        RECT 2076.050 209.000 2076.370 209.060 ;
        RECT 2046.610 208.860 2076.370 209.000 ;
        RECT 2046.610 208.800 2046.930 208.860 ;
        RECT 2061.790 208.800 2062.110 208.860 ;
        RECT 2076.050 208.800 2076.370 208.860 ;
      LAYER via ;
        RECT 2046.640 208.800 2046.900 209.060 ;
        RECT 2061.820 208.800 2062.080 209.060 ;
        RECT 2076.080 208.800 2076.340 209.060 ;
      LAYER met2 ;
        RECT 2046.035 209.170 2046.315 210.965 ;
        RECT 2061.215 209.170 2061.495 210.965 ;
        RECT 2076.855 209.170 2077.135 210.965 ;
        RECT 2046.035 209.090 2046.840 209.170 ;
        RECT 2061.215 209.090 2062.020 209.170 ;
        RECT 2076.140 209.090 2077.135 209.170 ;
        RECT 2046.035 209.030 2046.900 209.090 ;
        RECT 2046.035 208.565 2046.315 209.030 ;
        RECT 2046.640 208.770 2046.900 209.030 ;
        RECT 2061.215 209.030 2062.080 209.090 ;
        RECT 2061.215 208.565 2061.495 209.030 ;
        RECT 2061.820 208.770 2062.080 209.030 ;
        RECT 2076.080 209.030 2077.135 209.090 ;
        RECT 2076.080 208.770 2076.340 209.030 ;
        RECT 2076.855 208.565 2077.135 209.030 ;
    END
  END flash_io0_ieb_core
  PIN flash_io0_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.370 221.835 2055.650 222.205 ;
        RECT 2055.440 210.965 2055.580 221.835 ;
        RECT 2098.610 221.155 2098.890 221.525 ;
        RECT 2098.680 210.965 2098.820 221.155 ;
        RECT 2055.235 209.100 2055.580 210.965 ;
        RECT 2098.475 209.100 2098.820 210.965 ;
        RECT 2055.235 208.565 2055.515 209.100 ;
        RECT 2098.475 208.565 2098.755 209.100 ;
      LAYER via2 ;
        RECT 2055.370 221.880 2055.650 222.160 ;
        RECT 2098.610 221.200 2098.890 221.480 ;
      LAYER met3 ;
        RECT 2055.345 222.170 2055.675 222.185 ;
        RECT 2055.345 221.870 2097.750 222.170 ;
        RECT 2055.345 221.855 2055.675 221.870 ;
        RECT 2097.450 221.490 2097.750 221.870 ;
        RECT 2098.585 221.490 2098.915 221.505 ;
        RECT 2097.450 221.190 2098.915 221.490 ;
        RECT 2098.585 221.175 2098.915 221.190 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.900 95.440 ;
    END
  END flash_io1
  PIN flash_io1_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2320.770 209.000 2321.090 209.060 ;
        RECT 2335.950 209.000 2336.270 209.060 ;
        RECT 2350.210 209.000 2350.530 209.060 ;
        RECT 2320.770 208.860 2350.530 209.000 ;
        RECT 2320.770 208.800 2321.090 208.860 ;
        RECT 2335.950 208.800 2336.270 208.860 ;
        RECT 2350.210 208.800 2350.530 208.860 ;
      LAYER via ;
        RECT 2320.800 208.800 2321.060 209.060 ;
        RECT 2335.980 208.800 2336.240 209.060 ;
        RECT 2350.240 208.800 2350.500 209.060 ;
      LAYER met2 ;
        RECT 2320.035 209.170 2320.315 210.965 ;
        RECT 2335.215 209.170 2335.495 210.965 ;
        RECT 2350.855 209.170 2351.135 210.965 ;
        RECT 2320.035 209.090 2321.000 209.170 ;
        RECT 2335.215 209.090 2336.180 209.170 ;
        RECT 2350.300 209.090 2351.135 209.170 ;
        RECT 2320.035 209.030 2321.060 209.090 ;
        RECT 2320.035 208.565 2320.315 209.030 ;
        RECT 2320.800 208.770 2321.060 209.030 ;
        RECT 2335.215 209.030 2336.240 209.090 ;
        RECT 2335.215 208.565 2335.495 209.030 ;
        RECT 2335.980 208.770 2336.240 209.030 ;
        RECT 2350.240 209.030 2351.135 209.090 ;
        RECT 2350.240 208.770 2350.500 209.030 ;
        RECT 2350.855 208.565 2351.135 209.030 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.070 221.835 2329.350 222.205 ;
        RECT 2372.310 221.835 2372.590 222.205 ;
        RECT 2329.140 210.965 2329.280 221.835 ;
        RECT 2372.380 210.965 2372.520 221.835 ;
        RECT 2329.140 209.030 2329.515 210.965 ;
        RECT 2372.380 209.030 2372.755 210.965 ;
        RECT 2329.235 208.565 2329.515 209.030 ;
        RECT 2372.475 208.565 2372.755 209.030 ;
      LAYER via2 ;
        RECT 2329.070 221.880 2329.350 222.160 ;
        RECT 2372.310 221.880 2372.590 222.160 ;
      LAYER met3 ;
        RECT 2329.045 222.170 2329.375 222.185 ;
        RECT 2372.285 222.170 2372.615 222.185 ;
        RECT 2329.045 221.870 2372.615 222.170 ;
        RECT 2329.045 221.855 2329.375 221.870 ;
        RECT 2372.285 221.855 2372.615 221.870 ;
    END
  END flash_io1_oeb_core
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.900 95.440 ;
    END
  END gpio
  PIN gpio_in_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 221.155 2594.310 221.525 ;
        RECT 2624.850 221.155 2625.130 221.525 ;
        RECT 2594.100 210.965 2594.240 221.155 ;
        RECT 2624.920 210.965 2625.060 221.155 ;
        RECT 2594.035 208.565 2594.315 210.965 ;
        RECT 2624.855 208.565 2625.135 210.965 ;
      LAYER via2 ;
        RECT 2594.030 221.200 2594.310 221.480 ;
        RECT 2624.850 221.200 2625.130 221.480 ;
      LAYER met3 ;
        RECT 2594.005 221.490 2594.335 221.505 ;
        RECT 2624.825 221.490 2625.155 221.505 ;
        RECT 2594.005 221.190 2625.155 221.490 ;
        RECT 2594.005 221.175 2594.335 221.190 ;
        RECT 2624.825 221.175 2625.155 221.190 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.475 208.565 2646.755 210.965 ;
    END
  END gpio_outenb_core
  PIN vccd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd_pad
  PIN vdda_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda_pad
  PIN vddio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio_pad
  PIN vddio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4361.050 94.880 4421.890 ;
    END
  END vddio_pad2
  PIN vssa_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa_pad
  PIN vssd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd_pad
  PIN vssio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
  END vssio_pad
  PIN vssio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1704.050 5093.120 1764.890 5153.945 ;
    END
  END vssio_pad2
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 498.200 3555.010 560.900 ;
    END
  END mprj_io[0]
  PIN mprj_io_analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 521.015 3379.435 521.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 527.455 3379.435 527.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 542.635 3379.435 542.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 524.235 3379.435 524.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 515.035 3379.435 515.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 545.855 3379.435 546.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 549.075 3379.435 549.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 564.255 3379.435 564.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 530.215 3379.435 530.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 567.475 3379.435 567.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 551.835 3379.435 552.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 505.835 3379.435 506.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 561.035 3379.435 561.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 496.635 3379.435 496.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in_3v3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 570.235 3379.435 570.515 ;
    END
  END mprj_io_in_3v3[0]
  PIN mprj_gpio_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3372.055 3379.435 3372.335 ;
    END
  END mprj_gpio_analog[3]
  PIN mprj_gpio_noesd[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3381.255 3379.435 3381.535 ;
    END
  END mprj_gpio_noesd[3]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3361.200 3555.010 3423.900 ;
    END
  END mprj_io[10]
  PIN mprj_io_analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3384.015 3379.435 3384.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3390.455 3379.435 3390.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3405.635 3379.435 3405.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3387.235 3379.435 3387.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3378.035 3379.435 3378.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3408.855 3379.435 3409.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3412.075 3379.435 3412.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3427.255 3379.435 3427.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3393.215 3379.435 3393.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3430.475 3379.435 3430.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3414.835 3379.435 3415.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3368.835 3379.435 3369.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3424.035 3379.435 3424.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3359.635 3379.435 3359.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in_3v3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.235 3379.435 3433.515 ;
    END
  END mprj_io_in_3v3[10]
  PIN mprj_gpio_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3593.055 3379.435 3593.335 ;
    END
  END mprj_gpio_analog[4]
  PIN mprj_gpio_noesd[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3602.255 3379.435 3602.535 ;
    END
  END mprj_gpio_noesd[4]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3582.200 3555.010 3644.900 ;
    END
  END mprj_io[11]
  PIN mprj_io_analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3605.015 3379.435 3605.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3611.455 3379.435 3611.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3626.635 3379.435 3626.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3608.235 3379.435 3608.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3599.035 3379.435 3599.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3629.855 3379.435 3630.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3633.075 3379.435 3633.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3648.255 3379.435 3648.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3614.215 3379.435 3614.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3651.475 3379.435 3651.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3635.835 3379.435 3636.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3589.835 3379.435 3590.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.035 3379.435 3645.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3580.635 3379.435 3580.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in_3v3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.235 3379.435 3654.515 ;
    END
  END mprj_io_in_3v3[11]
  PIN mprj_gpio_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3815.055 3379.435 3815.335 ;
    END
  END mprj_gpio_analog[5]
  PIN mprj_gpio_noesd[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3824.255 3379.435 3824.535 ;
    END
  END mprj_gpio_noesd[5]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3804.200 3555.010 3866.900 ;
    END
  END mprj_io[12]
  PIN mprj_io_analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3827.015 3379.435 3827.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3833.455 3379.435 3833.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3848.635 3379.435 3848.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3830.235 3379.435 3830.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3821.035 3379.435 3821.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3851.855 3379.435 3852.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3855.075 3379.435 3855.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.255 3379.435 3870.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3836.215 3379.435 3836.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3873.475 3379.435 3873.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3857.835 3379.435 3858.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3811.835 3379.435 3812.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3867.035 3379.435 3867.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3802.635 3379.435 3802.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in_3v3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3876.235 3379.435 3876.515 ;
    END
  END mprj_io_in_3v3[12]
  PIN mprj_gpio_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4252.055 3379.435 4252.335 ;
    END
  END mprj_gpio_analog[6]
  PIN mprj_gpio_noesd[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4261.255 3379.435 4261.535 ;
    END
  END mprj_gpio_noesd[6]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4241.200 3555.010 4303.900 ;
    END
  END mprj_io[13]
  PIN mprj_io_analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4264.015 3379.435 4264.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4270.455 3379.435 4270.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4285.635 3379.435 4285.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4267.235 3379.435 4267.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4258.035 3379.435 4258.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4288.855 3379.435 4289.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4292.075 3379.435 4292.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4307.255 3379.435 4307.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4273.215 3379.435 4273.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4310.475 3379.435 4310.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4294.835 3379.435 4295.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4248.835 3379.435 4249.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4304.035 3379.435 4304.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4239.635 3379.435 4239.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in_3v3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4313.235 3379.435 4313.515 ;
    END
  END mprj_io_in_3v3[13]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 720.200 3555.010 782.900 ;
    END
  END mprj_io[1]
  PIN mprj_io_analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 743.015 3379.435 743.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.455 3379.435 749.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.635 3379.435 764.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 746.235 3379.435 746.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 737.035 3379.435 737.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 767.855 3379.435 768.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 771.075 3379.435 771.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 786.255 3379.435 786.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 752.215 3379.435 752.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 789.475 3379.435 789.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 773.835 3379.435 774.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 727.835 3379.435 728.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.035 3379.435 783.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 718.635 3379.435 718.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in_3v3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 792.235 3379.435 792.515 ;
    END
  END mprj_io_in_3v3[1]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 941.200 3555.010 1003.900 ;
    END
  END mprj_io[2]
  PIN mprj_io_analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.015 3379.435 964.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 970.455 3379.435 970.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 985.635 3379.435 985.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 967.235 3379.435 967.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 958.035 3379.435 958.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 988.855 3379.435 989.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 992.075 3379.435 992.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1007.255 3379.435 1007.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 973.215 3379.435 973.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.475 3379.435 1010.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 994.835 3379.435 995.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 948.835 3379.435 949.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.035 3379.435 1004.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 939.635 3379.435 939.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in_3v3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1013.235 3379.435 1013.515 ;
    END
  END mprj_io_in_3v3[2]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1162.200 3555.010 1224.900 ;
    END
  END mprj_io[3]
  PIN mprj_io_analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1185.015 3379.435 1185.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1191.455 3379.435 1191.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.635 3379.435 1206.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1179.035 3379.435 1179.315 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.855 3379.435 1210.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1188.235 3379.435 1188.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1213.075 3379.435 1213.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1228.255 3379.435 1228.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1194.215 3379.435 1194.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1231.475 3379.435 1231.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.835 3379.435 1216.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1169.835 3379.435 1170.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1225.035 3379.435 1225.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1160.635 3379.435 1160.915 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in_3v3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.235 3379.435 1234.515 ;
    END
  END mprj_io_in_3v3[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1384.200 3555.010 1446.900 ;
    END
  END mprj_io[4]
  PIN mprj_io_analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1407.015 3379.435 1407.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1413.455 3379.435 1413.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1428.635 3379.435 1428.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1410.235 3379.435 1410.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1401.035 3379.435 1401.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.855 3379.435 1432.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1435.075 3379.435 1435.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1450.255 3379.435 1450.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1416.215 3379.435 1416.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1453.475 3379.435 1453.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.835 3379.435 1438.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1391.835 3379.435 1392.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1447.035 3379.435 1447.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1382.635 3379.435 1382.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in_3v3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1456.235 3379.435 1456.515 ;
    END
  END mprj_io_in_3v3[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1605.200 3555.010 1667.900 ;
    END
  END mprj_io[5]
  PIN mprj_io_analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1628.015 3379.435 1628.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1634.455 3379.435 1634.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1649.635 3379.435 1649.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.235 3379.435 1631.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1622.035 3379.435 1622.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1652.855 3379.435 1653.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.075 3379.435 1656.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1671.255 3379.435 1671.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1637.215 3379.435 1637.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1674.475 3379.435 1674.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1658.835 3379.435 1659.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1612.835 3379.435 1613.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1668.035 3379.435 1668.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1603.635 3379.435 1603.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in_3v3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.235 3379.435 1677.515 ;
    END
  END mprj_io_in_3v3[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1826.200 3555.010 1888.900 ;
    END
  END mprj_io[6]
  PIN mprj_io_analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1849.015 3379.435 1849.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1855.455 3379.435 1855.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1870.635 3379.435 1870.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1852.235 3379.435 1852.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1843.035 3379.435 1843.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1873.855 3379.435 1874.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1877.075 3379.435 1877.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1892.255 3379.435 1892.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1858.215 3379.435 1858.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1895.475 3379.435 1895.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1879.835 3379.435 1880.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1833.835 3379.435 1834.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1889.035 3379.435 1889.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1824.635 3379.435 1824.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in_3v3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1898.235 3379.435 1898.515 ;
    END
  END mprj_io_in_3v3[6]
  PIN mprj_gpio_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2708.055 3379.435 2708.335 ;
    END
  END mprj_gpio_analog[0]
  PIN mprj_gpio_noesd[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2717.255 3379.435 2717.535 ;
    END
  END mprj_gpio_noesd[0]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2697.200 3555.010 2759.900 ;
    END
  END mprj_io[7]
  PIN mprj_io_analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2720.015 3379.435 2720.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2726.455 3379.435 2726.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2741.635 3379.435 2741.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2723.235 3379.435 2723.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2714.035 3379.435 2714.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2744.855 3379.435 2745.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2748.075 3379.435 2748.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2763.255 3379.435 2763.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2729.215 3379.435 2729.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2766.475 3379.435 2766.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2750.835 3379.435 2751.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2704.835 3379.435 2705.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2760.035 3379.435 2760.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2695.635 3379.435 2695.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in_3v3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2769.235 3379.435 2769.515 ;
    END
  END mprj_io_in_3v3[7]
  PIN mprj_gpio_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2929.055 3379.435 2929.335 ;
    END
  END mprj_gpio_analog[1]
  PIN mprj_gpio_noesd[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2938.255 3379.435 2938.535 ;
    END
  END mprj_gpio_noesd[1]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2918.200 3555.010 2980.900 ;
    END
  END mprj_io[8]
  PIN mprj_io_analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2941.015 3379.435 2941.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2947.455 3379.435 2947.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2962.635 3379.435 2962.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2944.235 3379.435 2944.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2935.035 3379.435 2935.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2965.855 3379.435 2966.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.075 3379.435 2969.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2984.255 3379.435 2984.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2950.215 3379.435 2950.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2987.475 3379.435 2987.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2971.835 3379.435 2972.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2925.835 3379.435 2926.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2981.035 3379.435 2981.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2916.635 3379.435 2916.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in_3v3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2990.235 3379.435 2990.515 ;
    END
  END mprj_io_in_3v3[8]
  PIN mprj_gpio_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3151.055 3379.435 3151.335 ;
    END
  END mprj_gpio_analog[2]
  PIN mprj_gpio_noesd[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3160.255 3379.435 3160.535 ;
    END
  END mprj_gpio_noesd[2]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3140.200 3555.010 3202.900 ;
    END
  END mprj_io[9]
  PIN mprj_io_analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3163.015 3379.435 3163.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3169.455 3379.435 3169.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3184.635 3379.435 3184.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3166.235 3379.435 3166.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3157.035 3379.435 3157.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3187.855 3379.435 3188.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3191.075 3379.435 3191.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3206.255 3379.435 3206.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3172.215 3379.435 3172.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3209.475 3379.435 3209.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3193.835 3379.435 3194.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3147.835 3379.435 3148.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.035 3379.435 3203.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3138.635 3379.435 3138.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_in_3v3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3212.235 3379.435 3212.515 ;
    END
  END mprj_io_in_3v3[9]
  PIN mprj_gpio_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3988.665 210.965 3988.945 ;
    END
  END mprj_gpio_analog[7]
  PIN mprj_gpio_noesd[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3979.465 210.965 3979.745 ;
    END
  END mprj_gpio_noesd[7]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3937.100 95.440 3999.800 ;
    END
  END mprj_io[25]
  PIN mprj_io_analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3976.705 210.965 3976.985 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3970.265 210.965 3970.545 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3955.085 210.965 3955.365 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3973.485 210.965 3973.765 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3982.685 210.965 3982.965 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.865 210.965 3952.145 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3948.645 210.965 3948.925 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3933.465 210.965 3933.745 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3967.505 210.965 3967.785 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3930.245 210.965 3930.525 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3945.885 210.965 3946.165 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3991.885 210.965 3992.165 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3936.685 210.965 3936.965 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4001.085 210.965 4001.365 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in_3v3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3927.485 210.965 3927.765 ;
    END
  END mprj_io_in_3v3[14]
  PIN mprj_gpio_analog[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1403.665 210.965 1403.945 ;
    END
  END mprj_gpio_analog[17]
  PIN mprj_gpio_noesd[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1394.465 210.965 1394.745 ;
    END
  END mprj_gpio_noesd[17]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1352.100 95.440 1414.800 ;
    END
  END mprj_io[35]
  PIN mprj_io_analog_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1391.705 210.965 1391.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1385.265 210.965 1385.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1370.085 210.965 1370.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1388.485 210.965 1388.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1397.685 210.965 1397.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1366.865 210.965 1367.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_holdover[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1363.645 210.965 1363.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1348.465 210.965 1348.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1382.505 210.965 1382.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1345.245 210.965 1345.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1360.885 210.965 1361.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_slow_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1406.885 210.965 1407.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1351.685 210.965 1351.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1416.085 210.965 1416.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in_3v3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1342.485 210.965 1342.765 ;
    END
  END mprj_io_in_3v3[24]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1136.100 95.440 1198.800 ;
    END
  END mprj_io[36]
  PIN mprj_io_analog_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1175.705 210.965 1175.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1169.265 210.965 1169.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1154.085 210.965 1154.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1172.485 210.965 1172.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1181.685 210.965 1181.965 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1150.865 210.965 1151.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_holdover[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1147.645 210.965 1147.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1132.465 210.965 1132.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1166.505 210.965 1166.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1129.245 210.965 1129.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1144.885 210.965 1145.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1190.885 210.965 1191.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1135.685 210.965 1135.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1200.085 210.965 1200.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in_3v3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1126.485 210.965 1126.765 ;
    END
  END mprj_io_in_3v3[25]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 920.100 95.440 982.800 ;
    END
  END mprj_io[37]
  PIN mprj_io_analog_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 959.705 210.965 959.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 953.265 210.965 953.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 938.085 210.965 938.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 956.485 210.965 956.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 965.685 210.965 965.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 934.865 210.965 935.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_holdover[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 931.645 210.965 931.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 916.465 210.965 916.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 950.505 210.965 950.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 913.245 210.965 913.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 928.885 210.965 929.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 974.885 210.965 975.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 919.685 210.965 919.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 984.085 210.965 984.365 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in_3v3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 910.485 210.965 910.765 ;
    END
  END mprj_io_in_3v3[26]
  PIN mprj_gpio_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3772.665 210.965 3772.945 ;
    END
  END mprj_gpio_analog[8]
  PIN mprj_gpio_noesd[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3763.465 210.965 3763.745 ;
    END
  END mprj_gpio_noesd[8]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3721.100 95.440 3783.800 ;
    END
  END mprj_io[26]
  PIN mprj_io_analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3760.705 210.965 3760.985 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3754.265 210.965 3754.545 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3739.085 210.965 3739.365 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3757.485 210.965 3757.765 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3766.685 210.965 3766.965 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.865 210.965 3736.145 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3732.645 210.965 3732.925 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3717.465 210.965 3717.745 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3751.505 210.965 3751.785 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3714.245 210.965 3714.525 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3729.885 210.965 3730.165 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3775.885 210.965 3776.165 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3720.685 210.965 3720.965 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3785.085 210.965 3785.365 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in_3v3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3711.485 210.965 3711.765 ;
    END
  END mprj_io_in_3v3[15]
  PIN mprj_gpio_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3556.665 210.965 3556.945 ;
    END
  END mprj_gpio_analog[9]
  PIN mprj_gpio_noesd[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3547.465 210.965 3547.745 ;
    END
  END mprj_gpio_noesd[9]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3505.100 95.440 3567.800 ;
    END
  END mprj_io[27]
  PIN mprj_io_analog_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3544.705 210.965 3544.985 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3538.265 210.965 3538.545 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3523.085 210.965 3523.365 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3541.485 210.965 3541.765 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3550.685 210.965 3550.965 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.865 210.965 3520.145 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_holdover[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3516.645 210.965 3516.925 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3501.465 210.965 3501.745 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3535.505 210.965 3535.785 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3498.245 210.965 3498.525 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3513.885 210.965 3514.165 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3559.885 210.965 3560.165 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3504.685 210.965 3504.965 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3569.085 210.965 3569.365 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in_3v3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3495.485 210.965 3495.765 ;
    END
  END mprj_io_in_3v3[16]
  PIN mprj_gpio_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.665 210.965 3339.945 ;
    END
  END mprj_gpio_analog[10]
  PIN mprj_gpio_noesd[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.465 210.965 3330.745 ;
    END
  END mprj_gpio_noesd[10]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3288.100 95.440 3350.800 ;
    END
  END mprj_io[28]
  PIN mprj_io_analog_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3327.705 210.965 3327.985 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.265 210.965 3321.545 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3306.085 210.965 3306.365 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.485 210.965 3324.765 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3333.685 210.965 3333.965 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3302.865 210.965 3303.145 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_holdover[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.645 210.965 3299.925 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.465 210.965 3284.745 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.505 210.965 3318.785 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.245 210.965 3281.525 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.885 210.965 3297.165 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3342.885 210.965 3343.165 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3287.685 210.965 3287.965 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3352.085 210.965 3352.365 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in_3v3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.485 210.965 3278.765 ;
    END
  END mprj_io_in_3v3[17]
  PIN mprj_gpio_analog[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.665 210.965 3123.945 ;
    END
  END mprj_gpio_analog[11]
  PIN mprj_gpio_noesd[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.465 210.965 3114.745 ;
    END
  END mprj_gpio_noesd[11]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3072.100 95.440 3134.800 ;
    END
  END mprj_io[29]
  PIN mprj_io_analog_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3111.705 210.965 3111.985 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.265 210.965 3105.545 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3090.085 210.965 3090.365 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.485 210.965 3108.765 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3117.685 210.965 3117.965 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3086.865 210.965 3087.145 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_holdover[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.645 210.965 3083.925 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.465 210.965 3068.745 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.505 210.965 3102.785 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.245 210.965 3065.525 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.885 210.965 3081.165 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3126.885 210.965 3127.165 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3071.685 210.965 3071.965 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3136.085 210.965 3136.365 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in_3v3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.485 210.965 3062.765 ;
    END
  END mprj_io_in_3v3[18]
  PIN mprj_gpio_analog[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.665 210.965 2907.945 ;
    END
  END mprj_gpio_analog[12]
  PIN mprj_gpio_noesd[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.465 210.965 2898.745 ;
    END
  END mprj_gpio_noesd[12]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2856.100 95.440 2918.800 ;
    END
  END mprj_io[30]
  PIN mprj_io_analog_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2895.705 210.965 2895.985 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.265 210.965 2889.545 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2874.085 210.965 2874.365 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.485 210.965 2892.765 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2901.685 210.965 2901.965 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2870.865 210.965 2871.145 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_holdover[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.645 210.965 2867.925 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.465 210.965 2852.745 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.505 210.965 2886.785 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.245 210.965 2849.525 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.885 210.965 2865.165 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2910.885 210.965 2911.165 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2855.685 210.965 2855.965 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2920.085 210.965 2920.365 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in_3v3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.485 210.965 2846.765 ;
    END
  END mprj_io_in_3v3[19]
  PIN mprj_gpio_analog[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.665 210.965 2691.945 ;
    END
  END mprj_gpio_analog[13]
  PIN mprj_gpio_noesd[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.465 210.965 2682.745 ;
    END
  END mprj_gpio_noesd[13]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2640.100 95.440 2702.800 ;
    END
  END mprj_io[31]
  PIN mprj_io_analog_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2679.705 210.965 2679.985 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.265 210.965 2673.545 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2658.085 210.965 2658.365 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.485 210.965 2676.765 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2685.685 210.965 2685.965 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2654.865 210.965 2655.145 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_holdover[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.645 210.965 2651.925 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.465 210.965 2636.745 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.505 210.965 2670.785 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.245 210.965 2633.525 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.885 210.965 2649.165 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2694.885 210.965 2695.165 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2639.685 210.965 2639.965 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2704.085 210.965 2704.365 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in_3v3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.485 210.965 2630.765 ;
    END
  END mprj_io_in_3v3[20]
  PIN mprj_gpio_analog[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2052.665 210.965 2052.945 ;
    END
  END mprj_gpio_analog[14]
  PIN mprj_gpio_noesd[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2043.465 210.965 2043.745 ;
    END
  END mprj_gpio_noesd[14]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2001.100 95.440 2063.800 ;
    END
  END mprj_io[32]
  PIN mprj_io_analog_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2040.705 210.965 2040.985 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2034.265 210.965 2034.545 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2019.085 210.965 2019.365 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2037.485 210.965 2037.765 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2046.685 210.965 2046.965 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2015.865 210.965 2016.145 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_holdover[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2012.645 210.965 2012.925 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1997.465 210.965 1997.745 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2031.505 210.965 2031.785 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1994.245 210.965 1994.525 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2009.885 210.965 2010.165 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2055.885 210.965 2056.165 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2000.685 210.965 2000.965 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2065.085 210.965 2065.365 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in_3v3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1991.485 210.965 1991.765 ;
    END
  END mprj_io_in_3v3[21]
  PIN mprj_gpio_analog[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1836.665 210.965 1836.945 ;
    END
  END mprj_gpio_analog[15]
  PIN mprj_gpio_noesd[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1827.465 210.965 1827.745 ;
    END
  END mprj_gpio_noesd[15]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1785.100 95.440 1847.800 ;
    END
  END mprj_io[33]
  PIN mprj_io_analog_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1824.705 210.965 1824.985 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1818.265 210.965 1818.545 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1803.085 210.965 1803.365 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1821.485 210.965 1821.765 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1830.685 210.965 1830.965 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1799.865 210.965 1800.145 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_holdover[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1796.645 210.965 1796.925 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1781.465 210.965 1781.745 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1815.505 210.965 1815.785 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1778.245 210.965 1778.525 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1793.885 210.965 1794.165 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1839.885 210.965 1840.165 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1784.685 210.965 1784.965 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1849.085 210.965 1849.365 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in_3v3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1775.485 210.965 1775.765 ;
    END
  END mprj_io_in_3v3[22]
  PIN mprj_gpio_analog[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1619.665 210.965 1619.945 ;
    END
  END mprj_gpio_analog[16]
  PIN mprj_gpio_noesd[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1610.465 210.965 1610.745 ;
    END
  END mprj_gpio_noesd[16]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1568.100 95.440 1630.800 ;
    END
  END mprj_io[34]
  PIN mprj_io_analog_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1607.705 210.965 1607.985 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1601.265 210.965 1601.545 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1586.085 210.965 1586.365 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1604.485 210.965 1604.765 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1613.685 210.965 1613.965 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1582.865 210.965 1583.145 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_holdover[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1579.645 210.965 1579.925 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1564.465 210.965 1564.745 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1598.505 210.965 1598.785 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1561.245 210.965 1561.525 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1576.885 210.965 1577.165 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1622.885 210.965 1623.165 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1567.685 210.965 1567.965 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1632.085 210.965 1632.365 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in_3v3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1558.485 210.965 1558.765 ;
    END
  END mprj_io_in_3v3[23]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3368.650 4277.100 3368.970 4277.160 ;
        RECT 3376.930 4277.100 3377.250 4277.160 ;
        RECT 3368.650 4276.960 3377.250 4277.100 ;
        RECT 3368.650 4276.900 3368.970 4276.960 ;
        RECT 3376.930 4276.900 3377.250 4276.960 ;
        RECT 211.210 3940.160 211.530 3940.220 ;
        RECT 212.130 3940.160 212.450 3940.220 ;
        RECT 211.210 3940.020 212.450 3940.160 ;
        RECT 211.210 3939.960 211.530 3940.020 ;
        RECT 212.130 3939.960 212.450 3940.020 ;
        RECT 3368.650 3866.720 3368.970 3866.780 ;
        RECT 3376.010 3866.720 3376.330 3866.780 ;
        RECT 3376.930 3866.720 3377.250 3866.780 ;
        RECT 3368.650 3866.580 3377.250 3866.720 ;
        RECT 3368.650 3866.520 3368.970 3866.580 ;
        RECT 3376.010 3866.520 3376.330 3866.580 ;
        RECT 3376.930 3866.520 3377.250 3866.580 ;
        RECT 3368.650 3845.640 3368.970 3845.700 ;
        RECT 3376.010 3845.640 3376.330 3845.700 ;
        RECT 3376.930 3845.640 3377.250 3845.700 ;
        RECT 3368.650 3845.500 3377.250 3845.640 ;
        RECT 3368.650 3845.440 3368.970 3845.500 ;
        RECT 3376.010 3845.440 3376.330 3845.500 ;
        RECT 3376.930 3845.440 3377.250 3845.500 ;
        RECT 3368.650 3643.000 3368.970 3643.060 ;
        RECT 3376.930 3643.000 3377.250 3643.060 ;
        RECT 3368.650 3642.860 3377.250 3643.000 ;
        RECT 3368.650 3642.800 3368.970 3642.860 ;
        RECT 3376.930 3642.800 3377.250 3642.860 ;
        RECT 3367.270 3620.220 3367.590 3620.280 ;
        RECT 3376.930 3620.220 3377.250 3620.280 ;
        RECT 3367.270 3620.080 3377.250 3620.220 ;
        RECT 3367.270 3620.020 3367.590 3620.080 ;
        RECT 3376.930 3620.020 3377.250 3620.080 ;
        RECT 3367.270 3421.660 3367.590 3421.720 ;
        RECT 3376.470 3421.660 3376.790 3421.720 ;
        RECT 3367.270 3421.520 3376.790 3421.660 ;
        RECT 3367.270 3421.460 3367.590 3421.520 ;
        RECT 3376.470 3421.460 3376.790 3421.520 ;
        RECT 3369.110 3400.580 3369.430 3400.640 ;
        RECT 3376.930 3400.580 3377.250 3400.640 ;
        RECT 3369.110 3400.440 3377.250 3400.580 ;
        RECT 3369.110 3400.380 3369.430 3400.440 ;
        RECT 3376.930 3400.380 3377.250 3400.440 ;
        RECT 3369.110 3200.660 3369.430 3200.720 ;
        RECT 3376.470 3200.660 3376.790 3200.720 ;
        RECT 3369.110 3200.520 3376.790 3200.660 ;
        RECT 3369.110 3200.460 3369.430 3200.520 ;
        RECT 3376.470 3200.460 3376.790 3200.520 ;
        RECT 3368.650 3178.900 3368.970 3178.960 ;
        RECT 3376.470 3178.900 3376.790 3178.960 ;
        RECT 3368.650 3178.760 3376.790 3178.900 ;
        RECT 3368.650 3178.700 3368.970 3178.760 ;
        RECT 3376.470 3178.700 3376.790 3178.760 ;
        RECT 3368.650 2980.680 3368.970 2980.740 ;
        RECT 3376.010 2980.680 3376.330 2980.740 ;
        RECT 3376.930 2980.680 3377.250 2980.740 ;
        RECT 3368.650 2980.540 3377.250 2980.680 ;
        RECT 3368.650 2980.480 3368.970 2980.540 ;
        RECT 3376.010 2980.480 3376.330 2980.540 ;
        RECT 3376.930 2980.480 3377.250 2980.540 ;
        RECT 3368.650 2954.160 3368.970 2954.220 ;
        RECT 3376.010 2954.160 3376.330 2954.220 ;
        RECT 3376.930 2954.160 3377.250 2954.220 ;
        RECT 3368.650 2954.020 3377.250 2954.160 ;
        RECT 3368.650 2953.960 3368.970 2954.020 ;
        RECT 3376.010 2953.960 3376.330 2954.020 ;
        RECT 3376.930 2953.960 3377.250 2954.020 ;
        RECT 208.910 2882.760 209.230 2882.820 ;
        RECT 211.210 2882.760 211.530 2882.820 ;
        RECT 212.130 2882.760 212.450 2882.820 ;
        RECT 208.910 2882.620 212.450 2882.760 ;
        RECT 208.910 2882.560 209.230 2882.620 ;
        RECT 211.210 2882.560 211.530 2882.620 ;
        RECT 212.130 2882.560 212.450 2882.620 ;
        RECT 3368.650 2757.640 3368.970 2757.700 ;
        RECT 3376.010 2757.640 3376.330 2757.700 ;
        RECT 3368.650 2757.500 3376.330 2757.640 ;
        RECT 3368.650 2757.440 3368.970 2757.500 ;
        RECT 3376.010 2757.440 3376.330 2757.500 ;
        RECT 3367.270 2735.200 3367.590 2735.260 ;
        RECT 3376.010 2735.200 3376.330 2735.260 ;
        RECT 3376.930 2735.200 3377.250 2735.260 ;
        RECT 3367.270 2735.060 3377.250 2735.200 ;
        RECT 3367.270 2735.000 3367.590 2735.060 ;
        RECT 3376.010 2735.000 3376.330 2735.060 ;
        RECT 3376.930 2735.000 3377.250 2735.060 ;
        RECT 3367.730 1864.120 3368.050 1864.180 ;
        RECT 3376.930 1864.120 3377.250 1864.180 ;
        RECT 3367.730 1863.980 3377.250 1864.120 ;
        RECT 3367.730 1863.920 3368.050 1863.980 ;
        RECT 3376.930 1863.920 3377.250 1863.980 ;
        RECT 3367.730 1665.560 3368.050 1665.620 ;
        RECT 3376.470 1665.560 3376.790 1665.620 ;
        RECT 3367.730 1665.420 3376.790 1665.560 ;
        RECT 3367.730 1665.360 3368.050 1665.420 ;
        RECT 3376.470 1665.360 3376.790 1665.420 ;
        RECT 3368.650 1641.420 3368.970 1641.480 ;
        RECT 3376.930 1641.420 3377.250 1641.480 ;
        RECT 3368.650 1641.280 3377.250 1641.420 ;
        RECT 3368.650 1641.220 3368.970 1641.280 ;
        RECT 3376.930 1641.220 3377.250 1641.280 ;
        RECT 211.210 1565.600 211.530 1565.660 ;
        RECT 211.210 1565.460 211.900 1565.600 ;
        RECT 211.210 1565.400 211.530 1565.460 ;
        RECT 211.760 1564.640 211.900 1565.460 ;
        RECT 211.670 1564.380 211.990 1564.640 ;
        RECT 3368.650 1446.600 3368.970 1446.660 ;
        RECT 3376.930 1446.600 3377.250 1446.660 ;
        RECT 3368.650 1446.460 3377.250 1446.600 ;
        RECT 3368.650 1446.400 3368.970 1446.460 ;
        RECT 3376.930 1446.400 3377.250 1446.460 ;
        RECT 211.670 1420.560 211.990 1420.820 ;
        RECT 211.760 1419.800 211.900 1420.560 ;
        RECT 3368.650 1420.420 3368.970 1420.480 ;
        RECT 3376.930 1420.420 3377.250 1420.480 ;
        RECT 3368.650 1420.280 3377.250 1420.420 ;
        RECT 3368.650 1420.220 3368.970 1420.280 ;
        RECT 3376.930 1420.220 3377.250 1420.280 ;
        RECT 211.670 1419.540 211.990 1419.800 ;
        RECT 3368.650 1223.220 3368.970 1223.280 ;
        RECT 3376.930 1223.220 3377.250 1223.280 ;
        RECT 3368.650 1223.080 3377.250 1223.220 ;
        RECT 3368.650 1223.020 3368.970 1223.080 ;
        RECT 3376.930 1223.020 3377.250 1223.080 ;
        RECT 3368.650 1198.400 3368.970 1198.460 ;
        RECT 3376.930 1198.400 3377.250 1198.460 ;
        RECT 3368.650 1198.260 3377.250 1198.400 ;
        RECT 3368.650 1198.200 3368.970 1198.260 ;
        RECT 3376.930 1198.200 3377.250 1198.260 ;
        RECT 3368.650 1002.220 3368.970 1002.280 ;
        RECT 3376.930 1002.220 3377.250 1002.280 ;
        RECT 3368.650 1002.080 3377.250 1002.220 ;
        RECT 3368.650 1002.020 3368.970 1002.080 ;
        RECT 3376.930 1002.020 3377.250 1002.080 ;
        RECT 3368.650 979.100 3368.970 979.160 ;
        RECT 3376.930 979.100 3377.250 979.160 ;
        RECT 3368.650 978.960 3377.250 979.100 ;
        RECT 3368.650 978.900 3368.970 978.960 ;
        RECT 3376.930 978.900 3377.250 978.960 ;
        RECT 3368.650 781.560 3368.970 781.620 ;
        RECT 3376.930 781.560 3377.250 781.620 ;
        RECT 3368.650 781.420 3377.250 781.560 ;
        RECT 3368.650 781.360 3368.970 781.420 ;
        RECT 3376.930 781.360 3377.250 781.420 ;
        RECT 3369.110 758.780 3369.430 758.840 ;
        RECT 3376.470 758.780 3376.790 758.840 ;
        RECT 3369.110 758.640 3376.790 758.780 ;
        RECT 3369.110 758.580 3369.430 758.640 ;
        RECT 3376.470 758.580 3376.790 758.640 ;
        RECT 3369.110 559.200 3369.430 559.260 ;
        RECT 3376.930 559.200 3377.250 559.260 ;
        RECT 3369.110 559.060 3377.250 559.200 ;
        RECT 3369.110 559.000 3369.430 559.060 ;
        RECT 3376.930 559.000 3377.250 559.060 ;
        RECT 3368.190 536.760 3368.510 536.820 ;
        RECT 3376.470 536.760 3376.790 536.820 ;
        RECT 3368.190 536.620 3376.790 536.760 ;
        RECT 3368.190 536.560 3368.510 536.620 ;
        RECT 3376.470 536.560 3376.790 536.620 ;
        RECT 3368.190 234.840 3368.510 234.900 ;
        RECT 2637.340 234.700 3368.510 234.840 ;
        RECT 2637.340 234.560 2637.480 234.700 ;
        RECT 3368.190 234.640 3368.510 234.700 ;
        RECT 2637.250 234.300 2637.570 234.560 ;
        RECT 211.670 228.040 211.990 228.100 ;
        RECT 718.130 228.040 718.450 228.100 ;
        RECT 211.670 227.900 718.450 228.040 ;
        RECT 211.670 227.840 211.990 227.900 ;
        RECT 718.130 227.840 718.450 227.900 ;
        RECT 1815.230 221.580 1815.550 221.640 ;
        RECT 2067.770 221.580 2068.090 221.640 ;
        RECT 2089.390 221.580 2089.710 221.640 ;
        RECT 2341.470 221.580 2341.790 221.640 ;
        RECT 2363.090 221.580 2363.410 221.640 ;
        RECT 1517.930 221.440 1519.680 221.580 ;
        RECT 999.190 221.240 999.510 221.300 ;
        RECT 1517.930 221.240 1518.070 221.440 ;
        RECT 1519.540 221.300 1519.680 221.440 ;
        RECT 1807.730 221.440 2615.860 221.580 ;
        RECT 999.190 221.100 1518.070 221.240 ;
        RECT 1519.450 221.240 1519.770 221.300 ;
        RECT 1541.070 221.240 1541.390 221.300 ;
        RECT 1793.610 221.240 1793.930 221.300 ;
        RECT 1807.730 221.240 1807.870 221.440 ;
        RECT 1815.230 221.380 1815.550 221.440 ;
        RECT 2067.770 221.380 2068.090 221.440 ;
        RECT 2089.390 221.380 2089.710 221.440 ;
        RECT 2341.470 221.380 2341.790 221.440 ;
        RECT 2363.090 221.380 2363.410 221.440 ;
        RECT 1519.450 221.100 1807.870 221.240 ;
        RECT 999.190 221.040 999.510 221.100 ;
        RECT 1519.450 221.040 1519.770 221.100 ;
        RECT 1541.070 221.040 1541.390 221.100 ;
        RECT 1793.610 221.040 1793.930 221.100 ;
        RECT 2615.720 220.960 2615.860 221.440 ;
        RECT 718.130 220.900 718.450 220.960 ;
        RECT 725.490 220.900 725.810 220.960 ;
        RECT 976.650 220.900 976.970 220.960 ;
        RECT 998.270 220.900 998.590 220.960 ;
        RECT 718.130 220.760 998.590 220.900 ;
        RECT 718.130 220.700 718.450 220.760 ;
        RECT 725.490 220.700 725.810 220.760 ;
        RECT 976.650 220.700 976.970 220.760 ;
        RECT 998.270 220.700 998.590 220.760 ;
        RECT 2615.630 220.900 2615.950 220.960 ;
        RECT 2637.250 220.900 2637.570 220.960 ;
        RECT 2615.630 220.760 2637.570 220.900 ;
        RECT 2615.630 220.700 2615.950 220.760 ;
        RECT 2637.250 220.700 2637.570 220.760 ;
      LAYER via ;
        RECT 3368.680 4276.900 3368.940 4277.160 ;
        RECT 3376.960 4276.900 3377.220 4277.160 ;
        RECT 211.240 3939.960 211.500 3940.220 ;
        RECT 212.160 3939.960 212.420 3940.220 ;
        RECT 3368.680 3866.520 3368.940 3866.780 ;
        RECT 3376.040 3866.520 3376.300 3866.780 ;
        RECT 3376.960 3866.520 3377.220 3866.780 ;
        RECT 3368.680 3845.440 3368.940 3845.700 ;
        RECT 3376.040 3845.440 3376.300 3845.700 ;
        RECT 3376.960 3845.440 3377.220 3845.700 ;
        RECT 3368.680 3642.800 3368.940 3643.060 ;
        RECT 3376.960 3642.800 3377.220 3643.060 ;
        RECT 3367.300 3620.020 3367.560 3620.280 ;
        RECT 3376.960 3620.020 3377.220 3620.280 ;
        RECT 3367.300 3421.460 3367.560 3421.720 ;
        RECT 3376.500 3421.460 3376.760 3421.720 ;
        RECT 3369.140 3400.380 3369.400 3400.640 ;
        RECT 3376.960 3400.380 3377.220 3400.640 ;
        RECT 3369.140 3200.460 3369.400 3200.720 ;
        RECT 3376.500 3200.460 3376.760 3200.720 ;
        RECT 3368.680 3178.700 3368.940 3178.960 ;
        RECT 3376.500 3178.700 3376.760 3178.960 ;
        RECT 3368.680 2980.480 3368.940 2980.740 ;
        RECT 3376.040 2980.480 3376.300 2980.740 ;
        RECT 3376.960 2980.480 3377.220 2980.740 ;
        RECT 3368.680 2953.960 3368.940 2954.220 ;
        RECT 3376.040 2953.960 3376.300 2954.220 ;
        RECT 3376.960 2953.960 3377.220 2954.220 ;
        RECT 208.940 2882.560 209.200 2882.820 ;
        RECT 211.240 2882.560 211.500 2882.820 ;
        RECT 212.160 2882.560 212.420 2882.820 ;
        RECT 3368.680 2757.440 3368.940 2757.700 ;
        RECT 3376.040 2757.440 3376.300 2757.700 ;
        RECT 3367.300 2735.000 3367.560 2735.260 ;
        RECT 3376.040 2735.000 3376.300 2735.260 ;
        RECT 3376.960 2735.000 3377.220 2735.260 ;
        RECT 3367.760 1863.920 3368.020 1864.180 ;
        RECT 3376.960 1863.920 3377.220 1864.180 ;
        RECT 3367.760 1665.360 3368.020 1665.620 ;
        RECT 3376.500 1665.360 3376.760 1665.620 ;
        RECT 3368.680 1641.220 3368.940 1641.480 ;
        RECT 3376.960 1641.220 3377.220 1641.480 ;
        RECT 211.240 1565.400 211.500 1565.660 ;
        RECT 211.700 1564.380 211.960 1564.640 ;
        RECT 3368.680 1446.400 3368.940 1446.660 ;
        RECT 3376.960 1446.400 3377.220 1446.660 ;
        RECT 211.700 1420.560 211.960 1420.820 ;
        RECT 3368.680 1420.220 3368.940 1420.480 ;
        RECT 3376.960 1420.220 3377.220 1420.480 ;
        RECT 211.700 1419.540 211.960 1419.800 ;
        RECT 3368.680 1223.020 3368.940 1223.280 ;
        RECT 3376.960 1223.020 3377.220 1223.280 ;
        RECT 3368.680 1198.200 3368.940 1198.460 ;
        RECT 3376.960 1198.200 3377.220 1198.460 ;
        RECT 3368.680 1002.020 3368.940 1002.280 ;
        RECT 3376.960 1002.020 3377.220 1002.280 ;
        RECT 3368.680 978.900 3368.940 979.160 ;
        RECT 3376.960 978.900 3377.220 979.160 ;
        RECT 3368.680 781.360 3368.940 781.620 ;
        RECT 3376.960 781.360 3377.220 781.620 ;
        RECT 3369.140 758.580 3369.400 758.840 ;
        RECT 3376.500 758.580 3376.760 758.840 ;
        RECT 3369.140 559.000 3369.400 559.260 ;
        RECT 3376.960 559.000 3377.220 559.260 ;
        RECT 3368.220 536.560 3368.480 536.820 ;
        RECT 3376.500 536.560 3376.760 536.820 ;
        RECT 3368.220 234.640 3368.480 234.900 ;
        RECT 2637.280 234.300 2637.540 234.560 ;
        RECT 211.700 227.840 211.960 228.100 ;
        RECT 718.160 227.840 718.420 228.100 ;
        RECT 999.220 221.040 999.480 221.300 ;
        RECT 1519.480 221.040 1519.740 221.300 ;
        RECT 1541.100 221.040 1541.360 221.300 ;
        RECT 1793.640 221.040 1793.900 221.300 ;
        RECT 1815.260 221.380 1815.520 221.640 ;
        RECT 2067.800 221.380 2068.060 221.640 ;
        RECT 2089.420 221.380 2089.680 221.640 ;
        RECT 2341.500 221.380 2341.760 221.640 ;
        RECT 2363.120 221.380 2363.380 221.640 ;
        RECT 718.160 220.700 718.420 220.960 ;
        RECT 725.520 220.700 725.780 220.960 ;
        RECT 976.680 220.700 976.940 220.960 ;
        RECT 998.300 220.700 998.560 220.960 ;
        RECT 2615.660 220.700 2615.920 220.960 ;
        RECT 2637.280 220.700 2637.540 220.960 ;
      LAYER met2 ;
        RECT 3377.035 4301.410 3379.435 4301.555 ;
        RECT 3376.560 4301.275 3379.435 4301.410 ;
        RECT 3376.560 4301.270 3377.090 4301.275 ;
        RECT 3376.560 4279.865 3376.700 4301.270 ;
        RECT 3377.035 4279.865 3379.435 4279.935 ;
        RECT 3376.560 4279.725 3379.435 4279.865 ;
        RECT 3377.020 4279.655 3379.435 4279.725 ;
        RECT 3377.020 4277.190 3377.160 4279.655 ;
        RECT 3368.680 4276.870 3368.940 4277.190 ;
        RECT 3376.960 4276.870 3377.220 4277.190 ;
        RECT 208.610 3961.345 211.440 3961.410 ;
        RECT 208.565 3961.270 211.440 3961.345 ;
        RECT 208.565 3961.065 210.965 3961.270 ;
        RECT 211.300 3940.330 211.440 3961.270 ;
        RECT 209.460 3940.250 211.440 3940.330 ;
        RECT 209.460 3940.190 211.500 3940.250 ;
        RECT 209.460 3939.725 209.600 3940.190 ;
        RECT 211.240 3939.930 211.500 3940.190 ;
        RECT 212.160 3939.930 212.420 3940.250 ;
        RECT 211.300 3939.775 211.440 3939.930 ;
        RECT 208.565 3939.445 210.965 3939.725 ;
        RECT 212.220 3747.890 212.360 3939.930 ;
        RECT 3368.740 3866.810 3368.880 4276.870 ;
        RECT 3368.680 3866.490 3368.940 3866.810 ;
        RECT 3376.040 3866.490 3376.300 3866.810 ;
        RECT 3376.960 3866.490 3377.220 3866.810 ;
        RECT 3376.100 3845.730 3376.240 3866.490 ;
        RECT 3377.020 3864.555 3377.160 3866.490 ;
        RECT 3377.020 3864.415 3379.435 3864.555 ;
        RECT 3377.035 3864.275 3379.435 3864.415 ;
        RECT 3368.680 3845.410 3368.940 3845.730 ;
        RECT 3376.040 3845.410 3376.300 3845.730 ;
        RECT 3376.960 3845.410 3377.220 3845.730 ;
        RECT 209.000 3747.750 212.360 3747.890 ;
        RECT 209.000 3745.345 209.140 3747.750 ;
        RECT 208.565 3745.065 210.965 3745.345 ;
        RECT 208.610 3745.030 209.140 3745.065 ;
        RECT 208.565 3723.655 210.965 3723.725 ;
        RECT 211.300 3723.655 211.440 3747.750 ;
        RECT 208.565 3723.515 211.440 3723.655 ;
        RECT 208.565 3723.445 210.965 3723.515 ;
        RECT 211.300 3643.270 211.440 3723.515 ;
        RECT 211.300 3643.130 211.900 3643.270 ;
        RECT 208.565 3529.275 210.965 3529.345 ;
        RECT 211.760 3529.275 211.900 3643.130 ;
        RECT 3368.740 3643.090 3368.880 3845.410 ;
        RECT 3377.020 3842.935 3377.160 3845.410 ;
        RECT 3377.020 3842.795 3379.435 3842.935 ;
        RECT 3377.035 3842.655 3379.435 3842.795 ;
        RECT 3368.680 3642.770 3368.940 3643.090 ;
        RECT 3376.960 3642.770 3377.220 3643.090 ;
        RECT 3377.020 3642.555 3377.160 3642.770 ;
        RECT 3377.020 3642.490 3379.435 3642.555 ;
        RECT 3376.560 3642.350 3379.435 3642.490 ;
        RECT 3376.560 3623.450 3376.700 3642.350 ;
        RECT 3377.035 3642.275 3379.435 3642.350 ;
        RECT 3376.560 3623.310 3377.160 3623.450 ;
        RECT 3377.020 3620.935 3377.160 3623.310 ;
        RECT 3377.020 3620.655 3379.435 3620.935 ;
        RECT 3377.020 3620.310 3377.160 3620.655 ;
        RECT 3367.300 3619.990 3367.560 3620.310 ;
        RECT 3376.960 3619.990 3377.220 3620.310 ;
        RECT 208.565 3529.135 211.900 3529.275 ;
        RECT 208.565 3529.065 210.965 3529.135 ;
        RECT 208.565 3507.445 210.965 3507.725 ;
        RECT 209.460 3507.170 209.600 3507.445 ;
        RECT 211.300 3507.170 211.440 3529.135 ;
        RECT 209.460 3507.030 211.440 3507.170 ;
        RECT 211.300 3450.070 211.440 3507.030 ;
        RECT 211.300 3449.930 211.900 3450.070 ;
        RECT 211.760 3312.690 211.900 3449.930 ;
        RECT 3367.360 3421.750 3367.500 3619.990 ;
        RECT 3376.560 3421.750 3376.700 3421.905 ;
        RECT 3367.300 3421.430 3367.560 3421.750 ;
        RECT 3376.500 3421.490 3376.760 3421.750 ;
        RECT 3377.035 3421.490 3379.435 3421.555 ;
        RECT 3376.500 3421.430 3379.435 3421.490 ;
        RECT 3376.560 3421.350 3379.435 3421.430 ;
        RECT 3376.560 3401.770 3376.700 3421.350 ;
        RECT 3377.035 3421.275 3379.435 3421.350 ;
        RECT 3376.560 3401.630 3377.160 3401.770 ;
        RECT 3377.020 3400.670 3377.160 3401.630 ;
        RECT 3369.140 3400.350 3369.400 3400.670 ;
        RECT 3376.960 3400.350 3377.220 3400.670 ;
        RECT 209.460 3312.550 211.900 3312.690 ;
        RECT 209.460 3312.345 209.600 3312.550 ;
        RECT 208.565 3312.065 210.965 3312.345 ;
        RECT 208.565 3290.655 210.965 3290.725 ;
        RECT 211.300 3290.655 211.440 3312.550 ;
        RECT 208.565 3290.515 211.440 3290.655 ;
        RECT 208.565 3290.445 210.965 3290.515 ;
        RECT 211.300 3256.870 211.440 3290.515 ;
        RECT 211.300 3256.730 211.900 3256.870 ;
        RECT 208.565 3096.065 210.965 3096.345 ;
        RECT 209.460 3095.770 209.600 3096.065 ;
        RECT 211.760 3095.770 211.900 3256.730 ;
        RECT 3369.200 3200.750 3369.340 3400.350 ;
        RECT 3377.020 3399.935 3377.160 3400.350 ;
        RECT 3377.020 3399.660 3379.435 3399.935 ;
        RECT 3377.035 3399.655 3379.435 3399.660 ;
        RECT 3376.560 3200.750 3376.700 3200.905 ;
        RECT 3369.140 3200.430 3369.400 3200.750 ;
        RECT 3376.500 3200.490 3376.760 3200.750 ;
        RECT 3377.035 3200.490 3379.435 3200.555 ;
        RECT 3376.500 3200.430 3379.435 3200.490 ;
        RECT 3376.560 3200.350 3379.435 3200.430 ;
        RECT 3376.560 3179.410 3376.700 3200.350 ;
        RECT 3377.035 3200.275 3379.435 3200.350 ;
        RECT 3376.560 3179.270 3377.160 3179.410 ;
        RECT 3376.560 3178.990 3376.700 3179.270 ;
        RECT 3368.680 3178.670 3368.940 3178.990 ;
        RECT 3376.500 3178.670 3376.760 3178.990 ;
        RECT 3377.020 3178.935 3377.160 3179.270 ;
        RECT 209.460 3095.630 211.900 3095.770 ;
        RECT 208.565 3074.445 210.965 3074.725 ;
        RECT 209.000 3074.010 209.140 3074.445 ;
        RECT 211.300 3074.010 211.440 3095.630 ;
        RECT 209.000 3073.870 211.900 3074.010 ;
        RECT 211.760 3022.270 211.900 3073.870 ;
        RECT 211.760 3022.130 212.360 3022.270 ;
        RECT 212.220 2882.850 212.360 3022.130 ;
        RECT 3368.740 2980.770 3368.880 3178.670 ;
        RECT 3377.020 3178.660 3379.435 3178.935 ;
        RECT 3377.035 3178.655 3379.435 3178.660 ;
        RECT 3368.680 2980.450 3368.940 2980.770 ;
        RECT 3376.040 2980.450 3376.300 2980.770 ;
        RECT 3376.960 2980.450 3377.220 2980.770 ;
        RECT 3376.100 2954.250 3376.240 2980.450 ;
        RECT 3377.020 2978.555 3377.160 2980.450 ;
        RECT 3377.020 2978.415 3379.435 2978.555 ;
        RECT 3377.035 2978.275 3379.435 2978.415 ;
        RECT 3377.035 2956.795 3379.435 2956.935 ;
        RECT 3377.020 2956.655 3379.435 2956.795 ;
        RECT 3377.020 2954.250 3377.160 2956.655 ;
        RECT 3368.680 2953.930 3368.940 2954.250 ;
        RECT 3376.040 2953.930 3376.300 2954.250 ;
        RECT 3376.960 2953.930 3377.220 2954.250 ;
        RECT 208.940 2882.530 209.200 2882.850 ;
        RECT 211.240 2882.530 211.500 2882.850 ;
        RECT 212.160 2882.530 212.420 2882.850 ;
        RECT 209.000 2880.345 209.140 2882.530 ;
        RECT 208.565 2880.065 210.965 2880.345 ;
        RECT 208.565 2858.655 210.965 2858.725 ;
        RECT 211.300 2858.655 211.440 2882.530 ;
        RECT 208.565 2858.515 211.900 2858.655 ;
        RECT 208.565 2858.445 210.965 2858.515 ;
        RECT 208.565 2664.275 210.965 2664.345 ;
        RECT 211.760 2664.275 211.900 2858.515 ;
        RECT 3368.740 2757.730 3368.880 2953.930 ;
        RECT 3376.100 2757.730 3376.240 2757.900 ;
        RECT 3368.680 2757.410 3368.940 2757.730 ;
        RECT 3376.040 2757.485 3376.300 2757.730 ;
        RECT 3377.035 2757.485 3379.435 2757.555 ;
        RECT 3376.040 2757.410 3379.435 2757.485 ;
        RECT 3376.100 2757.345 3379.435 2757.410 ;
        RECT 3376.100 2735.290 3376.240 2757.345 ;
        RECT 3377.035 2757.275 3379.435 2757.345 ;
        RECT 3377.035 2735.795 3379.435 2735.935 ;
        RECT 3377.020 2735.655 3379.435 2735.795 ;
        RECT 3377.020 2735.290 3377.160 2735.655 ;
        RECT 3367.300 2734.970 3367.560 2735.290 ;
        RECT 3376.040 2734.970 3376.300 2735.290 ;
        RECT 3376.960 2734.970 3377.220 2735.290 ;
        RECT 208.565 2664.135 211.900 2664.275 ;
        RECT 208.565 2664.065 210.965 2664.135 ;
        RECT 208.565 2642.445 210.965 2642.725 ;
        RECT 209.460 2642.210 209.600 2642.445 ;
        RECT 211.300 2642.210 211.440 2664.135 ;
        RECT 209.460 2642.070 211.440 2642.210 ;
        RECT 211.300 2097.670 211.440 2642.070 ;
        RECT 211.300 2097.530 211.900 2097.670 ;
        RECT 211.760 2027.490 211.900 2097.530 ;
        RECT 209.000 2027.350 211.900 2027.490 ;
        RECT 209.000 2025.345 209.140 2027.350 ;
        RECT 208.565 2025.065 210.965 2025.345 ;
        RECT 208.565 2003.690 210.965 2003.725 ;
        RECT 211.300 2003.690 211.440 2027.350 ;
        RECT 208.565 2003.550 211.440 2003.690 ;
        RECT 208.565 2003.445 210.965 2003.550 ;
        RECT 211.300 1904.470 211.440 2003.550 ;
        RECT 3367.360 1904.470 3367.500 2734.970 ;
        RECT 211.300 1904.330 211.900 1904.470 ;
        RECT 3367.360 1904.330 3367.960 1904.470 ;
        RECT 208.565 1809.065 210.965 1809.345 ;
        RECT 209.000 1807.870 209.140 1809.065 ;
        RECT 211.760 1807.870 211.900 1904.330 ;
        RECT 3367.820 1864.210 3367.960 1904.330 ;
        RECT 3377.035 1886.485 3379.435 1886.555 ;
        RECT 3376.560 1886.345 3379.435 1886.485 ;
        RECT 3376.560 1864.290 3376.700 1886.345 ;
        RECT 3377.035 1886.275 3379.435 1886.345 ;
        RECT 3377.035 1864.900 3379.435 1864.935 ;
        RECT 3377.020 1864.655 3379.435 1864.900 ;
        RECT 3377.020 1864.290 3377.160 1864.655 ;
        RECT 3376.560 1864.210 3377.160 1864.290 ;
        RECT 3367.760 1863.890 3368.020 1864.210 ;
        RECT 3376.560 1864.150 3377.220 1864.210 ;
        RECT 3376.960 1863.890 3377.220 1864.150 ;
        RECT 209.000 1807.730 211.900 1807.870 ;
        RECT 208.565 1787.655 210.965 1787.725 ;
        RECT 211.300 1787.655 211.440 1807.730 ;
        RECT 208.565 1787.515 211.900 1787.655 ;
        RECT 208.565 1787.445 210.965 1787.515 ;
        RECT 208.565 1592.065 210.965 1592.345 ;
        RECT 209.460 1591.610 209.600 1592.065 ;
        RECT 211.760 1591.610 211.900 1787.515 ;
        RECT 3367.820 1665.650 3367.960 1863.890 ;
        RECT 3376.560 1665.650 3376.700 1665.900 ;
        RECT 3367.760 1665.330 3368.020 1665.650 ;
        RECT 3376.500 1665.485 3376.760 1665.650 ;
        RECT 3377.035 1665.485 3379.435 1665.555 ;
        RECT 3376.500 1665.345 3379.435 1665.485 ;
        RECT 3376.500 1665.330 3376.760 1665.345 ;
        RECT 3376.560 1643.290 3376.700 1665.330 ;
        RECT 3377.035 1665.275 3379.435 1665.345 ;
        RECT 3377.035 1643.900 3379.435 1643.935 ;
        RECT 3377.020 1643.655 3379.435 1643.900 ;
        RECT 3377.020 1643.290 3377.160 1643.655 ;
        RECT 3376.560 1643.150 3377.160 1643.290 ;
        RECT 3377.020 1641.510 3377.160 1643.150 ;
        RECT 3368.680 1641.190 3368.940 1641.510 ;
        RECT 3376.960 1641.190 3377.220 1641.510 ;
        RECT 209.460 1591.470 211.900 1591.610 ;
        RECT 208.565 1570.445 210.965 1570.725 ;
        RECT 208.610 1570.390 209.600 1570.445 ;
        RECT 209.460 1569.850 209.600 1570.390 ;
        RECT 211.300 1569.850 211.440 1591.470 ;
        RECT 209.460 1569.710 211.440 1569.850 ;
        RECT 211.300 1565.690 211.440 1569.710 ;
        RECT 211.240 1565.370 211.500 1565.690 ;
        RECT 211.700 1564.350 211.960 1564.670 ;
        RECT 211.760 1420.850 211.900 1564.350 ;
        RECT 3368.740 1446.690 3368.880 1641.190 ;
        RECT 3368.680 1446.370 3368.940 1446.690 ;
        RECT 3376.960 1446.370 3377.220 1446.690 ;
        RECT 3377.020 1444.555 3377.160 1446.370 ;
        RECT 3377.020 1444.485 3379.435 1444.555 ;
        RECT 3376.560 1444.345 3379.435 1444.485 ;
        RECT 3376.560 1425.690 3376.700 1444.345 ;
        RECT 3377.035 1444.275 3379.435 1444.345 ;
        RECT 3376.560 1425.550 3377.160 1425.690 ;
        RECT 3377.020 1422.935 3377.160 1425.550 ;
        RECT 3377.020 1422.655 3379.435 1422.935 ;
        RECT 211.700 1420.530 211.960 1420.850 ;
        RECT 3377.020 1420.510 3377.160 1422.655 ;
        RECT 3368.680 1420.190 3368.940 1420.510 ;
        RECT 3376.960 1420.190 3377.220 1420.510 ;
        RECT 211.700 1419.510 211.960 1419.830 ;
        RECT 211.760 1376.730 211.900 1419.510 ;
        RECT 209.000 1376.590 211.900 1376.730 ;
        RECT 209.000 1376.345 209.140 1376.590 ;
        RECT 208.565 1376.065 210.965 1376.345 ;
        RECT 208.565 1354.655 210.965 1354.725 ;
        RECT 211.300 1354.655 211.440 1376.590 ;
        RECT 208.565 1354.515 211.440 1354.655 ;
        RECT 208.565 1354.445 210.965 1354.515 ;
        RECT 211.300 1324.870 211.440 1354.515 ;
        RECT 211.300 1324.730 211.900 1324.870 ;
        RECT 211.760 1162.530 211.900 1324.730 ;
        RECT 3368.740 1223.310 3368.880 1420.190 ;
        RECT 3368.680 1222.990 3368.940 1223.310 ;
        RECT 3376.960 1222.990 3377.220 1223.310 ;
        RECT 3377.020 1222.555 3377.160 1222.990 ;
        RECT 3377.020 1222.275 3379.435 1222.555 ;
        RECT 3377.020 1219.650 3377.160 1222.275 ;
        RECT 3376.560 1219.510 3377.160 1219.650 ;
        RECT 3376.560 1200.865 3376.700 1219.510 ;
        RECT 3377.035 1200.865 3379.435 1200.935 ;
        RECT 3376.560 1200.725 3379.435 1200.865 ;
        RECT 3377.020 1200.655 3379.435 1200.725 ;
        RECT 3377.020 1198.490 3377.160 1200.655 ;
        RECT 3368.680 1198.170 3368.940 1198.490 ;
        RECT 3376.960 1198.170 3377.220 1198.490 ;
        RECT 209.000 1162.390 211.900 1162.530 ;
        RECT 209.000 1160.345 209.140 1162.390 ;
        RECT 208.565 1160.065 210.965 1160.345 ;
        RECT 211.300 1139.410 211.440 1162.390 ;
        RECT 209.000 1139.270 211.440 1139.410 ;
        RECT 209.000 1138.730 209.140 1139.270 ;
        RECT 208.610 1138.725 209.140 1138.730 ;
        RECT 208.565 1138.445 210.965 1138.725 ;
        RECT 211.300 1131.670 211.440 1139.270 ;
        RECT 211.300 1131.530 211.900 1131.670 ;
        RECT 211.760 944.930 211.900 1131.530 ;
        RECT 3368.740 1002.310 3368.880 1198.170 ;
        RECT 3368.680 1001.990 3368.940 1002.310 ;
        RECT 3376.960 1001.990 3377.220 1002.310 ;
        RECT 3377.020 1001.555 3377.160 1001.990 ;
        RECT 3377.020 1001.275 3379.435 1001.555 ;
        RECT 3377.020 998.650 3377.160 1001.275 ;
        RECT 3376.560 998.510 3377.160 998.650 ;
        RECT 3376.560 979.865 3376.700 998.510 ;
        RECT 3377.035 979.865 3379.435 979.935 ;
        RECT 3376.560 979.725 3379.435 979.865 ;
        RECT 3377.020 979.655 3379.435 979.725 ;
        RECT 3377.020 979.190 3377.160 979.655 ;
        RECT 3368.680 978.870 3368.940 979.190 ;
        RECT 3376.960 978.870 3377.220 979.190 ;
        RECT 209.460 944.790 211.900 944.930 ;
        RECT 209.460 944.345 209.600 944.790 ;
        RECT 208.565 944.065 210.965 944.345 ;
        RECT 208.565 922.655 210.965 922.725 ;
        RECT 211.300 922.655 211.440 944.790 ;
        RECT 208.565 922.515 211.900 922.655 ;
        RECT 208.565 922.445 210.965 922.515 ;
        RECT 211.760 228.130 211.900 922.515 ;
        RECT 3368.740 781.650 3368.880 978.870 ;
        RECT 3368.680 781.330 3368.940 781.650 ;
        RECT 3376.960 781.330 3377.220 781.650 ;
        RECT 3377.020 781.050 3377.160 781.330 ;
        RECT 3376.560 780.910 3377.160 781.050 ;
        RECT 3376.560 758.870 3376.700 780.910 ;
        RECT 3377.020 780.555 3377.160 780.910 ;
        RECT 3377.020 780.300 3379.435 780.555 ;
        RECT 3377.035 780.275 3379.435 780.300 ;
        RECT 3369.140 758.550 3369.400 758.870 ;
        RECT 3376.500 758.865 3376.760 758.870 ;
        RECT 3377.035 758.865 3379.435 758.935 ;
        RECT 3376.500 758.725 3379.435 758.865 ;
        RECT 3376.500 758.550 3376.760 758.725 ;
        RECT 3377.035 758.655 3379.435 758.725 ;
        RECT 3369.200 559.290 3369.340 758.550 ;
        RECT 3376.560 758.310 3376.700 758.550 ;
        RECT 3369.140 558.970 3369.400 559.290 ;
        RECT 3376.960 558.970 3377.220 559.290 ;
        RECT 3377.020 558.555 3377.160 558.970 ;
        RECT 3377.020 558.485 3379.435 558.555 ;
        RECT 3376.560 558.345 3379.435 558.485 ;
        RECT 3376.560 536.930 3376.700 558.345 ;
        RECT 3377.035 558.275 3379.435 558.345 ;
        RECT 3377.035 536.930 3379.435 536.935 ;
        RECT 3376.560 536.850 3379.435 536.930 ;
        RECT 3368.220 536.530 3368.480 536.850 ;
        RECT 3376.500 536.790 3379.435 536.850 ;
        RECT 3376.500 536.530 3376.760 536.790 ;
        RECT 3377.035 536.655 3379.435 536.790 ;
        RECT 3368.280 234.930 3368.420 536.530 ;
        RECT 3376.560 536.375 3376.700 536.530 ;
        RECT 3368.220 234.610 3368.480 234.930 ;
        RECT 2637.280 234.270 2637.540 234.590 ;
        RECT 211.700 227.810 211.960 228.130 ;
        RECT 718.160 227.810 718.420 228.130 ;
        RECT 718.220 220.990 718.360 227.810 ;
        RECT 1815.260 221.350 1815.520 221.670 ;
        RECT 2067.800 221.350 2068.060 221.670 ;
        RECT 2089.420 221.350 2089.680 221.670 ;
        RECT 2341.500 221.350 2341.760 221.670 ;
        RECT 2363.120 221.350 2363.380 221.670 ;
        RECT 999.220 221.010 999.480 221.330 ;
        RECT 1519.480 221.010 1519.740 221.330 ;
        RECT 1541.100 221.010 1541.360 221.330 ;
        RECT 1793.640 221.010 1793.900 221.330 ;
        RECT 718.160 220.670 718.420 220.990 ;
        RECT 725.520 220.670 725.780 220.990 ;
        RECT 976.680 220.670 976.940 220.990 ;
        RECT 998.300 220.730 998.560 220.990 ;
        RECT 999.280 220.730 999.420 221.010 ;
        RECT 998.300 220.670 999.420 220.730 ;
        RECT 725.580 201.010 725.720 220.670 ;
        RECT 976.740 210.965 976.880 220.670 ;
        RECT 998.360 220.590 999.420 220.670 ;
        RECT 998.360 210.965 998.500 220.590 ;
        RECT 1519.540 210.965 1519.680 221.010 ;
        RECT 1541.160 210.965 1541.300 221.010 ;
        RECT 1793.700 210.965 1793.840 221.010 ;
        RECT 1815.320 210.965 1815.460 221.350 ;
        RECT 2067.860 210.965 2068.000 221.350 ;
        RECT 2089.480 210.965 2089.620 221.350 ;
        RECT 976.655 208.565 976.935 210.965 ;
        RECT 998.275 208.565 998.555 210.965 ;
        RECT 1519.540 209.030 1519.935 210.965 ;
        RECT 1541.160 209.030 1541.555 210.965 ;
        RECT 1519.655 208.565 1519.935 209.030 ;
        RECT 1541.275 208.565 1541.555 209.030 ;
        RECT 1793.655 208.565 1793.935 210.965 ;
        RECT 1815.275 208.565 1815.555 210.965 ;
        RECT 2067.655 209.100 2068.000 210.965 ;
        RECT 2089.275 209.100 2089.620 210.965 ;
        RECT 2341.560 210.965 2341.700 221.350 ;
        RECT 2363.180 210.965 2363.320 221.350 ;
        RECT 2637.340 220.990 2637.480 234.270 ;
        RECT 2615.660 220.670 2615.920 220.990 ;
        RECT 2637.280 220.670 2637.540 220.990 ;
        RECT 2615.720 210.965 2615.860 220.670 ;
        RECT 2637.340 210.965 2637.480 220.670 ;
        RECT 2067.655 208.565 2067.935 209.100 ;
        RECT 2089.275 208.565 2089.555 209.100 ;
        RECT 2341.560 209.030 2341.935 210.965 ;
        RECT 2363.180 209.030 2363.555 210.965 ;
        RECT 2341.655 208.565 2341.935 209.030 ;
        RECT 2363.275 208.565 2363.555 209.030 ;
        RECT 2615.655 208.565 2615.935 210.965 ;
        RECT 2637.275 208.565 2637.555 210.965 ;
        RECT 725.515 200.870 725.720 201.010 ;
        RECT 725.515 200.000 725.655 200.870 ;
        RECT 725.455 198.530 725.715 200.000 ;
    END
  END porb_h
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 708.335 190.155 709.065 200.000 ;
        RECT 708.335 189.855 709.365 190.155 ;
        RECT 708.335 189.555 709.100 189.855 ;
        RECT 709.365 189.555 709.830 189.855 ;
        RECT 708.335 189.090 709.830 189.555 ;
        RECT 709.100 185.230 709.830 189.090 ;
    END
  END resetb_core_h
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 468.035 181.615 663.965 185.065 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 143.265 964.910 143.595 ;
    END
  END vssa
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 158.370 664.270 158.415 ;
        RECT 467.730 153.810 664.345 158.370 ;
        RECT 467.730 153.765 664.270 153.810 ;
    END
  END vssd
  PIN mprj_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3159.720 4988.000 3184.720 5070.350 ;
    END
  END mprj_analog[1]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3142.050 5093.120 3202.890 5153.945 ;
    END
  END mprj_io[15]
  PIN mprj_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2653.720 4988.000 2678.720 5070.350 ;
    END
  END mprj_analog[2]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2636.050 5093.120 2696.890 5153.945 ;
    END
  END mprj_io[16]
  PIN mprj_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2395.720 4988.000 2420.720 5070.350 ;
    END
  END mprj_analog[3]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2378.050 5093.120 2438.890 5153.945 ;
    END
  END mprj_io[17]
  PIN mprj_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2148.720 4988.000 2173.720 5070.350 ;
    END
  END mprj_analog[4]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2131.050 5093.120 2191.890 5153.945 ;
    END
  END mprj_io[18]
  PIN mprj_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3388.000 4673.000 3403.685 4744.610 ;
    END
  END mprj_analog[0]
  PIN mprj_clamp_high[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3388.000 4720.710 3413.660 4744.610 ;
    END
  END mprj_clamp_high[0]
  PIN mprj_clamp_low[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3388.000 4770.605 3390.055 4794.505 ;
    END
  END mprj_clamp_low[0]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4727.110 3553.945 4787.950 ;
    END
  END mprj_io[14]
  PIN vccd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 4467.330 3557.165 4521.730 ;
    END
  END vccd1_pad
  PIN vdda1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4026.110 3553.945 4086.950 ;
    END
  END vdda1_pad
  PIN vdda1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2482.110 3553.945 2542.950 ;
    END
  END vdda1_pad2
  PIN vssa1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1_pad
  PIN vssa1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2049.110 3553.945 2109.950 ;
    END
  END vssa1_pad2
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3396.885 2115.730 3401.535 2259.270 ;
    END
  END vccd1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 2116.035 3406.385 2258.965 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3444.405 2115.730 3444.735 2723.910 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 2308.500 3429.600 2332.500 ;
    END
  END vssd1
  PIN vssd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 2268.330 3557.165 2322.730 ;
    END
  END vssd1_pad
  PIN mprj_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 879.720 4988.000 904.720 5070.350 ;
    END
  END mprj_analog[7]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 862.050 5093.120 922.890 5153.945 ;
    END
  END mprj_io[21]
  PIN mprj_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 639.720 4988.000 664.720 5070.350 ;
    END
  END mprj_analog[8]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 622.050 5093.120 682.890 5153.945 ;
    END
  END mprj_io[22]
  PIN mprj_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.720 4988.000 424.720 5070.350 ;
    END
  END mprj_analog[9]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 382.050 5093.120 442.890 5153.945 ;
    END
  END mprj_io[23]
  PIN mprj_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.650 4800.720 200.000 4825.720 ;
    END
  END mprj_analog[10]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4783.050 94.880 4843.890 ;
    END
  END mprj_io[24]
  PIN mprj_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1454.390 4988.000 1526.000 5003.685 ;
    END
  END mprj_analog[5]
  PIN mprj_clamp_high[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.390 4988.000 1478.290 5013.660 ;
    END
  END mprj_clamp_high[1]
  PIN mprj_clamp_low[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.495 4988.000 1428.395 4990.055 ;
    END
  END mprj_clamp_low[1]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1411.050 5093.120 1471.890 5153.945 ;
    END
  END mprj_io[19]
  PIN mprj_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1197.390 4988.000 1269.000 5003.685 ;
    END
  END mprj_analog[6]
  PIN mprj_clamp_high[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.390 4988.000 1221.290 5013.660 ;
    END
  END mprj_clamp_high[2]
  PIN mprj_clamp_low[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.495 4988.000 1171.395 4990.055 ;
    END
  END mprj_clamp_low[2]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1154.050 5093.120 1214.890 5153.945 ;
    END
  END mprj_io[20]
  PIN vccd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 4575.270 98.100 4629.670 ;
    END
  END vccd2_pad
  PIN vdda2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 2424.050 94.880 2484.890 ;
    END
  END vdda2_pad
  PIN vssa2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4149.050 94.880 4209.890 ;
    END
  END vssa2_pad
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 192.515 2279.730 197.965 2418.270 ;
    END
  END vccd
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 2279.730 191.115 2418.270 ;
    END
  END vccd2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2280.035 185.065 2417.965 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 164.665 2279.730 168.115 2418.270 ;
    END
  END vddio
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 2037.090 143.595 2631.610 ;
    END
  END vssa2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.400 2206.500 198.000 2230.500 ;
    END
  END vssd2
  PIN vssd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 2216.270 98.100 2270.670 ;
    END
  END vssd2_pad
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.035 2281.000 24.215 2282.465 ;
        RECT 0.000 2279.730 24.215 2281.000 ;
    END
  END vssio
  OBS
      LAYER pwell ;
        RECT 1150.495 4988.935 1158.285 5011.790 ;
      LAYER nwell ;
        RECT 1158.860 4988.685 1217.965 4990.205 ;
      LAYER pwell ;
        RECT 1407.495 4988.935 1415.285 5011.790 ;
      LAYER nwell ;
        RECT 1415.860 4988.685 1474.965 4990.205 ;
        RECT 1708.860 4988.685 1767.965 4990.205 ;
        RECT 2889.860 4988.685 2948.965 4990.205 ;
      LAYER pwell ;
        RECT 3388.935 4783.715 3411.790 4791.505 ;
      LAYER nwell ;
        RECT 3388.685 4724.035 3390.205 4783.140 ;
        RECT 197.795 4365.860 199.315 4424.965 ;
      LAYER pwell ;
        RECT 176.210 4357.495 199.065 4365.285 ;
      LAYER nwell ;
        RECT 3393.665 4311.890 3397.325 4315.415 ;
        RECT 3444.590 4314.285 3469.235 4315.715 ;
        RECT 3476.485 4315.120 3480.400 4315.415 ;
        RECT 3407.155 4250.170 3411.080 4310.420 ;
        RECT 3444.590 4291.485 3446.020 4314.285 ;
        RECT 3448.180 4311.190 3450.340 4314.285 ;
        RECT 3448.180 4304.540 3449.020 4311.190 ;
        RECT 3448.770 4301.465 3449.020 4304.540 ;
        RECT 3467.805 4290.185 3469.235 4314.285 ;
        RECT 3473.580 4312.205 3480.400 4315.120 ;
        RECT 3473.580 4310.470 3479.820 4312.205 ;
        RECT 3474.660 4309.025 3479.820 4310.470 ;
      LAYER pwell ;
        RECT 3480.935 4309.785 3518.355 4315.215 ;
      LAYER nwell ;
        RECT 3474.660 4306.580 3476.280 4309.025 ;
        RECT 3474.660 4306.505 3475.740 4306.580 ;
      LAYER pwell ;
        RECT 3480.935 4305.700 3484.255 4309.785 ;
        RECT 3482.955 4275.615 3484.255 4305.700 ;
        RECT 3489.965 4309.265 3518.355 4309.785 ;
        RECT 3489.965 4275.615 3491.550 4309.265 ;
        RECT 3482.955 4269.160 3485.985 4275.615 ;
        RECT 3482.955 4268.410 3483.260 4269.160 ;
      LAYER nwell ;
        RECT 3422.265 4256.725 3424.055 4266.085 ;
        RECT 3420.410 4250.170 3424.055 4256.725 ;
        RECT 3407.155 4234.550 3413.345 4250.170 ;
        RECT 3417.785 4234.550 3424.055 4250.170 ;
        RECT 3460.595 4252.350 3461.265 4268.060 ;
        RECT 3438.620 4235.875 3440.050 4244.665 ;
        RECT 3453.195 4235.875 3454.045 4244.665 ;
        RECT 3460.595 4235.875 3461.775 4252.350 ;
        RECT 3438.620 4235.760 3461.775 4235.875 ;
        RECT 3471.165 4235.760 3472.345 4268.060 ;
        RECT 3482.245 4252.350 3483.165 4268.060 ;
        RECT 3481.735 4235.760 3483.165 4252.350 ;
        RECT 3438.620 4234.330 3483.165 4235.760 ;
      LAYER pwell ;
        RECT 3483.975 4238.230 3485.985 4269.160 ;
        RECT 3488.820 4262.120 3491.550 4275.615 ;
        RECT 3487.520 4238.230 3491.550 4262.120 ;
        RECT 3483.975 4237.135 3491.550 4238.230 ;
        RECT 3513.135 4274.755 3518.355 4309.265 ;
        RECT 3513.135 4248.090 3517.315 4274.755 ;
      LAYER nwell ;
        RECT 3518.665 4268.960 3528.380 4315.415 ;
      LAYER pwell ;
        RECT 3513.135 4237.135 3518.355 4248.090 ;
        RECT 3483.975 4234.710 3518.355 4237.135 ;
      LAYER nwell ;
        RECT 3518.665 4234.560 3528.385 4268.960 ;
      LAYER pwell ;
        RECT 3528.685 4234.710 3532.565 4315.290 ;
      LAYER nwell ;
        RECT 3532.880 4308.615 3566.975 4315.415 ;
        RECT 3532.880 4236.370 3534.690 4308.615 ;
        RECT 3556.515 4307.485 3566.975 4308.615 ;
        RECT 3556.515 4248.030 3558.475 4307.485 ;
        RECT 3561.545 4248.030 3566.975 4307.485 ;
        RECT 3556.515 4236.370 3566.975 4248.030 ;
        RECT 3532.880 4234.565 3566.975 4236.370 ;
        RECT 3532.880 4234.560 3558.230 4234.565 ;
        RECT 197.795 4153.860 199.315 4212.965 ;
      LAYER pwell ;
        RECT 3388.935 4082.715 3411.790 4090.505 ;
      LAYER nwell ;
        RECT 3388.685 4023.035 3390.205 4082.140 ;
        RECT 29.770 4006.435 55.120 4006.440 ;
        RECT 21.025 4004.630 55.120 4006.435 ;
        RECT 21.025 3992.970 31.485 4004.630 ;
        RECT 21.025 3933.515 26.455 3992.970 ;
        RECT 29.525 3933.515 31.485 3992.970 ;
        RECT 21.025 3932.385 31.485 3933.515 ;
        RECT 53.310 3932.385 55.120 4004.630 ;
        RECT 21.025 3925.585 55.120 3932.385 ;
      LAYER pwell ;
        RECT 55.435 3925.710 59.315 4006.290 ;
      LAYER nwell ;
        RECT 59.615 3972.040 69.335 4006.440 ;
      LAYER pwell ;
        RECT 69.645 4003.865 104.025 4006.290 ;
        RECT 69.645 3992.910 74.865 4003.865 ;
      LAYER nwell ;
        RECT 59.620 3925.585 69.335 3972.040 ;
      LAYER pwell ;
        RECT 70.685 3966.245 74.865 3992.910 ;
        RECT 69.645 3931.735 74.865 3966.245 ;
        RECT 96.450 4002.770 104.025 4003.865 ;
        RECT 96.450 3978.880 100.480 4002.770 ;
        RECT 96.450 3965.385 99.180 3978.880 ;
        RECT 102.015 3971.840 104.025 4002.770 ;
      LAYER nwell ;
        RECT 104.835 4005.240 149.380 4006.670 ;
        RECT 104.835 3988.650 106.265 4005.240 ;
        RECT 104.835 3972.940 105.755 3988.650 ;
        RECT 115.655 3972.940 116.835 4005.240 ;
        RECT 126.225 4005.125 149.380 4005.240 ;
        RECT 126.225 3988.650 127.405 4005.125 ;
        RECT 133.955 3996.335 134.805 4005.125 ;
        RECT 147.950 3996.335 149.380 4005.125 ;
        RECT 126.735 3972.940 127.405 3988.650 ;
        RECT 163.945 3990.830 170.215 4006.450 ;
        RECT 174.655 3990.830 180.845 4006.450 ;
        RECT 163.945 3984.275 167.590 3990.830 ;
        RECT 163.945 3974.915 165.735 3984.275 ;
      LAYER pwell ;
        RECT 104.740 3971.840 105.045 3972.590 ;
        RECT 102.015 3965.385 105.045 3971.840 ;
        RECT 96.450 3931.735 98.035 3965.385 ;
        RECT 69.645 3931.215 98.035 3931.735 ;
        RECT 103.745 3935.300 105.045 3965.385 ;
        RECT 103.745 3931.215 107.065 3935.300 ;
      LAYER nwell ;
        RECT 112.260 3934.420 113.340 3934.495 ;
        RECT 111.720 3931.975 113.340 3934.420 ;
      LAYER pwell ;
        RECT 69.645 3925.785 107.065 3931.215 ;
      LAYER nwell ;
        RECT 108.180 3930.530 113.340 3931.975 ;
        RECT 108.180 3928.795 114.420 3930.530 ;
        RECT 107.600 3925.880 114.420 3928.795 ;
        RECT 118.765 3926.715 120.195 3950.815 ;
        RECT 138.980 3936.460 139.230 3939.535 ;
        RECT 138.980 3929.810 139.820 3936.460 ;
        RECT 137.660 3926.715 139.820 3929.810 ;
        RECT 141.980 3926.715 143.410 3949.515 ;
        RECT 176.920 3930.580 180.845 3990.830 ;
        RECT 107.600 3925.585 111.515 3925.880 ;
        RECT 118.765 3925.285 143.410 3926.715 ;
        RECT 190.675 3925.585 194.335 3929.110 ;
        RECT 3393.665 3874.890 3397.325 3878.415 ;
        RECT 3444.590 3877.285 3469.235 3878.715 ;
        RECT 3476.485 3878.120 3480.400 3878.415 ;
        RECT 3407.155 3813.170 3411.080 3873.420 ;
        RECT 3444.590 3854.485 3446.020 3877.285 ;
        RECT 3448.180 3874.190 3450.340 3877.285 ;
        RECT 3448.180 3867.540 3449.020 3874.190 ;
        RECT 3448.770 3864.465 3449.020 3867.540 ;
        RECT 3467.805 3853.185 3469.235 3877.285 ;
        RECT 3473.580 3875.205 3480.400 3878.120 ;
        RECT 3473.580 3873.470 3479.820 3875.205 ;
        RECT 3474.660 3872.025 3479.820 3873.470 ;
      LAYER pwell ;
        RECT 3480.935 3872.785 3518.355 3878.215 ;
      LAYER nwell ;
        RECT 3474.660 3869.580 3476.280 3872.025 ;
        RECT 3474.660 3869.505 3475.740 3869.580 ;
      LAYER pwell ;
        RECT 3480.935 3868.700 3484.255 3872.785 ;
        RECT 3482.955 3838.615 3484.255 3868.700 ;
        RECT 3489.965 3872.265 3518.355 3872.785 ;
        RECT 3489.965 3838.615 3491.550 3872.265 ;
        RECT 3482.955 3832.160 3485.985 3838.615 ;
        RECT 3482.955 3831.410 3483.260 3832.160 ;
      LAYER nwell ;
        RECT 3422.265 3819.725 3424.055 3829.085 ;
        RECT 3420.410 3813.170 3424.055 3819.725 ;
        RECT 3407.155 3797.550 3413.345 3813.170 ;
        RECT 3417.785 3797.550 3424.055 3813.170 ;
        RECT 3460.595 3815.350 3461.265 3831.060 ;
        RECT 3438.620 3798.875 3440.050 3807.665 ;
        RECT 3453.195 3798.875 3454.045 3807.665 ;
        RECT 3460.595 3798.875 3461.775 3815.350 ;
        RECT 3438.620 3798.760 3461.775 3798.875 ;
        RECT 3471.165 3798.760 3472.345 3831.060 ;
        RECT 3482.245 3815.350 3483.165 3831.060 ;
        RECT 3481.735 3798.760 3483.165 3815.350 ;
        RECT 3438.620 3797.330 3483.165 3798.760 ;
      LAYER pwell ;
        RECT 3483.975 3801.230 3485.985 3832.160 ;
        RECT 3488.820 3825.120 3491.550 3838.615 ;
        RECT 3487.520 3801.230 3491.550 3825.120 ;
        RECT 3483.975 3800.135 3491.550 3801.230 ;
        RECT 3513.135 3837.755 3518.355 3872.265 ;
        RECT 3513.135 3811.090 3517.315 3837.755 ;
      LAYER nwell ;
        RECT 3518.665 3831.960 3528.380 3878.415 ;
      LAYER pwell ;
        RECT 3513.135 3800.135 3518.355 3811.090 ;
        RECT 3483.975 3797.710 3518.355 3800.135 ;
      LAYER nwell ;
        RECT 3518.665 3797.560 3528.385 3831.960 ;
      LAYER pwell ;
        RECT 3528.685 3797.710 3532.565 3878.290 ;
      LAYER nwell ;
        RECT 3532.880 3871.615 3566.975 3878.415 ;
        RECT 3532.880 3799.370 3534.690 3871.615 ;
        RECT 3556.515 3870.485 3566.975 3871.615 ;
        RECT 3556.515 3811.030 3558.475 3870.485 ;
        RECT 3561.545 3811.030 3566.975 3870.485 ;
        RECT 3556.515 3799.370 3566.975 3811.030 ;
        RECT 3532.880 3797.565 3566.975 3799.370 ;
        RECT 3532.880 3797.560 3558.230 3797.565 ;
        RECT 29.770 3790.435 55.120 3790.440 ;
        RECT 21.025 3788.630 55.120 3790.435 ;
        RECT 21.025 3776.970 31.485 3788.630 ;
        RECT 21.025 3717.515 26.455 3776.970 ;
        RECT 29.525 3717.515 31.485 3776.970 ;
        RECT 21.025 3716.385 31.485 3717.515 ;
        RECT 53.310 3716.385 55.120 3788.630 ;
        RECT 21.025 3709.585 55.120 3716.385 ;
      LAYER pwell ;
        RECT 55.435 3709.710 59.315 3790.290 ;
      LAYER nwell ;
        RECT 59.615 3756.040 69.335 3790.440 ;
      LAYER pwell ;
        RECT 69.645 3787.865 104.025 3790.290 ;
        RECT 69.645 3776.910 74.865 3787.865 ;
      LAYER nwell ;
        RECT 59.620 3709.585 69.335 3756.040 ;
      LAYER pwell ;
        RECT 70.685 3750.245 74.865 3776.910 ;
        RECT 69.645 3715.735 74.865 3750.245 ;
        RECT 96.450 3786.770 104.025 3787.865 ;
        RECT 96.450 3762.880 100.480 3786.770 ;
        RECT 96.450 3749.385 99.180 3762.880 ;
        RECT 102.015 3755.840 104.025 3786.770 ;
      LAYER nwell ;
        RECT 104.835 3789.240 149.380 3790.670 ;
        RECT 104.835 3772.650 106.265 3789.240 ;
        RECT 104.835 3756.940 105.755 3772.650 ;
        RECT 115.655 3756.940 116.835 3789.240 ;
        RECT 126.225 3789.125 149.380 3789.240 ;
        RECT 126.225 3772.650 127.405 3789.125 ;
        RECT 133.955 3780.335 134.805 3789.125 ;
        RECT 147.950 3780.335 149.380 3789.125 ;
        RECT 126.735 3756.940 127.405 3772.650 ;
        RECT 163.945 3774.830 170.215 3790.450 ;
        RECT 174.655 3774.830 180.845 3790.450 ;
        RECT 163.945 3768.275 167.590 3774.830 ;
        RECT 163.945 3758.915 165.735 3768.275 ;
      LAYER pwell ;
        RECT 104.740 3755.840 105.045 3756.590 ;
        RECT 102.015 3749.385 105.045 3755.840 ;
        RECT 96.450 3715.735 98.035 3749.385 ;
        RECT 69.645 3715.215 98.035 3715.735 ;
        RECT 103.745 3719.300 105.045 3749.385 ;
        RECT 103.745 3715.215 107.065 3719.300 ;
      LAYER nwell ;
        RECT 112.260 3718.420 113.340 3718.495 ;
        RECT 111.720 3715.975 113.340 3718.420 ;
      LAYER pwell ;
        RECT 69.645 3709.785 107.065 3715.215 ;
      LAYER nwell ;
        RECT 108.180 3714.530 113.340 3715.975 ;
        RECT 108.180 3712.795 114.420 3714.530 ;
        RECT 107.600 3709.880 114.420 3712.795 ;
        RECT 118.765 3710.715 120.195 3734.815 ;
        RECT 138.980 3720.460 139.230 3723.535 ;
        RECT 138.980 3713.810 139.820 3720.460 ;
        RECT 137.660 3710.715 139.820 3713.810 ;
        RECT 141.980 3710.715 143.410 3733.515 ;
        RECT 176.920 3714.580 180.845 3774.830 ;
        RECT 107.600 3709.585 111.515 3709.880 ;
        RECT 118.765 3709.285 143.410 3710.715 ;
        RECT 190.675 3709.585 194.335 3713.110 ;
        RECT 3393.665 3652.890 3397.325 3656.415 ;
        RECT 3444.590 3655.285 3469.235 3656.715 ;
        RECT 3476.485 3656.120 3480.400 3656.415 ;
        RECT 3407.155 3591.170 3411.080 3651.420 ;
        RECT 3444.590 3632.485 3446.020 3655.285 ;
        RECT 3448.180 3652.190 3450.340 3655.285 ;
        RECT 3448.180 3645.540 3449.020 3652.190 ;
        RECT 3448.770 3642.465 3449.020 3645.540 ;
        RECT 3467.805 3631.185 3469.235 3655.285 ;
        RECT 3473.580 3653.205 3480.400 3656.120 ;
        RECT 3473.580 3651.470 3479.820 3653.205 ;
        RECT 3474.660 3650.025 3479.820 3651.470 ;
      LAYER pwell ;
        RECT 3480.935 3650.785 3518.355 3656.215 ;
      LAYER nwell ;
        RECT 3474.660 3647.580 3476.280 3650.025 ;
        RECT 3474.660 3647.505 3475.740 3647.580 ;
      LAYER pwell ;
        RECT 3480.935 3646.700 3484.255 3650.785 ;
        RECT 3482.955 3616.615 3484.255 3646.700 ;
        RECT 3489.965 3650.265 3518.355 3650.785 ;
        RECT 3489.965 3616.615 3491.550 3650.265 ;
        RECT 3482.955 3610.160 3485.985 3616.615 ;
        RECT 3482.955 3609.410 3483.260 3610.160 ;
      LAYER nwell ;
        RECT 3422.265 3597.725 3424.055 3607.085 ;
        RECT 3420.410 3591.170 3424.055 3597.725 ;
        RECT 3407.155 3575.550 3413.345 3591.170 ;
        RECT 3417.785 3575.550 3424.055 3591.170 ;
        RECT 3460.595 3593.350 3461.265 3609.060 ;
        RECT 3438.620 3576.875 3440.050 3585.665 ;
        RECT 3453.195 3576.875 3454.045 3585.665 ;
        RECT 3460.595 3576.875 3461.775 3593.350 ;
        RECT 3438.620 3576.760 3461.775 3576.875 ;
        RECT 3471.165 3576.760 3472.345 3609.060 ;
        RECT 3482.245 3593.350 3483.165 3609.060 ;
        RECT 3481.735 3576.760 3483.165 3593.350 ;
        RECT 3438.620 3575.330 3483.165 3576.760 ;
      LAYER pwell ;
        RECT 3483.975 3579.230 3485.985 3610.160 ;
        RECT 3488.820 3603.120 3491.550 3616.615 ;
        RECT 3487.520 3579.230 3491.550 3603.120 ;
        RECT 3483.975 3578.135 3491.550 3579.230 ;
        RECT 3513.135 3615.755 3518.355 3650.265 ;
        RECT 3513.135 3589.090 3517.315 3615.755 ;
      LAYER nwell ;
        RECT 3518.665 3609.960 3528.380 3656.415 ;
      LAYER pwell ;
        RECT 3513.135 3578.135 3518.355 3589.090 ;
        RECT 3483.975 3575.710 3518.355 3578.135 ;
      LAYER nwell ;
        RECT 3518.665 3575.560 3528.385 3609.960 ;
      LAYER pwell ;
        RECT 3528.685 3575.710 3532.565 3656.290 ;
      LAYER nwell ;
        RECT 3532.880 3649.615 3566.975 3656.415 ;
        RECT 3532.880 3577.370 3534.690 3649.615 ;
        RECT 3556.515 3648.485 3566.975 3649.615 ;
        RECT 3556.515 3589.030 3558.475 3648.485 ;
        RECT 3561.545 3589.030 3566.975 3648.485 ;
        RECT 3556.515 3577.370 3566.975 3589.030 ;
        RECT 3532.880 3575.565 3566.975 3577.370 ;
        RECT 3532.880 3575.560 3558.230 3575.565 ;
        RECT 29.770 3574.435 55.120 3574.440 ;
        RECT 21.025 3572.630 55.120 3574.435 ;
        RECT 21.025 3560.970 31.485 3572.630 ;
        RECT 21.025 3501.515 26.455 3560.970 ;
        RECT 29.525 3501.515 31.485 3560.970 ;
        RECT 21.025 3500.385 31.485 3501.515 ;
        RECT 53.310 3500.385 55.120 3572.630 ;
        RECT 21.025 3493.585 55.120 3500.385 ;
      LAYER pwell ;
        RECT 55.435 3493.710 59.315 3574.290 ;
      LAYER nwell ;
        RECT 59.615 3540.040 69.335 3574.440 ;
      LAYER pwell ;
        RECT 69.645 3571.865 104.025 3574.290 ;
        RECT 69.645 3560.910 74.865 3571.865 ;
      LAYER nwell ;
        RECT 59.620 3493.585 69.335 3540.040 ;
      LAYER pwell ;
        RECT 70.685 3534.245 74.865 3560.910 ;
        RECT 69.645 3499.735 74.865 3534.245 ;
        RECT 96.450 3570.770 104.025 3571.865 ;
        RECT 96.450 3546.880 100.480 3570.770 ;
        RECT 96.450 3533.385 99.180 3546.880 ;
        RECT 102.015 3539.840 104.025 3570.770 ;
      LAYER nwell ;
        RECT 104.835 3573.240 149.380 3574.670 ;
        RECT 104.835 3556.650 106.265 3573.240 ;
        RECT 104.835 3540.940 105.755 3556.650 ;
        RECT 115.655 3540.940 116.835 3573.240 ;
        RECT 126.225 3573.125 149.380 3573.240 ;
        RECT 126.225 3556.650 127.405 3573.125 ;
        RECT 133.955 3564.335 134.805 3573.125 ;
        RECT 147.950 3564.335 149.380 3573.125 ;
        RECT 126.735 3540.940 127.405 3556.650 ;
        RECT 163.945 3558.830 170.215 3574.450 ;
        RECT 174.655 3558.830 180.845 3574.450 ;
        RECT 163.945 3552.275 167.590 3558.830 ;
        RECT 163.945 3542.915 165.735 3552.275 ;
      LAYER pwell ;
        RECT 104.740 3539.840 105.045 3540.590 ;
        RECT 102.015 3533.385 105.045 3539.840 ;
        RECT 96.450 3499.735 98.035 3533.385 ;
        RECT 69.645 3499.215 98.035 3499.735 ;
        RECT 103.745 3503.300 105.045 3533.385 ;
        RECT 103.745 3499.215 107.065 3503.300 ;
      LAYER nwell ;
        RECT 112.260 3502.420 113.340 3502.495 ;
        RECT 111.720 3499.975 113.340 3502.420 ;
      LAYER pwell ;
        RECT 69.645 3493.785 107.065 3499.215 ;
      LAYER nwell ;
        RECT 108.180 3498.530 113.340 3499.975 ;
        RECT 108.180 3496.795 114.420 3498.530 ;
        RECT 107.600 3493.880 114.420 3496.795 ;
        RECT 118.765 3494.715 120.195 3518.815 ;
        RECT 138.980 3504.460 139.230 3507.535 ;
        RECT 138.980 3497.810 139.820 3504.460 ;
        RECT 137.660 3494.715 139.820 3497.810 ;
        RECT 141.980 3494.715 143.410 3517.515 ;
        RECT 176.920 3498.580 180.845 3558.830 ;
        RECT 107.600 3493.585 111.515 3493.880 ;
        RECT 118.765 3493.285 143.410 3494.715 ;
        RECT 190.675 3493.585 194.335 3497.110 ;
        RECT 3393.665 3431.890 3397.325 3435.415 ;
        RECT 3444.590 3434.285 3469.235 3435.715 ;
        RECT 3476.485 3435.120 3480.400 3435.415 ;
        RECT 3407.155 3370.170 3411.080 3430.420 ;
        RECT 3444.590 3411.485 3446.020 3434.285 ;
        RECT 3448.180 3431.190 3450.340 3434.285 ;
        RECT 3448.180 3424.540 3449.020 3431.190 ;
        RECT 3448.770 3421.465 3449.020 3424.540 ;
        RECT 3467.805 3410.185 3469.235 3434.285 ;
        RECT 3473.580 3432.205 3480.400 3435.120 ;
        RECT 3473.580 3430.470 3479.820 3432.205 ;
        RECT 3474.660 3429.025 3479.820 3430.470 ;
      LAYER pwell ;
        RECT 3480.935 3429.785 3518.355 3435.215 ;
      LAYER nwell ;
        RECT 3474.660 3426.580 3476.280 3429.025 ;
        RECT 3474.660 3426.505 3475.740 3426.580 ;
      LAYER pwell ;
        RECT 3480.935 3425.700 3484.255 3429.785 ;
        RECT 3482.955 3395.615 3484.255 3425.700 ;
        RECT 3489.965 3429.265 3518.355 3429.785 ;
        RECT 3489.965 3395.615 3491.550 3429.265 ;
        RECT 3482.955 3389.160 3485.985 3395.615 ;
        RECT 3482.955 3388.410 3483.260 3389.160 ;
      LAYER nwell ;
        RECT 3422.265 3376.725 3424.055 3386.085 ;
        RECT 3420.410 3370.170 3424.055 3376.725 ;
        RECT 29.770 3357.435 55.120 3357.440 ;
        RECT 21.025 3355.630 55.120 3357.435 ;
        RECT 21.025 3343.970 31.485 3355.630 ;
        RECT 21.025 3284.515 26.455 3343.970 ;
        RECT 29.525 3284.515 31.485 3343.970 ;
        RECT 21.025 3283.385 31.485 3284.515 ;
        RECT 53.310 3283.385 55.120 3355.630 ;
        RECT 21.025 3276.585 55.120 3283.385 ;
      LAYER pwell ;
        RECT 55.435 3276.710 59.315 3357.290 ;
      LAYER nwell ;
        RECT 59.615 3323.040 69.335 3357.440 ;
      LAYER pwell ;
        RECT 69.645 3354.865 104.025 3357.290 ;
        RECT 69.645 3343.910 74.865 3354.865 ;
      LAYER nwell ;
        RECT 59.620 3276.585 69.335 3323.040 ;
      LAYER pwell ;
        RECT 70.685 3317.245 74.865 3343.910 ;
        RECT 69.645 3282.735 74.865 3317.245 ;
        RECT 96.450 3353.770 104.025 3354.865 ;
        RECT 96.450 3329.880 100.480 3353.770 ;
        RECT 96.450 3316.385 99.180 3329.880 ;
        RECT 102.015 3322.840 104.025 3353.770 ;
      LAYER nwell ;
        RECT 104.835 3356.240 149.380 3357.670 ;
        RECT 104.835 3339.650 106.265 3356.240 ;
        RECT 104.835 3323.940 105.755 3339.650 ;
        RECT 115.655 3323.940 116.835 3356.240 ;
        RECT 126.225 3356.125 149.380 3356.240 ;
        RECT 126.225 3339.650 127.405 3356.125 ;
        RECT 133.955 3347.335 134.805 3356.125 ;
        RECT 147.950 3347.335 149.380 3356.125 ;
        RECT 126.735 3323.940 127.405 3339.650 ;
        RECT 163.945 3341.830 170.215 3357.450 ;
        RECT 174.655 3341.830 180.845 3357.450 ;
        RECT 3407.155 3354.550 3413.345 3370.170 ;
        RECT 3417.785 3354.550 3424.055 3370.170 ;
        RECT 3460.595 3372.350 3461.265 3388.060 ;
        RECT 3438.620 3355.875 3440.050 3364.665 ;
        RECT 3453.195 3355.875 3454.045 3364.665 ;
        RECT 3460.595 3355.875 3461.775 3372.350 ;
        RECT 3438.620 3355.760 3461.775 3355.875 ;
        RECT 3471.165 3355.760 3472.345 3388.060 ;
        RECT 3482.245 3372.350 3483.165 3388.060 ;
        RECT 3481.735 3355.760 3483.165 3372.350 ;
        RECT 3438.620 3354.330 3483.165 3355.760 ;
      LAYER pwell ;
        RECT 3483.975 3358.230 3485.985 3389.160 ;
        RECT 3488.820 3382.120 3491.550 3395.615 ;
        RECT 3487.520 3358.230 3491.550 3382.120 ;
        RECT 3483.975 3357.135 3491.550 3358.230 ;
        RECT 3513.135 3394.755 3518.355 3429.265 ;
        RECT 3513.135 3368.090 3517.315 3394.755 ;
      LAYER nwell ;
        RECT 3518.665 3388.960 3528.380 3435.415 ;
      LAYER pwell ;
        RECT 3513.135 3357.135 3518.355 3368.090 ;
        RECT 3483.975 3354.710 3518.355 3357.135 ;
      LAYER nwell ;
        RECT 3518.665 3354.560 3528.385 3388.960 ;
      LAYER pwell ;
        RECT 3528.685 3354.710 3532.565 3435.290 ;
      LAYER nwell ;
        RECT 3532.880 3428.615 3566.975 3435.415 ;
        RECT 3532.880 3356.370 3534.690 3428.615 ;
        RECT 3556.515 3427.485 3566.975 3428.615 ;
        RECT 3556.515 3368.030 3558.475 3427.485 ;
        RECT 3561.545 3368.030 3566.975 3427.485 ;
        RECT 3556.515 3356.370 3566.975 3368.030 ;
        RECT 3532.880 3354.565 3566.975 3356.370 ;
        RECT 3532.880 3354.560 3558.230 3354.565 ;
        RECT 163.945 3335.275 167.590 3341.830 ;
        RECT 163.945 3325.915 165.735 3335.275 ;
      LAYER pwell ;
        RECT 104.740 3322.840 105.045 3323.590 ;
        RECT 102.015 3316.385 105.045 3322.840 ;
        RECT 96.450 3282.735 98.035 3316.385 ;
        RECT 69.645 3282.215 98.035 3282.735 ;
        RECT 103.745 3286.300 105.045 3316.385 ;
        RECT 103.745 3282.215 107.065 3286.300 ;
      LAYER nwell ;
        RECT 112.260 3285.420 113.340 3285.495 ;
        RECT 111.720 3282.975 113.340 3285.420 ;
      LAYER pwell ;
        RECT 69.645 3276.785 107.065 3282.215 ;
      LAYER nwell ;
        RECT 108.180 3281.530 113.340 3282.975 ;
        RECT 108.180 3279.795 114.420 3281.530 ;
        RECT 107.600 3276.880 114.420 3279.795 ;
        RECT 118.765 3277.715 120.195 3301.815 ;
        RECT 138.980 3287.460 139.230 3290.535 ;
        RECT 138.980 3280.810 139.820 3287.460 ;
        RECT 137.660 3277.715 139.820 3280.810 ;
        RECT 141.980 3277.715 143.410 3300.515 ;
        RECT 176.920 3281.580 180.845 3341.830 ;
        RECT 107.600 3276.585 111.515 3276.880 ;
        RECT 118.765 3276.285 143.410 3277.715 ;
        RECT 190.675 3276.585 194.335 3280.110 ;
        RECT 3393.665 3210.890 3397.325 3214.415 ;
        RECT 3444.590 3213.285 3469.235 3214.715 ;
        RECT 3476.485 3214.120 3480.400 3214.415 ;
        RECT 3407.155 3149.170 3411.080 3209.420 ;
        RECT 3444.590 3190.485 3446.020 3213.285 ;
        RECT 3448.180 3210.190 3450.340 3213.285 ;
        RECT 3448.180 3203.540 3449.020 3210.190 ;
        RECT 3448.770 3200.465 3449.020 3203.540 ;
        RECT 3467.805 3189.185 3469.235 3213.285 ;
        RECT 3473.580 3211.205 3480.400 3214.120 ;
        RECT 3473.580 3209.470 3479.820 3211.205 ;
        RECT 3474.660 3208.025 3479.820 3209.470 ;
      LAYER pwell ;
        RECT 3480.935 3208.785 3518.355 3214.215 ;
      LAYER nwell ;
        RECT 3474.660 3205.580 3476.280 3208.025 ;
        RECT 3474.660 3205.505 3475.740 3205.580 ;
      LAYER pwell ;
        RECT 3480.935 3204.700 3484.255 3208.785 ;
        RECT 3482.955 3174.615 3484.255 3204.700 ;
        RECT 3489.965 3208.265 3518.355 3208.785 ;
        RECT 3489.965 3174.615 3491.550 3208.265 ;
        RECT 3482.955 3168.160 3485.985 3174.615 ;
        RECT 3482.955 3167.410 3483.260 3168.160 ;
      LAYER nwell ;
        RECT 3422.265 3155.725 3424.055 3165.085 ;
        RECT 3420.410 3149.170 3424.055 3155.725 ;
        RECT 29.770 3141.435 55.120 3141.440 ;
        RECT 21.025 3139.630 55.120 3141.435 ;
        RECT 21.025 3127.970 31.485 3139.630 ;
        RECT 21.025 3068.515 26.455 3127.970 ;
        RECT 29.525 3068.515 31.485 3127.970 ;
        RECT 21.025 3067.385 31.485 3068.515 ;
        RECT 53.310 3067.385 55.120 3139.630 ;
        RECT 21.025 3060.585 55.120 3067.385 ;
      LAYER pwell ;
        RECT 55.435 3060.710 59.315 3141.290 ;
      LAYER nwell ;
        RECT 59.615 3107.040 69.335 3141.440 ;
      LAYER pwell ;
        RECT 69.645 3138.865 104.025 3141.290 ;
        RECT 69.645 3127.910 74.865 3138.865 ;
      LAYER nwell ;
        RECT 59.620 3060.585 69.335 3107.040 ;
      LAYER pwell ;
        RECT 70.685 3101.245 74.865 3127.910 ;
        RECT 69.645 3066.735 74.865 3101.245 ;
        RECT 96.450 3137.770 104.025 3138.865 ;
        RECT 96.450 3113.880 100.480 3137.770 ;
        RECT 96.450 3100.385 99.180 3113.880 ;
        RECT 102.015 3106.840 104.025 3137.770 ;
      LAYER nwell ;
        RECT 104.835 3140.240 149.380 3141.670 ;
        RECT 104.835 3123.650 106.265 3140.240 ;
        RECT 104.835 3107.940 105.755 3123.650 ;
        RECT 115.655 3107.940 116.835 3140.240 ;
        RECT 126.225 3140.125 149.380 3140.240 ;
        RECT 126.225 3123.650 127.405 3140.125 ;
        RECT 133.955 3131.335 134.805 3140.125 ;
        RECT 147.950 3131.335 149.380 3140.125 ;
        RECT 126.735 3107.940 127.405 3123.650 ;
        RECT 163.945 3125.830 170.215 3141.450 ;
        RECT 174.655 3125.830 180.845 3141.450 ;
        RECT 3407.155 3133.550 3413.345 3149.170 ;
        RECT 3417.785 3133.550 3424.055 3149.170 ;
        RECT 3460.595 3151.350 3461.265 3167.060 ;
        RECT 3438.620 3134.875 3440.050 3143.665 ;
        RECT 3453.195 3134.875 3454.045 3143.665 ;
        RECT 3460.595 3134.875 3461.775 3151.350 ;
        RECT 3438.620 3134.760 3461.775 3134.875 ;
        RECT 3471.165 3134.760 3472.345 3167.060 ;
        RECT 3482.245 3151.350 3483.165 3167.060 ;
        RECT 3481.735 3134.760 3483.165 3151.350 ;
        RECT 3438.620 3133.330 3483.165 3134.760 ;
      LAYER pwell ;
        RECT 3483.975 3137.230 3485.985 3168.160 ;
        RECT 3488.820 3161.120 3491.550 3174.615 ;
        RECT 3487.520 3137.230 3491.550 3161.120 ;
        RECT 3483.975 3136.135 3491.550 3137.230 ;
        RECT 3513.135 3173.755 3518.355 3208.265 ;
        RECT 3513.135 3147.090 3517.315 3173.755 ;
      LAYER nwell ;
        RECT 3518.665 3167.960 3528.380 3214.415 ;
      LAYER pwell ;
        RECT 3513.135 3136.135 3518.355 3147.090 ;
        RECT 3483.975 3133.710 3518.355 3136.135 ;
      LAYER nwell ;
        RECT 3518.665 3133.560 3528.385 3167.960 ;
      LAYER pwell ;
        RECT 3528.685 3133.710 3532.565 3214.290 ;
      LAYER nwell ;
        RECT 3532.880 3207.615 3566.975 3214.415 ;
        RECT 3532.880 3135.370 3534.690 3207.615 ;
        RECT 3556.515 3206.485 3566.975 3207.615 ;
        RECT 3556.515 3147.030 3558.475 3206.485 ;
        RECT 3561.545 3147.030 3566.975 3206.485 ;
        RECT 3556.515 3135.370 3566.975 3147.030 ;
        RECT 3532.880 3133.565 3566.975 3135.370 ;
        RECT 3532.880 3133.560 3558.230 3133.565 ;
        RECT 163.945 3119.275 167.590 3125.830 ;
        RECT 163.945 3109.915 165.735 3119.275 ;
      LAYER pwell ;
        RECT 104.740 3106.840 105.045 3107.590 ;
        RECT 102.015 3100.385 105.045 3106.840 ;
        RECT 96.450 3066.735 98.035 3100.385 ;
        RECT 69.645 3066.215 98.035 3066.735 ;
        RECT 103.745 3070.300 105.045 3100.385 ;
        RECT 103.745 3066.215 107.065 3070.300 ;
      LAYER nwell ;
        RECT 112.260 3069.420 113.340 3069.495 ;
        RECT 111.720 3066.975 113.340 3069.420 ;
      LAYER pwell ;
        RECT 69.645 3060.785 107.065 3066.215 ;
      LAYER nwell ;
        RECT 108.180 3065.530 113.340 3066.975 ;
        RECT 108.180 3063.795 114.420 3065.530 ;
        RECT 107.600 3060.880 114.420 3063.795 ;
        RECT 118.765 3061.715 120.195 3085.815 ;
        RECT 138.980 3071.460 139.230 3074.535 ;
        RECT 138.980 3064.810 139.820 3071.460 ;
        RECT 137.660 3061.715 139.820 3064.810 ;
        RECT 141.980 3061.715 143.410 3084.515 ;
        RECT 176.920 3065.580 180.845 3125.830 ;
        RECT 107.600 3060.585 111.515 3060.880 ;
        RECT 118.765 3060.285 143.410 3061.715 ;
        RECT 190.675 3060.585 194.335 3064.110 ;
        RECT 3393.665 2988.890 3397.325 2992.415 ;
        RECT 3444.590 2991.285 3469.235 2992.715 ;
        RECT 3476.485 2992.120 3480.400 2992.415 ;
        RECT 3407.155 2927.170 3411.080 2987.420 ;
        RECT 3444.590 2968.485 3446.020 2991.285 ;
        RECT 3448.180 2988.190 3450.340 2991.285 ;
        RECT 3448.180 2981.540 3449.020 2988.190 ;
        RECT 3448.770 2978.465 3449.020 2981.540 ;
        RECT 3467.805 2967.185 3469.235 2991.285 ;
        RECT 3473.580 2989.205 3480.400 2992.120 ;
        RECT 3473.580 2987.470 3479.820 2989.205 ;
        RECT 3474.660 2986.025 3479.820 2987.470 ;
      LAYER pwell ;
        RECT 3480.935 2986.785 3518.355 2992.215 ;
      LAYER nwell ;
        RECT 3474.660 2983.580 3476.280 2986.025 ;
        RECT 3474.660 2983.505 3475.740 2983.580 ;
      LAYER pwell ;
        RECT 3480.935 2982.700 3484.255 2986.785 ;
        RECT 3482.955 2952.615 3484.255 2982.700 ;
        RECT 3489.965 2986.265 3518.355 2986.785 ;
        RECT 3489.965 2952.615 3491.550 2986.265 ;
        RECT 3482.955 2946.160 3485.985 2952.615 ;
        RECT 3482.955 2945.410 3483.260 2946.160 ;
      LAYER nwell ;
        RECT 3422.265 2933.725 3424.055 2943.085 ;
        RECT 3420.410 2927.170 3424.055 2933.725 ;
        RECT 29.770 2925.435 55.120 2925.440 ;
        RECT 21.025 2923.630 55.120 2925.435 ;
        RECT 21.025 2911.970 31.485 2923.630 ;
        RECT 21.025 2852.515 26.455 2911.970 ;
        RECT 29.525 2852.515 31.485 2911.970 ;
        RECT 21.025 2851.385 31.485 2852.515 ;
        RECT 53.310 2851.385 55.120 2923.630 ;
        RECT 21.025 2844.585 55.120 2851.385 ;
      LAYER pwell ;
        RECT 55.435 2844.710 59.315 2925.290 ;
      LAYER nwell ;
        RECT 59.615 2891.040 69.335 2925.440 ;
      LAYER pwell ;
        RECT 69.645 2922.865 104.025 2925.290 ;
        RECT 69.645 2911.910 74.865 2922.865 ;
      LAYER nwell ;
        RECT 59.620 2844.585 69.335 2891.040 ;
      LAYER pwell ;
        RECT 70.685 2885.245 74.865 2911.910 ;
        RECT 69.645 2850.735 74.865 2885.245 ;
        RECT 96.450 2921.770 104.025 2922.865 ;
        RECT 96.450 2897.880 100.480 2921.770 ;
        RECT 96.450 2884.385 99.180 2897.880 ;
        RECT 102.015 2890.840 104.025 2921.770 ;
      LAYER nwell ;
        RECT 104.835 2924.240 149.380 2925.670 ;
        RECT 104.835 2907.650 106.265 2924.240 ;
        RECT 104.835 2891.940 105.755 2907.650 ;
        RECT 115.655 2891.940 116.835 2924.240 ;
        RECT 126.225 2924.125 149.380 2924.240 ;
        RECT 126.225 2907.650 127.405 2924.125 ;
        RECT 133.955 2915.335 134.805 2924.125 ;
        RECT 147.950 2915.335 149.380 2924.125 ;
        RECT 126.735 2891.940 127.405 2907.650 ;
        RECT 163.945 2909.830 170.215 2925.450 ;
        RECT 174.655 2909.830 180.845 2925.450 ;
        RECT 3407.155 2911.550 3413.345 2927.170 ;
        RECT 3417.785 2911.550 3424.055 2927.170 ;
        RECT 3460.595 2929.350 3461.265 2945.060 ;
        RECT 3438.620 2912.875 3440.050 2921.665 ;
        RECT 3453.195 2912.875 3454.045 2921.665 ;
        RECT 3460.595 2912.875 3461.775 2929.350 ;
        RECT 3438.620 2912.760 3461.775 2912.875 ;
        RECT 3471.165 2912.760 3472.345 2945.060 ;
        RECT 3482.245 2929.350 3483.165 2945.060 ;
        RECT 3481.735 2912.760 3483.165 2929.350 ;
        RECT 3438.620 2911.330 3483.165 2912.760 ;
      LAYER pwell ;
        RECT 3483.975 2915.230 3485.985 2946.160 ;
        RECT 3488.820 2939.120 3491.550 2952.615 ;
        RECT 3487.520 2915.230 3491.550 2939.120 ;
        RECT 3483.975 2914.135 3491.550 2915.230 ;
        RECT 3513.135 2951.755 3518.355 2986.265 ;
        RECT 3513.135 2925.090 3517.315 2951.755 ;
      LAYER nwell ;
        RECT 3518.665 2945.960 3528.380 2992.415 ;
      LAYER pwell ;
        RECT 3513.135 2914.135 3518.355 2925.090 ;
        RECT 3483.975 2911.710 3518.355 2914.135 ;
      LAYER nwell ;
        RECT 3518.665 2911.560 3528.385 2945.960 ;
      LAYER pwell ;
        RECT 3528.685 2911.710 3532.565 2992.290 ;
      LAYER nwell ;
        RECT 3532.880 2985.615 3566.975 2992.415 ;
        RECT 3532.880 2913.370 3534.690 2985.615 ;
        RECT 3556.515 2984.485 3566.975 2985.615 ;
        RECT 3556.515 2925.030 3558.475 2984.485 ;
        RECT 3561.545 2925.030 3566.975 2984.485 ;
        RECT 3556.515 2913.370 3566.975 2925.030 ;
        RECT 3532.880 2911.565 3566.975 2913.370 ;
        RECT 3532.880 2911.560 3558.230 2911.565 ;
        RECT 163.945 2903.275 167.590 2909.830 ;
        RECT 163.945 2893.915 165.735 2903.275 ;
      LAYER pwell ;
        RECT 104.740 2890.840 105.045 2891.590 ;
        RECT 102.015 2884.385 105.045 2890.840 ;
        RECT 96.450 2850.735 98.035 2884.385 ;
        RECT 69.645 2850.215 98.035 2850.735 ;
        RECT 103.745 2854.300 105.045 2884.385 ;
        RECT 103.745 2850.215 107.065 2854.300 ;
      LAYER nwell ;
        RECT 112.260 2853.420 113.340 2853.495 ;
        RECT 111.720 2850.975 113.340 2853.420 ;
      LAYER pwell ;
        RECT 69.645 2844.785 107.065 2850.215 ;
      LAYER nwell ;
        RECT 108.180 2849.530 113.340 2850.975 ;
        RECT 108.180 2847.795 114.420 2849.530 ;
        RECT 107.600 2844.880 114.420 2847.795 ;
        RECT 118.765 2845.715 120.195 2869.815 ;
        RECT 138.980 2855.460 139.230 2858.535 ;
        RECT 138.980 2848.810 139.820 2855.460 ;
        RECT 137.660 2845.715 139.820 2848.810 ;
        RECT 141.980 2845.715 143.410 2868.515 ;
        RECT 176.920 2849.580 180.845 2909.830 ;
        RECT 107.600 2844.585 111.515 2844.880 ;
        RECT 118.765 2844.285 143.410 2845.715 ;
        RECT 190.675 2844.585 194.335 2848.110 ;
        RECT 3393.665 2767.890 3397.325 2771.415 ;
        RECT 3444.590 2770.285 3469.235 2771.715 ;
        RECT 3476.485 2771.120 3480.400 2771.415 ;
        RECT 29.770 2709.435 55.120 2709.440 ;
        RECT 21.025 2707.630 55.120 2709.435 ;
        RECT 21.025 2695.970 31.485 2707.630 ;
        RECT 21.025 2636.515 26.455 2695.970 ;
        RECT 29.525 2636.515 31.485 2695.970 ;
        RECT 21.025 2635.385 31.485 2636.515 ;
        RECT 53.310 2635.385 55.120 2707.630 ;
        RECT 21.025 2628.585 55.120 2635.385 ;
      LAYER pwell ;
        RECT 55.435 2628.710 59.315 2709.290 ;
      LAYER nwell ;
        RECT 59.615 2675.040 69.335 2709.440 ;
      LAYER pwell ;
        RECT 69.645 2706.865 104.025 2709.290 ;
        RECT 69.645 2695.910 74.865 2706.865 ;
      LAYER nwell ;
        RECT 59.620 2628.585 69.335 2675.040 ;
      LAYER pwell ;
        RECT 70.685 2669.245 74.865 2695.910 ;
        RECT 69.645 2634.735 74.865 2669.245 ;
        RECT 96.450 2705.770 104.025 2706.865 ;
        RECT 96.450 2681.880 100.480 2705.770 ;
        RECT 96.450 2668.385 99.180 2681.880 ;
        RECT 102.015 2674.840 104.025 2705.770 ;
      LAYER nwell ;
        RECT 104.835 2708.240 149.380 2709.670 ;
        RECT 104.835 2691.650 106.265 2708.240 ;
        RECT 104.835 2675.940 105.755 2691.650 ;
        RECT 115.655 2675.940 116.835 2708.240 ;
        RECT 126.225 2708.125 149.380 2708.240 ;
        RECT 126.225 2691.650 127.405 2708.125 ;
        RECT 133.955 2699.335 134.805 2708.125 ;
        RECT 147.950 2699.335 149.380 2708.125 ;
        RECT 126.735 2675.940 127.405 2691.650 ;
        RECT 163.945 2693.830 170.215 2709.450 ;
        RECT 174.655 2693.830 180.845 2709.450 ;
        RECT 163.945 2687.275 167.590 2693.830 ;
        RECT 163.945 2677.915 165.735 2687.275 ;
      LAYER pwell ;
        RECT 104.740 2674.840 105.045 2675.590 ;
        RECT 102.015 2668.385 105.045 2674.840 ;
        RECT 96.450 2634.735 98.035 2668.385 ;
        RECT 69.645 2634.215 98.035 2634.735 ;
        RECT 103.745 2638.300 105.045 2668.385 ;
        RECT 103.745 2634.215 107.065 2638.300 ;
      LAYER nwell ;
        RECT 112.260 2637.420 113.340 2637.495 ;
        RECT 111.720 2634.975 113.340 2637.420 ;
      LAYER pwell ;
        RECT 69.645 2628.785 107.065 2634.215 ;
      LAYER nwell ;
        RECT 108.180 2633.530 113.340 2634.975 ;
        RECT 108.180 2631.795 114.420 2633.530 ;
        RECT 107.600 2628.880 114.420 2631.795 ;
        RECT 118.765 2629.715 120.195 2653.815 ;
        RECT 138.980 2639.460 139.230 2642.535 ;
        RECT 138.980 2632.810 139.820 2639.460 ;
        RECT 137.660 2629.715 139.820 2632.810 ;
        RECT 141.980 2629.715 143.410 2652.515 ;
        RECT 176.920 2633.580 180.845 2693.830 ;
        RECT 3407.155 2706.170 3411.080 2766.420 ;
        RECT 3444.590 2747.485 3446.020 2770.285 ;
        RECT 3448.180 2767.190 3450.340 2770.285 ;
        RECT 3448.180 2760.540 3449.020 2767.190 ;
        RECT 3448.770 2757.465 3449.020 2760.540 ;
        RECT 3467.805 2746.185 3469.235 2770.285 ;
        RECT 3473.580 2768.205 3480.400 2771.120 ;
        RECT 3473.580 2766.470 3479.820 2768.205 ;
        RECT 3474.660 2765.025 3479.820 2766.470 ;
      LAYER pwell ;
        RECT 3480.935 2765.785 3518.355 2771.215 ;
      LAYER nwell ;
        RECT 3474.660 2762.580 3476.280 2765.025 ;
        RECT 3474.660 2762.505 3475.740 2762.580 ;
      LAYER pwell ;
        RECT 3480.935 2761.700 3484.255 2765.785 ;
        RECT 3482.955 2731.615 3484.255 2761.700 ;
        RECT 3489.965 2765.265 3518.355 2765.785 ;
        RECT 3489.965 2731.615 3491.550 2765.265 ;
        RECT 3482.955 2725.160 3485.985 2731.615 ;
        RECT 3482.955 2724.410 3483.260 2725.160 ;
      LAYER nwell ;
        RECT 3422.265 2712.725 3424.055 2722.085 ;
        RECT 3420.410 2706.170 3424.055 2712.725 ;
        RECT 3407.155 2690.550 3413.345 2706.170 ;
        RECT 3417.785 2690.550 3424.055 2706.170 ;
        RECT 3460.595 2708.350 3461.265 2724.060 ;
        RECT 3438.620 2691.875 3440.050 2700.665 ;
        RECT 3453.195 2691.875 3454.045 2700.665 ;
        RECT 3460.595 2691.875 3461.775 2708.350 ;
        RECT 3438.620 2691.760 3461.775 2691.875 ;
        RECT 3471.165 2691.760 3472.345 2724.060 ;
        RECT 3482.245 2708.350 3483.165 2724.060 ;
        RECT 3481.735 2691.760 3483.165 2708.350 ;
        RECT 3438.620 2690.330 3483.165 2691.760 ;
      LAYER pwell ;
        RECT 3483.975 2694.230 3485.985 2725.160 ;
        RECT 3488.820 2718.120 3491.550 2731.615 ;
        RECT 3487.520 2694.230 3491.550 2718.120 ;
        RECT 3483.975 2693.135 3491.550 2694.230 ;
        RECT 3513.135 2730.755 3518.355 2765.265 ;
        RECT 3513.135 2704.090 3517.315 2730.755 ;
      LAYER nwell ;
        RECT 3518.665 2724.960 3528.380 2771.415 ;
      LAYER pwell ;
        RECT 3513.135 2693.135 3518.355 2704.090 ;
        RECT 3483.975 2690.710 3518.355 2693.135 ;
      LAYER nwell ;
        RECT 3518.665 2690.560 3528.385 2724.960 ;
      LAYER pwell ;
        RECT 3528.685 2690.710 3532.565 2771.290 ;
      LAYER nwell ;
        RECT 3532.880 2764.615 3566.975 2771.415 ;
        RECT 3532.880 2692.370 3534.690 2764.615 ;
        RECT 3556.515 2763.485 3566.975 2764.615 ;
        RECT 3556.515 2704.030 3558.475 2763.485 ;
        RECT 3561.545 2704.030 3566.975 2763.485 ;
        RECT 3556.515 2692.370 3566.975 2704.030 ;
        RECT 3532.880 2690.565 3566.975 2692.370 ;
        RECT 3532.880 2690.560 3558.230 2690.565 ;
        RECT 107.600 2628.585 111.515 2628.880 ;
        RECT 118.765 2628.285 143.410 2629.715 ;
        RECT 190.675 2628.585 194.335 2632.110 ;
      LAYER pwell ;
        RECT 3388.935 2538.715 3411.790 2546.505 ;
      LAYER nwell ;
        RECT 197.795 2428.860 199.315 2487.965 ;
        RECT 3388.685 2479.035 3390.205 2538.140 ;
      LAYER pwell ;
        RECT 176.210 2420.495 199.065 2428.285 ;
      LAYER nwell ;
        RECT 29.770 2070.435 55.120 2070.440 ;
        RECT 21.025 2068.630 55.120 2070.435 ;
        RECT 21.025 2056.970 31.485 2068.630 ;
        RECT 21.025 1997.515 26.455 2056.970 ;
        RECT 29.525 1997.515 31.485 2056.970 ;
        RECT 21.025 1996.385 31.485 1997.515 ;
        RECT 53.310 1996.385 55.120 2068.630 ;
        RECT 21.025 1989.585 55.120 1996.385 ;
      LAYER pwell ;
        RECT 55.435 1989.710 59.315 2070.290 ;
      LAYER nwell ;
        RECT 59.615 2036.040 69.335 2070.440 ;
      LAYER pwell ;
        RECT 69.645 2067.865 104.025 2070.290 ;
        RECT 69.645 2056.910 74.865 2067.865 ;
      LAYER nwell ;
        RECT 59.620 1989.585 69.335 2036.040 ;
      LAYER pwell ;
        RECT 70.685 2030.245 74.865 2056.910 ;
        RECT 69.645 1995.735 74.865 2030.245 ;
        RECT 96.450 2066.770 104.025 2067.865 ;
        RECT 96.450 2042.880 100.480 2066.770 ;
        RECT 96.450 2029.385 99.180 2042.880 ;
        RECT 102.015 2035.840 104.025 2066.770 ;
      LAYER nwell ;
        RECT 104.835 2069.240 149.380 2070.670 ;
        RECT 104.835 2052.650 106.265 2069.240 ;
        RECT 104.835 2036.940 105.755 2052.650 ;
        RECT 115.655 2036.940 116.835 2069.240 ;
        RECT 126.225 2069.125 149.380 2069.240 ;
        RECT 126.225 2052.650 127.405 2069.125 ;
        RECT 133.955 2060.335 134.805 2069.125 ;
        RECT 147.950 2060.335 149.380 2069.125 ;
        RECT 126.735 2036.940 127.405 2052.650 ;
        RECT 163.945 2054.830 170.215 2070.450 ;
        RECT 174.655 2054.830 180.845 2070.450 ;
        RECT 163.945 2048.275 167.590 2054.830 ;
        RECT 163.945 2038.915 165.735 2048.275 ;
      LAYER pwell ;
        RECT 104.740 2035.840 105.045 2036.590 ;
        RECT 102.015 2029.385 105.045 2035.840 ;
        RECT 96.450 1995.735 98.035 2029.385 ;
        RECT 69.645 1995.215 98.035 1995.735 ;
        RECT 103.745 1999.300 105.045 2029.385 ;
        RECT 103.745 1995.215 107.065 1999.300 ;
      LAYER nwell ;
        RECT 112.260 1998.420 113.340 1998.495 ;
        RECT 111.720 1995.975 113.340 1998.420 ;
      LAYER pwell ;
        RECT 69.645 1989.785 107.065 1995.215 ;
      LAYER nwell ;
        RECT 108.180 1994.530 113.340 1995.975 ;
        RECT 108.180 1992.795 114.420 1994.530 ;
        RECT 107.600 1989.880 114.420 1992.795 ;
        RECT 118.765 1990.715 120.195 2014.815 ;
        RECT 138.980 2000.460 139.230 2003.535 ;
        RECT 138.980 1993.810 139.820 2000.460 ;
        RECT 137.660 1990.715 139.820 1993.810 ;
        RECT 141.980 1990.715 143.410 2013.515 ;
        RECT 176.920 1994.580 180.845 2054.830 ;
        RECT 3388.685 2046.035 3390.205 2105.140 ;
        RECT 107.600 1989.585 111.515 1989.880 ;
        RECT 118.765 1989.285 143.410 1990.715 ;
        RECT 190.675 1989.585 194.335 1993.110 ;
        RECT 3393.665 1896.890 3397.325 1900.415 ;
        RECT 3444.590 1899.285 3469.235 1900.715 ;
        RECT 3476.485 1900.120 3480.400 1900.415 ;
        RECT 29.770 1854.435 55.120 1854.440 ;
        RECT 21.025 1852.630 55.120 1854.435 ;
        RECT 21.025 1840.970 31.485 1852.630 ;
        RECT 21.025 1781.515 26.455 1840.970 ;
        RECT 29.525 1781.515 31.485 1840.970 ;
        RECT 21.025 1780.385 31.485 1781.515 ;
        RECT 53.310 1780.385 55.120 1852.630 ;
        RECT 21.025 1773.585 55.120 1780.385 ;
      LAYER pwell ;
        RECT 55.435 1773.710 59.315 1854.290 ;
      LAYER nwell ;
        RECT 59.615 1820.040 69.335 1854.440 ;
      LAYER pwell ;
        RECT 69.645 1851.865 104.025 1854.290 ;
        RECT 69.645 1840.910 74.865 1851.865 ;
      LAYER nwell ;
        RECT 59.620 1773.585 69.335 1820.040 ;
      LAYER pwell ;
        RECT 70.685 1814.245 74.865 1840.910 ;
        RECT 69.645 1779.735 74.865 1814.245 ;
        RECT 96.450 1850.770 104.025 1851.865 ;
        RECT 96.450 1826.880 100.480 1850.770 ;
        RECT 96.450 1813.385 99.180 1826.880 ;
        RECT 102.015 1819.840 104.025 1850.770 ;
      LAYER nwell ;
        RECT 104.835 1853.240 149.380 1854.670 ;
        RECT 104.835 1836.650 106.265 1853.240 ;
        RECT 104.835 1820.940 105.755 1836.650 ;
        RECT 115.655 1820.940 116.835 1853.240 ;
        RECT 126.225 1853.125 149.380 1853.240 ;
        RECT 126.225 1836.650 127.405 1853.125 ;
        RECT 133.955 1844.335 134.805 1853.125 ;
        RECT 147.950 1844.335 149.380 1853.125 ;
        RECT 126.735 1820.940 127.405 1836.650 ;
        RECT 163.945 1838.830 170.215 1854.450 ;
        RECT 174.655 1838.830 180.845 1854.450 ;
        RECT 163.945 1832.275 167.590 1838.830 ;
        RECT 163.945 1822.915 165.735 1832.275 ;
      LAYER pwell ;
        RECT 104.740 1819.840 105.045 1820.590 ;
        RECT 102.015 1813.385 105.045 1819.840 ;
        RECT 96.450 1779.735 98.035 1813.385 ;
        RECT 69.645 1779.215 98.035 1779.735 ;
        RECT 103.745 1783.300 105.045 1813.385 ;
        RECT 103.745 1779.215 107.065 1783.300 ;
      LAYER nwell ;
        RECT 112.260 1782.420 113.340 1782.495 ;
        RECT 111.720 1779.975 113.340 1782.420 ;
      LAYER pwell ;
        RECT 69.645 1773.785 107.065 1779.215 ;
      LAYER nwell ;
        RECT 108.180 1778.530 113.340 1779.975 ;
        RECT 108.180 1776.795 114.420 1778.530 ;
        RECT 107.600 1773.880 114.420 1776.795 ;
        RECT 118.765 1774.715 120.195 1798.815 ;
        RECT 138.980 1784.460 139.230 1787.535 ;
        RECT 138.980 1777.810 139.820 1784.460 ;
        RECT 137.660 1774.715 139.820 1777.810 ;
        RECT 141.980 1774.715 143.410 1797.515 ;
        RECT 176.920 1778.580 180.845 1838.830 ;
        RECT 3407.155 1835.170 3411.080 1895.420 ;
        RECT 3444.590 1876.485 3446.020 1899.285 ;
        RECT 3448.180 1896.190 3450.340 1899.285 ;
        RECT 3448.180 1889.540 3449.020 1896.190 ;
        RECT 3448.770 1886.465 3449.020 1889.540 ;
        RECT 3467.805 1875.185 3469.235 1899.285 ;
        RECT 3473.580 1897.205 3480.400 1900.120 ;
        RECT 3473.580 1895.470 3479.820 1897.205 ;
        RECT 3474.660 1894.025 3479.820 1895.470 ;
      LAYER pwell ;
        RECT 3480.935 1894.785 3518.355 1900.215 ;
      LAYER nwell ;
        RECT 3474.660 1891.580 3476.280 1894.025 ;
        RECT 3474.660 1891.505 3475.740 1891.580 ;
      LAYER pwell ;
        RECT 3480.935 1890.700 3484.255 1894.785 ;
        RECT 3482.955 1860.615 3484.255 1890.700 ;
        RECT 3489.965 1894.265 3518.355 1894.785 ;
        RECT 3489.965 1860.615 3491.550 1894.265 ;
        RECT 3482.955 1854.160 3485.985 1860.615 ;
        RECT 3482.955 1853.410 3483.260 1854.160 ;
      LAYER nwell ;
        RECT 3422.265 1841.725 3424.055 1851.085 ;
        RECT 3420.410 1835.170 3424.055 1841.725 ;
        RECT 3407.155 1819.550 3413.345 1835.170 ;
        RECT 3417.785 1819.550 3424.055 1835.170 ;
        RECT 3460.595 1837.350 3461.265 1853.060 ;
        RECT 3438.620 1820.875 3440.050 1829.665 ;
        RECT 3453.195 1820.875 3454.045 1829.665 ;
        RECT 3460.595 1820.875 3461.775 1837.350 ;
        RECT 3438.620 1820.760 3461.775 1820.875 ;
        RECT 3471.165 1820.760 3472.345 1853.060 ;
        RECT 3482.245 1837.350 3483.165 1853.060 ;
        RECT 3481.735 1820.760 3483.165 1837.350 ;
        RECT 3438.620 1819.330 3483.165 1820.760 ;
      LAYER pwell ;
        RECT 3483.975 1823.230 3485.985 1854.160 ;
        RECT 3488.820 1847.120 3491.550 1860.615 ;
        RECT 3487.520 1823.230 3491.550 1847.120 ;
        RECT 3483.975 1822.135 3491.550 1823.230 ;
        RECT 3513.135 1859.755 3518.355 1894.265 ;
        RECT 3513.135 1833.090 3517.315 1859.755 ;
      LAYER nwell ;
        RECT 3518.665 1853.960 3528.380 1900.415 ;
      LAYER pwell ;
        RECT 3513.135 1822.135 3518.355 1833.090 ;
        RECT 3483.975 1819.710 3518.355 1822.135 ;
      LAYER nwell ;
        RECT 3518.665 1819.560 3528.385 1853.960 ;
      LAYER pwell ;
        RECT 3528.685 1819.710 3532.565 1900.290 ;
      LAYER nwell ;
        RECT 3532.880 1893.615 3566.975 1900.415 ;
        RECT 3532.880 1821.370 3534.690 1893.615 ;
        RECT 3556.515 1892.485 3566.975 1893.615 ;
        RECT 3556.515 1833.030 3558.475 1892.485 ;
        RECT 3561.545 1833.030 3566.975 1892.485 ;
        RECT 3556.515 1821.370 3566.975 1833.030 ;
        RECT 3532.880 1819.565 3566.975 1821.370 ;
        RECT 3532.880 1819.560 3558.230 1819.565 ;
        RECT 107.600 1773.585 111.515 1773.880 ;
        RECT 118.765 1773.285 143.410 1774.715 ;
        RECT 190.675 1773.585 194.335 1777.110 ;
        RECT 3393.665 1675.890 3397.325 1679.415 ;
        RECT 3444.590 1678.285 3469.235 1679.715 ;
        RECT 3476.485 1679.120 3480.400 1679.415 ;
        RECT 29.770 1637.435 55.120 1637.440 ;
        RECT 21.025 1635.630 55.120 1637.435 ;
        RECT 21.025 1623.970 31.485 1635.630 ;
        RECT 21.025 1564.515 26.455 1623.970 ;
        RECT 29.525 1564.515 31.485 1623.970 ;
        RECT 21.025 1563.385 31.485 1564.515 ;
        RECT 53.310 1563.385 55.120 1635.630 ;
        RECT 21.025 1556.585 55.120 1563.385 ;
      LAYER pwell ;
        RECT 55.435 1556.710 59.315 1637.290 ;
      LAYER nwell ;
        RECT 59.615 1603.040 69.335 1637.440 ;
      LAYER pwell ;
        RECT 69.645 1634.865 104.025 1637.290 ;
        RECT 69.645 1623.910 74.865 1634.865 ;
      LAYER nwell ;
        RECT 59.620 1556.585 69.335 1603.040 ;
      LAYER pwell ;
        RECT 70.685 1597.245 74.865 1623.910 ;
        RECT 69.645 1562.735 74.865 1597.245 ;
        RECT 96.450 1633.770 104.025 1634.865 ;
        RECT 96.450 1609.880 100.480 1633.770 ;
        RECT 96.450 1596.385 99.180 1609.880 ;
        RECT 102.015 1602.840 104.025 1633.770 ;
      LAYER nwell ;
        RECT 104.835 1636.240 149.380 1637.670 ;
        RECT 104.835 1619.650 106.265 1636.240 ;
        RECT 104.835 1603.940 105.755 1619.650 ;
        RECT 115.655 1603.940 116.835 1636.240 ;
        RECT 126.225 1636.125 149.380 1636.240 ;
        RECT 126.225 1619.650 127.405 1636.125 ;
        RECT 133.955 1627.335 134.805 1636.125 ;
        RECT 147.950 1627.335 149.380 1636.125 ;
        RECT 126.735 1603.940 127.405 1619.650 ;
        RECT 163.945 1621.830 170.215 1637.450 ;
        RECT 174.655 1621.830 180.845 1637.450 ;
        RECT 163.945 1615.275 167.590 1621.830 ;
        RECT 163.945 1605.915 165.735 1615.275 ;
      LAYER pwell ;
        RECT 104.740 1602.840 105.045 1603.590 ;
        RECT 102.015 1596.385 105.045 1602.840 ;
        RECT 96.450 1562.735 98.035 1596.385 ;
        RECT 69.645 1562.215 98.035 1562.735 ;
        RECT 103.745 1566.300 105.045 1596.385 ;
        RECT 103.745 1562.215 107.065 1566.300 ;
      LAYER nwell ;
        RECT 112.260 1565.420 113.340 1565.495 ;
        RECT 111.720 1562.975 113.340 1565.420 ;
      LAYER pwell ;
        RECT 69.645 1556.785 107.065 1562.215 ;
      LAYER nwell ;
        RECT 108.180 1561.530 113.340 1562.975 ;
        RECT 108.180 1559.795 114.420 1561.530 ;
        RECT 107.600 1556.880 114.420 1559.795 ;
        RECT 118.765 1557.715 120.195 1581.815 ;
        RECT 138.980 1567.460 139.230 1570.535 ;
        RECT 138.980 1560.810 139.820 1567.460 ;
        RECT 137.660 1557.715 139.820 1560.810 ;
        RECT 141.980 1557.715 143.410 1580.515 ;
        RECT 176.920 1561.580 180.845 1621.830 ;
        RECT 3407.155 1614.170 3411.080 1674.420 ;
        RECT 3444.590 1655.485 3446.020 1678.285 ;
        RECT 3448.180 1675.190 3450.340 1678.285 ;
        RECT 3448.180 1668.540 3449.020 1675.190 ;
        RECT 3448.770 1665.465 3449.020 1668.540 ;
        RECT 3467.805 1654.185 3469.235 1678.285 ;
        RECT 3473.580 1676.205 3480.400 1679.120 ;
        RECT 3473.580 1674.470 3479.820 1676.205 ;
        RECT 3474.660 1673.025 3479.820 1674.470 ;
      LAYER pwell ;
        RECT 3480.935 1673.785 3518.355 1679.215 ;
      LAYER nwell ;
        RECT 3474.660 1670.580 3476.280 1673.025 ;
        RECT 3474.660 1670.505 3475.740 1670.580 ;
      LAYER pwell ;
        RECT 3480.935 1669.700 3484.255 1673.785 ;
        RECT 3482.955 1639.615 3484.255 1669.700 ;
        RECT 3489.965 1673.265 3518.355 1673.785 ;
        RECT 3489.965 1639.615 3491.550 1673.265 ;
        RECT 3482.955 1633.160 3485.985 1639.615 ;
        RECT 3482.955 1632.410 3483.260 1633.160 ;
      LAYER nwell ;
        RECT 3422.265 1620.725 3424.055 1630.085 ;
        RECT 3420.410 1614.170 3424.055 1620.725 ;
        RECT 3407.155 1598.550 3413.345 1614.170 ;
        RECT 3417.785 1598.550 3424.055 1614.170 ;
        RECT 3460.595 1616.350 3461.265 1632.060 ;
        RECT 3438.620 1599.875 3440.050 1608.665 ;
        RECT 3453.195 1599.875 3454.045 1608.665 ;
        RECT 3460.595 1599.875 3461.775 1616.350 ;
        RECT 3438.620 1599.760 3461.775 1599.875 ;
        RECT 3471.165 1599.760 3472.345 1632.060 ;
        RECT 3482.245 1616.350 3483.165 1632.060 ;
        RECT 3481.735 1599.760 3483.165 1616.350 ;
        RECT 3438.620 1598.330 3483.165 1599.760 ;
      LAYER pwell ;
        RECT 3483.975 1602.230 3485.985 1633.160 ;
        RECT 3488.820 1626.120 3491.550 1639.615 ;
        RECT 3487.520 1602.230 3491.550 1626.120 ;
        RECT 3483.975 1601.135 3491.550 1602.230 ;
        RECT 3513.135 1638.755 3518.355 1673.265 ;
        RECT 3513.135 1612.090 3517.315 1638.755 ;
      LAYER nwell ;
        RECT 3518.665 1632.960 3528.380 1679.415 ;
      LAYER pwell ;
        RECT 3513.135 1601.135 3518.355 1612.090 ;
        RECT 3483.975 1598.710 3518.355 1601.135 ;
      LAYER nwell ;
        RECT 3518.665 1598.560 3528.385 1632.960 ;
      LAYER pwell ;
        RECT 3528.685 1598.710 3532.565 1679.290 ;
      LAYER nwell ;
        RECT 3532.880 1672.615 3566.975 1679.415 ;
        RECT 3532.880 1600.370 3534.690 1672.615 ;
        RECT 3556.515 1671.485 3566.975 1672.615 ;
        RECT 3556.515 1612.030 3558.475 1671.485 ;
        RECT 3561.545 1612.030 3566.975 1671.485 ;
        RECT 3556.515 1600.370 3566.975 1612.030 ;
        RECT 3532.880 1598.565 3566.975 1600.370 ;
        RECT 3532.880 1598.560 3558.230 1598.565 ;
        RECT 107.600 1556.585 111.515 1556.880 ;
        RECT 118.765 1556.285 143.410 1557.715 ;
        RECT 190.675 1556.585 194.335 1560.110 ;
        RECT 3393.665 1454.890 3397.325 1458.415 ;
        RECT 3444.590 1457.285 3469.235 1458.715 ;
        RECT 3476.485 1458.120 3480.400 1458.415 ;
        RECT 29.770 1421.435 55.120 1421.440 ;
        RECT 21.025 1419.630 55.120 1421.435 ;
        RECT 21.025 1407.970 31.485 1419.630 ;
        RECT 21.025 1348.515 26.455 1407.970 ;
        RECT 29.525 1348.515 31.485 1407.970 ;
        RECT 21.025 1347.385 31.485 1348.515 ;
        RECT 53.310 1347.385 55.120 1419.630 ;
        RECT 21.025 1340.585 55.120 1347.385 ;
      LAYER pwell ;
        RECT 55.435 1340.710 59.315 1421.290 ;
      LAYER nwell ;
        RECT 59.615 1387.040 69.335 1421.440 ;
      LAYER pwell ;
        RECT 69.645 1418.865 104.025 1421.290 ;
        RECT 69.645 1407.910 74.865 1418.865 ;
      LAYER nwell ;
        RECT 59.620 1340.585 69.335 1387.040 ;
      LAYER pwell ;
        RECT 70.685 1381.245 74.865 1407.910 ;
        RECT 69.645 1346.735 74.865 1381.245 ;
        RECT 96.450 1417.770 104.025 1418.865 ;
        RECT 96.450 1393.880 100.480 1417.770 ;
        RECT 96.450 1380.385 99.180 1393.880 ;
        RECT 102.015 1386.840 104.025 1417.770 ;
      LAYER nwell ;
        RECT 104.835 1420.240 149.380 1421.670 ;
        RECT 104.835 1403.650 106.265 1420.240 ;
        RECT 104.835 1387.940 105.755 1403.650 ;
        RECT 115.655 1387.940 116.835 1420.240 ;
        RECT 126.225 1420.125 149.380 1420.240 ;
        RECT 126.225 1403.650 127.405 1420.125 ;
        RECT 133.955 1411.335 134.805 1420.125 ;
        RECT 147.950 1411.335 149.380 1420.125 ;
        RECT 126.735 1387.940 127.405 1403.650 ;
        RECT 163.945 1405.830 170.215 1421.450 ;
        RECT 174.655 1405.830 180.845 1421.450 ;
        RECT 163.945 1399.275 167.590 1405.830 ;
        RECT 163.945 1389.915 165.735 1399.275 ;
      LAYER pwell ;
        RECT 104.740 1386.840 105.045 1387.590 ;
        RECT 102.015 1380.385 105.045 1386.840 ;
        RECT 96.450 1346.735 98.035 1380.385 ;
        RECT 69.645 1346.215 98.035 1346.735 ;
        RECT 103.745 1350.300 105.045 1380.385 ;
        RECT 103.745 1346.215 107.065 1350.300 ;
      LAYER nwell ;
        RECT 112.260 1349.420 113.340 1349.495 ;
        RECT 111.720 1346.975 113.340 1349.420 ;
      LAYER pwell ;
        RECT 69.645 1340.785 107.065 1346.215 ;
      LAYER nwell ;
        RECT 108.180 1345.530 113.340 1346.975 ;
        RECT 108.180 1343.795 114.420 1345.530 ;
        RECT 107.600 1340.880 114.420 1343.795 ;
        RECT 118.765 1341.715 120.195 1365.815 ;
        RECT 138.980 1351.460 139.230 1354.535 ;
        RECT 138.980 1344.810 139.820 1351.460 ;
        RECT 137.660 1341.715 139.820 1344.810 ;
        RECT 141.980 1341.715 143.410 1364.515 ;
        RECT 176.920 1345.580 180.845 1405.830 ;
        RECT 3407.155 1393.170 3411.080 1453.420 ;
        RECT 3444.590 1434.485 3446.020 1457.285 ;
        RECT 3448.180 1454.190 3450.340 1457.285 ;
        RECT 3448.180 1447.540 3449.020 1454.190 ;
        RECT 3448.770 1444.465 3449.020 1447.540 ;
        RECT 3467.805 1433.185 3469.235 1457.285 ;
        RECT 3473.580 1455.205 3480.400 1458.120 ;
        RECT 3473.580 1453.470 3479.820 1455.205 ;
        RECT 3474.660 1452.025 3479.820 1453.470 ;
      LAYER pwell ;
        RECT 3480.935 1452.785 3518.355 1458.215 ;
      LAYER nwell ;
        RECT 3474.660 1449.580 3476.280 1452.025 ;
        RECT 3474.660 1449.505 3475.740 1449.580 ;
      LAYER pwell ;
        RECT 3480.935 1448.700 3484.255 1452.785 ;
        RECT 3482.955 1418.615 3484.255 1448.700 ;
        RECT 3489.965 1452.265 3518.355 1452.785 ;
        RECT 3489.965 1418.615 3491.550 1452.265 ;
        RECT 3482.955 1412.160 3485.985 1418.615 ;
        RECT 3482.955 1411.410 3483.260 1412.160 ;
      LAYER nwell ;
        RECT 3422.265 1399.725 3424.055 1409.085 ;
        RECT 3420.410 1393.170 3424.055 1399.725 ;
        RECT 3407.155 1377.550 3413.345 1393.170 ;
        RECT 3417.785 1377.550 3424.055 1393.170 ;
        RECT 3460.595 1395.350 3461.265 1411.060 ;
        RECT 3438.620 1378.875 3440.050 1387.665 ;
        RECT 3453.195 1378.875 3454.045 1387.665 ;
        RECT 3460.595 1378.875 3461.775 1395.350 ;
        RECT 3438.620 1378.760 3461.775 1378.875 ;
        RECT 3471.165 1378.760 3472.345 1411.060 ;
        RECT 3482.245 1395.350 3483.165 1411.060 ;
        RECT 3481.735 1378.760 3483.165 1395.350 ;
        RECT 3438.620 1377.330 3483.165 1378.760 ;
      LAYER pwell ;
        RECT 3483.975 1381.230 3485.985 1412.160 ;
        RECT 3488.820 1405.120 3491.550 1418.615 ;
        RECT 3487.520 1381.230 3491.550 1405.120 ;
        RECT 3483.975 1380.135 3491.550 1381.230 ;
        RECT 3513.135 1417.755 3518.355 1452.265 ;
        RECT 3513.135 1391.090 3517.315 1417.755 ;
      LAYER nwell ;
        RECT 3518.665 1411.960 3528.380 1458.415 ;
      LAYER pwell ;
        RECT 3513.135 1380.135 3518.355 1391.090 ;
        RECT 3483.975 1377.710 3518.355 1380.135 ;
      LAYER nwell ;
        RECT 3518.665 1377.560 3528.385 1411.960 ;
      LAYER pwell ;
        RECT 3528.685 1377.710 3532.565 1458.290 ;
      LAYER nwell ;
        RECT 3532.880 1451.615 3566.975 1458.415 ;
        RECT 3532.880 1379.370 3534.690 1451.615 ;
        RECT 3556.515 1450.485 3566.975 1451.615 ;
        RECT 3556.515 1391.030 3558.475 1450.485 ;
        RECT 3561.545 1391.030 3566.975 1450.485 ;
        RECT 3556.515 1379.370 3566.975 1391.030 ;
        RECT 3532.880 1377.565 3566.975 1379.370 ;
        RECT 3532.880 1377.560 3558.230 1377.565 ;
        RECT 107.600 1340.585 111.515 1340.880 ;
        RECT 118.765 1340.285 143.410 1341.715 ;
        RECT 190.675 1340.585 194.335 1344.110 ;
        RECT 3393.665 1232.890 3397.325 1236.415 ;
        RECT 3444.590 1235.285 3469.235 1236.715 ;
        RECT 3476.485 1236.120 3480.400 1236.415 ;
        RECT 29.770 1205.435 55.120 1205.440 ;
        RECT 21.025 1203.630 55.120 1205.435 ;
        RECT 21.025 1191.970 31.485 1203.630 ;
        RECT 21.025 1132.515 26.455 1191.970 ;
        RECT 29.525 1132.515 31.485 1191.970 ;
        RECT 21.025 1131.385 31.485 1132.515 ;
        RECT 53.310 1131.385 55.120 1203.630 ;
        RECT 21.025 1124.585 55.120 1131.385 ;
      LAYER pwell ;
        RECT 55.435 1124.710 59.315 1205.290 ;
      LAYER nwell ;
        RECT 59.615 1171.040 69.335 1205.440 ;
      LAYER pwell ;
        RECT 69.645 1202.865 104.025 1205.290 ;
        RECT 69.645 1191.910 74.865 1202.865 ;
      LAYER nwell ;
        RECT 59.620 1124.585 69.335 1171.040 ;
      LAYER pwell ;
        RECT 70.685 1165.245 74.865 1191.910 ;
        RECT 69.645 1130.735 74.865 1165.245 ;
        RECT 96.450 1201.770 104.025 1202.865 ;
        RECT 96.450 1177.880 100.480 1201.770 ;
        RECT 96.450 1164.385 99.180 1177.880 ;
        RECT 102.015 1170.840 104.025 1201.770 ;
      LAYER nwell ;
        RECT 104.835 1204.240 149.380 1205.670 ;
        RECT 104.835 1187.650 106.265 1204.240 ;
        RECT 104.835 1171.940 105.755 1187.650 ;
        RECT 115.655 1171.940 116.835 1204.240 ;
        RECT 126.225 1204.125 149.380 1204.240 ;
        RECT 126.225 1187.650 127.405 1204.125 ;
        RECT 133.955 1195.335 134.805 1204.125 ;
        RECT 147.950 1195.335 149.380 1204.125 ;
        RECT 126.735 1171.940 127.405 1187.650 ;
        RECT 163.945 1189.830 170.215 1205.450 ;
        RECT 174.655 1189.830 180.845 1205.450 ;
        RECT 163.945 1183.275 167.590 1189.830 ;
        RECT 163.945 1173.915 165.735 1183.275 ;
      LAYER pwell ;
        RECT 104.740 1170.840 105.045 1171.590 ;
        RECT 102.015 1164.385 105.045 1170.840 ;
        RECT 96.450 1130.735 98.035 1164.385 ;
        RECT 69.645 1130.215 98.035 1130.735 ;
        RECT 103.745 1134.300 105.045 1164.385 ;
        RECT 103.745 1130.215 107.065 1134.300 ;
      LAYER nwell ;
        RECT 112.260 1133.420 113.340 1133.495 ;
        RECT 111.720 1130.975 113.340 1133.420 ;
      LAYER pwell ;
        RECT 69.645 1124.785 107.065 1130.215 ;
      LAYER nwell ;
        RECT 108.180 1129.530 113.340 1130.975 ;
        RECT 108.180 1127.795 114.420 1129.530 ;
        RECT 107.600 1124.880 114.420 1127.795 ;
        RECT 118.765 1125.715 120.195 1149.815 ;
        RECT 138.980 1135.460 139.230 1138.535 ;
        RECT 138.980 1128.810 139.820 1135.460 ;
        RECT 137.660 1125.715 139.820 1128.810 ;
        RECT 141.980 1125.715 143.410 1148.515 ;
        RECT 176.920 1129.580 180.845 1189.830 ;
        RECT 3407.155 1171.170 3411.080 1231.420 ;
        RECT 3444.590 1212.485 3446.020 1235.285 ;
        RECT 3448.180 1232.190 3450.340 1235.285 ;
        RECT 3448.180 1225.540 3449.020 1232.190 ;
        RECT 3448.770 1222.465 3449.020 1225.540 ;
        RECT 3467.805 1211.185 3469.235 1235.285 ;
        RECT 3473.580 1233.205 3480.400 1236.120 ;
        RECT 3473.580 1231.470 3479.820 1233.205 ;
        RECT 3474.660 1230.025 3479.820 1231.470 ;
      LAYER pwell ;
        RECT 3480.935 1230.785 3518.355 1236.215 ;
      LAYER nwell ;
        RECT 3474.660 1227.580 3476.280 1230.025 ;
        RECT 3474.660 1227.505 3475.740 1227.580 ;
      LAYER pwell ;
        RECT 3480.935 1226.700 3484.255 1230.785 ;
        RECT 3482.955 1196.615 3484.255 1226.700 ;
        RECT 3489.965 1230.265 3518.355 1230.785 ;
        RECT 3489.965 1196.615 3491.550 1230.265 ;
        RECT 3482.955 1190.160 3485.985 1196.615 ;
        RECT 3482.955 1189.410 3483.260 1190.160 ;
      LAYER nwell ;
        RECT 3422.265 1177.725 3424.055 1187.085 ;
        RECT 3420.410 1171.170 3424.055 1177.725 ;
        RECT 3407.155 1155.550 3413.345 1171.170 ;
        RECT 3417.785 1155.550 3424.055 1171.170 ;
        RECT 3460.595 1173.350 3461.265 1189.060 ;
        RECT 3438.620 1156.875 3440.050 1165.665 ;
        RECT 3453.195 1156.875 3454.045 1165.665 ;
        RECT 3460.595 1156.875 3461.775 1173.350 ;
        RECT 3438.620 1156.760 3461.775 1156.875 ;
        RECT 3471.165 1156.760 3472.345 1189.060 ;
        RECT 3482.245 1173.350 3483.165 1189.060 ;
        RECT 3481.735 1156.760 3483.165 1173.350 ;
        RECT 3438.620 1155.330 3483.165 1156.760 ;
      LAYER pwell ;
        RECT 3483.975 1159.230 3485.985 1190.160 ;
        RECT 3488.820 1183.120 3491.550 1196.615 ;
        RECT 3487.520 1159.230 3491.550 1183.120 ;
        RECT 3483.975 1158.135 3491.550 1159.230 ;
        RECT 3513.135 1195.755 3518.355 1230.265 ;
        RECT 3513.135 1169.090 3517.315 1195.755 ;
      LAYER nwell ;
        RECT 3518.665 1189.960 3528.380 1236.415 ;
      LAYER pwell ;
        RECT 3513.135 1158.135 3518.355 1169.090 ;
        RECT 3483.975 1155.710 3518.355 1158.135 ;
      LAYER nwell ;
        RECT 3518.665 1155.560 3528.385 1189.960 ;
      LAYER pwell ;
        RECT 3528.685 1155.710 3532.565 1236.290 ;
      LAYER nwell ;
        RECT 3532.880 1229.615 3566.975 1236.415 ;
        RECT 3532.880 1157.370 3534.690 1229.615 ;
        RECT 3556.515 1228.485 3566.975 1229.615 ;
        RECT 3556.515 1169.030 3558.475 1228.485 ;
        RECT 3561.545 1169.030 3566.975 1228.485 ;
        RECT 3556.515 1157.370 3566.975 1169.030 ;
        RECT 3532.880 1155.565 3566.975 1157.370 ;
        RECT 3532.880 1155.560 3558.230 1155.565 ;
        RECT 107.600 1124.585 111.515 1124.880 ;
        RECT 118.765 1124.285 143.410 1125.715 ;
        RECT 190.675 1124.585 194.335 1128.110 ;
        RECT 3393.665 1011.890 3397.325 1015.415 ;
        RECT 3444.590 1014.285 3469.235 1015.715 ;
        RECT 3476.485 1015.120 3480.400 1015.415 ;
        RECT 29.770 989.435 55.120 989.440 ;
        RECT 21.025 987.630 55.120 989.435 ;
        RECT 21.025 975.970 31.485 987.630 ;
        RECT 21.025 916.515 26.455 975.970 ;
        RECT 29.525 916.515 31.485 975.970 ;
        RECT 21.025 915.385 31.485 916.515 ;
        RECT 53.310 915.385 55.120 987.630 ;
        RECT 21.025 908.585 55.120 915.385 ;
      LAYER pwell ;
        RECT 55.435 908.710 59.315 989.290 ;
      LAYER nwell ;
        RECT 59.615 955.040 69.335 989.440 ;
      LAYER pwell ;
        RECT 69.645 986.865 104.025 989.290 ;
        RECT 69.645 975.910 74.865 986.865 ;
      LAYER nwell ;
        RECT 59.620 908.585 69.335 955.040 ;
      LAYER pwell ;
        RECT 70.685 949.245 74.865 975.910 ;
        RECT 69.645 914.735 74.865 949.245 ;
        RECT 96.450 985.770 104.025 986.865 ;
        RECT 96.450 961.880 100.480 985.770 ;
        RECT 96.450 948.385 99.180 961.880 ;
        RECT 102.015 954.840 104.025 985.770 ;
      LAYER nwell ;
        RECT 104.835 988.240 149.380 989.670 ;
        RECT 104.835 971.650 106.265 988.240 ;
        RECT 104.835 955.940 105.755 971.650 ;
        RECT 115.655 955.940 116.835 988.240 ;
        RECT 126.225 988.125 149.380 988.240 ;
        RECT 126.225 971.650 127.405 988.125 ;
        RECT 133.955 979.335 134.805 988.125 ;
        RECT 147.950 979.335 149.380 988.125 ;
        RECT 126.735 955.940 127.405 971.650 ;
        RECT 163.945 973.830 170.215 989.450 ;
        RECT 174.655 973.830 180.845 989.450 ;
        RECT 163.945 967.275 167.590 973.830 ;
        RECT 163.945 957.915 165.735 967.275 ;
      LAYER pwell ;
        RECT 104.740 954.840 105.045 955.590 ;
        RECT 102.015 948.385 105.045 954.840 ;
        RECT 96.450 914.735 98.035 948.385 ;
        RECT 69.645 914.215 98.035 914.735 ;
        RECT 103.745 918.300 105.045 948.385 ;
        RECT 103.745 914.215 107.065 918.300 ;
      LAYER nwell ;
        RECT 112.260 917.420 113.340 917.495 ;
        RECT 111.720 914.975 113.340 917.420 ;
      LAYER pwell ;
        RECT 69.645 908.785 107.065 914.215 ;
      LAYER nwell ;
        RECT 108.180 913.530 113.340 914.975 ;
        RECT 108.180 911.795 114.420 913.530 ;
        RECT 107.600 908.880 114.420 911.795 ;
        RECT 118.765 909.715 120.195 933.815 ;
        RECT 138.980 919.460 139.230 922.535 ;
        RECT 138.980 912.810 139.820 919.460 ;
        RECT 137.660 909.715 139.820 912.810 ;
        RECT 141.980 909.715 143.410 932.515 ;
        RECT 176.920 913.580 180.845 973.830 ;
        RECT 3407.155 950.170 3411.080 1010.420 ;
        RECT 3444.590 991.485 3446.020 1014.285 ;
        RECT 3448.180 1011.190 3450.340 1014.285 ;
        RECT 3448.180 1004.540 3449.020 1011.190 ;
        RECT 3448.770 1001.465 3449.020 1004.540 ;
        RECT 3467.805 990.185 3469.235 1014.285 ;
        RECT 3473.580 1012.205 3480.400 1015.120 ;
        RECT 3473.580 1010.470 3479.820 1012.205 ;
        RECT 3474.660 1009.025 3479.820 1010.470 ;
      LAYER pwell ;
        RECT 3480.935 1009.785 3518.355 1015.215 ;
      LAYER nwell ;
        RECT 3474.660 1006.580 3476.280 1009.025 ;
        RECT 3474.660 1006.505 3475.740 1006.580 ;
      LAYER pwell ;
        RECT 3480.935 1005.700 3484.255 1009.785 ;
        RECT 3482.955 975.615 3484.255 1005.700 ;
        RECT 3489.965 1009.265 3518.355 1009.785 ;
        RECT 3489.965 975.615 3491.550 1009.265 ;
        RECT 3482.955 969.160 3485.985 975.615 ;
        RECT 3482.955 968.410 3483.260 969.160 ;
      LAYER nwell ;
        RECT 3422.265 956.725 3424.055 966.085 ;
        RECT 3420.410 950.170 3424.055 956.725 ;
        RECT 3407.155 934.550 3413.345 950.170 ;
        RECT 3417.785 934.550 3424.055 950.170 ;
        RECT 3460.595 952.350 3461.265 968.060 ;
        RECT 3438.620 935.875 3440.050 944.665 ;
        RECT 3453.195 935.875 3454.045 944.665 ;
        RECT 3460.595 935.875 3461.775 952.350 ;
        RECT 3438.620 935.760 3461.775 935.875 ;
        RECT 3471.165 935.760 3472.345 968.060 ;
        RECT 3482.245 952.350 3483.165 968.060 ;
        RECT 3481.735 935.760 3483.165 952.350 ;
        RECT 3438.620 934.330 3483.165 935.760 ;
      LAYER pwell ;
        RECT 3483.975 938.230 3485.985 969.160 ;
        RECT 3488.820 962.120 3491.550 975.615 ;
        RECT 3487.520 938.230 3491.550 962.120 ;
        RECT 3483.975 937.135 3491.550 938.230 ;
        RECT 3513.135 974.755 3518.355 1009.265 ;
        RECT 3513.135 948.090 3517.315 974.755 ;
      LAYER nwell ;
        RECT 3518.665 968.960 3528.380 1015.415 ;
      LAYER pwell ;
        RECT 3513.135 937.135 3518.355 948.090 ;
        RECT 3483.975 934.710 3518.355 937.135 ;
      LAYER nwell ;
        RECT 3518.665 934.560 3528.385 968.960 ;
      LAYER pwell ;
        RECT 3528.685 934.710 3532.565 1015.290 ;
      LAYER nwell ;
        RECT 3532.880 1008.615 3566.975 1015.415 ;
        RECT 3532.880 936.370 3534.690 1008.615 ;
        RECT 3556.515 1007.485 3566.975 1008.615 ;
        RECT 3556.515 948.030 3558.475 1007.485 ;
        RECT 3561.545 948.030 3566.975 1007.485 ;
        RECT 3556.515 936.370 3566.975 948.030 ;
        RECT 3532.880 934.565 3566.975 936.370 ;
        RECT 3532.880 934.560 3558.230 934.565 ;
        RECT 107.600 908.585 111.515 908.880 ;
        RECT 118.765 908.285 143.410 909.715 ;
        RECT 190.675 908.585 194.335 912.110 ;
        RECT 3393.665 790.890 3397.325 794.415 ;
        RECT 3444.590 793.285 3469.235 794.715 ;
        RECT 3476.485 794.120 3480.400 794.415 ;
        RECT 3407.155 729.170 3411.080 789.420 ;
        RECT 3444.590 770.485 3446.020 793.285 ;
        RECT 3448.180 790.190 3450.340 793.285 ;
        RECT 3448.180 783.540 3449.020 790.190 ;
        RECT 3448.770 780.465 3449.020 783.540 ;
        RECT 3467.805 769.185 3469.235 793.285 ;
        RECT 3473.580 791.205 3480.400 794.120 ;
        RECT 3473.580 789.470 3479.820 791.205 ;
        RECT 3474.660 788.025 3479.820 789.470 ;
      LAYER pwell ;
        RECT 3480.935 788.785 3518.355 794.215 ;
      LAYER nwell ;
        RECT 3474.660 785.580 3476.280 788.025 ;
        RECT 3474.660 785.505 3475.740 785.580 ;
      LAYER pwell ;
        RECT 3480.935 784.700 3484.255 788.785 ;
        RECT 3482.955 754.615 3484.255 784.700 ;
        RECT 3489.965 788.265 3518.355 788.785 ;
        RECT 3489.965 754.615 3491.550 788.265 ;
        RECT 3482.955 748.160 3485.985 754.615 ;
        RECT 3482.955 747.410 3483.260 748.160 ;
      LAYER nwell ;
        RECT 3422.265 735.725 3424.055 745.085 ;
        RECT 3420.410 729.170 3424.055 735.725 ;
        RECT 3407.155 713.550 3413.345 729.170 ;
        RECT 3417.785 713.550 3424.055 729.170 ;
        RECT 3460.595 731.350 3461.265 747.060 ;
        RECT 3438.620 714.875 3440.050 723.665 ;
        RECT 3453.195 714.875 3454.045 723.665 ;
        RECT 3460.595 714.875 3461.775 731.350 ;
        RECT 3438.620 714.760 3461.775 714.875 ;
        RECT 3471.165 714.760 3472.345 747.060 ;
        RECT 3482.245 731.350 3483.165 747.060 ;
        RECT 3481.735 714.760 3483.165 731.350 ;
        RECT 3438.620 713.330 3483.165 714.760 ;
      LAYER pwell ;
        RECT 3483.975 717.230 3485.985 748.160 ;
        RECT 3488.820 741.120 3491.550 754.615 ;
        RECT 3487.520 717.230 3491.550 741.120 ;
        RECT 3483.975 716.135 3491.550 717.230 ;
        RECT 3513.135 753.755 3518.355 788.265 ;
        RECT 3513.135 727.090 3517.315 753.755 ;
      LAYER nwell ;
        RECT 3518.665 747.960 3528.380 794.415 ;
      LAYER pwell ;
        RECT 3513.135 716.135 3518.355 727.090 ;
        RECT 3483.975 713.710 3518.355 716.135 ;
      LAYER nwell ;
        RECT 3518.665 713.560 3528.385 747.960 ;
      LAYER pwell ;
        RECT 3528.685 713.710 3532.565 794.290 ;
      LAYER nwell ;
        RECT 3532.880 787.615 3566.975 794.415 ;
        RECT 3532.880 715.370 3534.690 787.615 ;
        RECT 3556.515 786.485 3566.975 787.615 ;
        RECT 3556.515 727.030 3558.475 786.485 ;
        RECT 3561.545 727.030 3566.975 786.485 ;
        RECT 3556.515 715.370 3566.975 727.030 ;
        RECT 3532.880 713.565 3566.975 715.370 ;
        RECT 3532.880 713.560 3558.230 713.565 ;
        RECT 197.795 562.860 199.315 621.965 ;
        RECT 3393.665 568.890 3397.325 572.415 ;
        RECT 3444.590 571.285 3469.235 572.715 ;
        RECT 3476.485 572.120 3480.400 572.415 ;
      LAYER pwell ;
        RECT 176.210 554.495 199.065 562.285 ;
      LAYER nwell ;
        RECT 3407.155 507.170 3411.080 567.420 ;
        RECT 3444.590 548.485 3446.020 571.285 ;
        RECT 3448.180 568.190 3450.340 571.285 ;
        RECT 3448.180 561.540 3449.020 568.190 ;
        RECT 3448.770 558.465 3449.020 561.540 ;
        RECT 3467.805 547.185 3469.235 571.285 ;
        RECT 3473.580 569.205 3480.400 572.120 ;
        RECT 3473.580 567.470 3479.820 569.205 ;
        RECT 3474.660 566.025 3479.820 567.470 ;
      LAYER pwell ;
        RECT 3480.935 566.785 3518.355 572.215 ;
      LAYER nwell ;
        RECT 3474.660 563.580 3476.280 566.025 ;
        RECT 3474.660 563.505 3475.740 563.580 ;
      LAYER pwell ;
        RECT 3480.935 562.700 3484.255 566.785 ;
        RECT 3482.955 532.615 3484.255 562.700 ;
        RECT 3489.965 566.265 3518.355 566.785 ;
        RECT 3489.965 532.615 3491.550 566.265 ;
        RECT 3482.955 526.160 3485.985 532.615 ;
        RECT 3482.955 525.410 3483.260 526.160 ;
      LAYER nwell ;
        RECT 3422.265 513.725 3424.055 523.085 ;
        RECT 3420.410 507.170 3424.055 513.725 ;
        RECT 3407.155 491.550 3413.345 507.170 ;
        RECT 3417.785 491.550 3424.055 507.170 ;
        RECT 3460.595 509.350 3461.265 525.060 ;
        RECT 3438.620 492.875 3440.050 501.665 ;
        RECT 3453.195 492.875 3454.045 501.665 ;
        RECT 3460.595 492.875 3461.775 509.350 ;
        RECT 3438.620 492.760 3461.775 492.875 ;
        RECT 3471.165 492.760 3472.345 525.060 ;
        RECT 3482.245 509.350 3483.165 525.060 ;
        RECT 3481.735 492.760 3483.165 509.350 ;
        RECT 3438.620 491.330 3483.165 492.760 ;
      LAYER pwell ;
        RECT 3483.975 495.230 3485.985 526.160 ;
        RECT 3488.820 519.120 3491.550 532.615 ;
        RECT 3487.520 495.230 3491.550 519.120 ;
        RECT 3483.975 494.135 3491.550 495.230 ;
        RECT 3513.135 531.755 3518.355 566.265 ;
        RECT 3513.135 505.090 3517.315 531.755 ;
      LAYER nwell ;
        RECT 3518.665 525.960 3528.380 572.415 ;
      LAYER pwell ;
        RECT 3513.135 494.135 3518.355 505.090 ;
        RECT 3483.975 491.710 3518.355 494.135 ;
      LAYER nwell ;
        RECT 3518.665 491.560 3528.385 525.960 ;
      LAYER pwell ;
        RECT 3528.685 491.710 3532.565 572.290 ;
      LAYER nwell ;
        RECT 3532.880 565.615 3566.975 572.415 ;
        RECT 3532.880 493.370 3534.690 565.615 ;
        RECT 3556.515 564.485 3566.975 565.615 ;
        RECT 3556.515 505.030 3558.475 564.485 ;
        RECT 3561.545 505.030 3566.975 564.485 ;
        RECT 3556.515 493.370 3566.975 505.030 ;
        RECT 3532.880 491.565 3566.975 493.370 ;
        RECT 3532.880 491.560 3558.230 491.565 ;
        RECT 398.035 197.795 457.140 199.315 ;
        RECT 2849.035 197.795 2908.140 199.315 ;
        RECT 3118.035 197.795 3177.140 199.315 ;
        RECT 1008.890 190.675 1012.415 194.335 ;
        RECT 1551.890 190.675 1555.415 194.335 ;
        RECT 1825.890 190.675 1829.415 194.335 ;
        RECT 2099.890 190.675 2103.415 194.335 ;
        RECT 2373.890 190.675 2377.415 194.335 ;
        RECT 2647.890 190.675 2651.415 194.335 ;
        RECT 931.550 176.920 1007.420 180.845 ;
        RECT 1474.550 176.920 1550.420 180.845 ;
        RECT 1748.550 176.920 1824.420 180.845 ;
        RECT 2022.550 176.920 2098.420 180.845 ;
        RECT 2296.550 176.920 2372.420 180.845 ;
        RECT 2570.550 176.920 2646.420 180.845 ;
        RECT 931.550 174.655 947.170 176.920 ;
        RECT 1474.550 174.655 1490.170 176.920 ;
        RECT 1748.550 174.655 1764.170 176.920 ;
        RECT 2022.550 174.655 2038.170 176.920 ;
        RECT 2296.550 174.655 2312.170 176.920 ;
        RECT 2570.550 174.655 2586.170 176.920 ;
      LAYER pwell ;
        RECT 3177.715 176.210 3185.505 199.065 ;
      LAYER nwell ;
        RECT 931.550 167.590 947.170 170.215 ;
        RECT 1474.550 167.590 1490.170 170.215 ;
        RECT 1748.550 167.590 1764.170 170.215 ;
        RECT 2022.550 167.590 2038.170 170.215 ;
        RECT 2296.550 167.590 2312.170 170.215 ;
        RECT 2570.550 167.590 2586.170 170.215 ;
        RECT 931.550 165.735 953.725 167.590 ;
        RECT 1474.550 165.735 1496.725 167.590 ;
        RECT 1748.550 165.735 1770.725 167.590 ;
        RECT 2022.550 165.735 2044.725 167.590 ;
        RECT 2296.550 165.735 2318.725 167.590 ;
        RECT 2570.550 165.735 2592.725 167.590 ;
        RECT 931.550 163.945 963.085 165.735 ;
        RECT 1474.550 163.945 1506.085 165.735 ;
        RECT 1748.550 163.945 1780.085 165.735 ;
        RECT 2022.550 163.945 2054.085 165.735 ;
        RECT 2296.550 163.945 2328.085 165.735 ;
        RECT 2570.550 163.945 2602.085 165.735 ;
        RECT 931.330 147.950 941.665 149.380 ;
        RECT 1474.330 147.950 1484.665 149.380 ;
        RECT 1748.330 147.950 1758.665 149.380 ;
        RECT 2022.330 147.950 2032.665 149.380 ;
        RECT 2296.330 147.950 2306.665 149.380 ;
        RECT 2570.330 147.950 2580.665 149.380 ;
        RECT 931.330 134.805 932.875 147.950 ;
        RECT 988.485 141.980 1012.715 143.410 ;
        RECT 1011.285 139.820 1012.715 141.980 ;
        RECT 1001.540 139.230 1012.715 139.820 ;
        RECT 998.465 138.980 1012.715 139.230 ;
        RECT 1008.190 137.660 1012.715 138.980 ;
        RECT 931.330 133.955 941.665 134.805 ;
        RECT 931.330 127.405 932.875 133.955 ;
        RECT 931.330 126.735 965.060 127.405 ;
        RECT 931.330 126.225 949.350 126.735 ;
        RECT 931.330 116.835 932.760 126.225 ;
        RECT 1011.285 120.195 1012.715 137.660 ;
        RECT 987.185 118.765 1012.715 120.195 ;
        RECT 1474.330 134.805 1475.875 147.950 ;
        RECT 1531.485 141.980 1555.715 143.410 ;
        RECT 1554.285 139.820 1555.715 141.980 ;
        RECT 1544.540 139.230 1555.715 139.820 ;
        RECT 1541.465 138.980 1555.715 139.230 ;
        RECT 1551.190 137.660 1555.715 138.980 ;
        RECT 1474.330 133.955 1484.665 134.805 ;
        RECT 1474.330 127.405 1475.875 133.955 ;
        RECT 1474.330 126.735 1508.060 127.405 ;
        RECT 1474.330 126.225 1492.350 126.735 ;
        RECT 1474.330 116.835 1475.760 126.225 ;
        RECT 1554.285 120.195 1555.715 137.660 ;
        RECT 1530.185 118.765 1555.715 120.195 ;
        RECT 1748.330 134.805 1749.875 147.950 ;
        RECT 1805.485 141.980 1829.715 143.410 ;
        RECT 1828.285 139.820 1829.715 141.980 ;
        RECT 1818.540 139.230 1829.715 139.820 ;
        RECT 1815.465 138.980 1829.715 139.230 ;
        RECT 1825.190 137.660 1829.715 138.980 ;
        RECT 1748.330 133.955 1758.665 134.805 ;
        RECT 1748.330 127.405 1749.875 133.955 ;
        RECT 1748.330 126.735 1782.060 127.405 ;
        RECT 1748.330 126.225 1766.350 126.735 ;
        RECT 1748.330 116.835 1749.760 126.225 ;
        RECT 1828.285 120.195 1829.715 137.660 ;
        RECT 1804.185 118.765 1829.715 120.195 ;
        RECT 2022.330 134.805 2023.875 147.950 ;
        RECT 2079.485 141.980 2103.715 143.410 ;
        RECT 2102.285 139.820 2103.715 141.980 ;
        RECT 2092.540 139.230 2103.715 139.820 ;
        RECT 2089.465 138.980 2103.715 139.230 ;
        RECT 2099.190 137.660 2103.715 138.980 ;
        RECT 2022.330 133.955 2032.665 134.805 ;
        RECT 2022.330 127.405 2023.875 133.955 ;
        RECT 2022.330 126.735 2056.060 127.405 ;
        RECT 2022.330 126.225 2040.350 126.735 ;
        RECT 2022.330 116.835 2023.760 126.225 ;
        RECT 2102.285 120.195 2103.715 137.660 ;
        RECT 2078.185 118.765 2103.715 120.195 ;
        RECT 2296.330 134.805 2297.875 147.950 ;
        RECT 2353.485 141.980 2377.715 143.410 ;
        RECT 2376.285 139.820 2377.715 141.980 ;
        RECT 2366.540 139.230 2377.715 139.820 ;
        RECT 2363.465 138.980 2377.715 139.230 ;
        RECT 2373.190 137.660 2377.715 138.980 ;
        RECT 2296.330 133.955 2306.665 134.805 ;
        RECT 2296.330 127.405 2297.875 133.955 ;
        RECT 2296.330 126.735 2330.060 127.405 ;
        RECT 2296.330 126.225 2314.350 126.735 ;
        RECT 2296.330 116.835 2297.760 126.225 ;
        RECT 2376.285 120.195 2377.715 137.660 ;
        RECT 2352.185 118.765 2377.715 120.195 ;
        RECT 2570.330 134.805 2571.875 147.950 ;
        RECT 2627.485 141.980 2651.715 143.410 ;
        RECT 2650.285 139.820 2651.715 141.980 ;
        RECT 2640.540 139.230 2651.715 139.820 ;
        RECT 2637.465 138.980 2651.715 139.230 ;
        RECT 2647.190 137.660 2651.715 138.980 ;
        RECT 2570.330 133.955 2580.665 134.805 ;
        RECT 2570.330 127.405 2571.875 133.955 ;
        RECT 2570.330 126.735 2604.060 127.405 ;
        RECT 2570.330 126.225 2588.350 126.735 ;
        RECT 2570.330 116.835 2571.760 126.225 ;
        RECT 2650.285 120.195 2651.715 137.660 ;
        RECT 2626.185 118.765 2651.715 120.195 ;
        RECT 931.330 115.655 965.060 116.835 ;
        RECT 1474.330 115.655 1508.060 116.835 ;
        RECT 1748.330 115.655 1782.060 116.835 ;
        RECT 2022.330 115.655 2056.060 116.835 ;
        RECT 2296.330 115.655 2330.060 116.835 ;
        RECT 2570.330 115.655 2604.060 116.835 ;
        RECT 931.330 106.265 932.760 115.655 ;
        RECT 1007.470 113.340 1012.120 114.420 ;
        RECT 1003.505 112.260 1012.120 113.340 ;
        RECT 1003.580 111.720 1012.120 112.260 ;
        RECT 1006.025 111.515 1012.120 111.720 ;
        RECT 1006.025 108.180 1012.415 111.515 ;
        RECT 1009.205 107.600 1012.415 108.180 ;
        RECT 931.330 105.755 949.350 106.265 ;
        RECT 931.330 104.835 965.060 105.755 ;
      LAYER pwell ;
        RECT 1002.700 105.045 1012.215 107.065 ;
        RECT 965.410 104.740 1012.215 105.045 ;
      LAYER nwell ;
        RECT 1474.330 106.265 1475.760 115.655 ;
        RECT 1550.470 113.340 1555.120 114.420 ;
        RECT 1546.505 112.260 1555.120 113.340 ;
        RECT 1546.580 111.720 1555.120 112.260 ;
        RECT 1549.025 111.515 1555.120 111.720 ;
        RECT 1549.025 108.180 1555.415 111.515 ;
        RECT 1552.205 107.600 1555.415 108.180 ;
        RECT 1474.330 105.755 1492.350 106.265 ;
        RECT 1474.330 104.835 1508.060 105.755 ;
      LAYER pwell ;
        RECT 1545.700 105.045 1555.215 107.065 ;
        RECT 1508.410 104.740 1555.215 105.045 ;
      LAYER nwell ;
        RECT 1748.330 106.265 1749.760 115.655 ;
        RECT 1824.470 113.340 1829.120 114.420 ;
        RECT 1820.505 112.260 1829.120 113.340 ;
        RECT 1820.580 111.720 1829.120 112.260 ;
        RECT 1823.025 111.515 1829.120 111.720 ;
        RECT 1823.025 108.180 1829.415 111.515 ;
        RECT 1826.205 107.600 1829.415 108.180 ;
        RECT 1748.330 105.755 1766.350 106.265 ;
        RECT 1748.330 104.835 1782.060 105.755 ;
      LAYER pwell ;
        RECT 1819.700 105.045 1829.215 107.065 ;
        RECT 1782.410 104.740 1829.215 105.045 ;
      LAYER nwell ;
        RECT 2022.330 106.265 2023.760 115.655 ;
        RECT 2098.470 113.340 2103.120 114.420 ;
        RECT 2094.505 112.260 2103.120 113.340 ;
        RECT 2094.580 111.720 2103.120 112.260 ;
        RECT 2097.025 111.515 2103.120 111.720 ;
        RECT 2097.025 108.180 2103.415 111.515 ;
        RECT 2100.205 107.600 2103.415 108.180 ;
        RECT 2022.330 105.755 2040.350 106.265 ;
        RECT 2022.330 104.835 2056.060 105.755 ;
      LAYER pwell ;
        RECT 2093.700 105.045 2103.215 107.065 ;
        RECT 2056.410 104.740 2103.215 105.045 ;
      LAYER nwell ;
        RECT 2296.330 106.265 2297.760 115.655 ;
        RECT 2372.470 113.340 2377.120 114.420 ;
        RECT 2368.505 112.260 2377.120 113.340 ;
        RECT 2368.580 111.720 2377.120 112.260 ;
        RECT 2371.025 111.515 2377.120 111.720 ;
        RECT 2371.025 108.180 2377.415 111.515 ;
        RECT 2374.205 107.600 2377.415 108.180 ;
        RECT 2296.330 105.755 2314.350 106.265 ;
        RECT 2296.330 104.835 2330.060 105.755 ;
      LAYER pwell ;
        RECT 2367.700 105.045 2377.215 107.065 ;
        RECT 2330.410 104.740 2377.215 105.045 ;
      LAYER nwell ;
        RECT 2570.330 106.265 2571.760 115.655 ;
        RECT 2646.470 113.340 2651.120 114.420 ;
        RECT 2642.505 112.260 2651.120 113.340 ;
        RECT 2642.580 111.720 2651.120 112.260 ;
        RECT 2645.025 111.515 2651.120 111.720 ;
        RECT 2645.025 108.180 2651.415 111.515 ;
        RECT 2648.205 107.600 2651.415 108.180 ;
        RECT 2570.330 105.755 2588.350 106.265 ;
        RECT 2570.330 104.835 2604.060 105.755 ;
      LAYER pwell ;
        RECT 2641.700 105.045 2651.215 107.065 ;
        RECT 2604.410 104.740 2651.215 105.045 ;
        RECT 966.160 104.025 1012.215 104.740 ;
        RECT 1509.160 104.025 1555.215 104.740 ;
        RECT 1783.160 104.025 1829.215 104.740 ;
        RECT 2057.160 104.025 2103.215 104.740 ;
        RECT 2331.160 104.025 2377.215 104.740 ;
        RECT 2605.160 104.025 2651.215 104.740 ;
        RECT 931.710 103.745 1012.215 104.025 ;
        RECT 679.530 103.265 738.130 103.270 ;
        RECT 662.870 102.005 738.130 103.265 ;
        RECT 662.870 100.770 666.070 102.005 ;
        RECT 679.530 100.770 738.130 102.005 ;
        RECT 662.870 97.475 738.130 100.770 ;
        RECT 662.870 75.865 664.440 97.475 ;
        RECT 736.565 75.865 738.130 97.475 ;
        RECT 662.870 70.685 738.130 75.865 ;
        RECT 662.870 69.645 676.090 70.685 ;
        RECT 696.250 69.645 738.130 70.685 ;
        RECT 931.710 102.015 972.615 103.745 ;
        RECT 931.710 100.480 935.230 102.015 ;
        RECT 931.710 99.180 959.120 100.480 ;
        RECT 931.710 98.035 972.615 99.180 ;
        RECT 1006.785 98.035 1012.215 103.745 ;
        RECT 931.710 96.450 1012.215 98.035 ;
        RECT 931.710 74.865 934.135 96.450 ;
        RECT 1006.265 74.865 1012.215 96.450 ;
        RECT 931.710 70.685 1012.215 74.865 ;
        RECT 931.710 69.645 945.090 70.685 ;
        RECT 971.755 69.645 1012.215 70.685 ;
        RECT 1474.710 103.745 1555.215 104.025 ;
        RECT 1474.710 102.015 1515.615 103.745 ;
        RECT 1474.710 100.480 1478.230 102.015 ;
        RECT 1474.710 99.180 1502.120 100.480 ;
        RECT 1474.710 98.035 1515.615 99.180 ;
        RECT 1549.785 98.035 1555.215 103.745 ;
        RECT 1474.710 96.450 1555.215 98.035 ;
        RECT 1474.710 74.865 1477.135 96.450 ;
        RECT 1549.265 74.865 1555.215 96.450 ;
        RECT 1474.710 70.685 1555.215 74.865 ;
        RECT 1474.710 69.645 1488.090 70.685 ;
        RECT 1514.755 69.645 1555.215 70.685 ;
        RECT 1748.710 103.745 1829.215 104.025 ;
        RECT 1748.710 102.015 1789.615 103.745 ;
        RECT 1748.710 100.480 1752.230 102.015 ;
        RECT 1748.710 99.180 1776.120 100.480 ;
        RECT 1748.710 98.035 1789.615 99.180 ;
        RECT 1823.785 98.035 1829.215 103.745 ;
        RECT 1748.710 96.450 1829.215 98.035 ;
        RECT 1748.710 74.865 1751.135 96.450 ;
        RECT 1823.265 74.865 1829.215 96.450 ;
        RECT 1748.710 70.685 1829.215 74.865 ;
        RECT 1748.710 69.645 1762.090 70.685 ;
        RECT 1788.755 69.645 1829.215 70.685 ;
        RECT 2022.710 103.745 2103.215 104.025 ;
        RECT 2022.710 102.015 2063.615 103.745 ;
        RECT 2022.710 100.480 2026.230 102.015 ;
        RECT 2022.710 99.180 2050.120 100.480 ;
        RECT 2022.710 98.035 2063.615 99.180 ;
        RECT 2097.785 98.035 2103.215 103.745 ;
        RECT 2022.710 96.450 2103.215 98.035 ;
        RECT 2022.710 74.865 2025.135 96.450 ;
        RECT 2097.265 74.865 2103.215 96.450 ;
        RECT 2022.710 70.685 2103.215 74.865 ;
        RECT 2022.710 69.645 2036.090 70.685 ;
        RECT 2062.755 69.645 2103.215 70.685 ;
        RECT 2296.710 103.745 2377.215 104.025 ;
        RECT 2296.710 102.015 2337.615 103.745 ;
        RECT 2296.710 100.480 2300.230 102.015 ;
        RECT 2296.710 99.180 2324.120 100.480 ;
        RECT 2296.710 98.035 2337.615 99.180 ;
        RECT 2371.785 98.035 2377.215 103.745 ;
        RECT 2296.710 96.450 2377.215 98.035 ;
        RECT 2296.710 74.865 2299.135 96.450 ;
        RECT 2371.265 74.865 2377.215 96.450 ;
        RECT 2296.710 70.685 2377.215 74.865 ;
        RECT 2296.710 69.645 2310.090 70.685 ;
        RECT 2336.755 69.645 2377.215 70.685 ;
        RECT 2570.710 103.745 2651.215 104.025 ;
        RECT 2570.710 102.015 2611.615 103.745 ;
        RECT 2570.710 100.480 2574.230 102.015 ;
        RECT 2570.710 99.180 2598.120 100.480 ;
        RECT 2570.710 98.035 2611.615 99.180 ;
        RECT 2645.785 98.035 2651.215 103.745 ;
        RECT 2570.710 96.450 2651.215 98.035 ;
        RECT 2570.710 74.865 2573.135 96.450 ;
        RECT 2645.265 74.865 2651.215 96.450 ;
        RECT 2570.710 70.685 2651.215 74.865 ;
        RECT 2570.710 69.645 2584.090 70.685 ;
        RECT 2610.755 69.645 2651.215 70.685 ;
      LAYER nwell ;
        RECT 662.670 59.620 738.330 69.335 ;
        RECT 931.560 59.620 1012.415 69.335 ;
        RECT 1474.560 59.620 1555.415 69.335 ;
        RECT 1748.560 59.620 1829.415 69.335 ;
        RECT 2022.560 59.620 2103.415 69.335 ;
        RECT 2296.560 59.620 2377.415 69.335 ;
        RECT 2570.560 59.620 2651.415 69.335 ;
        RECT 931.560 59.615 965.960 59.620 ;
        RECT 1474.560 59.615 1508.960 59.620 ;
        RECT 1748.560 59.615 1782.960 59.620 ;
        RECT 2022.560 59.615 2056.960 59.620 ;
        RECT 2296.560 59.615 2330.960 59.620 ;
        RECT 2570.560 59.615 2604.960 59.620 ;
      LAYER pwell ;
        RECT 662.710 55.435 738.290 59.315 ;
        RECT 931.710 55.435 1012.290 59.315 ;
        RECT 1474.710 55.435 1555.290 59.315 ;
        RECT 1748.710 55.435 1829.290 59.315 ;
        RECT 2022.710 55.435 2103.290 59.315 ;
        RECT 2296.710 55.435 2377.290 59.315 ;
        RECT 2570.710 55.435 2651.290 59.315 ;
      LAYER nwell ;
        RECT 662.380 53.310 738.515 55.120 ;
        RECT 662.380 31.485 664.905 53.310 ;
        RECT 736.325 31.485 738.515 53.310 ;
        RECT 662.380 29.790 738.515 31.485 ;
        RECT 931.560 53.310 1012.415 55.120 ;
        RECT 931.560 31.485 933.370 53.310 ;
        RECT 1005.615 31.485 1012.415 53.310 ;
        RECT 931.560 29.770 1012.415 31.485 ;
        RECT 1474.560 53.310 1555.415 55.120 ;
        RECT 1474.560 31.485 1476.370 53.310 ;
        RECT 1548.615 31.485 1555.415 53.310 ;
        RECT 1474.560 29.770 1555.415 31.485 ;
        RECT 1748.560 53.310 1829.415 55.120 ;
        RECT 1748.560 31.485 1750.370 53.310 ;
        RECT 1822.615 31.485 1829.415 53.310 ;
        RECT 1748.560 29.770 1829.415 31.485 ;
        RECT 2022.560 53.310 2103.415 55.120 ;
        RECT 2022.560 31.485 2024.370 53.310 ;
        RECT 2096.615 31.485 2103.415 53.310 ;
        RECT 2022.560 29.770 2103.415 31.485 ;
        RECT 2296.560 53.310 2377.415 55.120 ;
        RECT 2296.560 31.485 2298.370 53.310 ;
        RECT 2370.615 31.485 2377.415 53.310 ;
        RECT 2296.560 29.770 2377.415 31.485 ;
        RECT 2570.560 53.310 2651.415 55.120 ;
        RECT 2570.560 31.485 2572.370 53.310 ;
        RECT 2644.615 31.485 2651.415 53.310 ;
        RECT 2570.560 29.770 2651.415 31.485 ;
        RECT 931.565 29.525 1012.415 29.770 ;
        RECT 931.565 26.455 945.030 29.525 ;
        RECT 1004.485 26.455 1012.415 29.525 ;
        RECT 931.565 21.025 1012.415 26.455 ;
        RECT 1474.565 29.525 1555.415 29.770 ;
        RECT 1474.565 26.455 1488.030 29.525 ;
        RECT 1547.485 26.455 1555.415 29.525 ;
        RECT 1474.565 21.025 1555.415 26.455 ;
        RECT 1748.565 29.525 1829.415 29.770 ;
        RECT 1748.565 26.455 1762.030 29.525 ;
        RECT 1821.485 26.455 1829.415 29.525 ;
        RECT 1748.565 21.025 1829.415 26.455 ;
        RECT 2022.565 29.525 2103.415 29.770 ;
        RECT 2022.565 26.455 2036.030 29.525 ;
        RECT 2095.485 26.455 2103.415 29.525 ;
        RECT 2022.565 21.025 2103.415 26.455 ;
        RECT 2296.565 29.525 2377.415 29.770 ;
        RECT 2296.565 26.455 2310.030 29.525 ;
        RECT 2369.485 26.455 2377.415 29.525 ;
        RECT 2296.565 21.025 2377.415 26.455 ;
        RECT 2570.565 29.525 2651.415 29.770 ;
        RECT 2570.565 26.455 2584.030 29.525 ;
        RECT 2643.485 26.455 2651.415 29.525 ;
        RECT 2570.565 21.025 2651.415 26.455 ;
      LAYER li1 ;
        RECT 377.905 5036.265 447.045 5169.100 ;
        RECT 617.905 5036.265 687.045 5169.100 ;
        RECT 857.905 5036.265 927.045 5169.100 ;
        RECT 1147.610 4990.035 1219.855 5187.695 ;
        RECT 1404.610 4990.035 1476.855 5187.695 ;
        RECT 1698.070 4990.035 1769.775 5187.695 ;
        RECT 2126.905 5036.265 2196.045 5169.100 ;
        RECT 2373.905 5036.265 2443.045 5169.100 ;
        RECT 2631.905 5036.265 2701.045 5169.100 ;
        RECT 2879.070 4990.035 2950.775 5187.695 ;
        RECT 3137.905 5036.265 3207.045 5169.100 ;
        RECT 1147.610 4989.065 1158.155 4990.035 ;
        RECT 1159.035 4989.920 1160.045 4990.035 ;
        RECT 1216.730 4989.920 1217.680 4990.035 ;
        RECT 1159.035 4988.970 1217.680 4989.920 ;
        RECT 1404.610 4989.065 1415.155 4990.035 ;
        RECT 1416.035 4989.920 1417.045 4990.035 ;
        RECT 1473.730 4989.920 1474.680 4990.035 ;
        RECT 1416.035 4988.970 1474.680 4989.920 ;
        RECT 1709.065 4989.890 1710.045 4990.035 ;
        RECT 1766.760 4989.890 1767.650 4990.035 ;
        RECT 1709.065 4989.000 1767.650 4989.890 ;
        RECT 2890.065 4989.890 2891.045 4990.035 ;
        RECT 2947.760 4989.890 2948.650 4990.035 ;
        RECT 2890.065 4989.000 2948.650 4989.890 ;
        RECT 18.900 4778.905 151.735 4848.045 ;
        RECT 3389.065 4783.845 3587.695 4794.390 ;
        RECT 3390.035 4782.965 3587.695 4783.845 ;
        RECT 3388.970 4781.955 3587.695 4782.965 ;
        RECT 3388.970 4725.270 3389.920 4781.955 ;
        RECT 3390.035 4725.270 3587.695 4781.955 ;
        RECT 3388.970 4724.320 3587.695 4725.270 ;
        RECT 3390.035 4722.145 3587.695 4724.320 ;
        RECT 0.220 4565.240 196.980 4639.755 ;
        RECT 3391.020 4457.245 3587.780 4531.760 ;
        RECT 0.305 4424.680 197.965 4426.855 ;
        RECT 0.305 4423.730 199.030 4424.680 ;
        RECT 0.305 4367.045 197.965 4423.730 ;
        RECT 198.080 4367.045 199.030 4423.730 ;
        RECT 0.305 4366.035 199.030 4367.045 ;
        RECT 0.305 4365.155 197.965 4366.035 ;
        RECT 0.305 4354.610 198.935 4365.155 ;
        RECT 3483.895 4315.085 3518.220 4315.115 ;
        RECT 3519.275 4315.085 3528.150 4315.115 ;
        RECT 3393.995 4315.000 3396.995 4315.085 ;
        RECT 3445.220 4315.000 3468.605 4315.085 ;
        RECT 3476.815 4315.000 3480.070 4315.085 ;
        RECT 3481.065 4315.000 3518.225 4315.085 ;
        RECT 3518.995 4315.000 3528.150 4315.085 ;
        RECT 3528.815 4315.000 3532.435 4315.160 ;
        RECT 3533.155 4315.085 3558.090 4315.115 ;
        RECT 3533.155 4315.000 3566.645 4315.085 ;
        RECT 3388.230 4235.000 3587.705 4315.000 ;
        RECT 3407.485 4234.880 3413.015 4235.000 ;
        RECT 3418.115 4234.880 3423.725 4235.000 ;
        RECT 3439.250 4234.915 3482.580 4235.000 ;
        RECT 3484.105 4234.840 3518.225 4235.000 ;
        RECT 3518.995 4234.915 3528.055 4235.000 ;
        RECT 3528.815 4234.840 3532.435 4235.000 ;
        RECT 3533.215 4234.895 3566.645 4235.000 ;
        RECT 0.305 4212.650 197.965 4214.775 ;
        RECT 0.305 4211.760 199.000 4212.650 ;
        RECT 0.305 4155.045 197.965 4211.760 ;
        RECT 198.110 4155.045 199.000 4211.760 ;
        RECT 0.305 4154.065 199.000 4155.045 ;
        RECT 0.305 4143.070 197.965 4154.065 ;
        RECT 3389.065 4082.845 3587.695 4093.390 ;
        RECT 3390.035 4081.965 3587.695 4082.845 ;
        RECT 3388.970 4080.955 3587.695 4081.965 ;
        RECT 3388.970 4024.270 3389.920 4080.955 ;
        RECT 3390.035 4024.270 3587.695 4080.955 ;
        RECT 3388.970 4023.320 3587.695 4024.270 ;
        RECT 3390.035 4021.145 3587.695 4023.320 ;
        RECT 21.355 4006.000 54.785 4006.105 ;
        RECT 55.565 4006.000 59.185 4006.160 ;
        RECT 59.945 4006.000 69.005 4006.085 ;
        RECT 69.775 4006.000 103.895 4006.160 ;
        RECT 105.420 4006.000 148.750 4006.085 ;
        RECT 164.275 4006.000 169.885 4006.120 ;
        RECT 174.985 4006.000 180.515 4006.120 ;
        RECT 0.295 3926.000 199.770 4006.000 ;
        RECT 21.355 3925.915 54.845 3926.000 ;
        RECT 29.910 3925.885 54.845 3925.915 ;
        RECT 55.565 3925.840 59.185 3926.000 ;
        RECT 59.850 3925.915 69.005 3926.000 ;
        RECT 69.775 3925.915 106.935 3926.000 ;
        RECT 107.930 3925.915 111.185 3926.000 ;
        RECT 119.395 3925.915 142.780 3926.000 ;
        RECT 191.005 3925.915 194.005 3926.000 ;
        RECT 59.850 3925.885 68.725 3925.915 ;
        RECT 69.780 3925.885 104.105 3925.915 ;
        RECT 3483.895 3878.085 3518.220 3878.115 ;
        RECT 3519.275 3878.085 3528.150 3878.115 ;
        RECT 3393.995 3878.000 3396.995 3878.085 ;
        RECT 3445.220 3878.000 3468.605 3878.085 ;
        RECT 3476.815 3878.000 3480.070 3878.085 ;
        RECT 3481.065 3878.000 3518.225 3878.085 ;
        RECT 3518.995 3878.000 3528.150 3878.085 ;
        RECT 3528.815 3878.000 3532.435 3878.160 ;
        RECT 3533.155 3878.085 3558.090 3878.115 ;
        RECT 3533.155 3878.000 3566.645 3878.085 ;
        RECT 3388.230 3798.000 3587.705 3878.000 ;
        RECT 3407.485 3797.880 3413.015 3798.000 ;
        RECT 3418.115 3797.880 3423.725 3798.000 ;
        RECT 3439.250 3797.915 3482.580 3798.000 ;
        RECT 3484.105 3797.840 3518.225 3798.000 ;
        RECT 3518.995 3797.915 3528.055 3798.000 ;
        RECT 3528.815 3797.840 3532.435 3798.000 ;
        RECT 3533.215 3797.895 3566.645 3798.000 ;
        RECT 21.355 3790.000 54.785 3790.105 ;
        RECT 55.565 3790.000 59.185 3790.160 ;
        RECT 59.945 3790.000 69.005 3790.085 ;
        RECT 69.775 3790.000 103.895 3790.160 ;
        RECT 105.420 3790.000 148.750 3790.085 ;
        RECT 164.275 3790.000 169.885 3790.120 ;
        RECT 174.985 3790.000 180.515 3790.120 ;
        RECT 0.295 3710.000 199.770 3790.000 ;
        RECT 21.355 3709.915 54.845 3710.000 ;
        RECT 29.910 3709.885 54.845 3709.915 ;
        RECT 55.565 3709.840 59.185 3710.000 ;
        RECT 59.850 3709.915 69.005 3710.000 ;
        RECT 69.775 3709.915 106.935 3710.000 ;
        RECT 107.930 3709.915 111.185 3710.000 ;
        RECT 119.395 3709.915 142.780 3710.000 ;
        RECT 191.005 3709.915 194.005 3710.000 ;
        RECT 59.850 3709.885 68.725 3709.915 ;
        RECT 69.780 3709.885 104.105 3709.915 ;
        RECT 3483.895 3656.085 3518.220 3656.115 ;
        RECT 3519.275 3656.085 3528.150 3656.115 ;
        RECT 3393.995 3656.000 3396.995 3656.085 ;
        RECT 3445.220 3656.000 3468.605 3656.085 ;
        RECT 3476.815 3656.000 3480.070 3656.085 ;
        RECT 3481.065 3656.000 3518.225 3656.085 ;
        RECT 3518.995 3656.000 3528.150 3656.085 ;
        RECT 3528.815 3656.000 3532.435 3656.160 ;
        RECT 3533.155 3656.085 3558.090 3656.115 ;
        RECT 3533.155 3656.000 3566.645 3656.085 ;
        RECT 3388.230 3576.000 3587.705 3656.000 ;
        RECT 3407.485 3575.880 3413.015 3576.000 ;
        RECT 3418.115 3575.880 3423.725 3576.000 ;
        RECT 3439.250 3575.915 3482.580 3576.000 ;
        RECT 3484.105 3575.840 3518.225 3576.000 ;
        RECT 3518.995 3575.915 3528.055 3576.000 ;
        RECT 3528.815 3575.840 3532.435 3576.000 ;
        RECT 3533.215 3575.895 3566.645 3576.000 ;
        RECT 21.355 3574.000 54.785 3574.105 ;
        RECT 55.565 3574.000 59.185 3574.160 ;
        RECT 59.945 3574.000 69.005 3574.085 ;
        RECT 69.775 3574.000 103.895 3574.160 ;
        RECT 105.420 3574.000 148.750 3574.085 ;
        RECT 164.275 3574.000 169.885 3574.120 ;
        RECT 174.985 3574.000 180.515 3574.120 ;
        RECT 0.295 3494.000 199.770 3574.000 ;
        RECT 21.355 3493.915 54.845 3494.000 ;
        RECT 29.910 3493.885 54.845 3493.915 ;
        RECT 55.565 3493.840 59.185 3494.000 ;
        RECT 59.850 3493.915 69.005 3494.000 ;
        RECT 69.775 3493.915 106.935 3494.000 ;
        RECT 107.930 3493.915 111.185 3494.000 ;
        RECT 119.395 3493.915 142.780 3494.000 ;
        RECT 191.005 3493.915 194.005 3494.000 ;
        RECT 59.850 3493.885 68.725 3493.915 ;
        RECT 69.780 3493.885 104.105 3493.915 ;
        RECT 3483.895 3435.085 3518.220 3435.115 ;
        RECT 3519.275 3435.085 3528.150 3435.115 ;
        RECT 3393.995 3435.000 3396.995 3435.085 ;
        RECT 3445.220 3435.000 3468.605 3435.085 ;
        RECT 3476.815 3435.000 3480.070 3435.085 ;
        RECT 3481.065 3435.000 3518.225 3435.085 ;
        RECT 3518.995 3435.000 3528.150 3435.085 ;
        RECT 3528.815 3435.000 3532.435 3435.160 ;
        RECT 3533.155 3435.085 3558.090 3435.115 ;
        RECT 3533.155 3435.000 3566.645 3435.085 ;
        RECT 21.355 3357.000 54.785 3357.105 ;
        RECT 55.565 3357.000 59.185 3357.160 ;
        RECT 59.945 3357.000 69.005 3357.085 ;
        RECT 69.775 3357.000 103.895 3357.160 ;
        RECT 105.420 3357.000 148.750 3357.085 ;
        RECT 164.275 3357.000 169.885 3357.120 ;
        RECT 174.985 3357.000 180.515 3357.120 ;
        RECT 0.295 3277.000 199.770 3357.000 ;
        RECT 3388.230 3355.000 3587.705 3435.000 ;
        RECT 3407.485 3354.880 3413.015 3355.000 ;
        RECT 3418.115 3354.880 3423.725 3355.000 ;
        RECT 3439.250 3354.915 3482.580 3355.000 ;
        RECT 3484.105 3354.840 3518.225 3355.000 ;
        RECT 3518.995 3354.915 3528.055 3355.000 ;
        RECT 3528.815 3354.840 3532.435 3355.000 ;
        RECT 3533.215 3354.895 3566.645 3355.000 ;
        RECT 21.355 3276.915 54.845 3277.000 ;
        RECT 29.910 3276.885 54.845 3276.915 ;
        RECT 55.565 3276.840 59.185 3277.000 ;
        RECT 59.850 3276.915 69.005 3277.000 ;
        RECT 69.775 3276.915 106.935 3277.000 ;
        RECT 107.930 3276.915 111.185 3277.000 ;
        RECT 119.395 3276.915 142.780 3277.000 ;
        RECT 191.005 3276.915 194.005 3277.000 ;
        RECT 59.850 3276.885 68.725 3276.915 ;
        RECT 69.780 3276.885 104.105 3276.915 ;
        RECT 3483.895 3214.085 3518.220 3214.115 ;
        RECT 3519.275 3214.085 3528.150 3214.115 ;
        RECT 3393.995 3214.000 3396.995 3214.085 ;
        RECT 3445.220 3214.000 3468.605 3214.085 ;
        RECT 3476.815 3214.000 3480.070 3214.085 ;
        RECT 3481.065 3214.000 3518.225 3214.085 ;
        RECT 3518.995 3214.000 3528.150 3214.085 ;
        RECT 3528.815 3214.000 3532.435 3214.160 ;
        RECT 3533.155 3214.085 3558.090 3214.115 ;
        RECT 3533.155 3214.000 3566.645 3214.085 ;
        RECT 21.355 3141.000 54.785 3141.105 ;
        RECT 55.565 3141.000 59.185 3141.160 ;
        RECT 59.945 3141.000 69.005 3141.085 ;
        RECT 69.775 3141.000 103.895 3141.160 ;
        RECT 105.420 3141.000 148.750 3141.085 ;
        RECT 164.275 3141.000 169.885 3141.120 ;
        RECT 174.985 3141.000 180.515 3141.120 ;
        RECT 0.295 3061.000 199.770 3141.000 ;
        RECT 3388.230 3134.000 3587.705 3214.000 ;
        RECT 3407.485 3133.880 3413.015 3134.000 ;
        RECT 3418.115 3133.880 3423.725 3134.000 ;
        RECT 3439.250 3133.915 3482.580 3134.000 ;
        RECT 3484.105 3133.840 3518.225 3134.000 ;
        RECT 3518.995 3133.915 3528.055 3134.000 ;
        RECT 3528.815 3133.840 3532.435 3134.000 ;
        RECT 3533.215 3133.895 3566.645 3134.000 ;
        RECT 21.355 3060.915 54.845 3061.000 ;
        RECT 29.910 3060.885 54.845 3060.915 ;
        RECT 55.565 3060.840 59.185 3061.000 ;
        RECT 59.850 3060.915 69.005 3061.000 ;
        RECT 69.775 3060.915 106.935 3061.000 ;
        RECT 107.930 3060.915 111.185 3061.000 ;
        RECT 119.395 3060.915 142.780 3061.000 ;
        RECT 191.005 3060.915 194.005 3061.000 ;
        RECT 59.850 3060.885 68.725 3060.915 ;
        RECT 69.780 3060.885 104.105 3060.915 ;
        RECT 3483.895 2992.085 3518.220 2992.115 ;
        RECT 3519.275 2992.085 3528.150 2992.115 ;
        RECT 3393.995 2992.000 3396.995 2992.085 ;
        RECT 3445.220 2992.000 3468.605 2992.085 ;
        RECT 3476.815 2992.000 3480.070 2992.085 ;
        RECT 3481.065 2992.000 3518.225 2992.085 ;
        RECT 3518.995 2992.000 3528.150 2992.085 ;
        RECT 3528.815 2992.000 3532.435 2992.160 ;
        RECT 3533.155 2992.085 3558.090 2992.115 ;
        RECT 3533.155 2992.000 3566.645 2992.085 ;
        RECT 21.355 2925.000 54.785 2925.105 ;
        RECT 55.565 2925.000 59.185 2925.160 ;
        RECT 59.945 2925.000 69.005 2925.085 ;
        RECT 69.775 2925.000 103.895 2925.160 ;
        RECT 105.420 2925.000 148.750 2925.085 ;
        RECT 164.275 2925.000 169.885 2925.120 ;
        RECT 174.985 2925.000 180.515 2925.120 ;
        RECT 0.295 2845.000 199.770 2925.000 ;
        RECT 3388.230 2912.000 3587.705 2992.000 ;
        RECT 3407.485 2911.880 3413.015 2912.000 ;
        RECT 3418.115 2911.880 3423.725 2912.000 ;
        RECT 3439.250 2911.915 3482.580 2912.000 ;
        RECT 3484.105 2911.840 3518.225 2912.000 ;
        RECT 3518.995 2911.915 3528.055 2912.000 ;
        RECT 3528.815 2911.840 3532.435 2912.000 ;
        RECT 3533.215 2911.895 3566.645 2912.000 ;
        RECT 21.355 2844.915 54.845 2845.000 ;
        RECT 29.910 2844.885 54.845 2844.915 ;
        RECT 55.565 2844.840 59.185 2845.000 ;
        RECT 59.850 2844.915 69.005 2845.000 ;
        RECT 69.775 2844.915 106.935 2845.000 ;
        RECT 107.930 2844.915 111.185 2845.000 ;
        RECT 119.395 2844.915 142.780 2845.000 ;
        RECT 191.005 2844.915 194.005 2845.000 ;
        RECT 59.850 2844.885 68.725 2844.915 ;
        RECT 69.780 2844.885 104.105 2844.915 ;
        RECT 3483.895 2771.085 3518.220 2771.115 ;
        RECT 3519.275 2771.085 3528.150 2771.115 ;
        RECT 3393.995 2771.000 3396.995 2771.085 ;
        RECT 3445.220 2771.000 3468.605 2771.085 ;
        RECT 3476.815 2771.000 3480.070 2771.085 ;
        RECT 3481.065 2771.000 3518.225 2771.085 ;
        RECT 3518.995 2771.000 3528.150 2771.085 ;
        RECT 3528.815 2771.000 3532.435 2771.160 ;
        RECT 3533.155 2771.085 3558.090 2771.115 ;
        RECT 3533.155 2771.000 3566.645 2771.085 ;
        RECT 21.355 2709.000 54.785 2709.105 ;
        RECT 55.565 2709.000 59.185 2709.160 ;
        RECT 59.945 2709.000 69.005 2709.085 ;
        RECT 69.775 2709.000 103.895 2709.160 ;
        RECT 105.420 2709.000 148.750 2709.085 ;
        RECT 164.275 2709.000 169.885 2709.120 ;
        RECT 174.985 2709.000 180.515 2709.120 ;
        RECT 0.295 2629.000 199.770 2709.000 ;
        RECT 3388.230 2691.000 3587.705 2771.000 ;
        RECT 3407.485 2690.880 3413.015 2691.000 ;
        RECT 3418.115 2690.880 3423.725 2691.000 ;
        RECT 3439.250 2690.915 3482.580 2691.000 ;
        RECT 3484.105 2690.840 3518.225 2691.000 ;
        RECT 3518.995 2690.915 3528.055 2691.000 ;
        RECT 3528.815 2690.840 3532.435 2691.000 ;
        RECT 3533.215 2690.895 3566.645 2691.000 ;
        RECT 21.355 2628.915 54.845 2629.000 ;
        RECT 29.910 2628.885 54.845 2628.915 ;
        RECT 55.565 2628.840 59.185 2629.000 ;
        RECT 59.850 2628.915 69.005 2629.000 ;
        RECT 69.775 2628.915 106.935 2629.000 ;
        RECT 107.930 2628.915 111.185 2629.000 ;
        RECT 119.395 2628.915 142.780 2629.000 ;
        RECT 191.005 2628.915 194.005 2629.000 ;
        RECT 59.850 2628.885 68.725 2628.915 ;
        RECT 69.780 2628.885 104.105 2628.915 ;
        RECT 3389.065 2538.845 3587.695 2549.390 ;
        RECT 3390.035 2537.965 3587.695 2538.845 ;
        RECT 3388.970 2536.955 3587.695 2537.965 ;
        RECT 0.305 2487.680 197.965 2489.855 ;
        RECT 0.305 2486.730 199.030 2487.680 ;
        RECT 0.305 2430.045 197.965 2486.730 ;
        RECT 198.080 2430.045 199.030 2486.730 ;
        RECT 3388.970 2480.270 3389.920 2536.955 ;
        RECT 3390.035 2480.270 3587.695 2536.955 ;
        RECT 3388.970 2479.320 3587.695 2480.270 ;
        RECT 3390.035 2477.145 3587.695 2479.320 ;
        RECT 0.305 2429.035 199.030 2430.045 ;
        RECT 0.305 2428.155 197.965 2429.035 ;
        RECT 0.305 2417.610 198.935 2428.155 ;
        RECT 0.220 2206.240 196.980 2280.755 ;
        RECT 3391.020 2258.245 3587.780 2332.760 ;
        RECT 3390.035 2104.935 3587.695 2115.930 ;
        RECT 3389.000 2103.955 3587.695 2104.935 ;
        RECT 21.355 2070.000 54.785 2070.105 ;
        RECT 55.565 2070.000 59.185 2070.160 ;
        RECT 59.945 2070.000 69.005 2070.085 ;
        RECT 69.775 2070.000 103.895 2070.160 ;
        RECT 105.420 2070.000 148.750 2070.085 ;
        RECT 164.275 2070.000 169.885 2070.120 ;
        RECT 174.985 2070.000 180.515 2070.120 ;
        RECT 0.295 1990.000 199.770 2070.000 ;
        RECT 3389.000 2047.240 3389.890 2103.955 ;
        RECT 3390.035 2047.240 3587.695 2103.955 ;
        RECT 3389.000 2046.350 3587.695 2047.240 ;
        RECT 3390.035 2044.225 3587.695 2046.350 ;
        RECT 21.355 1989.915 54.845 1990.000 ;
        RECT 29.910 1989.885 54.845 1989.915 ;
        RECT 55.565 1989.840 59.185 1990.000 ;
        RECT 59.850 1989.915 69.005 1990.000 ;
        RECT 69.775 1989.915 106.935 1990.000 ;
        RECT 107.930 1989.915 111.185 1990.000 ;
        RECT 119.395 1989.915 142.780 1990.000 ;
        RECT 191.005 1989.915 194.005 1990.000 ;
        RECT 59.850 1989.885 68.725 1989.915 ;
        RECT 69.780 1989.885 104.105 1989.915 ;
        RECT 3483.895 1900.085 3518.220 1900.115 ;
        RECT 3519.275 1900.085 3528.150 1900.115 ;
        RECT 3393.995 1900.000 3396.995 1900.085 ;
        RECT 3445.220 1900.000 3468.605 1900.085 ;
        RECT 3476.815 1900.000 3480.070 1900.085 ;
        RECT 3481.065 1900.000 3518.225 1900.085 ;
        RECT 3518.995 1900.000 3528.150 1900.085 ;
        RECT 3528.815 1900.000 3532.435 1900.160 ;
        RECT 3533.155 1900.085 3558.090 1900.115 ;
        RECT 3533.155 1900.000 3566.645 1900.085 ;
        RECT 21.355 1854.000 54.785 1854.105 ;
        RECT 55.565 1854.000 59.185 1854.160 ;
        RECT 59.945 1854.000 69.005 1854.085 ;
        RECT 69.775 1854.000 103.895 1854.160 ;
        RECT 105.420 1854.000 148.750 1854.085 ;
        RECT 164.275 1854.000 169.885 1854.120 ;
        RECT 174.985 1854.000 180.515 1854.120 ;
        RECT 0.295 1774.000 199.770 1854.000 ;
        RECT 3388.230 1820.000 3587.705 1900.000 ;
        RECT 3407.485 1819.880 3413.015 1820.000 ;
        RECT 3418.115 1819.880 3423.725 1820.000 ;
        RECT 3439.250 1819.915 3482.580 1820.000 ;
        RECT 3484.105 1819.840 3518.225 1820.000 ;
        RECT 3518.995 1819.915 3528.055 1820.000 ;
        RECT 3528.815 1819.840 3532.435 1820.000 ;
        RECT 3533.215 1819.895 3566.645 1820.000 ;
        RECT 21.355 1773.915 54.845 1774.000 ;
        RECT 29.910 1773.885 54.845 1773.915 ;
        RECT 55.565 1773.840 59.185 1774.000 ;
        RECT 59.850 1773.915 69.005 1774.000 ;
        RECT 69.775 1773.915 106.935 1774.000 ;
        RECT 107.930 1773.915 111.185 1774.000 ;
        RECT 119.395 1773.915 142.780 1774.000 ;
        RECT 191.005 1773.915 194.005 1774.000 ;
        RECT 59.850 1773.885 68.725 1773.915 ;
        RECT 69.780 1773.885 104.105 1773.915 ;
        RECT 3483.895 1679.085 3518.220 1679.115 ;
        RECT 3519.275 1679.085 3528.150 1679.115 ;
        RECT 3393.995 1679.000 3396.995 1679.085 ;
        RECT 3445.220 1679.000 3468.605 1679.085 ;
        RECT 3476.815 1679.000 3480.070 1679.085 ;
        RECT 3481.065 1679.000 3518.225 1679.085 ;
        RECT 3518.995 1679.000 3528.150 1679.085 ;
        RECT 3528.815 1679.000 3532.435 1679.160 ;
        RECT 3533.155 1679.085 3558.090 1679.115 ;
        RECT 3533.155 1679.000 3566.645 1679.085 ;
        RECT 21.355 1637.000 54.785 1637.105 ;
        RECT 55.565 1637.000 59.185 1637.160 ;
        RECT 59.945 1637.000 69.005 1637.085 ;
        RECT 69.775 1637.000 103.895 1637.160 ;
        RECT 105.420 1637.000 148.750 1637.085 ;
        RECT 164.275 1637.000 169.885 1637.120 ;
        RECT 174.985 1637.000 180.515 1637.120 ;
        RECT 0.295 1557.000 199.770 1637.000 ;
        RECT 3388.230 1599.000 3587.705 1679.000 ;
        RECT 3407.485 1598.880 3413.015 1599.000 ;
        RECT 3418.115 1598.880 3423.725 1599.000 ;
        RECT 3439.250 1598.915 3482.580 1599.000 ;
        RECT 3484.105 1598.840 3518.225 1599.000 ;
        RECT 3518.995 1598.915 3528.055 1599.000 ;
        RECT 3528.815 1598.840 3532.435 1599.000 ;
        RECT 3533.215 1598.895 3566.645 1599.000 ;
        RECT 21.355 1556.915 54.845 1557.000 ;
        RECT 29.910 1556.885 54.845 1556.915 ;
        RECT 55.565 1556.840 59.185 1557.000 ;
        RECT 59.850 1556.915 69.005 1557.000 ;
        RECT 69.775 1556.915 106.935 1557.000 ;
        RECT 107.930 1556.915 111.185 1557.000 ;
        RECT 119.395 1556.915 142.780 1557.000 ;
        RECT 191.005 1556.915 194.005 1557.000 ;
        RECT 59.850 1556.885 68.725 1556.915 ;
        RECT 69.780 1556.885 104.105 1556.915 ;
        RECT 3483.895 1458.085 3518.220 1458.115 ;
        RECT 3519.275 1458.085 3528.150 1458.115 ;
        RECT 3393.995 1458.000 3396.995 1458.085 ;
        RECT 3445.220 1458.000 3468.605 1458.085 ;
        RECT 3476.815 1458.000 3480.070 1458.085 ;
        RECT 3481.065 1458.000 3518.225 1458.085 ;
        RECT 3518.995 1458.000 3528.150 1458.085 ;
        RECT 3528.815 1458.000 3532.435 1458.160 ;
        RECT 3533.155 1458.085 3558.090 1458.115 ;
        RECT 3533.155 1458.000 3566.645 1458.085 ;
        RECT 21.355 1421.000 54.785 1421.105 ;
        RECT 55.565 1421.000 59.185 1421.160 ;
        RECT 59.945 1421.000 69.005 1421.085 ;
        RECT 69.775 1421.000 103.895 1421.160 ;
        RECT 105.420 1421.000 148.750 1421.085 ;
        RECT 164.275 1421.000 169.885 1421.120 ;
        RECT 174.985 1421.000 180.515 1421.120 ;
        RECT 0.295 1341.000 199.770 1421.000 ;
        RECT 3388.230 1378.000 3587.705 1458.000 ;
        RECT 3407.485 1377.880 3413.015 1378.000 ;
        RECT 3418.115 1377.880 3423.725 1378.000 ;
        RECT 3439.250 1377.915 3482.580 1378.000 ;
        RECT 3484.105 1377.840 3518.225 1378.000 ;
        RECT 3518.995 1377.915 3528.055 1378.000 ;
        RECT 3528.815 1377.840 3532.435 1378.000 ;
        RECT 3533.215 1377.895 3566.645 1378.000 ;
        RECT 21.355 1340.915 54.845 1341.000 ;
        RECT 29.910 1340.885 54.845 1340.915 ;
        RECT 55.565 1340.840 59.185 1341.000 ;
        RECT 59.850 1340.915 69.005 1341.000 ;
        RECT 69.775 1340.915 106.935 1341.000 ;
        RECT 107.930 1340.915 111.185 1341.000 ;
        RECT 119.395 1340.915 142.780 1341.000 ;
        RECT 191.005 1340.915 194.005 1341.000 ;
        RECT 59.850 1340.885 68.725 1340.915 ;
        RECT 69.780 1340.885 104.105 1340.915 ;
        RECT 3483.895 1236.085 3518.220 1236.115 ;
        RECT 3519.275 1236.085 3528.150 1236.115 ;
        RECT 3393.995 1236.000 3396.995 1236.085 ;
        RECT 3445.220 1236.000 3468.605 1236.085 ;
        RECT 3476.815 1236.000 3480.070 1236.085 ;
        RECT 3481.065 1236.000 3518.225 1236.085 ;
        RECT 3518.995 1236.000 3528.150 1236.085 ;
        RECT 3528.815 1236.000 3532.435 1236.160 ;
        RECT 3533.155 1236.085 3558.090 1236.115 ;
        RECT 3533.155 1236.000 3566.645 1236.085 ;
        RECT 21.355 1205.000 54.785 1205.105 ;
        RECT 55.565 1205.000 59.185 1205.160 ;
        RECT 59.945 1205.000 69.005 1205.085 ;
        RECT 69.775 1205.000 103.895 1205.160 ;
        RECT 105.420 1205.000 148.750 1205.085 ;
        RECT 164.275 1205.000 169.885 1205.120 ;
        RECT 174.985 1205.000 180.515 1205.120 ;
        RECT 0.295 1125.000 199.770 1205.000 ;
        RECT 3388.230 1156.000 3587.705 1236.000 ;
        RECT 3407.485 1155.880 3413.015 1156.000 ;
        RECT 3418.115 1155.880 3423.725 1156.000 ;
        RECT 3439.250 1155.915 3482.580 1156.000 ;
        RECT 3484.105 1155.840 3518.225 1156.000 ;
        RECT 3518.995 1155.915 3528.055 1156.000 ;
        RECT 3528.815 1155.840 3532.435 1156.000 ;
        RECT 3533.215 1155.895 3566.645 1156.000 ;
        RECT 21.355 1124.915 54.845 1125.000 ;
        RECT 29.910 1124.885 54.845 1124.915 ;
        RECT 55.565 1124.840 59.185 1125.000 ;
        RECT 59.850 1124.915 69.005 1125.000 ;
        RECT 69.775 1124.915 106.935 1125.000 ;
        RECT 107.930 1124.915 111.185 1125.000 ;
        RECT 119.395 1124.915 142.780 1125.000 ;
        RECT 191.005 1124.915 194.005 1125.000 ;
        RECT 59.850 1124.885 68.725 1124.915 ;
        RECT 69.780 1124.885 104.105 1124.915 ;
        RECT 3483.895 1015.085 3518.220 1015.115 ;
        RECT 3519.275 1015.085 3528.150 1015.115 ;
        RECT 3393.995 1015.000 3396.995 1015.085 ;
        RECT 3445.220 1015.000 3468.605 1015.085 ;
        RECT 3476.815 1015.000 3480.070 1015.085 ;
        RECT 3481.065 1015.000 3518.225 1015.085 ;
        RECT 3518.995 1015.000 3528.150 1015.085 ;
        RECT 3528.815 1015.000 3532.435 1015.160 ;
        RECT 3533.155 1015.085 3558.090 1015.115 ;
        RECT 3533.155 1015.000 3566.645 1015.085 ;
        RECT 21.355 989.000 54.785 989.105 ;
        RECT 55.565 989.000 59.185 989.160 ;
        RECT 59.945 989.000 69.005 989.085 ;
        RECT 69.775 989.000 103.895 989.160 ;
        RECT 105.420 989.000 148.750 989.085 ;
        RECT 164.275 989.000 169.885 989.120 ;
        RECT 174.985 989.000 180.515 989.120 ;
        RECT 0.295 909.000 199.770 989.000 ;
        RECT 3388.230 935.000 3587.705 1015.000 ;
        RECT 3407.485 934.880 3413.015 935.000 ;
        RECT 3418.115 934.880 3423.725 935.000 ;
        RECT 3439.250 934.915 3482.580 935.000 ;
        RECT 3484.105 934.840 3518.225 935.000 ;
        RECT 3518.995 934.915 3528.055 935.000 ;
        RECT 3528.815 934.840 3532.435 935.000 ;
        RECT 3533.215 934.895 3566.645 935.000 ;
        RECT 21.355 908.915 54.845 909.000 ;
        RECT 29.910 908.885 54.845 908.915 ;
        RECT 55.565 908.840 59.185 909.000 ;
        RECT 59.850 908.915 69.005 909.000 ;
        RECT 69.775 908.915 106.935 909.000 ;
        RECT 107.930 908.915 111.185 909.000 ;
        RECT 119.395 908.915 142.780 909.000 ;
        RECT 191.005 908.915 194.005 909.000 ;
        RECT 59.850 908.885 68.725 908.915 ;
        RECT 69.780 908.885 104.105 908.915 ;
        RECT 3483.895 794.085 3518.220 794.115 ;
        RECT 3519.275 794.085 3528.150 794.115 ;
        RECT 3393.995 794.000 3396.995 794.085 ;
        RECT 3445.220 794.000 3468.605 794.085 ;
        RECT 3476.815 794.000 3480.070 794.085 ;
        RECT 3481.065 794.000 3518.225 794.085 ;
        RECT 3518.995 794.000 3528.150 794.085 ;
        RECT 3528.815 794.000 3532.435 794.160 ;
        RECT 3533.155 794.085 3558.090 794.115 ;
        RECT 3533.155 794.000 3566.645 794.085 ;
        RECT 3388.230 714.000 3587.705 794.000 ;
        RECT 3407.485 713.880 3413.015 714.000 ;
        RECT 3418.115 713.880 3423.725 714.000 ;
        RECT 3439.250 713.915 3482.580 714.000 ;
        RECT 3484.105 713.840 3518.225 714.000 ;
        RECT 3518.995 713.915 3528.055 714.000 ;
        RECT 3528.815 713.840 3532.435 714.000 ;
        RECT 3533.215 713.895 3566.645 714.000 ;
        RECT 0.305 621.680 197.965 623.855 ;
        RECT 0.305 620.730 199.030 621.680 ;
        RECT 0.305 564.045 197.965 620.730 ;
        RECT 198.080 564.045 199.030 620.730 ;
        RECT 3483.895 572.085 3518.220 572.115 ;
        RECT 3519.275 572.085 3528.150 572.115 ;
        RECT 3393.995 572.000 3396.995 572.085 ;
        RECT 3445.220 572.000 3468.605 572.085 ;
        RECT 3476.815 572.000 3480.070 572.085 ;
        RECT 3481.065 572.000 3518.225 572.085 ;
        RECT 3518.995 572.000 3528.150 572.085 ;
        RECT 3528.815 572.000 3532.435 572.160 ;
        RECT 3533.155 572.085 3558.090 572.115 ;
        RECT 3533.155 572.000 3566.645 572.085 ;
        RECT 0.305 563.035 199.030 564.045 ;
        RECT 0.305 562.155 197.965 563.035 ;
        RECT 0.305 551.610 198.935 562.155 ;
        RECT 3388.230 492.000 3587.705 572.000 ;
        RECT 3407.485 491.880 3413.015 492.000 ;
        RECT 3418.115 491.880 3423.725 492.000 ;
        RECT 3439.250 491.915 3482.580 492.000 ;
        RECT 3484.105 491.840 3518.225 492.000 ;
        RECT 3518.995 491.915 3528.055 492.000 ;
        RECT 3528.815 491.840 3532.435 492.000 ;
        RECT 3533.215 491.895 3566.645 492.000 ;
        RECT 0.220 340.240 196.980 414.755 ;
        RECT 398.350 198.110 456.935 199.000 ;
        RECT 398.350 197.965 399.240 198.110 ;
        RECT 455.955 197.965 456.935 198.110 ;
        RECT 396.225 0.305 467.930 197.965 ;
        RECT 663.000 98.605 738.000 199.815 ;
        RECT 932.000 194.005 1012.000 199.770 ;
        RECT 932.000 191.005 1012.085 194.005 ;
        RECT 932.000 180.515 1012.000 191.005 ;
        RECT 931.880 174.985 1012.000 180.515 ;
        RECT 932.000 169.885 1012.000 174.985 ;
        RECT 931.880 164.275 1012.000 169.885 ;
        RECT 932.000 148.750 1012.000 164.275 ;
        RECT 931.915 142.780 1012.000 148.750 ;
        RECT 931.915 119.395 1012.085 142.780 ;
        RECT 931.915 111.185 1012.000 119.395 ;
        RECT 931.915 107.930 1012.085 111.185 ;
        RECT 931.915 106.935 1012.000 107.930 ;
        RECT 931.915 105.420 1012.085 106.935 ;
        RECT 932.000 104.105 1012.085 105.420 ;
        RECT 932.000 103.895 1012.115 104.105 ;
        RECT 663.000 69.775 738.265 98.605 ;
        RECT 931.840 69.780 1012.115 103.895 ;
        RECT 931.840 69.775 1012.085 69.780 ;
        RECT 663.000 59.185 738.000 69.775 ;
        RECT 932.000 69.005 1012.000 69.775 ;
        RECT 931.915 68.725 1012.085 69.005 ;
        RECT 931.915 59.945 1012.115 68.725 ;
        RECT 932.000 59.850 1012.115 59.945 ;
        RECT 932.000 59.185 1012.000 59.850 ;
        RECT 662.840 55.565 738.160 59.185 ;
        RECT 931.840 55.565 1012.160 59.185 ;
        RECT 663.000 0.780 738.000 55.565 ;
        RECT 932.000 54.845 1012.000 55.565 ;
        RECT 932.000 54.785 1012.115 54.845 ;
        RECT 931.895 29.910 1012.115 54.785 ;
        RECT 931.895 21.355 1012.085 29.910 ;
        RECT 932.000 0.295 1012.000 21.355 ;
        RECT 1206.245 0.220 1280.760 196.980 ;
        RECT 1475.000 194.005 1555.000 199.770 ;
        RECT 1749.000 194.005 1829.000 199.770 ;
        RECT 2023.000 194.005 2103.000 199.770 ;
        RECT 2297.000 194.005 2377.000 199.770 ;
        RECT 2571.000 194.005 2651.000 199.770 ;
        RECT 2849.350 198.110 2907.935 199.000 ;
        RECT 2849.350 197.965 2850.240 198.110 ;
        RECT 2906.955 197.965 2907.935 198.110 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.270 198.080 ;
        RECT 3175.955 197.965 3176.965 198.080 ;
        RECT 3177.845 197.965 3188.390 198.935 ;
        RECT 1475.000 191.005 1555.085 194.005 ;
        RECT 1749.000 191.005 1829.085 194.005 ;
        RECT 2023.000 191.005 2103.085 194.005 ;
        RECT 2297.000 191.005 2377.085 194.005 ;
        RECT 2571.000 191.005 2651.085 194.005 ;
        RECT 1475.000 180.515 1555.000 191.005 ;
        RECT 1749.000 180.515 1829.000 191.005 ;
        RECT 2023.000 180.515 2103.000 191.005 ;
        RECT 2297.000 180.515 2377.000 191.005 ;
        RECT 2571.000 180.515 2651.000 191.005 ;
        RECT 1474.880 174.985 1555.000 180.515 ;
        RECT 1748.880 174.985 1829.000 180.515 ;
        RECT 2022.880 174.985 2103.000 180.515 ;
        RECT 2296.880 174.985 2377.000 180.515 ;
        RECT 2570.880 174.985 2651.000 180.515 ;
        RECT 1475.000 169.885 1555.000 174.985 ;
        RECT 1749.000 169.885 1829.000 174.985 ;
        RECT 2023.000 169.885 2103.000 174.985 ;
        RECT 2297.000 169.885 2377.000 174.985 ;
        RECT 2571.000 169.885 2651.000 174.985 ;
        RECT 1474.880 164.275 1555.000 169.885 ;
        RECT 1748.880 164.275 1829.000 169.885 ;
        RECT 2022.880 164.275 2103.000 169.885 ;
        RECT 2296.880 164.275 2377.000 169.885 ;
        RECT 2570.880 164.275 2651.000 169.885 ;
        RECT 1475.000 148.750 1555.000 164.275 ;
        RECT 1749.000 148.750 1829.000 164.275 ;
        RECT 2023.000 148.750 2103.000 164.275 ;
        RECT 2297.000 148.750 2377.000 164.275 ;
        RECT 2571.000 148.750 2651.000 164.275 ;
        RECT 1474.915 142.780 1555.000 148.750 ;
        RECT 1748.915 142.780 1829.000 148.750 ;
        RECT 2022.915 142.780 2103.000 148.750 ;
        RECT 2296.915 142.780 2377.000 148.750 ;
        RECT 2570.915 142.780 2651.000 148.750 ;
        RECT 1474.915 119.395 1555.085 142.780 ;
        RECT 1748.915 119.395 1829.085 142.780 ;
        RECT 2022.915 119.395 2103.085 142.780 ;
        RECT 2296.915 119.395 2377.085 142.780 ;
        RECT 2570.915 119.395 2651.085 142.780 ;
        RECT 1474.915 111.185 1555.000 119.395 ;
        RECT 1748.915 111.185 1829.000 119.395 ;
        RECT 2022.915 111.185 2103.000 119.395 ;
        RECT 2296.915 111.185 2377.000 119.395 ;
        RECT 2570.915 111.185 2651.000 119.395 ;
        RECT 1474.915 107.930 1555.085 111.185 ;
        RECT 1748.915 107.930 1829.085 111.185 ;
        RECT 2022.915 107.930 2103.085 111.185 ;
        RECT 2296.915 107.930 2377.085 111.185 ;
        RECT 2570.915 107.930 2651.085 111.185 ;
        RECT 1474.915 106.935 1555.000 107.930 ;
        RECT 1748.915 106.935 1829.000 107.930 ;
        RECT 2022.915 106.935 2103.000 107.930 ;
        RECT 2296.915 106.935 2377.000 107.930 ;
        RECT 2570.915 106.935 2651.000 107.930 ;
        RECT 1474.915 105.420 1555.085 106.935 ;
        RECT 1748.915 105.420 1829.085 106.935 ;
        RECT 2022.915 105.420 2103.085 106.935 ;
        RECT 2296.915 105.420 2377.085 106.935 ;
        RECT 2570.915 105.420 2651.085 106.935 ;
        RECT 1475.000 104.105 1555.085 105.420 ;
        RECT 1749.000 104.105 1829.085 105.420 ;
        RECT 2023.000 104.105 2103.085 105.420 ;
        RECT 2297.000 104.105 2377.085 105.420 ;
        RECT 2571.000 104.105 2651.085 105.420 ;
        RECT 1475.000 103.895 1555.115 104.105 ;
        RECT 1749.000 103.895 1829.115 104.105 ;
        RECT 2023.000 103.895 2103.115 104.105 ;
        RECT 2297.000 103.895 2377.115 104.105 ;
        RECT 2571.000 103.895 2651.115 104.105 ;
        RECT 1474.840 69.780 1555.115 103.895 ;
        RECT 1748.840 69.780 1829.115 103.895 ;
        RECT 2022.840 69.780 2103.115 103.895 ;
        RECT 2296.840 69.780 2377.115 103.895 ;
        RECT 2570.840 69.780 2651.115 103.895 ;
        RECT 1474.840 69.775 1555.085 69.780 ;
        RECT 1748.840 69.775 1829.085 69.780 ;
        RECT 2022.840 69.775 2103.085 69.780 ;
        RECT 2296.840 69.775 2377.085 69.780 ;
        RECT 2570.840 69.775 2651.085 69.780 ;
        RECT 1475.000 69.005 1555.000 69.775 ;
        RECT 1749.000 69.005 1829.000 69.775 ;
        RECT 2023.000 69.005 2103.000 69.775 ;
        RECT 2297.000 69.005 2377.000 69.775 ;
        RECT 2571.000 69.005 2651.000 69.775 ;
        RECT 1474.915 68.725 1555.085 69.005 ;
        RECT 1748.915 68.725 1829.085 69.005 ;
        RECT 2022.915 68.725 2103.085 69.005 ;
        RECT 2296.915 68.725 2377.085 69.005 ;
        RECT 2570.915 68.725 2651.085 69.005 ;
        RECT 1474.915 59.945 1555.115 68.725 ;
        RECT 1748.915 59.945 1829.115 68.725 ;
        RECT 2022.915 59.945 2103.115 68.725 ;
        RECT 2296.915 59.945 2377.115 68.725 ;
        RECT 2570.915 59.945 2651.115 68.725 ;
        RECT 1475.000 59.850 1555.115 59.945 ;
        RECT 1749.000 59.850 1829.115 59.945 ;
        RECT 2023.000 59.850 2103.115 59.945 ;
        RECT 2297.000 59.850 2377.115 59.945 ;
        RECT 2571.000 59.850 2651.115 59.945 ;
        RECT 1475.000 59.185 1555.000 59.850 ;
        RECT 1749.000 59.185 1829.000 59.850 ;
        RECT 2023.000 59.185 2103.000 59.850 ;
        RECT 2297.000 59.185 2377.000 59.850 ;
        RECT 2571.000 59.185 2651.000 59.850 ;
        RECT 1474.840 55.565 1555.160 59.185 ;
        RECT 1748.840 55.565 1829.160 59.185 ;
        RECT 2022.840 55.565 2103.160 59.185 ;
        RECT 2296.840 55.565 2377.160 59.185 ;
        RECT 2570.840 55.565 2651.160 59.185 ;
        RECT 1475.000 54.845 1555.000 55.565 ;
        RECT 1749.000 54.845 1829.000 55.565 ;
        RECT 2023.000 54.845 2103.000 55.565 ;
        RECT 2297.000 54.845 2377.000 55.565 ;
        RECT 2571.000 54.845 2651.000 55.565 ;
        RECT 1475.000 54.785 1555.115 54.845 ;
        RECT 1749.000 54.785 1829.115 54.845 ;
        RECT 2023.000 54.785 2103.115 54.845 ;
        RECT 2297.000 54.785 2377.115 54.845 ;
        RECT 2571.000 54.785 2651.115 54.845 ;
        RECT 1474.895 29.910 1555.115 54.785 ;
        RECT 1748.895 29.910 1829.115 54.785 ;
        RECT 2022.895 29.910 2103.115 54.785 ;
        RECT 2296.895 29.910 2377.115 54.785 ;
        RECT 2570.895 29.910 2651.115 54.785 ;
        RECT 1474.895 21.355 1555.085 29.910 ;
        RECT 1748.895 21.355 1829.085 29.910 ;
        RECT 2022.895 21.355 2103.085 29.910 ;
        RECT 2296.895 21.355 2377.085 29.910 ;
        RECT 2570.895 21.355 2651.085 29.910 ;
        RECT 1475.000 0.295 1555.000 21.355 ;
        RECT 1749.000 0.295 1829.000 21.355 ;
        RECT 2023.000 0.295 2103.000 21.355 ;
        RECT 2297.000 0.295 2377.000 21.355 ;
        RECT 2571.000 0.295 2651.000 21.355 ;
        RECT 2847.225 0.305 2918.930 197.965 ;
        RECT 3116.145 0.305 3188.390 197.965 ;
      LAYER met1 ;
        RECT 379.250 5034.255 445.440 5036.855 ;
        RECT 619.250 5034.255 685.440 5036.855 ;
        RECT 859.250 5034.255 925.440 5036.855 ;
        RECT 1147.185 4990.035 1219.915 5187.725 ;
        RECT 1404.185 4990.035 1476.915 5187.725 ;
        RECT 1697.185 4990.035 1770.620 5187.725 ;
        RECT 2128.250 5034.255 2194.440 5036.855 ;
        RECT 2375.250 5034.255 2441.440 5036.855 ;
        RECT 2633.250 5034.255 2699.440 5036.855 ;
        RECT 2878.185 4990.035 2951.620 5187.725 ;
        RECT 3139.250 5034.255 3205.440 5036.855 ;
        RECT 1150.625 4989.130 1155.855 4990.035 ;
        RECT 1159.035 4989.920 1160.350 4990.035 ;
        POLYGON 1160.350 4990.035 1160.465 4989.920 1160.350 4989.920 ;
        POLYGON 1216.540 4990.035 1216.540 4989.920 1216.425 4989.920 ;
        RECT 1216.540 4989.920 1217.680 4990.035 ;
        RECT 1159.035 4988.970 1217.680 4989.920 ;
        RECT 1407.625 4989.130 1412.855 4990.035 ;
        RECT 1416.035 4989.920 1417.350 4990.035 ;
        POLYGON 1417.350 4990.035 1417.465 4989.920 1417.350 4989.920 ;
        POLYGON 1473.540 4990.035 1473.540 4989.920 1473.425 4989.920 ;
        RECT 1473.540 4989.920 1474.680 4990.035 ;
        RECT 1416.035 4988.970 1474.680 4989.920 ;
        RECT 1709.035 4989.920 1710.350 4990.035 ;
        POLYGON 1710.350 4990.035 1710.465 4989.920 1710.350 4989.920 ;
        POLYGON 1766.540 4990.035 1766.540 4989.920 1766.425 4989.920 ;
        RECT 1766.540 4989.920 1767.680 4990.035 ;
        RECT 1709.035 4988.970 1767.680 4989.920 ;
        RECT 2890.035 4989.920 2891.350 4990.035 ;
        POLYGON 2891.350 4990.035 2891.465 4989.920 2891.350 4989.920 ;
        POLYGON 2947.540 4990.035 2947.540 4989.920 2947.425 4989.920 ;
        RECT 2947.540 4989.920 2948.680 4990.035 ;
        RECT 2890.035 4988.970 2948.680 4989.920 ;
      LAYER met1 ;
        RECT 2928.890 4982.260 2929.210 4982.320 ;
        RECT 3373.710 4982.260 3374.030 4982.320 ;
        RECT 2928.890 4982.120 3374.030 4982.260 ;
        RECT 2928.890 4982.060 2929.210 4982.120 ;
        RECT 3373.710 4982.060 3374.030 4982.120 ;
        RECT 211.210 4981.920 211.530 4981.980 ;
        RECT 1697.470 4981.920 1697.790 4981.980 ;
        RECT 3367.730 4981.920 3368.050 4981.980 ;
        RECT 211.210 4981.780 3368.050 4981.920 ;
        RECT 211.210 4981.720 211.530 4981.780 ;
        RECT 1697.470 4981.720 1697.790 4981.780 ;
        RECT 3367.730 4981.720 3368.050 4981.780 ;
        RECT 224.550 4950.640 224.870 4950.700 ;
        RECT 3368.190 4950.640 3368.510 4950.700 ;
        RECT 224.550 4950.500 3368.510 4950.640 ;
        RECT 224.550 4950.440 224.870 4950.500 ;
        RECT 3368.190 4950.440 3368.510 4950.500 ;
        RECT 211.670 4950.300 211.990 4950.360 ;
        RECT 3367.270 4950.300 3367.590 4950.360 ;
        RECT 211.670 4950.160 3367.590 4950.300 ;
        RECT 211.670 4950.100 211.990 4950.160 ;
        RECT 3367.270 4950.100 3367.590 4950.160 ;
      LAYER met1 ;
        RECT 151.145 4780.250 153.745 4846.440 ;
        RECT 3390.035 4791.375 3587.725 4794.815 ;
        RECT 3389.130 4786.145 3587.725 4791.375 ;
        RECT 3390.035 4782.965 3587.725 4786.145 ;
        RECT 3388.970 4781.650 3587.725 4782.965 ;
        RECT 3388.970 4725.460 3389.920 4781.650 ;
        POLYGON 3389.920 4781.650 3390.035 4781.650 3389.920 4781.535 ;
        POLYGON 3389.920 4725.575 3390.035 4725.460 3389.920 4725.460 ;
        RECT 3390.035 4725.460 3587.725 4781.650 ;
        RECT 3388.970 4724.320 3587.725 4725.460 ;
        RECT 3390.035 4722.085 3587.725 4724.320 ;
        RECT 122.615 4646.935 204.885 4650.935 ;
        POLYGON 204.885 4650.935 208.885 4646.935 204.885 4646.935 ;
        RECT 122.615 4641.200 208.885 4646.935 ;
        RECT 0.160 4621.565 197.965 4640.000 ;
        RECT 198.780 4621.565 208.885 4641.200 ;
        RECT 0.160 4585.925 208.885 4621.565 ;
        RECT 0.160 4581.655 198.000 4585.925 ;
        RECT 0.160 4565.120 197.965 4581.655 ;
        RECT 3390.035 4515.345 3587.840 4531.880 ;
        RECT 3390.000 4511.075 3587.840 4515.345 ;
        RECT 3379.115 4475.435 3587.840 4511.075 ;
        RECT 3379.115 4455.800 3389.220 4475.435 ;
        RECT 3390.035 4457.000 3587.840 4475.435 ;
        RECT 3379.115 4450.065 3465.385 4455.800 ;
        POLYGON 3379.115 4450.065 3383.115 4450.065 3383.115 4446.065 ;
        RECT 3383.115 4446.065 3465.385 4450.065 ;
        RECT 0.275 4424.680 197.965 4426.915 ;
        RECT 0.275 4423.540 199.030 4424.680 ;
        RECT 0.275 4367.350 197.965 4423.540 ;
        POLYGON 197.965 4423.540 198.080 4423.540 198.080 4423.425 ;
        POLYGON 198.080 4367.465 198.080 4367.350 197.965 4367.350 ;
        RECT 198.080 4367.350 199.030 4423.540 ;
        RECT 0.275 4366.035 199.030 4367.350 ;
        RECT 0.275 4362.855 197.965 4366.035 ;
        RECT 0.275 4357.625 198.870 4362.855 ;
        RECT 0.275 4354.185 197.965 4357.625 ;
        RECT 3445.190 4315.000 3468.635 4315.115 ;
        RECT 3477.750 4315.000 3479.480 4315.145 ;
        RECT 3483.895 4315.000 3518.220 4315.115 ;
        RECT 3519.275 4315.000 3558.090 4315.115 ;
      LAYER met1 ;
        RECT 212.130 4306.000 212.450 4306.060 ;
        RECT 220.870 4306.000 221.190 4306.060 ;
        RECT 212.130 4305.860 221.190 4306.000 ;
        RECT 212.130 4305.800 212.450 4305.860 ;
        RECT 220.870 4305.800 221.190 4305.860 ;
        RECT 3367.730 4295.800 3368.050 4295.860 ;
        RECT 3376.930 4295.800 3377.250 4295.860 ;
        RECT 3367.730 4295.660 3377.250 4295.800 ;
        RECT 3367.730 4295.600 3368.050 4295.660 ;
        RECT 3376.930 4295.600 3377.250 4295.660 ;
        RECT 3368.190 4280.500 3368.510 4280.560 ;
        RECT 3376.930 4280.500 3377.250 4280.560 ;
        RECT 3368.190 4280.360 3377.250 4280.500 ;
        RECT 3368.190 4280.300 3368.510 4280.360 ;
        RECT 3376.930 4280.300 3377.250 4280.360 ;
        RECT 3367.270 4248.540 3367.590 4248.600 ;
        RECT 3376.930 4248.540 3377.250 4248.600 ;
        RECT 3367.270 4248.400 3377.250 4248.540 ;
        RECT 3367.270 4248.340 3367.590 4248.400 ;
        RECT 3376.930 4248.340 3377.250 4248.400 ;
      LAYER met1 ;
        RECT 3381.155 4235.000 3588.000 4315.000 ;
        RECT 3407.485 4234.885 3413.015 4235.000 ;
        RECT 3418.120 4234.885 3423.725 4235.000 ;
        RECT 3439.220 4234.940 3482.580 4235.000 ;
        RECT 3439.220 4234.885 3460.930 4234.940 ;
        POLYGON 3460.930 4234.940 3460.985 4234.940 3460.930 4234.885 ;
        RECT 3483.895 4234.855 3518.220 4235.000 ;
        RECT 3519.275 4234.855 3558.090 4235.000 ;
        RECT 3566.900 4234.980 3568.975 4235.000 ;
        RECT 0.275 4212.680 197.965 4215.620 ;
        RECT 0.275 4211.540 199.030 4212.680 ;
        RECT 0.275 4155.350 197.965 4211.540 ;
        POLYGON 197.965 4211.540 198.080 4211.540 198.080 4211.425 ;
        POLYGON 198.080 4155.465 198.080 4155.350 197.965 4155.350 ;
        RECT 198.080 4155.350 199.030 4211.540 ;
        RECT 0.275 4154.035 199.030 4155.350 ;
        RECT 0.275 4142.185 197.965 4154.035 ;
        RECT 3390.035 4090.375 3587.725 4093.815 ;
        RECT 3389.130 4085.145 3587.725 4090.375 ;
        RECT 3390.035 4081.965 3587.725 4085.145 ;
        RECT 3388.970 4080.650 3587.725 4081.965 ;
        RECT 3388.970 4024.460 3389.920 4080.650 ;
        POLYGON 3389.920 4080.650 3390.035 4080.650 3389.920 4080.535 ;
        POLYGON 3389.920 4024.575 3390.035 4024.460 3389.920 4024.460 ;
        RECT 3390.035 4024.460 3587.725 4080.650 ;
        RECT 3388.970 4023.320 3587.725 4024.460 ;
        RECT 3390.035 4021.085 3587.725 4023.320 ;
      LAYER met1 ;
        RECT 3376.470 4019.040 3376.790 4019.100 ;
        RECT 3387.970 4019.040 3388.290 4019.100 ;
        RECT 3376.470 4018.900 3388.290 4019.040 ;
        RECT 3376.470 4018.840 3376.790 4018.900 ;
        RECT 3387.970 4018.840 3388.290 4018.900 ;
      LAYER met1 ;
        RECT 19.025 4006.000 21.100 4006.020 ;
        RECT 29.910 4006.000 68.725 4006.145 ;
        RECT 69.780 4006.000 104.105 4006.145 ;
        POLYGON 127.070 4006.115 127.070 4006.060 127.015 4006.060 ;
        RECT 127.070 4006.060 148.780 4006.115 ;
        RECT 105.420 4006.000 148.780 4006.060 ;
        RECT 164.275 4006.000 169.880 4006.115 ;
        RECT 174.985 4006.000 180.515 4006.115 ;
        RECT 0.000 3926.000 206.845 4006.000 ;
      LAYER met1 ;
        RECT 211.210 4005.100 211.530 4005.160 ;
        RECT 213.050 4005.100 213.370 4005.160 ;
        RECT 211.210 4004.960 213.370 4005.100 ;
        RECT 211.210 4004.900 211.530 4004.960 ;
        RECT 213.050 4004.900 213.370 4004.960 ;
        RECT 208.910 3992.860 209.230 3992.920 ;
        RECT 211.670 3992.860 211.990 3992.920 ;
        RECT 208.910 3992.720 211.990 3992.860 ;
        RECT 208.910 3992.660 209.230 3992.720 ;
        RECT 211.670 3992.660 211.990 3992.720 ;
        RECT 208.910 3960.560 209.230 3960.620 ;
        RECT 212.130 3960.560 212.450 3960.620 ;
        RECT 208.910 3960.420 212.450 3960.560 ;
        RECT 208.910 3960.360 209.230 3960.420 ;
        RECT 212.130 3960.360 212.450 3960.420 ;
        RECT 208.910 3945.600 209.230 3945.660 ;
        RECT 213.050 3945.600 213.370 3945.660 ;
        RECT 208.910 3945.460 213.370 3945.600 ;
        RECT 208.910 3945.400 209.230 3945.460 ;
        RECT 213.050 3945.400 213.370 3945.460 ;
      LAYER met1 ;
        RECT 29.910 3925.885 68.725 3926.000 ;
        RECT 69.780 3925.885 104.105 3926.000 ;
        RECT 108.520 3925.855 110.250 3926.000 ;
        RECT 119.365 3925.885 142.810 3926.000 ;
        RECT 3445.190 3878.000 3468.635 3878.115 ;
        RECT 3477.750 3878.000 3479.480 3878.145 ;
        RECT 3483.895 3878.000 3518.220 3878.115 ;
        RECT 3519.275 3878.000 3558.090 3878.115 ;
      LAYER met1 ;
        RECT 3367.730 3864.000 3368.050 3864.060 ;
        RECT 3376.930 3864.000 3377.250 3864.060 ;
        RECT 3367.730 3863.860 3377.250 3864.000 ;
        RECT 3367.730 3863.800 3368.050 3863.860 ;
        RECT 3376.930 3863.800 3377.250 3863.860 ;
        RECT 3368.190 3848.360 3368.510 3848.420 ;
        RECT 3369.570 3848.360 3369.890 3848.420 ;
        RECT 3376.930 3848.360 3377.250 3848.420 ;
        RECT 3368.190 3848.220 3377.250 3848.360 ;
        RECT 3368.190 3848.160 3368.510 3848.220 ;
        RECT 3369.570 3848.160 3369.890 3848.220 ;
        RECT 3376.930 3848.160 3377.250 3848.220 ;
        RECT 3376.010 3838.160 3376.330 3838.220 ;
        RECT 3376.930 3838.160 3377.250 3838.220 ;
        RECT 3376.010 3838.020 3377.250 3838.160 ;
        RECT 3376.010 3837.960 3376.330 3838.020 ;
        RECT 3376.930 3837.960 3377.250 3838.020 ;
        RECT 3367.270 3806.540 3367.590 3806.600 ;
        RECT 3370.030 3806.540 3370.350 3806.600 ;
        RECT 3376.930 3806.540 3377.250 3806.600 ;
        RECT 3367.270 3806.400 3377.250 3806.540 ;
        RECT 3367.270 3806.340 3367.590 3806.400 ;
        RECT 3370.030 3806.340 3370.350 3806.400 ;
        RECT 3376.930 3806.340 3377.250 3806.400 ;
        RECT 3376.010 3801.100 3376.330 3801.160 ;
        RECT 3376.930 3801.100 3377.250 3801.160 ;
        RECT 3376.010 3800.960 3377.250 3801.100 ;
        RECT 3376.010 3800.900 3376.330 3800.960 ;
        RECT 3376.930 3800.900 3377.250 3800.960 ;
      LAYER met1 ;
        RECT 3381.155 3798.000 3588.000 3878.000 ;
        RECT 3407.485 3797.885 3413.015 3798.000 ;
        RECT 3418.120 3797.885 3423.725 3798.000 ;
        RECT 3439.220 3797.940 3482.580 3798.000 ;
        RECT 3439.220 3797.885 3460.930 3797.940 ;
        POLYGON 3460.930 3797.940 3460.985 3797.940 3460.930 3797.885 ;
        RECT 3483.895 3797.855 3518.220 3798.000 ;
        RECT 3519.275 3797.855 3558.090 3798.000 ;
        RECT 3566.900 3797.980 3568.975 3798.000 ;
        RECT 19.025 3790.000 21.100 3790.020 ;
        RECT 29.910 3790.000 68.725 3790.145 ;
        RECT 69.780 3790.000 104.105 3790.145 ;
        POLYGON 127.070 3790.115 127.070 3790.060 127.015 3790.060 ;
        RECT 127.070 3790.060 148.780 3790.115 ;
        RECT 105.420 3790.000 148.780 3790.060 ;
        RECT 164.275 3790.000 169.880 3790.115 ;
        RECT 174.985 3790.000 180.515 3790.115 ;
        RECT 0.000 3710.000 206.845 3790.000 ;
      LAYER met1 ;
        RECT 208.910 3781.380 209.230 3781.440 ;
        RECT 211.670 3781.380 211.990 3781.440 ;
        RECT 213.050 3781.380 213.370 3781.440 ;
        RECT 208.910 3781.240 213.370 3781.380 ;
        RECT 208.910 3781.180 209.230 3781.240 ;
        RECT 211.670 3781.180 211.990 3781.240 ;
        RECT 213.050 3781.180 213.370 3781.240 ;
        RECT 208.910 3741.600 209.230 3741.660 ;
        RECT 212.590 3741.600 212.910 3741.660 ;
        RECT 208.910 3741.460 212.910 3741.600 ;
        RECT 208.910 3741.400 209.230 3741.460 ;
        RECT 212.590 3741.400 212.910 3741.460 ;
        RECT 208.910 3724.260 209.230 3724.320 ;
        RECT 212.130 3724.260 212.450 3724.320 ;
        RECT 213.510 3724.260 213.830 3724.320 ;
        RECT 208.910 3724.120 213.830 3724.260 ;
        RECT 208.910 3724.060 209.230 3724.120 ;
        RECT 212.130 3724.060 212.450 3724.120 ;
        RECT 213.510 3724.060 213.830 3724.120 ;
      LAYER met1 ;
        RECT 29.910 3709.885 68.725 3710.000 ;
        RECT 69.780 3709.885 104.105 3710.000 ;
        RECT 108.520 3709.855 110.250 3710.000 ;
        RECT 119.365 3709.885 142.810 3710.000 ;
        RECT 3445.190 3656.000 3468.635 3656.115 ;
        RECT 3477.750 3656.000 3479.480 3656.145 ;
        RECT 3483.895 3656.000 3518.220 3656.115 ;
        RECT 3519.275 3656.000 3558.090 3656.115 ;
      LAYER met1 ;
        RECT 3367.730 3641.980 3368.050 3642.040 ;
        RECT 3376.930 3641.980 3377.250 3642.040 ;
        RECT 3367.730 3641.840 3377.250 3641.980 ;
        RECT 3367.730 3641.780 3368.050 3641.840 ;
        RECT 3376.930 3641.780 3377.250 3641.840 ;
        RECT 3369.570 3626.340 3369.890 3626.400 ;
        RECT 3376.930 3626.340 3377.250 3626.400 ;
        RECT 3369.570 3626.200 3377.250 3626.340 ;
        RECT 3369.570 3626.140 3369.890 3626.200 ;
        RECT 3376.930 3626.140 3377.250 3626.200 ;
        RECT 3368.190 3589.280 3368.510 3589.340 ;
        RECT 3370.030 3589.280 3370.350 3589.340 ;
        RECT 3376.930 3589.280 3377.250 3589.340 ;
        RECT 3368.190 3589.140 3377.250 3589.280 ;
        RECT 3368.190 3589.080 3368.510 3589.140 ;
        RECT 3370.030 3589.080 3370.350 3589.140 ;
        RECT 3376.930 3589.080 3377.250 3589.140 ;
      LAYER met1 ;
        RECT 3381.155 3576.000 3588.000 3656.000 ;
        RECT 3407.485 3575.885 3413.015 3576.000 ;
        RECT 3418.120 3575.885 3423.725 3576.000 ;
        RECT 3439.220 3575.940 3482.580 3576.000 ;
        RECT 3439.220 3575.885 3460.930 3575.940 ;
        POLYGON 3460.930 3575.940 3460.985 3575.940 3460.930 3575.885 ;
        RECT 3483.895 3575.855 3518.220 3576.000 ;
        RECT 3519.275 3575.855 3558.090 3576.000 ;
        RECT 3566.900 3575.980 3568.975 3576.000 ;
        RECT 19.025 3574.000 21.100 3574.020 ;
        RECT 29.910 3574.000 68.725 3574.145 ;
        RECT 69.780 3574.000 104.105 3574.145 ;
        POLYGON 127.070 3574.115 127.070 3574.060 127.015 3574.060 ;
        RECT 127.070 3574.060 148.780 3574.115 ;
        RECT 105.420 3574.000 148.780 3574.060 ;
        RECT 164.275 3574.000 169.880 3574.115 ;
        RECT 174.985 3574.000 180.515 3574.115 ;
        RECT 0.000 3494.000 206.845 3574.000 ;
      LAYER met1 ;
        RECT 208.910 3565.480 209.230 3565.540 ;
        RECT 213.050 3565.480 213.370 3565.540 ;
        RECT 208.910 3565.340 213.370 3565.480 ;
        RECT 208.910 3565.280 209.230 3565.340 ;
        RECT 213.050 3565.280 213.370 3565.340 ;
        RECT 208.910 3524.000 209.230 3524.060 ;
        RECT 212.590 3524.000 212.910 3524.060 ;
        RECT 208.910 3523.860 212.910 3524.000 ;
        RECT 208.910 3523.800 209.230 3523.860 ;
        RECT 212.590 3523.800 212.910 3523.860 ;
        RECT 208.910 3508.360 209.230 3508.420 ;
        RECT 212.130 3508.360 212.450 3508.420 ;
        RECT 208.910 3508.220 212.450 3508.360 ;
        RECT 208.910 3508.160 209.230 3508.220 ;
        RECT 212.130 3508.160 212.450 3508.220 ;
      LAYER met1 ;
        RECT 29.910 3493.885 68.725 3494.000 ;
        RECT 69.780 3493.885 104.105 3494.000 ;
        RECT 108.520 3493.855 110.250 3494.000 ;
        RECT 119.365 3493.885 142.810 3494.000 ;
        RECT 3445.190 3435.000 3468.635 3435.115 ;
        RECT 3477.750 3435.000 3479.480 3435.145 ;
        RECT 3483.895 3435.000 3518.220 3435.115 ;
        RECT 3519.275 3435.000 3558.090 3435.115 ;
      LAYER met1 ;
        RECT 3367.730 3415.540 3368.050 3415.600 ;
        RECT 3368.650 3415.540 3368.970 3415.600 ;
        RECT 3376.930 3415.540 3377.250 3415.600 ;
        RECT 3367.730 3415.400 3377.250 3415.540 ;
        RECT 3367.730 3415.340 3368.050 3415.400 ;
        RECT 3368.650 3415.340 3368.970 3415.400 ;
        RECT 3376.930 3415.340 3377.250 3415.400 ;
        RECT 3367.730 3402.280 3368.050 3402.340 ;
        RECT 3369.570 3402.280 3369.890 3402.340 ;
        RECT 3376.930 3402.280 3377.250 3402.340 ;
        RECT 3367.730 3402.140 3377.250 3402.280 ;
        RECT 3367.730 3402.080 3368.050 3402.140 ;
        RECT 3369.570 3402.080 3369.890 3402.140 ;
        RECT 3376.930 3402.080 3377.250 3402.140 ;
        RECT 3376.010 3394.120 3376.330 3394.180 ;
        RECT 3376.930 3394.120 3377.250 3394.180 ;
        RECT 3376.010 3393.980 3377.250 3394.120 ;
        RECT 3376.010 3393.920 3376.330 3393.980 ;
        RECT 3376.930 3393.920 3377.250 3393.980 ;
        RECT 3368.190 3368.280 3368.510 3368.340 ;
        RECT 3370.030 3368.280 3370.350 3368.340 ;
        RECT 3376.930 3368.280 3377.250 3368.340 ;
        RECT 3368.190 3368.140 3377.250 3368.280 ;
        RECT 3368.190 3368.080 3368.510 3368.140 ;
        RECT 3370.030 3368.080 3370.350 3368.140 ;
        RECT 3376.930 3368.080 3377.250 3368.140 ;
      LAYER met1 ;
        RECT 19.025 3357.000 21.100 3357.020 ;
        RECT 29.910 3357.000 68.725 3357.145 ;
        RECT 69.780 3357.000 104.105 3357.145 ;
        POLYGON 127.070 3357.115 127.070 3357.060 127.015 3357.060 ;
        RECT 127.070 3357.060 148.780 3357.115 ;
        RECT 105.420 3357.000 148.780 3357.060 ;
        RECT 164.275 3357.000 169.880 3357.115 ;
        RECT 174.985 3357.000 180.515 3357.115 ;
        RECT 0.000 3277.000 206.845 3357.000 ;
        RECT 3381.155 3355.000 3588.000 3435.000 ;
        RECT 3407.485 3354.885 3413.015 3355.000 ;
        RECT 3418.120 3354.885 3423.725 3355.000 ;
        RECT 3439.220 3354.940 3482.580 3355.000 ;
        RECT 3439.220 3354.885 3460.930 3354.940 ;
        POLYGON 3460.930 3354.940 3460.985 3354.940 3460.930 3354.885 ;
        RECT 3483.895 3354.855 3518.220 3355.000 ;
        RECT 3519.275 3354.855 3558.090 3355.000 ;
        RECT 3566.900 3354.980 3568.975 3355.000 ;
      LAYER met1 ;
        RECT 208.910 3343.800 209.230 3343.860 ;
        RECT 213.050 3343.800 213.370 3343.860 ;
        RECT 208.910 3343.660 213.370 3343.800 ;
        RECT 208.910 3343.600 209.230 3343.660 ;
        RECT 213.050 3343.600 213.370 3343.660 ;
        RECT 208.910 3306.740 209.230 3306.800 ;
        RECT 212.590 3306.740 212.910 3306.800 ;
        RECT 208.910 3306.600 212.910 3306.740 ;
        RECT 208.910 3306.540 209.230 3306.600 ;
        RECT 212.590 3306.540 212.910 3306.600 ;
        RECT 208.910 3296.540 209.230 3296.600 ;
        RECT 212.130 3296.540 212.450 3296.600 ;
        RECT 213.510 3296.540 213.830 3296.600 ;
        RECT 208.910 3296.400 213.830 3296.540 ;
        RECT 208.910 3296.340 209.230 3296.400 ;
        RECT 212.130 3296.340 212.450 3296.400 ;
        RECT 213.510 3296.340 213.830 3296.400 ;
      LAYER met1 ;
        RECT 29.910 3276.885 68.725 3277.000 ;
        RECT 69.780 3276.885 104.105 3277.000 ;
        RECT 108.520 3276.855 110.250 3277.000 ;
        RECT 119.365 3276.885 142.810 3277.000 ;
        RECT 3445.190 3214.000 3468.635 3214.115 ;
        RECT 3477.750 3214.000 3479.480 3214.145 ;
        RECT 3483.895 3214.000 3518.220 3214.115 ;
        RECT 3519.275 3214.000 3558.090 3214.115 ;
      LAYER met1 ;
        RECT 3368.190 3194.540 3368.510 3194.600 ;
        RECT 3376.930 3194.540 3377.250 3194.600 ;
        RECT 3368.190 3194.400 3377.250 3194.540 ;
        RECT 3368.190 3194.340 3368.510 3194.400 ;
        RECT 3376.930 3194.340 3377.250 3194.400 ;
        RECT 3367.730 3181.620 3368.050 3181.680 ;
        RECT 3376.930 3181.620 3377.250 3181.680 ;
        RECT 3367.730 3181.480 3377.250 3181.620 ;
        RECT 3367.730 3181.420 3368.050 3181.480 ;
        RECT 3376.930 3181.420 3377.250 3181.480 ;
        RECT 3376.010 3173.120 3376.330 3173.180 ;
        RECT 3376.930 3173.120 3377.250 3173.180 ;
        RECT 3376.010 3172.980 3377.250 3173.120 ;
        RECT 3376.010 3172.920 3376.330 3172.980 ;
        RECT 3376.930 3172.920 3377.250 3172.980 ;
        RECT 3367.270 3147.280 3367.590 3147.340 ;
        RECT 3370.030 3147.280 3370.350 3147.340 ;
        RECT 3376.930 3147.280 3377.250 3147.340 ;
        RECT 3367.270 3147.140 3377.250 3147.280 ;
        RECT 3367.270 3147.080 3367.590 3147.140 ;
        RECT 3370.030 3147.080 3370.350 3147.140 ;
        RECT 3376.930 3147.080 3377.250 3147.140 ;
      LAYER met1 ;
        RECT 19.025 3141.000 21.100 3141.020 ;
        RECT 29.910 3141.000 68.725 3141.145 ;
        RECT 69.780 3141.000 104.105 3141.145 ;
        POLYGON 127.070 3141.115 127.070 3141.060 127.015 3141.060 ;
        RECT 127.070 3141.060 148.780 3141.115 ;
        RECT 105.420 3141.000 148.780 3141.060 ;
        RECT 164.275 3141.000 169.880 3141.115 ;
        RECT 174.985 3141.000 180.515 3141.115 ;
        RECT 0.000 3061.000 206.845 3141.000 ;
        RECT 3381.155 3134.000 3588.000 3214.000 ;
        RECT 3407.485 3133.885 3413.015 3134.000 ;
        RECT 3418.120 3133.885 3423.725 3134.000 ;
        RECT 3439.220 3133.940 3482.580 3134.000 ;
        RECT 3439.220 3133.885 3460.930 3133.940 ;
        POLYGON 3460.930 3133.940 3460.985 3133.940 3460.930 3133.885 ;
        RECT 3483.895 3133.855 3518.220 3134.000 ;
        RECT 3519.275 3133.855 3558.090 3134.000 ;
        RECT 3566.900 3133.980 3568.975 3134.000 ;
      LAYER met1 ;
        RECT 208.910 3127.560 209.230 3127.620 ;
        RECT 213.050 3127.560 213.370 3127.620 ;
        RECT 208.910 3127.420 213.370 3127.560 ;
        RECT 208.910 3127.360 209.230 3127.420 ;
        RECT 213.050 3127.360 213.370 3127.420 ;
        RECT 208.910 3090.840 209.230 3090.900 ;
        RECT 212.590 3090.840 212.910 3090.900 ;
        RECT 208.910 3090.700 212.910 3090.840 ;
        RECT 208.910 3090.640 209.230 3090.700 ;
        RECT 212.590 3090.640 212.910 3090.700 ;
        RECT 208.910 3075.200 209.230 3075.260 ;
        RECT 213.510 3075.200 213.830 3075.260 ;
        RECT 208.910 3075.060 213.830 3075.200 ;
        RECT 208.910 3075.000 209.230 3075.060 ;
        RECT 211.300 3073.560 211.440 3075.060 ;
        RECT 213.510 3075.000 213.830 3075.060 ;
        RECT 211.210 3073.300 211.530 3073.560 ;
      LAYER met1 ;
        RECT 29.910 3060.885 68.725 3061.000 ;
        RECT 69.780 3060.885 104.105 3061.000 ;
        RECT 108.520 3060.855 110.250 3061.000 ;
        RECT 119.365 3060.885 142.810 3061.000 ;
        RECT 3445.190 2992.000 3468.635 2992.115 ;
        RECT 3477.750 2992.000 3479.480 2992.145 ;
        RECT 3483.895 2992.000 3518.220 2992.115 ;
        RECT 3519.275 2992.000 3558.090 2992.115 ;
      LAYER met1 ;
        RECT 3368.190 2975.920 3368.510 2975.980 ;
        RECT 3376.930 2975.920 3377.250 2975.980 ;
        RECT 3368.190 2975.780 3377.250 2975.920 ;
        RECT 3368.190 2975.720 3368.510 2975.780 ;
        RECT 3376.930 2975.720 3377.250 2975.780 ;
        RECT 3367.730 2959.600 3368.050 2959.660 ;
        RECT 3376.930 2959.600 3377.250 2959.660 ;
        RECT 3367.730 2959.460 3377.250 2959.600 ;
        RECT 3367.730 2959.400 3368.050 2959.460 ;
        RECT 3376.930 2959.400 3377.250 2959.460 ;
      LAYER met1 ;
        RECT 19.025 2925.000 21.100 2925.020 ;
        RECT 29.910 2925.000 68.725 2925.145 ;
        RECT 69.780 2925.000 104.105 2925.145 ;
        POLYGON 127.070 2925.115 127.070 2925.060 127.015 2925.060 ;
        RECT 127.070 2925.060 148.780 2925.115 ;
        RECT 105.420 2925.000 148.780 2925.060 ;
        RECT 164.275 2925.000 169.880 2925.115 ;
        RECT 174.985 2925.000 180.515 2925.115 ;
        RECT 0.000 2845.000 206.845 2925.000 ;
      LAYER met1 ;
        RECT 3367.270 2920.840 3367.590 2920.900 ;
        RECT 3369.570 2920.840 3369.890 2920.900 ;
        RECT 3376.930 2920.840 3377.250 2920.900 ;
        RECT 3367.270 2920.700 3377.250 2920.840 ;
        RECT 3367.270 2920.640 3367.590 2920.700 ;
        RECT 3369.570 2920.640 3369.890 2920.700 ;
        RECT 3376.930 2920.640 3377.250 2920.700 ;
        RECT 208.910 2916.420 209.230 2916.480 ;
        RECT 213.050 2916.420 213.370 2916.480 ;
        RECT 208.910 2916.280 213.370 2916.420 ;
        RECT 208.910 2916.220 209.230 2916.280 ;
        RECT 213.050 2916.220 213.370 2916.280 ;
      LAYER met1 ;
        RECT 3381.155 2912.000 3588.000 2992.000 ;
        RECT 3407.485 2911.885 3413.015 2912.000 ;
        RECT 3418.120 2911.885 3423.725 2912.000 ;
        RECT 3439.220 2911.940 3482.580 2912.000 ;
        RECT 3439.220 2911.885 3460.930 2911.940 ;
        POLYGON 3460.930 2911.940 3460.985 2911.940 3460.930 2911.885 ;
        RECT 3483.895 2911.855 3518.220 2912.000 ;
        RECT 3519.275 2911.855 3558.090 2912.000 ;
        RECT 3566.900 2911.980 3568.975 2912.000 ;
      LAYER met1 ;
        RECT 208.910 2879.700 209.230 2879.760 ;
        RECT 212.590 2879.700 212.910 2879.760 ;
        RECT 208.910 2879.560 212.910 2879.700 ;
        RECT 208.910 2879.500 209.230 2879.560 ;
        RECT 212.590 2879.500 212.910 2879.560 ;
        RECT 208.910 2859.300 209.230 2859.360 ;
        RECT 212.130 2859.300 212.450 2859.360 ;
        RECT 208.910 2859.160 212.450 2859.300 ;
        RECT 208.910 2859.100 209.230 2859.160 ;
        RECT 212.130 2859.100 212.450 2859.160 ;
      LAYER met1 ;
        RECT 29.910 2844.885 68.725 2845.000 ;
        RECT 69.780 2844.885 104.105 2845.000 ;
        RECT 108.520 2844.855 110.250 2845.000 ;
        RECT 119.365 2844.885 142.810 2845.000 ;
        RECT 3445.190 2771.000 3468.635 2771.115 ;
        RECT 3477.750 2771.000 3479.480 2771.145 ;
        RECT 3483.895 2771.000 3518.220 2771.115 ;
        RECT 3519.275 2771.000 3558.090 2771.115 ;
      LAYER met1 ;
        RECT 3368.190 2756.960 3368.510 2757.020 ;
        RECT 3376.930 2756.960 3377.250 2757.020 ;
        RECT 3368.190 2756.820 3377.250 2756.960 ;
        RECT 3368.190 2756.760 3368.510 2756.820 ;
        RECT 3376.930 2756.760 3377.250 2756.820 ;
        RECT 3367.730 2741.320 3368.050 2741.380 ;
        RECT 3376.930 2741.320 3377.250 2741.380 ;
        RECT 3367.730 2741.180 3377.250 2741.320 ;
        RECT 3367.730 2741.120 3368.050 2741.180 ;
        RECT 3376.930 2741.120 3377.250 2741.180 ;
      LAYER met1 ;
        RECT 19.025 2709.000 21.100 2709.020 ;
        RECT 29.910 2709.000 68.725 2709.145 ;
        RECT 69.780 2709.000 104.105 2709.145 ;
        POLYGON 127.070 2709.115 127.070 2709.060 127.015 2709.060 ;
        RECT 127.070 2709.060 148.780 2709.115 ;
        RECT 105.420 2709.000 148.780 2709.060 ;
        RECT 164.275 2709.000 169.880 2709.115 ;
        RECT 174.985 2709.000 180.515 2709.115 ;
        RECT 0.000 2629.000 206.845 2709.000 ;
      LAYER met1 ;
        RECT 3369.570 2704.600 3369.890 2704.660 ;
        RECT 3376.930 2704.600 3377.250 2704.660 ;
        RECT 3369.570 2704.460 3377.250 2704.600 ;
        RECT 3369.570 2704.400 3369.890 2704.460 ;
        RECT 3376.930 2704.400 3377.250 2704.460 ;
        RECT 208.910 2700.520 209.230 2700.580 ;
        RECT 213.050 2700.520 213.370 2700.580 ;
        RECT 208.910 2700.380 213.370 2700.520 ;
        RECT 208.910 2700.320 209.230 2700.380 ;
        RECT 213.050 2700.320 213.370 2700.380 ;
      LAYER met1 ;
        RECT 3381.155 2691.000 3588.000 2771.000 ;
        RECT 3407.485 2690.885 3413.015 2691.000 ;
        RECT 3418.120 2690.885 3423.725 2691.000 ;
        RECT 3439.220 2690.940 3482.580 2691.000 ;
        RECT 3439.220 2690.885 3460.930 2690.940 ;
        POLYGON 3460.930 2690.940 3460.985 2690.940 3460.930 2690.885 ;
        RECT 3483.895 2690.855 3518.220 2691.000 ;
        RECT 3519.275 2690.855 3558.090 2691.000 ;
        RECT 3566.900 2690.980 3568.975 2691.000 ;
      LAYER met1 ;
        RECT 208.910 2659.040 209.230 2659.100 ;
        RECT 212.590 2659.040 212.910 2659.100 ;
        RECT 213.510 2659.040 213.830 2659.100 ;
        RECT 208.910 2658.900 213.830 2659.040 ;
        RECT 208.910 2658.840 209.230 2658.900 ;
        RECT 212.590 2658.840 212.910 2658.900 ;
        RECT 213.510 2658.840 213.830 2658.900 ;
        RECT 208.910 2643.400 209.230 2643.460 ;
        RECT 212.130 2643.400 212.450 2643.460 ;
        RECT 208.910 2643.260 212.450 2643.400 ;
        RECT 208.910 2643.200 209.230 2643.260 ;
        RECT 212.130 2643.200 212.450 2643.260 ;
      LAYER met1 ;
        RECT 29.910 2628.885 68.725 2629.000 ;
        RECT 69.780 2628.885 104.105 2629.000 ;
        RECT 108.520 2628.855 110.250 2629.000 ;
        RECT 119.365 2628.885 142.810 2629.000 ;
        RECT 3390.035 2546.375 3587.725 2549.815 ;
        RECT 3389.130 2541.145 3587.725 2546.375 ;
        RECT 3390.035 2537.965 3587.725 2541.145 ;
        RECT 3388.970 2536.650 3587.725 2537.965 ;
      LAYER met1 ;
        RECT 3376.470 2497.540 3376.790 2497.600 ;
        RECT 3380.610 2497.540 3380.930 2497.600 ;
        RECT 3376.470 2497.400 3380.930 2497.540 ;
        RECT 3376.470 2497.340 3376.790 2497.400 ;
        RECT 3380.610 2497.340 3380.930 2497.400 ;
      LAYER met1 ;
        RECT 0.275 2487.680 197.965 2489.915 ;
        RECT 0.275 2486.540 199.030 2487.680 ;
        RECT 0.275 2430.350 197.965 2486.540 ;
        POLYGON 197.965 2486.540 198.080 2486.540 198.080 2486.425 ;
        POLYGON 198.080 2430.465 198.080 2430.350 197.965 2430.350 ;
        RECT 198.080 2430.350 199.030 2486.540 ;
        RECT 3388.970 2480.460 3389.920 2536.650 ;
        POLYGON 3389.920 2536.650 3390.035 2536.650 3389.920 2536.535 ;
        POLYGON 3389.920 2480.575 3390.035 2480.460 3389.920 2480.460 ;
        RECT 3390.035 2480.460 3587.725 2536.650 ;
        RECT 3388.970 2479.320 3587.725 2480.460 ;
        RECT 3390.035 2477.085 3587.725 2479.320 ;
      LAYER met1 ;
        RECT 3380.610 2474.420 3380.930 2474.480 ;
        RECT 3389.810 2474.420 3390.130 2474.480 ;
        RECT 3380.610 2474.280 3390.130 2474.420 ;
        RECT 3380.610 2474.220 3380.930 2474.280 ;
        RECT 3389.810 2474.220 3390.130 2474.280 ;
      LAYER met1 ;
        RECT 0.275 2429.035 199.030 2430.350 ;
        RECT 0.275 2425.855 197.965 2429.035 ;
        RECT 0.275 2420.625 198.870 2425.855 ;
        RECT 0.275 2417.185 197.965 2420.625 ;
        RECT 3390.035 2316.345 3587.840 2332.880 ;
        RECT 3390.000 2312.075 3587.840 2316.345 ;
        RECT 122.615 2287.935 204.885 2291.935 ;
        POLYGON 204.885 2291.935 208.885 2287.935 204.885 2287.935 ;
        RECT 122.615 2282.200 208.885 2287.935 ;
        RECT 0.160 2262.565 197.965 2281.000 ;
        RECT 198.780 2262.565 208.885 2282.200 ;
        RECT 0.160 2226.925 208.885 2262.565 ;
        RECT 3379.115 2276.435 3587.840 2312.075 ;
        RECT 3379.115 2256.800 3389.220 2276.435 ;
        RECT 3390.035 2258.000 3587.840 2276.435 ;
        RECT 3379.115 2251.065 3465.385 2256.800 ;
        POLYGON 3379.115 2251.065 3383.115 2251.065 3383.115 2247.065 ;
        RECT 3383.115 2247.065 3465.385 2251.065 ;
        RECT 0.160 2222.655 198.000 2226.925 ;
        RECT 0.160 2206.120 197.965 2222.655 ;
      LAYER met1 ;
        RECT 3370.030 2111.300 3370.350 2111.360 ;
        RECT 3373.710 2111.300 3374.030 2111.360 ;
        RECT 3370.030 2111.160 3374.030 2111.300 ;
        RECT 3370.030 2111.100 3370.350 2111.160 ;
        RECT 3373.710 2111.100 3374.030 2111.160 ;
      LAYER met1 ;
        RECT 3390.035 2104.965 3587.725 2116.815 ;
        RECT 3388.970 2103.650 3587.725 2104.965 ;
      LAYER met1 ;
        RECT 3370.030 2096.000 3370.350 2096.060 ;
        RECT 3387.510 2096.000 3387.830 2096.060 ;
        RECT 3370.030 2095.860 3387.830 2096.000 ;
        RECT 3370.030 2095.800 3370.350 2095.860 ;
        RECT 3387.510 2095.800 3387.830 2095.860 ;
      LAYER met1 ;
        RECT 19.025 2070.000 21.100 2070.020 ;
        RECT 29.910 2070.000 68.725 2070.145 ;
        RECT 69.780 2070.000 104.105 2070.145 ;
        POLYGON 127.070 2070.115 127.070 2070.060 127.015 2070.060 ;
        RECT 127.070 2070.060 148.780 2070.115 ;
        RECT 105.420 2070.000 148.780 2070.060 ;
        RECT 164.275 2070.000 169.880 2070.115 ;
        RECT 174.985 2070.000 180.515 2070.115 ;
        RECT 0.000 1990.000 206.845 2070.000 ;
      LAYER met1 ;
        RECT 208.910 2056.560 209.230 2056.620 ;
        RECT 212.590 2056.560 212.910 2056.620 ;
        RECT 208.910 2056.420 212.910 2056.560 ;
        RECT 208.910 2056.360 209.230 2056.420 ;
        RECT 212.590 2056.360 212.910 2056.420 ;
      LAYER met1 ;
        RECT 3388.970 2047.460 3389.920 2103.650 ;
        POLYGON 3389.920 2103.650 3390.035 2103.650 3389.920 2103.535 ;
        POLYGON 3389.920 2047.575 3390.035 2047.460 3389.920 2047.460 ;
        RECT 3390.035 2047.460 3587.725 2103.650 ;
        RECT 3388.970 2046.320 3587.725 2047.460 ;
        RECT 3390.035 2043.380 3587.725 2046.320 ;
      LAYER met1 ;
        RECT 208.910 2024.600 209.230 2024.660 ;
        RECT 213.510 2024.600 213.830 2024.660 ;
        RECT 208.910 2024.460 213.830 2024.600 ;
        RECT 208.910 2024.400 209.230 2024.460 ;
        RECT 213.510 2024.400 213.830 2024.460 ;
        RECT 208.910 2009.640 209.230 2009.700 ;
        RECT 212.130 2009.640 212.450 2009.700 ;
        RECT 208.910 2009.500 212.450 2009.640 ;
        RECT 208.910 2009.440 209.230 2009.500 ;
        RECT 212.130 2009.440 212.450 2009.500 ;
      LAYER met1 ;
        RECT 29.910 1989.885 68.725 1990.000 ;
        RECT 69.780 1989.885 104.105 1990.000 ;
        RECT 108.520 1989.855 110.250 1990.000 ;
        RECT 119.365 1989.885 142.810 1990.000 ;
        RECT 3445.190 1900.000 3468.635 1900.115 ;
        RECT 3477.750 1900.000 3479.480 1900.145 ;
        RECT 3483.895 1900.000 3518.220 1900.115 ;
        RECT 3519.275 1900.000 3558.090 1900.115 ;
      LAYER met1 ;
        RECT 3369.570 1880.780 3369.890 1880.840 ;
        RECT 3376.930 1880.780 3377.250 1880.840 ;
        RECT 3369.570 1880.640 3377.250 1880.780 ;
        RECT 3369.570 1880.580 3369.890 1880.640 ;
        RECT 3376.930 1880.580 3377.250 1880.640 ;
        RECT 3368.650 1865.480 3368.970 1865.540 ;
        RECT 3376.930 1865.480 3377.250 1865.540 ;
        RECT 3368.650 1865.340 3377.250 1865.480 ;
        RECT 3368.650 1865.280 3368.970 1865.340 ;
        RECT 3376.930 1865.280 3377.250 1865.340 ;
      LAYER met1 ;
        RECT 19.025 1854.000 21.100 1854.020 ;
        RECT 29.910 1854.000 68.725 1854.145 ;
        RECT 69.780 1854.000 104.105 1854.145 ;
        POLYGON 127.070 1854.115 127.070 1854.060 127.015 1854.060 ;
        RECT 127.070 1854.060 148.780 1854.115 ;
        RECT 105.420 1854.000 148.780 1854.060 ;
        RECT 164.275 1854.000 169.880 1854.115 ;
        RECT 174.985 1854.000 180.515 1854.115 ;
        RECT 0.000 1774.000 206.845 1854.000 ;
      LAYER met1 ;
        RECT 208.910 1845.420 209.230 1845.480 ;
        RECT 212.590 1845.420 212.910 1845.480 ;
        RECT 208.910 1845.280 212.910 1845.420 ;
        RECT 208.910 1845.220 209.230 1845.280 ;
        RECT 212.590 1845.220 212.910 1845.280 ;
        RECT 3370.030 1828.760 3370.350 1828.820 ;
        RECT 3376.930 1828.760 3377.250 1828.820 ;
        RECT 3370.030 1828.620 3377.250 1828.760 ;
        RECT 3370.030 1828.560 3370.350 1828.620 ;
        RECT 3376.930 1828.560 3377.250 1828.620 ;
      LAYER met1 ;
        RECT 3381.155 1820.000 3588.000 1900.000 ;
        RECT 3407.485 1819.885 3413.015 1820.000 ;
        RECT 3418.120 1819.885 3423.725 1820.000 ;
        RECT 3439.220 1819.940 3482.580 1820.000 ;
        RECT 3439.220 1819.885 3460.930 1819.940 ;
        POLYGON 3460.930 1819.940 3460.985 1819.940 3460.930 1819.885 ;
        RECT 3483.895 1819.855 3518.220 1820.000 ;
        RECT 3519.275 1819.855 3558.090 1820.000 ;
        RECT 3566.900 1819.980 3568.975 1820.000 ;
      LAYER met1 ;
        RECT 208.910 1806.660 209.230 1806.720 ;
        RECT 213.050 1806.660 213.370 1806.720 ;
        RECT 208.910 1806.520 213.370 1806.660 ;
        RECT 208.910 1806.460 209.230 1806.520 ;
        RECT 213.050 1806.460 213.370 1806.520 ;
        RECT 208.910 1788.300 209.230 1788.360 ;
        RECT 212.130 1788.300 212.450 1788.360 ;
        RECT 213.510 1788.300 213.830 1788.360 ;
        RECT 208.910 1788.160 213.830 1788.300 ;
        RECT 208.910 1788.100 209.230 1788.160 ;
        RECT 212.130 1788.100 212.450 1788.160 ;
        RECT 213.510 1788.100 213.830 1788.160 ;
      LAYER met1 ;
        RECT 29.910 1773.885 68.725 1774.000 ;
        RECT 69.780 1773.885 104.105 1774.000 ;
        RECT 108.520 1773.855 110.250 1774.000 ;
        RECT 119.365 1773.885 142.810 1774.000 ;
        RECT 3445.190 1679.000 3468.635 1679.115 ;
        RECT 3477.750 1679.000 3479.480 1679.145 ;
        RECT 3483.895 1679.000 3518.220 1679.115 ;
        RECT 3519.275 1679.000 3558.090 1679.115 ;
      LAYER met1 ;
        RECT 3368.650 1669.980 3368.970 1670.040 ;
        RECT 3376.010 1669.980 3376.330 1670.040 ;
        RECT 3368.650 1669.840 3376.330 1669.980 ;
        RECT 3368.650 1669.780 3368.970 1669.840 ;
        RECT 3376.010 1669.780 3376.330 1669.840 ;
        RECT 3367.270 1659.780 3367.590 1659.840 ;
        RECT 3369.570 1659.780 3369.890 1659.840 ;
        RECT 3376.930 1659.780 3377.250 1659.840 ;
        RECT 3367.270 1659.640 3377.250 1659.780 ;
        RECT 3367.270 1659.580 3367.590 1659.640 ;
        RECT 3369.570 1659.580 3369.890 1659.640 ;
        RECT 3376.930 1659.580 3377.250 1659.640 ;
        RECT 3367.730 1644.480 3368.050 1644.540 ;
        RECT 3376.010 1644.480 3376.330 1644.540 ;
        RECT 3376.930 1644.480 3377.250 1644.540 ;
        RECT 3367.730 1644.340 3377.250 1644.480 ;
        RECT 3367.730 1644.280 3368.050 1644.340 ;
        RECT 3376.010 1644.280 3376.330 1644.340 ;
        RECT 3376.930 1644.280 3377.250 1644.340 ;
      LAYER met1 ;
        RECT 19.025 1637.000 21.100 1637.020 ;
        RECT 29.910 1637.000 68.725 1637.145 ;
        RECT 69.780 1637.000 104.105 1637.145 ;
        POLYGON 127.070 1637.115 127.070 1637.060 127.015 1637.060 ;
        RECT 127.070 1637.060 148.780 1637.115 ;
        RECT 105.420 1637.000 148.780 1637.060 ;
        RECT 164.275 1637.000 169.880 1637.115 ;
        RECT 174.985 1637.000 180.515 1637.115 ;
        RECT 0.000 1557.000 206.845 1637.000 ;
      LAYER met1 ;
        RECT 208.910 1628.500 209.230 1628.560 ;
        RECT 212.590 1628.500 212.910 1628.560 ;
        RECT 208.910 1628.360 212.910 1628.500 ;
        RECT 208.910 1628.300 209.230 1628.360 ;
        RECT 212.590 1628.300 212.910 1628.360 ;
        RECT 3368.190 1612.520 3368.510 1612.580 ;
        RECT 3370.030 1612.520 3370.350 1612.580 ;
        RECT 3376.930 1612.520 3377.250 1612.580 ;
        RECT 3368.190 1612.380 3377.250 1612.520 ;
        RECT 3368.190 1612.320 3368.510 1612.380 ;
        RECT 3370.030 1612.320 3370.350 1612.380 ;
        RECT 3376.930 1612.320 3377.250 1612.380 ;
      LAYER met1 ;
        RECT 3381.155 1599.000 3588.000 1679.000 ;
        RECT 3407.485 1598.885 3413.015 1599.000 ;
        RECT 3418.120 1598.885 3423.725 1599.000 ;
        RECT 3439.220 1598.940 3482.580 1599.000 ;
        RECT 3439.220 1598.885 3460.930 1598.940 ;
        POLYGON 3460.930 1598.940 3460.985 1598.940 3460.930 1598.885 ;
        RECT 3483.895 1598.855 3518.220 1599.000 ;
        RECT 3519.275 1598.855 3558.090 1599.000 ;
        RECT 3566.900 1598.980 3568.975 1599.000 ;
      LAYER met1 ;
        RECT 208.910 1587.020 209.230 1587.080 ;
        RECT 213.050 1587.020 213.370 1587.080 ;
        RECT 208.910 1586.880 213.370 1587.020 ;
        RECT 208.910 1586.820 209.230 1586.880 ;
        RECT 213.050 1586.820 213.370 1586.880 ;
        RECT 208.910 1571.380 209.230 1571.440 ;
        RECT 212.590 1571.380 212.910 1571.440 ;
        RECT 213.510 1571.380 213.830 1571.440 ;
        RECT 208.910 1571.240 213.830 1571.380 ;
        RECT 208.910 1571.180 209.230 1571.240 ;
        RECT 212.590 1571.180 212.910 1571.240 ;
        RECT 213.510 1571.180 213.830 1571.240 ;
      LAYER met1 ;
        RECT 29.910 1556.885 68.725 1557.000 ;
        RECT 69.780 1556.885 104.105 1557.000 ;
        RECT 108.520 1556.855 110.250 1557.000 ;
        RECT 119.365 1556.885 142.810 1557.000 ;
        RECT 3445.190 1458.000 3468.635 1458.115 ;
        RECT 3477.750 1458.000 3479.480 1458.145 ;
        RECT 3483.895 1458.000 3518.220 1458.115 ;
        RECT 3519.275 1458.000 3558.090 1458.115 ;
      LAYER met1 ;
        RECT 3367.270 1443.880 3367.590 1443.940 ;
        RECT 3376.930 1443.880 3377.250 1443.940 ;
        RECT 3367.270 1443.740 3377.250 1443.880 ;
        RECT 3367.270 1443.680 3367.590 1443.740 ;
        RECT 3376.930 1443.680 3377.250 1443.740 ;
        RECT 3367.730 1426.540 3368.050 1426.600 ;
        RECT 3376.930 1426.540 3377.250 1426.600 ;
        RECT 3367.730 1426.400 3377.250 1426.540 ;
        RECT 3367.730 1426.340 3368.050 1426.400 ;
        RECT 3376.930 1426.340 3377.250 1426.400 ;
      LAYER met1 ;
        RECT 19.025 1421.000 21.100 1421.020 ;
        RECT 29.910 1421.000 68.725 1421.145 ;
        RECT 69.780 1421.000 104.105 1421.145 ;
        POLYGON 127.070 1421.115 127.070 1421.060 127.015 1421.060 ;
        RECT 127.070 1421.060 148.780 1421.115 ;
        RECT 105.420 1421.000 148.780 1421.060 ;
        RECT 164.275 1421.000 169.880 1421.115 ;
        RECT 174.985 1421.000 180.515 1421.115 ;
        RECT 0.000 1341.000 206.845 1421.000 ;
      LAYER met1 ;
        RECT 208.910 1407.840 209.230 1407.900 ;
        RECT 212.130 1407.840 212.450 1407.900 ;
        RECT 213.510 1407.840 213.830 1407.900 ;
        RECT 208.910 1407.700 213.830 1407.840 ;
        RECT 208.910 1407.640 209.230 1407.700 ;
        RECT 212.130 1407.640 212.450 1407.700 ;
        RECT 213.510 1407.640 213.830 1407.700 ;
        RECT 3368.190 1386.760 3368.510 1386.820 ;
        RECT 3376.930 1386.760 3377.250 1386.820 ;
        RECT 3368.190 1386.620 3377.250 1386.760 ;
        RECT 3368.190 1386.560 3368.510 1386.620 ;
        RECT 3376.930 1386.560 3377.250 1386.620 ;
      LAYER met1 ;
        RECT 3381.155 1378.000 3588.000 1458.000 ;
        RECT 3407.485 1377.885 3413.015 1378.000 ;
        RECT 3418.120 1377.885 3423.725 1378.000 ;
        RECT 3439.220 1377.940 3482.580 1378.000 ;
        RECT 3439.220 1377.885 3460.930 1377.940 ;
        POLYGON 3460.930 1377.940 3460.985 1377.940 3460.930 1377.885 ;
        RECT 3483.895 1377.855 3518.220 1378.000 ;
        RECT 3519.275 1377.855 3558.090 1378.000 ;
        RECT 3566.900 1377.980 3568.975 1378.000 ;
      LAYER met1 ;
        RECT 208.910 1373.500 209.230 1373.560 ;
        RECT 213.050 1373.500 213.370 1373.560 ;
        RECT 208.910 1373.360 213.370 1373.500 ;
        RECT 208.910 1373.300 209.230 1373.360 ;
        RECT 213.050 1373.300 213.370 1373.360 ;
        RECT 208.910 1360.580 209.230 1360.640 ;
        RECT 212.590 1360.580 212.910 1360.640 ;
        RECT 208.910 1360.440 212.910 1360.580 ;
        RECT 208.910 1360.380 209.230 1360.440 ;
        RECT 212.590 1360.380 212.910 1360.440 ;
      LAYER met1 ;
        RECT 29.910 1340.885 68.725 1341.000 ;
        RECT 69.780 1340.885 104.105 1341.000 ;
        RECT 108.520 1340.855 110.250 1341.000 ;
        RECT 119.365 1340.885 142.810 1341.000 ;
        RECT 3445.190 1236.000 3468.635 1236.115 ;
        RECT 3477.750 1236.000 3479.480 1236.145 ;
        RECT 3483.895 1236.000 3518.220 1236.115 ;
        RECT 3519.275 1236.000 3558.090 1236.115 ;
      LAYER met1 ;
        RECT 3367.270 1218.800 3367.590 1218.860 ;
        RECT 3376.930 1218.800 3377.250 1218.860 ;
        RECT 3367.270 1218.660 3377.250 1218.800 ;
        RECT 3367.270 1218.600 3367.590 1218.660 ;
        RECT 3376.930 1218.600 3377.250 1218.660 ;
      LAYER met1 ;
        RECT 19.025 1205.000 21.100 1205.020 ;
        RECT 29.910 1205.000 68.725 1205.145 ;
        RECT 69.780 1205.000 104.105 1205.145 ;
        POLYGON 127.070 1205.115 127.070 1205.060 127.015 1205.060 ;
        RECT 127.070 1205.060 148.780 1205.115 ;
        RECT 105.420 1205.000 148.780 1205.060 ;
        RECT 164.275 1205.000 169.880 1205.115 ;
        RECT 174.985 1205.000 180.515 1205.115 ;
        RECT 0.000 1125.000 206.845 1205.000 ;
      LAYER met1 ;
        RECT 3367.730 1201.460 3368.050 1201.520 ;
        RECT 3376.930 1201.460 3377.250 1201.520 ;
        RECT 3367.730 1201.320 3377.250 1201.460 ;
        RECT 3367.730 1201.260 3368.050 1201.320 ;
        RECT 3376.930 1201.260 3377.250 1201.320 ;
        RECT 208.910 1191.600 209.230 1191.660 ;
        RECT 212.130 1191.600 212.450 1191.660 ;
        RECT 213.510 1191.600 213.830 1191.660 ;
        RECT 208.910 1191.460 213.830 1191.600 ;
        RECT 208.910 1191.400 209.230 1191.460 ;
        RECT 212.130 1191.400 212.450 1191.460 ;
        RECT 213.510 1191.400 213.830 1191.460 ;
        RECT 3368.190 1169.500 3368.510 1169.560 ;
        RECT 3376.930 1169.500 3377.250 1169.560 ;
        RECT 3368.190 1169.360 3377.250 1169.500 ;
        RECT 3368.190 1169.300 3368.510 1169.360 ;
        RECT 3376.930 1169.300 3377.250 1169.360 ;
        RECT 208.910 1159.640 209.230 1159.700 ;
        RECT 213.050 1159.640 213.370 1159.700 ;
        RECT 208.910 1159.500 213.370 1159.640 ;
        RECT 208.910 1159.440 209.230 1159.500 ;
        RECT 213.050 1159.440 213.370 1159.500 ;
      LAYER met1 ;
        RECT 3381.155 1156.000 3588.000 1236.000 ;
        RECT 3407.485 1155.885 3413.015 1156.000 ;
        RECT 3418.120 1155.885 3423.725 1156.000 ;
        RECT 3439.220 1155.940 3482.580 1156.000 ;
        RECT 3439.220 1155.885 3460.930 1155.940 ;
        POLYGON 3460.930 1155.940 3460.985 1155.940 3460.930 1155.885 ;
        RECT 3483.895 1155.855 3518.220 1156.000 ;
        RECT 3519.275 1155.855 3558.090 1156.000 ;
        RECT 3566.900 1155.980 3568.975 1156.000 ;
      LAYER met1 ;
        RECT 208.910 1144.340 209.230 1144.400 ;
        RECT 212.590 1144.340 212.910 1144.400 ;
        RECT 208.910 1144.200 212.910 1144.340 ;
        RECT 208.910 1144.140 209.230 1144.200 ;
        RECT 212.590 1144.140 212.910 1144.200 ;
      LAYER met1 ;
        RECT 29.910 1124.885 68.725 1125.000 ;
        RECT 69.780 1124.885 104.105 1125.000 ;
        RECT 108.520 1124.855 110.250 1125.000 ;
        RECT 119.365 1124.885 142.810 1125.000 ;
        RECT 3445.190 1015.000 3468.635 1015.115 ;
        RECT 3477.750 1015.000 3479.480 1015.145 ;
        RECT 3483.895 1015.000 3518.220 1015.115 ;
        RECT 3519.275 1015.000 3558.090 1015.115 ;
      LAYER met1 ;
        RECT 3367.270 995.760 3367.590 995.820 ;
        RECT 3376.930 995.760 3377.250 995.820 ;
        RECT 3367.270 995.620 3377.250 995.760 ;
        RECT 3367.270 995.560 3367.590 995.620 ;
        RECT 3376.930 995.560 3377.250 995.620 ;
      LAYER met1 ;
        RECT 19.025 989.000 21.100 989.020 ;
        RECT 29.910 989.000 68.725 989.145 ;
        RECT 69.780 989.000 104.105 989.145 ;
        POLYGON 127.070 989.115 127.070 989.060 127.015 989.060 ;
        RECT 127.070 989.060 148.780 989.115 ;
        RECT 105.420 989.000 148.780 989.060 ;
        RECT 164.275 989.000 169.880 989.115 ;
        RECT 174.985 989.000 180.515 989.115 ;
        RECT 0.000 909.000 206.845 989.000 ;
      LAYER met1 ;
        RECT 3367.730 985.220 3368.050 985.280 ;
        RECT 3376.930 985.220 3377.250 985.280 ;
        RECT 3367.730 985.080 3377.250 985.220 ;
        RECT 3367.730 985.020 3368.050 985.080 ;
        RECT 3376.930 985.020 3377.250 985.080 ;
        RECT 208.910 975.700 209.230 975.760 ;
        RECT 212.130 975.700 212.450 975.760 ;
        RECT 208.910 975.560 212.450 975.700 ;
        RECT 208.910 975.500 209.230 975.560 ;
        RECT 212.130 975.500 212.450 975.560 ;
        RECT 3368.190 946.460 3368.510 946.520 ;
        RECT 3376.930 946.460 3377.250 946.520 ;
        RECT 3368.190 946.320 3377.250 946.460 ;
        RECT 3368.190 946.260 3368.510 946.320 ;
        RECT 3376.930 946.260 3377.250 946.320 ;
        RECT 208.910 943.740 209.230 943.800 ;
        RECT 212.590 943.740 212.910 943.800 ;
        RECT 213.970 943.740 214.290 943.800 ;
        RECT 208.910 943.600 214.290 943.740 ;
        RECT 208.910 943.540 209.230 943.600 ;
        RECT 212.590 943.540 212.910 943.600 ;
        RECT 213.970 943.540 214.290 943.600 ;
      LAYER met1 ;
        RECT 3381.155 935.000 3588.000 1015.000 ;
        RECT 3407.485 934.885 3413.015 935.000 ;
        RECT 3418.120 934.885 3423.725 935.000 ;
        RECT 3439.220 934.940 3482.580 935.000 ;
        RECT 3439.220 934.885 3460.930 934.940 ;
        POLYGON 3460.930 934.940 3460.985 934.940 3460.930 934.885 ;
        RECT 3483.895 934.855 3518.220 935.000 ;
        RECT 3519.275 934.855 3558.090 935.000 ;
        RECT 3566.900 934.980 3568.975 935.000 ;
      LAYER met1 ;
        RECT 208.910 928.440 209.230 928.500 ;
        RECT 213.510 928.440 213.830 928.500 ;
        RECT 208.910 928.300 213.830 928.440 ;
        RECT 208.910 928.240 209.230 928.300 ;
        RECT 213.510 928.240 213.830 928.300 ;
        RECT 211.210 921.980 211.530 922.040 ;
        RECT 213.510 921.980 213.830 922.040 ;
        RECT 211.210 921.840 213.830 921.980 ;
        RECT 211.210 921.780 211.530 921.840 ;
        RECT 213.510 921.780 213.830 921.840 ;
      LAYER met1 ;
        RECT 29.910 908.885 68.725 909.000 ;
        RECT 69.780 908.885 104.105 909.000 ;
        RECT 108.520 908.855 110.250 909.000 ;
        RECT 119.365 908.885 142.810 909.000 ;
        RECT 3445.190 794.000 3468.635 794.115 ;
        RECT 3477.750 794.000 3479.480 794.145 ;
        RECT 3483.895 794.000 3518.220 794.115 ;
        RECT 3519.275 794.000 3558.090 794.115 ;
      LAYER met1 ;
        RECT 3367.270 779.860 3367.590 779.920 ;
        RECT 3369.570 779.860 3369.890 779.920 ;
        RECT 3376.930 779.860 3377.250 779.920 ;
        RECT 3367.270 779.720 3377.250 779.860 ;
        RECT 3367.270 779.660 3367.590 779.720 ;
        RECT 3369.570 779.660 3369.890 779.720 ;
        RECT 3376.930 779.660 3377.250 779.720 ;
        RECT 3367.730 764.220 3368.050 764.280 ;
        RECT 3376.930 764.220 3377.250 764.280 ;
        RECT 3367.730 764.080 3377.250 764.220 ;
        RECT 3367.730 764.020 3368.050 764.080 ;
        RECT 3376.930 764.020 3377.250 764.080 ;
        RECT 3368.650 722.740 3368.970 722.800 ;
        RECT 3376.930 722.740 3377.250 722.800 ;
        RECT 3368.650 722.600 3377.250 722.740 ;
        RECT 3368.650 722.540 3368.970 722.600 ;
        RECT 3376.930 722.540 3377.250 722.600 ;
      LAYER met1 ;
        RECT 3381.155 714.000 3588.000 794.000 ;
        RECT 3407.485 713.885 3413.015 714.000 ;
        RECT 3418.120 713.885 3423.725 714.000 ;
        RECT 3439.220 713.940 3482.580 714.000 ;
        RECT 3439.220 713.885 3460.930 713.940 ;
        POLYGON 3460.930 713.940 3460.985 713.940 3460.930 713.885 ;
        RECT 3483.895 713.855 3518.220 714.000 ;
        RECT 3519.275 713.855 3558.090 714.000 ;
        RECT 3566.900 713.980 3568.975 714.000 ;
        RECT 0.275 621.680 197.965 623.915 ;
        RECT 0.275 620.540 199.030 621.680 ;
        RECT 0.275 564.350 197.965 620.540 ;
        POLYGON 197.965 620.540 198.080 620.540 198.080 620.425 ;
        POLYGON 198.080 564.465 198.080 564.350 197.965 564.350 ;
        RECT 198.080 564.350 199.030 620.540 ;
      LAYER met1 ;
        RECT 212.590 607.480 212.910 607.540 ;
        RECT 220.870 607.480 221.190 607.540 ;
        RECT 212.590 607.340 221.190 607.480 ;
        RECT 212.590 607.280 212.910 607.340 ;
        RECT 220.870 607.280 221.190 607.340 ;
      LAYER met1 ;
        RECT 3445.190 572.000 3468.635 572.115 ;
        RECT 3477.750 572.000 3479.480 572.145 ;
        RECT 3483.895 572.000 3518.220 572.115 ;
        RECT 3519.275 572.000 3558.090 572.115 ;
        RECT 0.275 563.035 199.030 564.350 ;
        RECT 0.275 559.855 197.965 563.035 ;
        RECT 0.275 554.625 198.870 559.855 ;
      LAYER met1 ;
        RECT 3367.270 557.840 3367.590 557.900 ;
        RECT 3369.570 557.840 3369.890 557.900 ;
        RECT 3376.930 557.840 3377.250 557.900 ;
        RECT 3367.270 557.700 3377.250 557.840 ;
        RECT 3367.270 557.640 3367.590 557.700 ;
        RECT 3369.570 557.640 3369.890 557.700 ;
        RECT 3376.930 557.640 3377.250 557.700 ;
      LAYER met1 ;
        RECT 0.275 551.185 197.965 554.625 ;
      LAYER met1 ;
        RECT 3367.730 542.200 3368.050 542.260 ;
        RECT 3376.930 542.200 3377.250 542.260 ;
        RECT 3367.730 542.060 3377.250 542.200 ;
        RECT 3367.730 542.000 3368.050 542.060 ;
        RECT 3376.930 542.000 3377.250 542.060 ;
        RECT 212.130 530.300 212.450 530.360 ;
        RECT 220.870 530.300 221.190 530.360 ;
        RECT 212.130 530.160 221.190 530.300 ;
        RECT 212.130 530.100 212.450 530.160 ;
        RECT 220.870 530.100 221.190 530.160 ;
      LAYER met1 ;
        RECT 3381.155 492.000 3588.000 572.000 ;
        RECT 3407.485 491.885 3413.015 492.000 ;
        RECT 3418.120 491.885 3423.725 492.000 ;
        RECT 3439.220 491.940 3482.580 492.000 ;
        RECT 3439.220 491.885 3460.930 491.940 ;
        POLYGON 3460.930 491.940 3460.985 491.940 3460.930 491.885 ;
        RECT 3483.895 491.855 3518.220 492.000 ;
        RECT 3519.275 491.855 3558.090 492.000 ;
        RECT 3566.900 491.980 3568.975 492.000 ;
        RECT 159.640 425.935 163.510 426.195 ;
        RECT 159.640 421.935 204.500 425.935 ;
        POLYGON 204.500 425.935 208.500 421.935 204.500 421.935 ;
        RECT 159.640 416.200 208.500 421.935 ;
        RECT 159.640 415.245 163.510 416.200 ;
        RECT 0.160 396.565 197.965 415.000 ;
        RECT 198.780 396.565 208.500 416.200 ;
        RECT 0.160 360.495 208.500 396.565 ;
        RECT 0.160 356.655 198.000 360.495 ;
        RECT 198.980 358.655 208.500 360.495 ;
        POLYGON 198.980 358.655 200.980 358.655 200.980 356.655 ;
        RECT 200.980 356.655 206.500 358.655 ;
        POLYGON 206.500 358.655 208.500 358.655 206.500 356.655 ;
        RECT 0.160 340.120 197.965 356.655 ;
      LAYER met1 ;
        RECT 224.090 234.640 224.410 234.900 ;
        RECT 1004.340 234.700 1488.860 234.840 ;
        RECT 224.180 234.500 224.320 234.640 ;
        RECT 1004.340 234.560 1004.480 234.700 ;
        RECT 717.670 234.500 717.990 234.560 ;
        RECT 224.180 234.360 717.990 234.500 ;
        RECT 717.670 234.300 717.990 234.360 ;
        RECT 1004.250 234.300 1004.570 234.560 ;
        RECT 1204.440 234.500 1204.580 234.700 ;
        RECT 1488.720 234.560 1488.860 234.700 ;
        RECT 1547.140 234.700 1763.020 234.840 ;
        RECT 1547.140 234.560 1547.280 234.700 ;
        RECT 1762.880 234.560 1763.020 234.700 ;
        RECT 1821.300 234.700 2037.180 234.840 ;
        RECT 1821.300 234.560 1821.440 234.700 ;
        RECT 2037.040 234.560 2037.180 234.700 ;
        RECT 2095.460 234.700 2310.880 234.840 ;
        RECT 2095.460 234.560 2095.600 234.700 ;
        RECT 2310.740 234.560 2310.880 234.700 ;
        RECT 2369.160 234.700 2585.040 234.840 ;
        RECT 2369.160 234.560 2369.300 234.700 ;
        RECT 2584.900 234.560 2585.040 234.700 ;
        RECT 1281.170 234.500 1281.490 234.560 ;
        RECT 1204.440 234.360 1281.490 234.500 ;
        RECT 1281.170 234.300 1281.490 234.360 ;
        RECT 1488.630 234.300 1488.950 234.560 ;
        RECT 1547.050 234.300 1547.370 234.560 ;
        RECT 1762.790 234.300 1763.110 234.560 ;
        RECT 1821.210 234.300 1821.530 234.560 ;
        RECT 2036.950 234.300 2037.270 234.560 ;
        RECT 2095.370 234.300 2095.690 234.560 ;
        RECT 2310.650 234.300 2310.970 234.560 ;
        RECT 2369.070 234.300 2369.390 234.560 ;
        RECT 2584.810 234.300 2585.130 234.560 ;
        RECT 211.210 228.380 211.530 228.440 ;
        RECT 704.790 228.380 705.110 228.440 ;
        RECT 211.210 228.240 705.110 228.380 ;
        RECT 211.210 228.180 211.530 228.240 ;
        RECT 704.790 228.180 705.110 228.240 ;
        RECT 933.410 228.040 933.730 228.100 ;
        RECT 973.430 228.040 973.750 228.100 ;
        RECT 933.410 227.900 973.750 228.040 ;
        RECT 933.410 227.840 933.730 227.900 ;
        RECT 973.430 227.840 973.750 227.900 ;
        RECT 2618.850 228.040 2619.170 228.100 ;
        RECT 3367.730 228.040 3368.050 228.100 ;
        RECT 2618.850 227.900 3368.050 228.040 ;
        RECT 2618.850 227.840 2619.170 227.900 ;
        RECT 3367.730 227.840 3368.050 227.900 ;
        RECT 224.550 227.700 224.870 227.760 ;
        RECT 979.870 227.700 980.190 227.760 ;
        RECT 224.550 227.560 980.190 227.700 ;
        RECT 224.550 227.500 224.870 227.560 ;
        RECT 979.870 227.500 980.190 227.560 ;
        RECT 2593.550 227.700 2593.870 227.760 ;
        RECT 3368.650 227.700 3368.970 227.760 ;
        RECT 2593.550 227.560 3368.970 227.700 ;
        RECT 2593.550 227.500 2593.870 227.560 ;
        RECT 3368.650 227.500 3368.970 227.560 ;
        RECT 1749.910 222.260 1750.230 222.320 ;
        RECT 1796.830 222.260 1797.150 222.320 ;
        RECT 2070.990 222.260 2071.310 222.320 ;
        RECT 1749.910 222.120 2071.310 222.260 ;
        RECT 1749.910 222.060 1750.230 222.120 ;
        RECT 1796.830 222.060 1797.150 222.120 ;
        RECT 2070.990 222.060 2071.310 222.120 ;
        RECT 942.610 221.920 942.930 221.980 ;
        RECT 964.230 221.920 964.550 221.980 ;
        RECT 1485.410 221.920 1485.730 221.980 ;
        RECT 1497.830 221.920 1498.150 221.980 ;
        RECT 1528.650 221.920 1528.970 221.980 ;
        RECT 2344.690 221.920 2345.010 221.980 ;
        RECT 2618.850 221.920 2619.170 221.980 ;
        RECT 942.610 221.780 1007.700 221.920 ;
        RECT 942.610 221.720 942.930 221.780 ;
        RECT 964.230 221.720 964.550 221.780 ;
        RECT 1007.560 221.640 1007.700 221.780 ;
        RECT 1421.330 221.780 1614.670 221.920 ;
        RECT 979.870 221.580 980.190 221.640 ;
        RECT 1007.470 221.580 1007.790 221.640 ;
        RECT 1421.330 221.580 1421.470 221.780 ;
        RECT 1485.410 221.720 1485.730 221.780 ;
        RECT 1497.830 221.720 1498.150 221.780 ;
        RECT 1528.650 221.720 1528.970 221.780 ;
        RECT 979.870 221.440 998.960 221.580 ;
        RECT 979.870 221.380 980.190 221.440 ;
        RECT 998.820 220.900 998.960 221.440 ;
        RECT 1007.470 221.440 1421.470 221.580 ;
        RECT 1476.210 221.580 1476.530 221.640 ;
        RECT 1516.230 221.580 1516.550 221.640 ;
        RECT 1476.210 221.440 1516.550 221.580 ;
        RECT 1614.530 221.580 1614.670 221.780 ;
        RECT 2344.690 221.780 2619.170 221.920 ;
        RECT 2344.690 221.720 2345.010 221.780 ;
        RECT 2618.850 221.720 2619.170 221.780 ;
        RECT 1759.570 221.580 1759.890 221.640 ;
        RECT 1771.990 221.580 1772.310 221.640 ;
        RECT 1802.810 221.580 1803.130 221.640 ;
        RECT 1614.530 221.440 1803.130 221.580 ;
        RECT 1007.470 221.380 1007.790 221.440 ;
        RECT 1476.210 221.380 1476.530 221.440 ;
        RECT 1516.230 221.380 1516.550 221.440 ;
        RECT 1759.570 221.380 1759.890 221.440 ;
        RECT 1771.990 221.380 1772.310 221.440 ;
        RECT 1802.810 221.380 1803.130 221.440 ;
        RECT 2033.730 221.240 2034.050 221.300 ;
        RECT 2307.430 221.240 2307.750 221.300 ;
        RECT 2581.590 221.240 2581.910 221.300 ;
        RECT 2593.550 221.240 2593.870 221.300 ;
        RECT 1904.330 221.100 2593.870 221.240 ;
        RECT 1522.670 220.900 1522.990 220.960 ;
        RECT 1749.910 220.900 1750.230 220.960 ;
        RECT 998.820 220.760 1750.230 220.900 ;
        RECT 1522.670 220.700 1522.990 220.760 ;
        RECT 1749.910 220.700 1750.230 220.760 ;
        RECT 1750.370 220.900 1750.690 220.960 ;
        RECT 1790.390 220.900 1790.710 220.960 ;
        RECT 1750.370 220.760 1790.710 220.900 ;
        RECT 1750.370 220.700 1750.690 220.760 ;
        RECT 1790.390 220.700 1790.710 220.760 ;
        RECT 1802.810 220.900 1803.130 220.960 ;
        RECT 1904.330 220.900 1904.470 221.100 ;
        RECT 2033.730 221.040 2034.050 221.100 ;
        RECT 2307.430 221.040 2307.750 221.100 ;
        RECT 2581.590 221.040 2581.910 221.100 ;
        RECT 2593.550 221.040 2593.870 221.100 ;
        RECT 1802.810 220.760 1904.470 220.900 ;
        RECT 2070.990 220.900 2071.310 220.960 ;
        RECT 2344.690 220.900 2345.010 220.960 ;
        RECT 2070.990 220.760 2345.010 220.900 ;
        RECT 1802.810 220.700 1803.130 220.760 ;
        RECT 2070.990 220.700 2071.310 220.760 ;
        RECT 2344.690 220.700 2345.010 220.760 ;
        RECT 2899.450 213.760 2899.770 213.820 ;
        RECT 3367.270 213.760 3367.590 213.820 ;
        RECT 2899.450 213.620 3367.590 213.760 ;
        RECT 2899.450 213.560 2899.770 213.620 ;
        RECT 3367.270 213.560 3367.590 213.620 ;
        RECT 946.290 209.680 946.610 209.740 ;
        RECT 955.490 209.680 955.810 209.740 ;
        RECT 961.470 209.680 961.790 209.740 ;
        RECT 967.910 209.680 968.230 209.740 ;
        RECT 982.170 209.680 982.490 209.740 ;
        RECT 946.290 209.540 982.490 209.680 ;
        RECT 946.290 209.480 946.610 209.540 ;
        RECT 955.490 209.480 955.810 209.540 ;
        RECT 961.470 209.480 961.790 209.540 ;
        RECT 967.910 209.480 968.230 209.540 ;
        RECT 982.170 209.480 982.490 209.540 ;
        RECT 992.290 209.680 992.610 209.740 ;
        RECT 1000.570 209.680 1000.890 209.740 ;
        RECT 992.290 209.540 1000.890 209.680 ;
        RECT 992.290 209.480 992.610 209.540 ;
        RECT 1000.570 209.480 1000.890 209.540 ;
        RECT 1489.550 209.680 1489.870 209.740 ;
        RECT 1503.350 209.680 1503.670 209.740 ;
        RECT 1489.550 209.540 1503.670 209.680 ;
        RECT 1489.550 209.480 1489.870 209.540 ;
        RECT 1503.350 209.480 1503.670 209.540 ;
        RECT 1511.170 209.680 1511.490 209.740 ;
        RECT 1526.350 209.680 1526.670 209.740 ;
        RECT 1532.790 209.680 1533.110 209.740 ;
        RECT 1543.370 209.680 1543.690 209.740 ;
        RECT 1511.170 209.540 1543.690 209.680 ;
        RECT 1511.170 209.480 1511.490 209.540 ;
        RECT 1526.350 209.480 1526.670 209.540 ;
        RECT 1532.790 209.480 1533.110 209.540 ;
        RECT 1543.370 209.480 1543.690 209.540 ;
        RECT 1763.250 209.680 1763.570 209.740 ;
        RECT 1777.510 209.680 1777.830 209.740 ;
        RECT 1763.250 209.540 1777.830 209.680 ;
        RECT 1763.250 209.480 1763.570 209.540 ;
        RECT 1777.510 209.480 1777.830 209.540 ;
        RECT 1784.870 209.680 1785.190 209.740 ;
        RECT 1799.130 209.680 1799.450 209.740 ;
        RECT 1805.570 209.680 1805.890 209.740 ;
        RECT 1817.530 209.680 1817.850 209.740 ;
        RECT 1784.870 209.540 1817.850 209.680 ;
        RECT 1784.870 209.480 1785.190 209.540 ;
        RECT 1799.130 209.480 1799.450 209.540 ;
        RECT 1805.570 209.480 1805.890 209.540 ;
        RECT 1817.530 209.480 1817.850 209.540 ;
        RECT 2037.410 209.680 2037.730 209.740 ;
        RECT 2051.210 209.680 2051.530 209.740 ;
        RECT 2057.650 209.680 2057.970 209.740 ;
        RECT 2072.830 209.680 2073.150 209.740 ;
        RECT 2079.270 209.680 2079.590 209.740 ;
        RECT 2091.230 209.680 2091.550 209.740 ;
        RECT 2037.410 209.540 2091.550 209.680 ;
        RECT 2037.410 209.480 2037.730 209.540 ;
        RECT 2051.210 209.480 2051.530 209.540 ;
        RECT 2057.650 209.480 2057.970 209.540 ;
        RECT 2072.830 209.480 2073.150 209.540 ;
        RECT 2079.270 209.480 2079.590 209.540 ;
        RECT 2091.230 209.480 2091.550 209.540 ;
        RECT 2311.570 209.680 2311.890 209.740 ;
        RECT 2325.370 209.680 2325.690 209.740 ;
        RECT 2331.810 209.680 2332.130 209.740 ;
        RECT 2346.990 209.680 2347.310 209.740 ;
        RECT 2353.430 209.680 2353.750 209.740 ;
        RECT 2365.390 209.680 2365.710 209.740 ;
        RECT 2311.570 209.540 2365.710 209.680 ;
        RECT 2311.570 209.480 2311.890 209.540 ;
        RECT 2325.370 209.480 2325.690 209.540 ;
        RECT 2331.810 209.480 2332.130 209.540 ;
        RECT 2346.990 209.480 2347.310 209.540 ;
        RECT 2353.430 209.480 2353.750 209.540 ;
        RECT 2365.390 209.480 2365.710 209.540 ;
        RECT 2585.270 209.680 2585.590 209.740 ;
        RECT 2599.530 209.680 2599.850 209.740 ;
        RECT 2605.970 209.680 2606.290 209.740 ;
        RECT 2621.150 209.680 2621.470 209.740 ;
        RECT 2627.590 209.680 2627.910 209.740 ;
        RECT 2639.550 209.680 2639.870 209.740 ;
        RECT 2585.270 209.540 2639.870 209.680 ;
        RECT 2585.270 209.480 2585.590 209.540 ;
        RECT 2599.530 209.480 2599.850 209.540 ;
        RECT 2605.970 209.480 2606.290 209.540 ;
        RECT 2621.150 209.480 2621.470 209.540 ;
        RECT 2627.590 209.480 2627.910 209.540 ;
        RECT 2639.550 209.480 2639.870 209.540 ;
        RECT 731.470 209.340 731.790 209.400 ;
        RECT 2844.250 209.340 2844.570 209.400 ;
        RECT 2899.450 209.340 2899.770 209.400 ;
        RECT 731.470 209.200 2899.770 209.340 ;
        RECT 731.470 209.140 731.790 209.200 ;
        RECT 2844.250 209.140 2844.570 209.200 ;
        RECT 2899.450 209.140 2899.770 209.200 ;
        RECT 994.590 209.000 994.910 209.060 ;
        RECT 1538.770 209.000 1539.090 209.060 ;
        RECT 1812.470 209.000 1812.790 209.060 ;
        RECT 2086.630 209.000 2086.950 209.060 ;
        RECT 2360.790 209.000 2361.110 209.060 ;
        RECT 2633.570 209.000 2633.890 209.060 ;
        RECT 841.730 208.860 1904.470 209.000 ;
        RECT 468.810 207.640 469.130 207.700 ;
        RECT 841.730 207.640 841.870 208.860 ;
        RECT 994.590 208.800 994.910 208.860 ;
        RECT 1538.770 208.800 1539.090 208.860 ;
        RECT 1812.470 208.800 1812.790 208.860 ;
        RECT 468.810 207.500 841.870 207.640 ;
      LAYER met1 ;
        POLYGON 1199.065 208.500 1199.065 207.500 1198.065 207.500 ;
        RECT 1199.065 207.500 1262.345 208.500 ;
      LAYER met1 ;
        RECT 468.810 207.440 469.130 207.500 ;
      LAYER met1 ;
        POLYGON 1198.065 207.500 1198.065 207.440 1198.005 207.440 ;
        RECT 1198.065 207.440 1262.345 207.500 ;
        POLYGON 1198.005 207.440 1198.005 206.845 1197.410 206.845 ;
        RECT 1198.005 206.845 1262.345 207.440 ;
      LAYER met1 ;
        RECT 675.810 201.180 676.130 201.240 ;
        RECT 717.670 201.180 717.990 201.240 ;
        RECT 675.810 201.040 717.990 201.180 ;
        RECT 675.810 200.980 676.130 201.040 ;
        RECT 717.670 200.980 717.990 201.040 ;
        RECT 704.950 200.500 705.270 200.560 ;
        RECT 715.330 200.500 715.650 200.560 ;
        RECT 722.730 200.500 723.050 200.560 ;
        RECT 731.470 200.500 731.790 200.560 ;
        RECT 704.950 200.360 731.790 200.500 ;
        RECT 704.950 200.300 705.270 200.360 ;
        RECT 712.930 200.000 713.070 200.360 ;
        RECT 715.330 200.300 715.650 200.360 ;
        RECT 722.730 200.300 723.050 200.360 ;
        RECT 731.470 200.300 731.790 200.360 ;
      LAYER met1 ;
        RECT 663.000 199.390 704.700 199.815 ;
      LAYER met1 ;
        RECT 704.980 199.670 705.240 200.000 ;
      LAYER met1 ;
        RECT 705.520 199.390 706.565 199.815 ;
      LAYER met1 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met1 ;
        RECT 707.775 199.390 709.490 199.815 ;
      LAYER met1 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met1 ;
        RECT 710.700 199.390 712.585 199.815 ;
        RECT 398.320 198.080 456.965 199.030 ;
        RECT 398.320 197.965 399.460 198.080 ;
        POLYGON 399.460 198.080 399.575 198.080 399.460 197.965 ;
        POLYGON 455.535 198.080 455.650 198.080 455.650 197.965 ;
        RECT 455.650 197.965 456.965 198.080 ;
        RECT 395.380 0.275 468.815 197.965 ;
        RECT 663.000 189.745 712.585 199.390 ;
      LAYER met1 ;
        RECT 712.865 190.025 713.095 200.000 ;
      LAYER met1 ;
        RECT 713.375 199.390 715.060 199.815 ;
      LAYER met1 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met1 ;
        RECT 715.920 199.390 722.585 199.815 ;
      LAYER met1 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met1 ;
        RECT 723.725 199.390 725.175 199.815 ;
      LAYER met1 ;
        RECT 725.455 199.670 725.715 200.000 ;
      LAYER met1 ;
        RECT 725.995 199.390 738.000 199.815 ;
        RECT 713.375 189.745 738.000 199.390 ;
        RECT 663.000 104.105 738.000 189.745 ;
        RECT 932.000 180.515 1012.000 206.845 ;
        RECT 931.885 174.985 1012.000 180.515 ;
        RECT 932.000 169.880 1012.000 174.985 ;
        RECT 931.885 164.275 1012.000 169.880 ;
        RECT 932.000 148.780 1012.000 164.275 ;
        POLYGON 1197.410 206.845 1197.410 204.500 1195.065 204.500 ;
        RECT 1197.410 206.500 1262.345 206.845 ;
        POLYGON 1262.345 208.500 1264.345 206.500 1262.345 206.500 ;
      LAYER met1 ;
        RECT 1904.330 207.640 1904.470 208.860 ;
        RECT 2086.260 208.860 2086.950 209.000 ;
        RECT 2086.260 207.640 2086.400 208.860 ;
        RECT 2086.630 208.800 2086.950 208.860 ;
        RECT 2360.420 208.860 2361.110 209.000 ;
        RECT 2360.420 207.640 2360.560 208.860 ;
        RECT 2360.790 208.800 2361.110 208.860 ;
        RECT 2580.530 208.860 2633.890 209.000 ;
        RECT 2580.530 207.640 2580.670 208.860 ;
        RECT 2633.570 208.800 2633.890 208.860 ;
        RECT 1904.330 207.500 2580.670 207.640 ;
      LAYER met1 ;
        RECT 1197.410 204.500 1264.345 206.500 ;
        RECT 1195.065 200.980 1264.345 204.500 ;
        RECT 1195.065 198.980 1262.345 200.980 ;
        POLYGON 1262.345 200.980 1264.345 200.980 1262.345 198.980 ;
        RECT 1195.065 198.780 1260.505 198.980 ;
        RECT 1195.065 163.510 1204.800 198.780 ;
        RECT 1224.435 198.000 1260.505 198.780 ;
        RECT 1224.435 197.965 1264.345 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 931.885 142.810 1012.000 148.780 ;
        RECT 931.885 127.070 1012.115 142.810 ;
        POLYGON 931.885 127.070 931.940 127.070 931.940 127.015 ;
        RECT 931.940 119.365 1012.115 127.070 ;
        RECT 931.940 110.250 1012.000 119.365 ;
        RECT 931.940 108.520 1012.145 110.250 ;
        RECT 931.940 105.420 1012.000 108.520 ;
        RECT 932.000 104.105 1012.000 105.420 ;
        RECT 662.855 69.780 738.145 104.105 ;
        RECT 931.855 69.780 1012.115 104.105 ;
        RECT 663.000 68.725 738.000 69.780 ;
        RECT 932.000 68.725 1012.000 69.780 ;
        RECT 662.855 29.910 738.145 68.725 ;
        RECT 931.855 29.910 1012.115 68.725 ;
        RECT 663.000 0.790 738.000 29.910 ;
        RECT 932.000 21.100 1012.000 29.910 ;
        RECT 931.980 19.025 1012.000 21.100 ;
        RECT 932.000 0.000 1012.000 19.025 ;
        RECT 1206.000 0.160 1280.880 197.965 ;
        RECT 1475.000 180.515 1555.000 206.845 ;
        RECT 1749.000 180.515 1829.000 206.845 ;
        RECT 2023.000 180.515 2103.000 206.845 ;
        RECT 2297.000 180.515 2377.000 206.845 ;
        RECT 2571.000 180.515 2651.000 206.845 ;
        RECT 2849.320 198.080 2907.965 199.030 ;
        RECT 2849.320 197.965 2850.460 198.080 ;
        POLYGON 2850.460 198.080 2850.575 198.080 2850.460 197.965 ;
        POLYGON 2906.535 198.080 2906.650 198.080 2906.650 197.965 ;
        RECT 2906.650 197.965 2907.965 198.080 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.460 198.080 ;
        POLYGON 3119.460 198.080 3119.575 198.080 3119.460 197.965 ;
        POLYGON 3175.535 198.080 3175.650 198.080 3175.650 197.965 ;
        RECT 3175.650 197.965 3176.965 198.080 ;
        RECT 3180.145 197.965 3185.375 198.870 ;
        RECT 1474.885 174.985 1555.000 180.515 ;
        RECT 1748.885 174.985 1829.000 180.515 ;
        RECT 2022.885 174.985 2103.000 180.515 ;
        RECT 2296.885 174.985 2377.000 180.515 ;
        RECT 2570.885 174.985 2651.000 180.515 ;
        RECT 1475.000 169.880 1555.000 174.985 ;
        RECT 1749.000 169.880 1829.000 174.985 ;
        RECT 2023.000 169.880 2103.000 174.985 ;
        RECT 2297.000 169.880 2377.000 174.985 ;
        RECT 2571.000 169.880 2651.000 174.985 ;
        RECT 1474.885 164.275 1555.000 169.880 ;
        RECT 1748.885 164.275 1829.000 169.880 ;
        RECT 2022.885 164.275 2103.000 169.880 ;
        RECT 2296.885 164.275 2377.000 169.880 ;
        RECT 2570.885 164.275 2651.000 169.880 ;
        RECT 1475.000 148.780 1555.000 164.275 ;
        RECT 1749.000 148.780 1829.000 164.275 ;
        RECT 2023.000 148.780 2103.000 164.275 ;
        RECT 2297.000 148.780 2377.000 164.275 ;
        RECT 2571.000 148.780 2651.000 164.275 ;
        RECT 1474.885 142.810 1555.000 148.780 ;
        RECT 1748.885 142.810 1829.000 148.780 ;
        RECT 2022.885 142.810 2103.000 148.780 ;
        RECT 2296.885 142.810 2377.000 148.780 ;
        RECT 2570.885 142.810 2651.000 148.780 ;
        RECT 1474.885 127.070 1555.115 142.810 ;
        POLYGON 1474.885 127.070 1474.940 127.070 1474.940 127.015 ;
        RECT 1474.940 119.365 1555.115 127.070 ;
        RECT 1748.885 127.070 1829.115 142.810 ;
        POLYGON 1748.885 127.070 1748.940 127.070 1748.940 127.015 ;
        RECT 1748.940 119.365 1829.115 127.070 ;
        RECT 2022.885 127.070 2103.115 142.810 ;
        POLYGON 2022.885 127.070 2022.940 127.070 2022.940 127.015 ;
        RECT 2022.940 119.365 2103.115 127.070 ;
        RECT 2296.885 127.070 2377.115 142.810 ;
        POLYGON 2296.885 127.070 2296.940 127.070 2296.940 127.015 ;
        RECT 2296.940 119.365 2377.115 127.070 ;
        RECT 2570.885 127.070 2651.115 142.810 ;
        POLYGON 2570.885 127.070 2570.940 127.070 2570.940 127.015 ;
        RECT 2570.940 119.365 2651.115 127.070 ;
        RECT 1474.940 110.250 1555.000 119.365 ;
        RECT 1748.940 110.250 1829.000 119.365 ;
        RECT 2022.940 110.250 2103.000 119.365 ;
        RECT 2296.940 110.250 2377.000 119.365 ;
        RECT 2570.940 110.250 2651.000 119.365 ;
        RECT 1474.940 108.520 1555.145 110.250 ;
        RECT 1748.940 108.520 1829.145 110.250 ;
        RECT 2022.940 108.520 2103.145 110.250 ;
        RECT 2296.940 108.520 2377.145 110.250 ;
        RECT 2570.940 108.520 2651.145 110.250 ;
        RECT 1474.940 105.420 1555.000 108.520 ;
        RECT 1748.940 105.420 1829.000 108.520 ;
        RECT 2022.940 105.420 2103.000 108.520 ;
        RECT 2296.940 105.420 2377.000 108.520 ;
        RECT 2570.940 105.420 2651.000 108.520 ;
        RECT 1475.000 104.105 1555.000 105.420 ;
        RECT 1749.000 104.105 1829.000 105.420 ;
        RECT 2023.000 104.105 2103.000 105.420 ;
        RECT 2297.000 104.105 2377.000 105.420 ;
        RECT 2571.000 104.105 2651.000 105.420 ;
        RECT 1474.855 69.780 1555.115 104.105 ;
        RECT 1748.855 69.780 1829.115 104.105 ;
        RECT 2022.855 69.780 2103.115 104.105 ;
        RECT 2296.855 69.780 2377.115 104.105 ;
        RECT 2570.855 69.780 2651.115 104.105 ;
        RECT 1475.000 68.725 1555.000 69.780 ;
        RECT 1749.000 68.725 1829.000 69.780 ;
        RECT 2023.000 68.725 2103.000 69.780 ;
        RECT 2297.000 68.725 2377.000 69.780 ;
        RECT 2571.000 68.725 2651.000 69.780 ;
        RECT 1474.855 29.910 1555.115 68.725 ;
        RECT 1748.855 29.910 1829.115 68.725 ;
        RECT 2022.855 29.910 2103.115 68.725 ;
        RECT 2296.855 29.910 2377.115 68.725 ;
        RECT 2570.855 29.910 2651.115 68.725 ;
        RECT 1475.000 21.100 1555.000 29.910 ;
        RECT 1749.000 21.100 1829.000 29.910 ;
        RECT 2023.000 21.100 2103.000 29.910 ;
        RECT 2297.000 21.100 2377.000 29.910 ;
        RECT 2571.000 21.100 2651.000 29.910 ;
        RECT 1474.980 19.025 1555.000 21.100 ;
        RECT 1748.980 19.025 1829.000 21.100 ;
        RECT 2022.980 19.025 2103.000 21.100 ;
        RECT 2296.980 19.025 2377.000 21.100 ;
        RECT 2570.980 19.025 2651.000 21.100 ;
        RECT 1475.000 0.000 1555.000 19.025 ;
        RECT 1749.000 0.000 1829.000 19.025 ;
        RECT 2023.000 0.000 2103.000 19.025 ;
        RECT 2297.000 0.000 2377.000 19.025 ;
        RECT 2571.000 0.000 2651.000 19.025 ;
        RECT 2846.380 0.275 2919.815 197.965 ;
        RECT 3116.085 0.275 3188.815 197.965 ;
      LAYER via ;
        RECT 2928.920 4982.060 2929.180 4982.320 ;
        RECT 3373.740 4982.060 3374.000 4982.320 ;
        RECT 211.240 4981.720 211.500 4981.980 ;
        RECT 1697.500 4981.720 1697.760 4981.980 ;
        RECT 3367.760 4981.720 3368.020 4981.980 ;
        RECT 224.580 4950.440 224.840 4950.700 ;
        RECT 3368.220 4950.440 3368.480 4950.700 ;
        RECT 211.700 4950.100 211.960 4950.360 ;
        RECT 3367.300 4950.100 3367.560 4950.360 ;
        RECT 212.160 4305.800 212.420 4306.060 ;
        RECT 220.900 4305.800 221.160 4306.060 ;
        RECT 3367.760 4295.600 3368.020 4295.860 ;
        RECT 3376.960 4295.600 3377.220 4295.860 ;
        RECT 3368.220 4280.300 3368.480 4280.560 ;
        RECT 3376.960 4280.300 3377.220 4280.560 ;
        RECT 3367.300 4248.340 3367.560 4248.600 ;
        RECT 3376.960 4248.340 3377.220 4248.600 ;
        RECT 3376.500 4018.840 3376.760 4019.100 ;
        RECT 3388.000 4018.840 3388.260 4019.100 ;
        RECT 211.240 4004.900 211.500 4005.160 ;
        RECT 213.080 4004.900 213.340 4005.160 ;
        RECT 208.940 3992.660 209.200 3992.920 ;
        RECT 211.700 3992.660 211.960 3992.920 ;
        RECT 208.940 3960.360 209.200 3960.620 ;
        RECT 212.160 3960.360 212.420 3960.620 ;
        RECT 208.940 3945.400 209.200 3945.660 ;
        RECT 213.080 3945.400 213.340 3945.660 ;
        RECT 3367.760 3863.800 3368.020 3864.060 ;
        RECT 3376.960 3863.800 3377.220 3864.060 ;
        RECT 3368.220 3848.160 3368.480 3848.420 ;
        RECT 3369.600 3848.160 3369.860 3848.420 ;
        RECT 3376.960 3848.160 3377.220 3848.420 ;
        RECT 3376.040 3837.960 3376.300 3838.220 ;
        RECT 3376.960 3837.960 3377.220 3838.220 ;
        RECT 3367.300 3806.340 3367.560 3806.600 ;
        RECT 3370.060 3806.340 3370.320 3806.600 ;
        RECT 3376.960 3806.340 3377.220 3806.600 ;
        RECT 3376.040 3800.900 3376.300 3801.160 ;
        RECT 3376.960 3800.900 3377.220 3801.160 ;
        RECT 208.940 3781.180 209.200 3781.440 ;
        RECT 211.700 3781.180 211.960 3781.440 ;
        RECT 213.080 3781.180 213.340 3781.440 ;
        RECT 208.940 3741.400 209.200 3741.660 ;
        RECT 212.620 3741.400 212.880 3741.660 ;
        RECT 208.940 3724.060 209.200 3724.320 ;
        RECT 212.160 3724.060 212.420 3724.320 ;
        RECT 213.540 3724.060 213.800 3724.320 ;
        RECT 3367.760 3641.780 3368.020 3642.040 ;
        RECT 3376.960 3641.780 3377.220 3642.040 ;
        RECT 3369.600 3626.140 3369.860 3626.400 ;
        RECT 3376.960 3626.140 3377.220 3626.400 ;
        RECT 3368.220 3589.080 3368.480 3589.340 ;
        RECT 3370.060 3589.080 3370.320 3589.340 ;
        RECT 3376.960 3589.080 3377.220 3589.340 ;
        RECT 208.940 3565.280 209.200 3565.540 ;
        RECT 213.080 3565.280 213.340 3565.540 ;
        RECT 208.940 3523.800 209.200 3524.060 ;
        RECT 212.620 3523.800 212.880 3524.060 ;
        RECT 208.940 3508.160 209.200 3508.420 ;
        RECT 212.160 3508.160 212.420 3508.420 ;
        RECT 3367.760 3415.340 3368.020 3415.600 ;
        RECT 3368.680 3415.340 3368.940 3415.600 ;
        RECT 3376.960 3415.340 3377.220 3415.600 ;
        RECT 3367.760 3402.080 3368.020 3402.340 ;
        RECT 3369.600 3402.080 3369.860 3402.340 ;
        RECT 3376.960 3402.080 3377.220 3402.340 ;
        RECT 3376.040 3393.920 3376.300 3394.180 ;
        RECT 3376.960 3393.920 3377.220 3394.180 ;
        RECT 3368.220 3368.080 3368.480 3368.340 ;
        RECT 3370.060 3368.080 3370.320 3368.340 ;
        RECT 3376.960 3368.080 3377.220 3368.340 ;
        RECT 208.940 3343.600 209.200 3343.860 ;
        RECT 213.080 3343.600 213.340 3343.860 ;
        RECT 208.940 3306.540 209.200 3306.800 ;
        RECT 212.620 3306.540 212.880 3306.800 ;
        RECT 208.940 3296.340 209.200 3296.600 ;
        RECT 212.160 3296.340 212.420 3296.600 ;
        RECT 213.540 3296.340 213.800 3296.600 ;
        RECT 3368.220 3194.340 3368.480 3194.600 ;
        RECT 3376.960 3194.340 3377.220 3194.600 ;
        RECT 3367.760 3181.420 3368.020 3181.680 ;
        RECT 3376.960 3181.420 3377.220 3181.680 ;
        RECT 3376.040 3172.920 3376.300 3173.180 ;
        RECT 3376.960 3172.920 3377.220 3173.180 ;
        RECT 3367.300 3147.080 3367.560 3147.340 ;
        RECT 3370.060 3147.080 3370.320 3147.340 ;
        RECT 3376.960 3147.080 3377.220 3147.340 ;
        RECT 208.940 3127.360 209.200 3127.620 ;
        RECT 213.080 3127.360 213.340 3127.620 ;
        RECT 208.940 3090.640 209.200 3090.900 ;
        RECT 212.620 3090.640 212.880 3090.900 ;
        RECT 208.940 3075.000 209.200 3075.260 ;
        RECT 213.540 3075.000 213.800 3075.260 ;
        RECT 211.240 3073.300 211.500 3073.560 ;
        RECT 3368.220 2975.720 3368.480 2975.980 ;
        RECT 3376.960 2975.720 3377.220 2975.980 ;
        RECT 3367.760 2959.400 3368.020 2959.660 ;
        RECT 3376.960 2959.400 3377.220 2959.660 ;
        RECT 3367.300 2920.640 3367.560 2920.900 ;
        RECT 3369.600 2920.640 3369.860 2920.900 ;
        RECT 3376.960 2920.640 3377.220 2920.900 ;
        RECT 208.940 2916.220 209.200 2916.480 ;
        RECT 213.080 2916.220 213.340 2916.480 ;
        RECT 208.940 2879.500 209.200 2879.760 ;
        RECT 212.620 2879.500 212.880 2879.760 ;
        RECT 208.940 2859.100 209.200 2859.360 ;
        RECT 212.160 2859.100 212.420 2859.360 ;
        RECT 3368.220 2756.760 3368.480 2757.020 ;
        RECT 3376.960 2756.760 3377.220 2757.020 ;
        RECT 3367.760 2741.120 3368.020 2741.380 ;
        RECT 3376.960 2741.120 3377.220 2741.380 ;
        RECT 3369.600 2704.400 3369.860 2704.660 ;
        RECT 3376.960 2704.400 3377.220 2704.660 ;
        RECT 208.940 2700.320 209.200 2700.580 ;
        RECT 213.080 2700.320 213.340 2700.580 ;
        RECT 208.940 2658.840 209.200 2659.100 ;
        RECT 212.620 2658.840 212.880 2659.100 ;
        RECT 213.540 2658.840 213.800 2659.100 ;
        RECT 208.940 2643.200 209.200 2643.460 ;
        RECT 212.160 2643.200 212.420 2643.460 ;
        RECT 3376.500 2497.340 3376.760 2497.600 ;
        RECT 3380.640 2497.340 3380.900 2497.600 ;
        RECT 3380.640 2474.220 3380.900 2474.480 ;
        RECT 3389.840 2474.220 3390.100 2474.480 ;
        RECT 3370.060 2111.100 3370.320 2111.360 ;
        RECT 3373.740 2111.100 3374.000 2111.360 ;
        RECT 3370.060 2095.800 3370.320 2096.060 ;
        RECT 3387.540 2095.800 3387.800 2096.060 ;
        RECT 208.940 2056.360 209.200 2056.620 ;
        RECT 212.620 2056.360 212.880 2056.620 ;
        RECT 208.940 2024.400 209.200 2024.660 ;
        RECT 213.540 2024.400 213.800 2024.660 ;
        RECT 208.940 2009.440 209.200 2009.700 ;
        RECT 212.160 2009.440 212.420 2009.700 ;
        RECT 3369.600 1880.580 3369.860 1880.840 ;
        RECT 3376.960 1880.580 3377.220 1880.840 ;
        RECT 3368.680 1865.280 3368.940 1865.540 ;
        RECT 3376.960 1865.280 3377.220 1865.540 ;
        RECT 208.940 1845.220 209.200 1845.480 ;
        RECT 212.620 1845.220 212.880 1845.480 ;
        RECT 3370.060 1828.560 3370.320 1828.820 ;
        RECT 3376.960 1828.560 3377.220 1828.820 ;
        RECT 208.940 1806.460 209.200 1806.720 ;
        RECT 213.080 1806.460 213.340 1806.720 ;
        RECT 208.940 1788.100 209.200 1788.360 ;
        RECT 212.160 1788.100 212.420 1788.360 ;
        RECT 213.540 1788.100 213.800 1788.360 ;
        RECT 3368.680 1669.780 3368.940 1670.040 ;
        RECT 3376.040 1669.780 3376.300 1670.040 ;
        RECT 3367.300 1659.580 3367.560 1659.840 ;
        RECT 3369.600 1659.580 3369.860 1659.840 ;
        RECT 3376.960 1659.580 3377.220 1659.840 ;
        RECT 3367.760 1644.280 3368.020 1644.540 ;
        RECT 3376.040 1644.280 3376.300 1644.540 ;
        RECT 3376.960 1644.280 3377.220 1644.540 ;
        RECT 208.940 1628.300 209.200 1628.560 ;
        RECT 212.620 1628.300 212.880 1628.560 ;
        RECT 3368.220 1612.320 3368.480 1612.580 ;
        RECT 3370.060 1612.320 3370.320 1612.580 ;
        RECT 3376.960 1612.320 3377.220 1612.580 ;
        RECT 208.940 1586.820 209.200 1587.080 ;
        RECT 213.080 1586.820 213.340 1587.080 ;
        RECT 208.940 1571.180 209.200 1571.440 ;
        RECT 212.620 1571.180 212.880 1571.440 ;
        RECT 213.540 1571.180 213.800 1571.440 ;
        RECT 3367.300 1443.680 3367.560 1443.940 ;
        RECT 3376.960 1443.680 3377.220 1443.940 ;
        RECT 3367.760 1426.340 3368.020 1426.600 ;
        RECT 3376.960 1426.340 3377.220 1426.600 ;
        RECT 208.940 1407.640 209.200 1407.900 ;
        RECT 212.160 1407.640 212.420 1407.900 ;
        RECT 213.540 1407.640 213.800 1407.900 ;
        RECT 3368.220 1386.560 3368.480 1386.820 ;
        RECT 3376.960 1386.560 3377.220 1386.820 ;
        RECT 208.940 1373.300 209.200 1373.560 ;
        RECT 213.080 1373.300 213.340 1373.560 ;
        RECT 208.940 1360.380 209.200 1360.640 ;
        RECT 212.620 1360.380 212.880 1360.640 ;
        RECT 3367.300 1218.600 3367.560 1218.860 ;
        RECT 3376.960 1218.600 3377.220 1218.860 ;
        RECT 3367.760 1201.260 3368.020 1201.520 ;
        RECT 3376.960 1201.260 3377.220 1201.520 ;
        RECT 208.940 1191.400 209.200 1191.660 ;
        RECT 212.160 1191.400 212.420 1191.660 ;
        RECT 213.540 1191.400 213.800 1191.660 ;
        RECT 3368.220 1169.300 3368.480 1169.560 ;
        RECT 3376.960 1169.300 3377.220 1169.560 ;
        RECT 208.940 1159.440 209.200 1159.700 ;
        RECT 213.080 1159.440 213.340 1159.700 ;
        RECT 208.940 1144.140 209.200 1144.400 ;
        RECT 212.620 1144.140 212.880 1144.400 ;
        RECT 3367.300 995.560 3367.560 995.820 ;
        RECT 3376.960 995.560 3377.220 995.820 ;
        RECT 3367.760 985.020 3368.020 985.280 ;
        RECT 3376.960 985.020 3377.220 985.280 ;
        RECT 208.940 975.500 209.200 975.760 ;
        RECT 212.160 975.500 212.420 975.760 ;
        RECT 3368.220 946.260 3368.480 946.520 ;
        RECT 3376.960 946.260 3377.220 946.520 ;
        RECT 208.940 943.540 209.200 943.800 ;
        RECT 212.620 943.540 212.880 943.800 ;
        RECT 214.000 943.540 214.260 943.800 ;
        RECT 208.940 928.240 209.200 928.500 ;
        RECT 213.540 928.240 213.800 928.500 ;
        RECT 211.240 921.780 211.500 922.040 ;
        RECT 213.540 921.780 213.800 922.040 ;
        RECT 3367.300 779.660 3367.560 779.920 ;
        RECT 3369.600 779.660 3369.860 779.920 ;
        RECT 3376.960 779.660 3377.220 779.920 ;
        RECT 3367.760 764.020 3368.020 764.280 ;
        RECT 3376.960 764.020 3377.220 764.280 ;
        RECT 3368.680 722.540 3368.940 722.800 ;
        RECT 3376.960 722.540 3377.220 722.800 ;
        RECT 212.620 607.280 212.880 607.540 ;
        RECT 220.900 607.280 221.160 607.540 ;
        RECT 3367.300 557.640 3367.560 557.900 ;
        RECT 3369.600 557.640 3369.860 557.900 ;
        RECT 3376.960 557.640 3377.220 557.900 ;
        RECT 3367.760 542.000 3368.020 542.260 ;
        RECT 3376.960 542.000 3377.220 542.260 ;
        RECT 212.160 530.100 212.420 530.360 ;
        RECT 220.900 530.100 221.160 530.360 ;
        RECT 224.120 234.640 224.380 234.900 ;
        RECT 717.700 234.300 717.960 234.560 ;
        RECT 1004.280 234.300 1004.540 234.560 ;
        RECT 1281.200 234.300 1281.460 234.560 ;
        RECT 1488.660 234.300 1488.920 234.560 ;
        RECT 1547.080 234.300 1547.340 234.560 ;
        RECT 1762.820 234.300 1763.080 234.560 ;
        RECT 1821.240 234.300 1821.500 234.560 ;
        RECT 2036.980 234.300 2037.240 234.560 ;
        RECT 2095.400 234.300 2095.660 234.560 ;
        RECT 2310.680 234.300 2310.940 234.560 ;
        RECT 2369.100 234.300 2369.360 234.560 ;
        RECT 2584.840 234.300 2585.100 234.560 ;
        RECT 211.240 228.180 211.500 228.440 ;
        RECT 704.820 228.180 705.080 228.440 ;
        RECT 933.440 227.840 933.700 228.100 ;
        RECT 973.460 227.840 973.720 228.100 ;
        RECT 2618.880 227.840 2619.140 228.100 ;
        RECT 3367.760 227.840 3368.020 228.100 ;
        RECT 224.580 227.500 224.840 227.760 ;
        RECT 979.900 227.500 980.160 227.760 ;
        RECT 2593.580 227.500 2593.840 227.760 ;
        RECT 3368.680 227.500 3368.940 227.760 ;
        RECT 1749.940 222.060 1750.200 222.320 ;
        RECT 1796.860 222.060 1797.120 222.320 ;
        RECT 2071.020 222.060 2071.280 222.320 ;
        RECT 942.640 221.720 942.900 221.980 ;
        RECT 964.260 221.720 964.520 221.980 ;
        RECT 979.900 221.380 980.160 221.640 ;
        RECT 1007.500 221.380 1007.760 221.640 ;
        RECT 1485.440 221.720 1485.700 221.980 ;
        RECT 1497.860 221.720 1498.120 221.980 ;
        RECT 1528.680 221.720 1528.940 221.980 ;
        RECT 1476.240 221.380 1476.500 221.640 ;
        RECT 1516.260 221.380 1516.520 221.640 ;
        RECT 2344.720 221.720 2344.980 221.980 ;
        RECT 2618.880 221.720 2619.140 221.980 ;
        RECT 1759.600 221.380 1759.860 221.640 ;
        RECT 1772.020 221.380 1772.280 221.640 ;
        RECT 1802.840 221.380 1803.100 221.640 ;
        RECT 1522.700 220.700 1522.960 220.960 ;
        RECT 1749.940 220.700 1750.200 220.960 ;
        RECT 1750.400 220.700 1750.660 220.960 ;
        RECT 1790.420 220.700 1790.680 220.960 ;
        RECT 1802.840 220.700 1803.100 220.960 ;
        RECT 2033.760 221.040 2034.020 221.300 ;
        RECT 2307.460 221.040 2307.720 221.300 ;
        RECT 2581.620 221.040 2581.880 221.300 ;
        RECT 2593.580 221.040 2593.840 221.300 ;
        RECT 2071.020 220.700 2071.280 220.960 ;
        RECT 2344.720 220.700 2344.980 220.960 ;
        RECT 2899.480 213.560 2899.740 213.820 ;
        RECT 3367.300 213.560 3367.560 213.820 ;
        RECT 946.320 209.480 946.580 209.740 ;
        RECT 955.520 209.480 955.780 209.740 ;
        RECT 961.500 209.480 961.760 209.740 ;
        RECT 967.940 209.480 968.200 209.740 ;
        RECT 982.200 209.480 982.460 209.740 ;
        RECT 992.320 209.480 992.580 209.740 ;
        RECT 1000.600 209.480 1000.860 209.740 ;
        RECT 1489.580 209.480 1489.840 209.740 ;
        RECT 1503.380 209.480 1503.640 209.740 ;
        RECT 1511.200 209.480 1511.460 209.740 ;
        RECT 1526.380 209.480 1526.640 209.740 ;
        RECT 1532.820 209.480 1533.080 209.740 ;
        RECT 1543.400 209.480 1543.660 209.740 ;
        RECT 1763.280 209.480 1763.540 209.740 ;
        RECT 1777.540 209.480 1777.800 209.740 ;
        RECT 1784.900 209.480 1785.160 209.740 ;
        RECT 1799.160 209.480 1799.420 209.740 ;
        RECT 1805.600 209.480 1805.860 209.740 ;
        RECT 1817.560 209.480 1817.820 209.740 ;
        RECT 2037.440 209.480 2037.700 209.740 ;
        RECT 2051.240 209.480 2051.500 209.740 ;
        RECT 2057.680 209.480 2057.940 209.740 ;
        RECT 2072.860 209.480 2073.120 209.740 ;
        RECT 2079.300 209.480 2079.560 209.740 ;
        RECT 2091.260 209.480 2091.520 209.740 ;
        RECT 2311.600 209.480 2311.860 209.740 ;
        RECT 2325.400 209.480 2325.660 209.740 ;
        RECT 2331.840 209.480 2332.100 209.740 ;
        RECT 2347.020 209.480 2347.280 209.740 ;
        RECT 2353.460 209.480 2353.720 209.740 ;
        RECT 2365.420 209.480 2365.680 209.740 ;
        RECT 2585.300 209.480 2585.560 209.740 ;
        RECT 2599.560 209.480 2599.820 209.740 ;
        RECT 2606.000 209.480 2606.260 209.740 ;
        RECT 2621.180 209.480 2621.440 209.740 ;
        RECT 2627.620 209.480 2627.880 209.740 ;
        RECT 2639.580 209.480 2639.840 209.740 ;
        RECT 731.500 209.140 731.760 209.400 ;
        RECT 2844.280 209.140 2844.540 209.400 ;
        RECT 2899.480 209.140 2899.740 209.400 ;
        RECT 468.840 207.440 469.100 207.700 ;
        RECT 994.620 208.800 994.880 209.060 ;
        RECT 1538.800 208.800 1539.060 209.060 ;
        RECT 1812.500 208.800 1812.760 209.060 ;
        RECT 675.840 200.980 676.100 201.240 ;
        RECT 717.700 200.980 717.960 201.240 ;
        RECT 704.980 200.300 705.240 200.560 ;
        RECT 715.360 200.300 715.620 200.560 ;
        RECT 722.760 200.300 723.020 200.560 ;
        RECT 731.500 200.300 731.760 200.560 ;
        RECT 2086.660 208.800 2086.920 209.060 ;
        RECT 2360.820 208.800 2361.080 209.060 ;
        RECT 2633.600 208.800 2633.860 209.060 ;
      LAYER met2 ;
        RECT 379.250 5034.255 445.440 5036.855 ;
        RECT 619.250 5034.255 685.440 5036.855 ;
        RECT 859.250 5034.255 925.440 5036.855 ;
        RECT 1147.265 5013.940 1221.290 5183.075 ;
        RECT 1404.265 5013.940 1478.290 5183.075 ;
        RECT 1147.265 4990.335 1197.110 5013.940 ;
        RECT 1404.265 4990.335 1454.110 5013.940 ;
        RECT 1171.675 4990.035 1197.110 4990.335 ;
        RECT 1428.675 4990.035 1454.110 4990.335 ;
        RECT 1697.265 4990.035 1771.290 5183.075 ;
        RECT 2128.250 5034.255 2194.440 5036.855 ;
        RECT 2375.250 5034.255 2441.440 5036.855 ;
        RECT 2633.250 5034.255 2699.440 5036.855 ;
        RECT 2878.265 4990.035 2952.290 5183.075 ;
        RECT 3139.250 5034.255 3205.440 5036.855 ;
        RECT 1172.895 4988.000 1174.895 4989.920 ;
        RECT 1429.895 4988.000 1431.895 4989.920 ;
        RECT 1697.495 4988.000 1721.395 4990.035 ;
        RECT 1722.895 4988.000 1724.895 4989.920 ;
        RECT 1747.390 4988.000 1771.290 4990.035 ;
        RECT 2878.495 4988.000 2902.395 4990.035 ;
        RECT 2903.895 4988.000 2905.895 4989.920 ;
        RECT 2928.390 4988.000 2952.290 4990.035 ;
      LAYER met2 ;
        RECT 2928.910 4987.275 2929.190 4987.645 ;
        RECT 1697.490 4985.235 1697.770 4985.605 ;
        RECT 1697.560 4982.010 1697.700 4985.235 ;
        RECT 2928.980 4982.350 2929.120 4987.275 ;
        RECT 2928.920 4982.030 2929.180 4982.350 ;
        RECT 3373.740 4982.030 3374.000 4982.350 ;
        RECT 211.240 4981.690 211.500 4982.010 ;
        RECT 1697.500 4981.690 1697.760 4982.010 ;
        RECT 3367.760 4981.690 3368.020 4982.010 ;
      LAYER met2 ;
        RECT 151.145 4780.250 153.745 4846.440 ;
        RECT 0.035 4641.200 151.405 4650.935 ;
        RECT 153.765 4640.000 158.415 4651.140 ;
        RECT 160.165 4641.200 174.575 4650.935 ;
        RECT 0.035 4639.700 197.965 4640.000 ;
        RECT 0.035 4619.095 198.000 4639.700 ;
        RECT 0.035 4618.535 197.965 4619.095 ;
        RECT 0.035 4585.925 198.000 4618.535 ;
        RECT 0.035 4585.495 197.965 4585.925 ;
        RECT 0.035 4565.500 198.000 4585.495 ;
        RECT 0.035 4565.000 197.965 4565.500 ;
        RECT 153.800 4554.025 158.450 4565.000 ;
        RECT 4.925 4404.390 200.000 4428.290 ;
        RECT 4.925 4378.395 197.965 4404.390 ;
        RECT 198.080 4379.895 200.000 4381.895 ;
        RECT 4.925 4354.495 200.000 4378.395 ;
        RECT 4.925 4354.265 197.965 4354.495 ;
        RECT 4.925 4192.390 200.000 4216.290 ;
        RECT 4.925 4166.395 197.965 4192.390 ;
        RECT 198.080 4167.895 200.000 4169.895 ;
        RECT 4.925 4142.495 200.000 4166.395 ;
        RECT 4.925 4142.265 197.965 4142.495 ;
        RECT 0.000 4004.865 208.565 4005.915 ;
      LAYER met2 ;
        RECT 211.300 4005.190 211.440 4981.690 ;
        RECT 224.580 4950.410 224.840 4950.730 ;
        RECT 211.700 4950.070 211.960 4950.390 ;
        RECT 211.240 4004.870 211.500 4005.190 ;
      LAYER met2 ;
        RECT 0.000 4004.025 208.285 4004.865 ;
      LAYER met2 ;
        RECT 208.565 4004.515 210.965 4004.585 ;
        RECT 208.565 4004.375 211.440 4004.515 ;
        RECT 208.565 4004.305 210.965 4004.375 ;
      LAYER met2 ;
        RECT 0.000 4001.645 208.565 4004.025 ;
        RECT 0.000 4000.805 208.285 4001.645 ;
        RECT 0.000 3998.425 208.565 4000.805 ;
        RECT 0.000 3997.585 208.285 3998.425 ;
      LAYER met2 ;
        RECT 208.565 3997.865 210.965 3998.145 ;
      LAYER met2 ;
        RECT 0.000 3995.665 208.565 3997.585 ;
        RECT 0.000 3994.825 208.285 3995.665 ;
      LAYER met2 ;
        RECT 208.610 3995.385 209.140 3995.410 ;
        RECT 208.565 3995.105 210.965 3995.385 ;
      LAYER met2 ;
        RECT 0.000 3992.445 208.565 3994.825 ;
      LAYER met2 ;
        RECT 209.000 3992.950 209.140 3995.105 ;
        RECT 208.940 3992.630 209.200 3992.950 ;
      LAYER met2 ;
        RECT 0.000 3991.605 208.285 3992.445 ;
        RECT 0.000 3989.225 208.565 3991.605 ;
        RECT 0.000 3988.385 208.285 3989.225 ;
        RECT 0.000 3986.465 208.565 3988.385 ;
        RECT 0.000 3985.625 208.285 3986.465 ;
      LAYER met2 ;
        RECT 208.565 3985.905 210.965 3986.185 ;
      LAYER met2 ;
        RECT 0.000 3983.245 208.565 3985.625 ;
        RECT 0.000 3982.405 208.285 3983.245 ;
        RECT 0.000 3980.025 208.565 3982.405 ;
        RECT 0.000 3979.185 208.285 3980.025 ;
        RECT 0.000 3977.265 208.565 3979.185 ;
        RECT 0.000 3976.425 208.285 3977.265 ;
        RECT 0.000 3974.045 208.565 3976.425 ;
        RECT 0.000 3973.205 208.285 3974.045 ;
        RECT 0.000 3970.825 208.565 3973.205 ;
        RECT 0.000 3969.985 208.285 3970.825 ;
        RECT 0.000 3968.065 208.565 3969.985 ;
        RECT 0.000 3967.225 208.285 3968.065 ;
        RECT 0.000 3964.845 208.565 3967.225 ;
      LAYER met2 ;
        RECT 211.300 3965.490 211.440 4004.375 ;
        RECT 211.760 3992.950 211.900 4950.070 ;
        RECT 224.640 4512.670 224.780 4950.410 ;
        RECT 3367.300 4950.070 3367.560 4950.390 ;
        RECT 224.180 4512.530 224.780 4512.670 ;
        RECT 224.180 4429.365 224.320 4512.530 ;
        RECT 220.890 4428.995 221.170 4429.365 ;
        RECT 224.110 4428.995 224.390 4429.365 ;
        RECT 220.960 4355.245 221.100 4428.995 ;
        RECT 220.890 4354.875 221.170 4355.245 ;
        RECT 220.960 4306.090 221.100 4354.875 ;
        RECT 212.160 4305.770 212.420 4306.090 ;
        RECT 220.900 4305.770 221.160 4306.090 ;
        RECT 211.700 3992.630 211.960 3992.950 ;
        RECT 209.000 3965.350 211.440 3965.490 ;
      LAYER met2 ;
        RECT 0.000 3964.005 208.285 3964.845 ;
      LAYER met2 ;
        RECT 209.000 3964.565 209.140 3965.350 ;
        RECT 208.565 3964.285 210.965 3964.565 ;
      LAYER met2 ;
        RECT 0.000 3961.625 208.565 3964.005 ;
        RECT 0.000 3960.785 208.285 3961.625 ;
        RECT 0.000 3958.405 208.565 3960.785 ;
      LAYER met2 ;
        RECT 208.940 3960.330 209.200 3960.650 ;
      LAYER met2 ;
        RECT 0.000 3957.565 208.285 3958.405 ;
      LAYER met2 ;
        RECT 209.000 3958.125 209.140 3960.330 ;
        RECT 208.565 3957.845 210.965 3958.125 ;
      LAYER met2 ;
        RECT 0.000 3955.645 208.565 3957.565 ;
        RECT 0.000 3954.805 208.285 3955.645 ;
        RECT 0.000 3952.425 208.565 3954.805 ;
        RECT 0.000 3951.585 208.285 3952.425 ;
        RECT 0.000 3949.205 208.565 3951.585 ;
        RECT 0.000 3948.365 208.285 3949.205 ;
        RECT 0.000 3946.445 208.565 3948.365 ;
        RECT 0.000 3945.605 208.285 3946.445 ;
        RECT 0.000 3943.225 208.565 3945.605 ;
      LAYER met2 ;
        RECT 208.940 3945.370 209.200 3945.690 ;
      LAYER met2 ;
        RECT 0.000 3942.385 208.285 3943.225 ;
      LAYER met2 ;
        RECT 209.000 3942.945 209.140 3945.370 ;
        RECT 208.565 3942.665 210.965 3942.945 ;
      LAYER met2 ;
        RECT 0.000 3940.005 208.565 3942.385 ;
        RECT 0.000 3939.165 208.285 3940.005 ;
        RECT 0.000 3937.245 208.565 3939.165 ;
        RECT 0.000 3936.405 208.285 3937.245 ;
        RECT 0.000 3934.025 208.565 3936.405 ;
        RECT 0.000 3933.185 208.285 3934.025 ;
        RECT 0.000 3930.805 208.565 3933.185 ;
        RECT 0.000 3929.965 208.285 3930.805 ;
        RECT 0.000 3928.045 208.565 3929.965 ;
        RECT 0.000 3927.205 208.285 3928.045 ;
        RECT 0.000 3926.210 208.565 3927.205 ;
        RECT 0.000 3788.865 208.565 3789.915 ;
        RECT 0.000 3788.025 208.285 3788.865 ;
      LAYER met2 ;
        RECT 208.565 3788.515 210.965 3788.585 ;
        RECT 208.565 3788.375 211.440 3788.515 ;
        RECT 208.565 3788.305 210.965 3788.375 ;
      LAYER met2 ;
        RECT 0.000 3785.645 208.565 3788.025 ;
        RECT 0.000 3784.805 208.285 3785.645 ;
        RECT 0.000 3782.425 208.565 3784.805 ;
        RECT 0.000 3781.585 208.285 3782.425 ;
      LAYER met2 ;
        RECT 208.565 3781.865 210.965 3782.145 ;
      LAYER met2 ;
        RECT 0.000 3779.665 208.565 3781.585 ;
      LAYER met2 ;
        RECT 208.940 3781.150 209.200 3781.470 ;
      LAYER met2 ;
        RECT 0.000 3778.825 208.285 3779.665 ;
      LAYER met2 ;
        RECT 209.000 3779.385 209.140 3781.150 ;
        RECT 208.565 3779.105 210.965 3779.385 ;
      LAYER met2 ;
        RECT 0.000 3776.445 208.565 3778.825 ;
        RECT 0.000 3775.605 208.285 3776.445 ;
        RECT 0.000 3773.225 208.565 3775.605 ;
        RECT 0.000 3772.385 208.285 3773.225 ;
        RECT 0.000 3770.465 208.565 3772.385 ;
        RECT 0.000 3769.625 208.285 3770.465 ;
      LAYER met2 ;
        RECT 208.565 3769.905 210.965 3770.185 ;
      LAYER met2 ;
        RECT 0.000 3767.245 208.565 3769.625 ;
        RECT 0.000 3766.405 208.285 3767.245 ;
        RECT 0.000 3764.025 208.565 3766.405 ;
        RECT 0.000 3763.185 208.285 3764.025 ;
        RECT 0.000 3761.265 208.565 3763.185 ;
        RECT 0.000 3760.425 208.285 3761.265 ;
        RECT 0.000 3758.045 208.565 3760.425 ;
        RECT 0.000 3757.205 208.285 3758.045 ;
        RECT 0.000 3754.825 208.565 3757.205 ;
        RECT 0.000 3753.985 208.285 3754.825 ;
        RECT 0.000 3752.065 208.565 3753.985 ;
        RECT 0.000 3751.225 208.285 3752.065 ;
        RECT 0.000 3748.845 208.565 3751.225 ;
      LAYER met2 ;
        RECT 211.300 3749.250 211.440 3788.375 ;
        RECT 211.760 3781.470 211.900 3992.630 ;
        RECT 212.220 3960.650 212.360 4305.770 ;
        RECT 3367.360 4248.630 3367.500 4950.070 ;
        RECT 3367.820 4295.890 3367.960 4981.690 ;
        RECT 3368.220 4950.410 3368.480 4950.730 ;
        RECT 3367.760 4295.570 3368.020 4295.890 ;
        RECT 3367.300 4248.310 3367.560 4248.630 ;
        RECT 213.080 4004.870 213.340 4005.190 ;
        RECT 212.160 3960.330 212.420 3960.650 ;
        RECT 212.220 3960.050 212.360 3960.330 ;
        RECT 212.220 3959.910 212.820 3960.050 ;
        RECT 211.700 3781.150 211.960 3781.470 ;
        RECT 209.000 3749.110 211.440 3749.250 ;
      LAYER met2 ;
        RECT 0.000 3748.005 208.285 3748.845 ;
      LAYER met2 ;
        RECT 209.000 3748.570 209.140 3749.110 ;
        RECT 208.610 3748.565 209.140 3748.570 ;
        RECT 208.565 3748.285 210.965 3748.565 ;
      LAYER met2 ;
        RECT 0.000 3745.625 208.565 3748.005 ;
        RECT 0.000 3744.785 208.285 3745.625 ;
        RECT 0.000 3742.405 208.565 3744.785 ;
        RECT 0.000 3741.565 208.285 3742.405 ;
      LAYER met2 ;
        RECT 208.565 3741.845 210.965 3742.125 ;
        RECT 209.000 3741.690 209.140 3741.845 ;
        RECT 212.680 3741.690 212.820 3959.910 ;
        RECT 213.140 3945.690 213.280 4004.870 ;
        RECT 213.080 3945.370 213.340 3945.690 ;
        RECT 213.140 3933.070 213.280 3945.370 ;
        RECT 213.140 3932.930 213.740 3933.070 ;
        RECT 213.080 3781.150 213.340 3781.470 ;
      LAYER met2 ;
        RECT 0.000 3739.645 208.565 3741.565 ;
      LAYER met2 ;
        RECT 208.940 3741.370 209.200 3741.690 ;
        RECT 212.620 3741.370 212.880 3741.690 ;
      LAYER met2 ;
        RECT 0.000 3738.805 208.285 3739.645 ;
        RECT 0.000 3736.425 208.565 3738.805 ;
        RECT 0.000 3735.585 208.285 3736.425 ;
        RECT 0.000 3733.205 208.565 3735.585 ;
        RECT 0.000 3732.365 208.285 3733.205 ;
        RECT 0.000 3730.445 208.565 3732.365 ;
        RECT 0.000 3729.605 208.285 3730.445 ;
        RECT 0.000 3727.225 208.565 3729.605 ;
        RECT 0.000 3726.385 208.285 3727.225 ;
      LAYER met2 ;
        RECT 208.565 3726.665 210.965 3726.945 ;
      LAYER met2 ;
        RECT 0.000 3724.005 208.565 3726.385 ;
      LAYER met2 ;
        RECT 209.000 3724.350 209.140 3726.665 ;
        RECT 208.940 3724.030 209.200 3724.350 ;
        RECT 212.160 3724.030 212.420 3724.350 ;
      LAYER met2 ;
        RECT 0.000 3723.165 208.285 3724.005 ;
        RECT 0.000 3721.245 208.565 3723.165 ;
        RECT 0.000 3720.405 208.285 3721.245 ;
        RECT 0.000 3718.025 208.565 3720.405 ;
        RECT 0.000 3717.185 208.285 3718.025 ;
        RECT 0.000 3714.805 208.565 3717.185 ;
        RECT 0.000 3713.965 208.285 3714.805 ;
        RECT 0.000 3712.045 208.565 3713.965 ;
        RECT 0.000 3711.205 208.285 3712.045 ;
        RECT 0.000 3710.210 208.565 3711.205 ;
        RECT 0.000 3572.865 208.565 3573.915 ;
        RECT 0.000 3572.025 208.285 3572.865 ;
      LAYER met2 ;
        RECT 208.565 3572.305 210.965 3572.585 ;
      LAYER met2 ;
        RECT 0.000 3569.645 208.565 3572.025 ;
      LAYER met2 ;
        RECT 209.460 3571.090 209.600 3572.305 ;
        RECT 209.460 3570.950 211.440 3571.090 ;
      LAYER met2 ;
        RECT 0.000 3568.805 208.285 3569.645 ;
        RECT 0.000 3566.425 208.565 3568.805 ;
        RECT 0.000 3565.585 208.285 3566.425 ;
      LAYER met2 ;
        RECT 208.565 3565.865 210.965 3566.145 ;
      LAYER met2 ;
        RECT 0.000 3563.665 208.565 3565.585 ;
      LAYER met2 ;
        RECT 208.940 3565.250 209.200 3565.570 ;
      LAYER met2 ;
        RECT 0.000 3562.825 208.285 3563.665 ;
      LAYER met2 ;
        RECT 209.000 3563.385 209.140 3565.250 ;
        RECT 208.565 3563.105 210.965 3563.385 ;
      LAYER met2 ;
        RECT 0.000 3560.445 208.565 3562.825 ;
        RECT 0.000 3559.605 208.285 3560.445 ;
        RECT 0.000 3557.225 208.565 3559.605 ;
        RECT 0.000 3556.385 208.285 3557.225 ;
        RECT 0.000 3554.465 208.565 3556.385 ;
        RECT 0.000 3553.625 208.285 3554.465 ;
      LAYER met2 ;
        RECT 208.565 3553.905 210.965 3554.185 ;
      LAYER met2 ;
        RECT 0.000 3551.245 208.565 3553.625 ;
        RECT 0.000 3550.405 208.285 3551.245 ;
        RECT 0.000 3548.025 208.565 3550.405 ;
        RECT 0.000 3547.185 208.285 3548.025 ;
        RECT 0.000 3545.265 208.565 3547.185 ;
        RECT 0.000 3544.425 208.285 3545.265 ;
        RECT 0.000 3542.045 208.565 3544.425 ;
        RECT 0.000 3541.205 208.285 3542.045 ;
        RECT 0.000 3538.825 208.565 3541.205 ;
        RECT 0.000 3537.985 208.285 3538.825 ;
        RECT 0.000 3536.065 208.565 3537.985 ;
        RECT 0.000 3535.225 208.285 3536.065 ;
        RECT 0.000 3532.845 208.565 3535.225 ;
        RECT 0.000 3532.005 208.285 3532.845 ;
      LAYER met2 ;
        RECT 208.565 3532.495 210.965 3532.565 ;
        RECT 211.300 3532.495 211.440 3570.950 ;
        RECT 208.565 3532.355 211.440 3532.495 ;
        RECT 208.565 3532.285 210.965 3532.355 ;
      LAYER met2 ;
        RECT 0.000 3529.625 208.565 3532.005 ;
        RECT 0.000 3528.785 208.285 3529.625 ;
        RECT 0.000 3526.405 208.565 3528.785 ;
        RECT 0.000 3525.565 208.285 3526.405 ;
      LAYER met2 ;
        RECT 208.565 3525.845 210.965 3526.125 ;
      LAYER met2 ;
        RECT 0.000 3523.645 208.565 3525.565 ;
      LAYER met2 ;
        RECT 209.000 3524.090 209.140 3525.845 ;
        RECT 208.940 3523.770 209.200 3524.090 ;
      LAYER met2 ;
        RECT 0.000 3522.805 208.285 3523.645 ;
        RECT 0.000 3520.425 208.565 3522.805 ;
        RECT 0.000 3519.585 208.285 3520.425 ;
        RECT 0.000 3517.205 208.565 3519.585 ;
        RECT 0.000 3516.365 208.285 3517.205 ;
        RECT 0.000 3514.445 208.565 3516.365 ;
        RECT 0.000 3513.605 208.285 3514.445 ;
        RECT 0.000 3511.225 208.565 3513.605 ;
        RECT 0.000 3510.385 208.285 3511.225 ;
      LAYER met2 ;
        RECT 208.565 3510.665 210.965 3510.945 ;
      LAYER met2 ;
        RECT 0.000 3508.005 208.565 3510.385 ;
      LAYER met2 ;
        RECT 209.000 3508.450 209.140 3510.665 ;
        RECT 212.220 3508.450 212.360 3724.030 ;
        RECT 212.680 3524.090 212.820 3741.370 ;
        RECT 213.140 3565.570 213.280 3781.150 ;
        RECT 213.600 3724.350 213.740 3932.930 ;
        RECT 3367.360 3806.630 3367.500 4248.310 ;
        RECT 3367.820 3864.090 3367.960 4295.570 ;
        RECT 3368.280 4280.590 3368.420 4950.410 ;
        RECT 3368.220 4280.270 3368.480 4280.590 ;
        RECT 3367.760 3863.770 3368.020 3864.090 ;
        RECT 3367.300 3806.310 3367.560 3806.630 ;
        RECT 213.540 3724.030 213.800 3724.350 ;
        RECT 3367.820 3642.070 3367.960 3863.770 ;
        RECT 3368.280 3848.450 3368.420 4280.270 ;
        RECT 3368.220 3848.130 3368.480 3848.450 ;
        RECT 3369.600 3848.130 3369.860 3848.450 ;
        RECT 3367.760 3641.750 3368.020 3642.070 ;
        RECT 213.080 3565.250 213.340 3565.570 ;
        RECT 212.620 3523.770 212.880 3524.090 ;
        RECT 208.940 3508.130 209.200 3508.450 ;
        RECT 212.160 3508.130 212.420 3508.450 ;
      LAYER met2 ;
        RECT 0.000 3507.165 208.285 3508.005 ;
        RECT 0.000 3505.245 208.565 3507.165 ;
        RECT 0.000 3504.405 208.285 3505.245 ;
        RECT 0.000 3502.025 208.565 3504.405 ;
        RECT 0.000 3501.185 208.285 3502.025 ;
        RECT 0.000 3498.805 208.565 3501.185 ;
        RECT 0.000 3497.965 208.285 3498.805 ;
        RECT 0.000 3496.045 208.565 3497.965 ;
        RECT 0.000 3495.205 208.285 3496.045 ;
        RECT 0.000 3494.210 208.565 3495.205 ;
        RECT 0.000 3355.865 208.565 3356.915 ;
        RECT 0.000 3355.025 208.285 3355.865 ;
      LAYER met2 ;
        RECT 208.565 3355.305 210.965 3355.585 ;
      LAYER met2 ;
        RECT 0.000 3352.645 208.565 3355.025 ;
      LAYER met2 ;
        RECT 209.000 3353.470 209.140 3355.305 ;
        RECT 209.000 3353.330 211.440 3353.470 ;
      LAYER met2 ;
        RECT 0.000 3351.805 208.285 3352.645 ;
        RECT 0.000 3349.425 208.565 3351.805 ;
        RECT 0.000 3348.585 208.285 3349.425 ;
      LAYER met2 ;
        RECT 208.565 3348.865 210.965 3349.145 ;
      LAYER met2 ;
        RECT 0.000 3346.665 208.565 3348.585 ;
        RECT 0.000 3345.825 208.285 3346.665 ;
      LAYER met2 ;
        RECT 208.565 3346.105 210.965 3346.385 ;
      LAYER met2 ;
        RECT 0.000 3343.445 208.565 3345.825 ;
      LAYER met2 ;
        RECT 209.000 3343.890 209.140 3346.105 ;
        RECT 208.940 3343.570 209.200 3343.890 ;
      LAYER met2 ;
        RECT 0.000 3342.605 208.285 3343.445 ;
        RECT 0.000 3340.225 208.565 3342.605 ;
        RECT 0.000 3339.385 208.285 3340.225 ;
        RECT 0.000 3337.465 208.565 3339.385 ;
        RECT 0.000 3336.625 208.285 3337.465 ;
      LAYER met2 ;
        RECT 208.565 3336.905 210.965 3337.185 ;
      LAYER met2 ;
        RECT 0.000 3334.245 208.565 3336.625 ;
        RECT 0.000 3333.405 208.285 3334.245 ;
        RECT 0.000 3331.025 208.565 3333.405 ;
        RECT 0.000 3330.185 208.285 3331.025 ;
        RECT 0.000 3328.265 208.565 3330.185 ;
        RECT 0.000 3327.425 208.285 3328.265 ;
        RECT 0.000 3325.045 208.565 3327.425 ;
        RECT 0.000 3324.205 208.285 3325.045 ;
        RECT 0.000 3321.825 208.565 3324.205 ;
        RECT 0.000 3320.985 208.285 3321.825 ;
        RECT 0.000 3319.065 208.565 3320.985 ;
        RECT 0.000 3318.225 208.285 3319.065 ;
        RECT 0.000 3315.845 208.565 3318.225 ;
      LAYER met2 ;
        RECT 211.300 3318.130 211.440 3353.330 ;
        RECT 209.460 3317.990 211.440 3318.130 ;
      LAYER met2 ;
        RECT 0.000 3315.005 208.285 3315.845 ;
      LAYER met2 ;
        RECT 209.460 3315.565 209.600 3317.990 ;
        RECT 208.565 3315.285 210.965 3315.565 ;
        RECT 208.610 3315.270 209.600 3315.285 ;
      LAYER met2 ;
        RECT 0.000 3312.625 208.565 3315.005 ;
        RECT 0.000 3311.785 208.285 3312.625 ;
        RECT 0.000 3309.405 208.565 3311.785 ;
        RECT 0.000 3308.565 208.285 3309.405 ;
      LAYER met2 ;
        RECT 208.565 3308.845 210.965 3309.125 ;
      LAYER met2 ;
        RECT 0.000 3306.645 208.565 3308.565 ;
      LAYER met2 ;
        RECT 209.000 3306.830 209.140 3308.845 ;
      LAYER met2 ;
        RECT 0.000 3305.805 208.285 3306.645 ;
      LAYER met2 ;
        RECT 208.940 3306.510 209.200 3306.830 ;
      LAYER met2 ;
        RECT 0.000 3303.425 208.565 3305.805 ;
        RECT 0.000 3302.585 208.285 3303.425 ;
        RECT 0.000 3300.205 208.565 3302.585 ;
        RECT 0.000 3299.365 208.285 3300.205 ;
        RECT 0.000 3297.445 208.565 3299.365 ;
        RECT 0.000 3296.605 208.285 3297.445 ;
      LAYER met2 ;
        RECT 212.220 3296.630 212.360 3508.130 ;
        RECT 212.680 3306.830 212.820 3523.770 ;
        RECT 213.140 3343.890 213.280 3565.250 ;
        RECT 3367.820 3415.630 3367.960 3641.750 ;
        RECT 3369.660 3626.430 3369.800 3848.130 ;
        RECT 3370.060 3806.310 3370.320 3806.630 ;
        RECT 3369.600 3626.110 3369.860 3626.430 ;
        RECT 3368.220 3589.050 3368.480 3589.370 ;
        RECT 3367.760 3415.310 3368.020 3415.630 ;
        RECT 3367.760 3402.050 3368.020 3402.370 ;
        RECT 213.080 3343.570 213.340 3343.890 ;
        RECT 212.620 3306.510 212.880 3306.830 ;
      LAYER met2 ;
        RECT 0.000 3294.225 208.565 3296.605 ;
      LAYER met2 ;
        RECT 208.940 3296.310 209.200 3296.630 ;
        RECT 212.160 3296.310 212.420 3296.630 ;
      LAYER met2 ;
        RECT 0.000 3293.385 208.285 3294.225 ;
      LAYER met2 ;
        RECT 209.000 3293.945 209.140 3296.310 ;
        RECT 208.565 3293.665 210.965 3293.945 ;
      LAYER met2 ;
        RECT 0.000 3291.005 208.565 3293.385 ;
        RECT 0.000 3290.165 208.285 3291.005 ;
        RECT 0.000 3288.245 208.565 3290.165 ;
        RECT 0.000 3287.405 208.285 3288.245 ;
        RECT 0.000 3285.025 208.565 3287.405 ;
        RECT 0.000 3284.185 208.285 3285.025 ;
        RECT 0.000 3281.805 208.565 3284.185 ;
        RECT 0.000 3280.965 208.285 3281.805 ;
        RECT 0.000 3279.045 208.565 3280.965 ;
        RECT 0.000 3278.205 208.285 3279.045 ;
        RECT 0.000 3277.210 208.565 3278.205 ;
        RECT 0.000 3139.865 208.565 3140.915 ;
        RECT 0.000 3139.025 208.285 3139.865 ;
      LAYER met2 ;
        RECT 208.565 3139.515 210.965 3139.585 ;
        RECT 208.565 3139.375 211.440 3139.515 ;
        RECT 208.565 3139.305 210.965 3139.375 ;
      LAYER met2 ;
        RECT 0.000 3136.645 208.565 3139.025 ;
        RECT 0.000 3135.805 208.285 3136.645 ;
        RECT 0.000 3133.425 208.565 3135.805 ;
        RECT 0.000 3132.585 208.285 3133.425 ;
      LAYER met2 ;
        RECT 208.565 3132.865 210.965 3133.145 ;
      LAYER met2 ;
        RECT 0.000 3130.665 208.565 3132.585 ;
        RECT 0.000 3129.825 208.285 3130.665 ;
      LAYER met2 ;
        RECT 208.610 3130.385 209.140 3130.450 ;
        RECT 208.565 3130.105 210.965 3130.385 ;
      LAYER met2 ;
        RECT 0.000 3127.445 208.565 3129.825 ;
      LAYER met2 ;
        RECT 209.000 3127.650 209.140 3130.105 ;
      LAYER met2 ;
        RECT 0.000 3126.605 208.285 3127.445 ;
      LAYER met2 ;
        RECT 208.940 3127.330 209.200 3127.650 ;
      LAYER met2 ;
        RECT 0.000 3124.225 208.565 3126.605 ;
        RECT 0.000 3123.385 208.285 3124.225 ;
        RECT 0.000 3121.465 208.565 3123.385 ;
        RECT 0.000 3120.625 208.285 3121.465 ;
      LAYER met2 ;
        RECT 208.565 3120.905 210.965 3121.185 ;
      LAYER met2 ;
        RECT 0.000 3118.245 208.565 3120.625 ;
        RECT 0.000 3117.405 208.285 3118.245 ;
        RECT 0.000 3115.025 208.565 3117.405 ;
        RECT 0.000 3114.185 208.285 3115.025 ;
        RECT 0.000 3112.265 208.565 3114.185 ;
        RECT 0.000 3111.425 208.285 3112.265 ;
        RECT 0.000 3109.045 208.565 3111.425 ;
        RECT 0.000 3108.205 208.285 3109.045 ;
        RECT 0.000 3105.825 208.565 3108.205 ;
        RECT 0.000 3104.985 208.285 3105.825 ;
        RECT 0.000 3103.065 208.565 3104.985 ;
        RECT 0.000 3102.225 208.285 3103.065 ;
        RECT 0.000 3099.845 208.565 3102.225 ;
      LAYER met2 ;
        RECT 211.300 3101.890 211.440 3139.375 ;
        RECT 209.460 3101.750 211.440 3101.890 ;
      LAYER met2 ;
        RECT 0.000 3099.005 208.285 3099.845 ;
      LAYER met2 ;
        RECT 209.460 3099.565 209.600 3101.750 ;
        RECT 208.565 3099.285 210.965 3099.565 ;
      LAYER met2 ;
        RECT 0.000 3096.625 208.565 3099.005 ;
        RECT 0.000 3095.785 208.285 3096.625 ;
        RECT 0.000 3093.405 208.565 3095.785 ;
        RECT 0.000 3092.565 208.285 3093.405 ;
      LAYER met2 ;
        RECT 208.565 3092.845 210.965 3093.125 ;
      LAYER met2 ;
        RECT 0.000 3090.645 208.565 3092.565 ;
      LAYER met2 ;
        RECT 209.000 3090.930 209.140 3092.845 ;
        RECT 212.680 3090.930 212.820 3306.510 ;
        RECT 213.140 3127.650 213.280 3343.570 ;
        RECT 213.540 3296.310 213.800 3296.630 ;
        RECT 213.080 3127.330 213.340 3127.650 ;
      LAYER met2 ;
        RECT 0.000 3089.805 208.285 3090.645 ;
      LAYER met2 ;
        RECT 208.940 3090.610 209.200 3090.930 ;
        RECT 212.620 3090.610 212.880 3090.930 ;
      LAYER met2 ;
        RECT 0.000 3087.425 208.565 3089.805 ;
        RECT 0.000 3086.585 208.285 3087.425 ;
        RECT 0.000 3084.205 208.565 3086.585 ;
        RECT 0.000 3083.365 208.285 3084.205 ;
        RECT 0.000 3081.445 208.565 3083.365 ;
        RECT 0.000 3080.605 208.285 3081.445 ;
        RECT 0.000 3078.225 208.565 3080.605 ;
        RECT 0.000 3077.385 208.285 3078.225 ;
      LAYER met2 ;
        RECT 208.565 3077.665 210.965 3077.945 ;
      LAYER met2 ;
        RECT 0.000 3075.005 208.565 3077.385 ;
      LAYER met2 ;
        RECT 209.000 3075.290 209.140 3077.665 ;
      LAYER met2 ;
        RECT 0.000 3074.165 208.285 3075.005 ;
      LAYER met2 ;
        RECT 208.940 3074.970 209.200 3075.290 ;
      LAYER met2 ;
        RECT 0.000 3072.245 208.565 3074.165 ;
      LAYER met2 ;
        RECT 211.240 3073.270 211.500 3073.590 ;
      LAYER met2 ;
        RECT 0.000 3071.405 208.285 3072.245 ;
        RECT 0.000 3069.025 208.565 3071.405 ;
        RECT 0.000 3068.185 208.285 3069.025 ;
        RECT 0.000 3065.805 208.565 3068.185 ;
        RECT 0.000 3064.965 208.285 3065.805 ;
        RECT 0.000 3063.045 208.565 3064.965 ;
        RECT 0.000 3062.205 208.285 3063.045 ;
        RECT 0.000 3061.210 208.565 3062.205 ;
        RECT 0.000 2923.865 208.565 2924.915 ;
      LAYER met2 ;
        RECT 211.300 2924.410 211.440 3073.270 ;
        RECT 211.300 2924.270 211.900 2924.410 ;
      LAYER met2 ;
        RECT 0.000 2923.025 208.285 2923.865 ;
      LAYER met2 ;
        RECT 208.565 2923.515 210.965 2923.585 ;
        RECT 208.565 2923.375 211.440 2923.515 ;
        RECT 208.565 2923.305 210.965 2923.375 ;
      LAYER met2 ;
        RECT 0.000 2920.645 208.565 2923.025 ;
        RECT 0.000 2919.805 208.285 2920.645 ;
        RECT 0.000 2917.425 208.565 2919.805 ;
        RECT 0.000 2916.585 208.285 2917.425 ;
      LAYER met2 ;
        RECT 208.565 2916.865 210.965 2917.145 ;
      LAYER met2 ;
        RECT 0.000 2914.665 208.565 2916.585 ;
      LAYER met2 ;
        RECT 208.940 2916.190 209.200 2916.510 ;
      LAYER met2 ;
        RECT 0.000 2913.825 208.285 2914.665 ;
      LAYER met2 ;
        RECT 209.000 2914.385 209.140 2916.190 ;
        RECT 208.565 2914.105 210.965 2914.385 ;
        RECT 208.610 2914.070 209.140 2914.105 ;
      LAYER met2 ;
        RECT 0.000 2911.445 208.565 2913.825 ;
        RECT 0.000 2910.605 208.285 2911.445 ;
        RECT 0.000 2908.225 208.565 2910.605 ;
        RECT 0.000 2907.385 208.285 2908.225 ;
        RECT 0.000 2905.465 208.565 2907.385 ;
        RECT 0.000 2904.625 208.285 2905.465 ;
      LAYER met2 ;
        RECT 208.565 2904.905 210.965 2905.185 ;
      LAYER met2 ;
        RECT 0.000 2902.245 208.565 2904.625 ;
        RECT 0.000 2901.405 208.285 2902.245 ;
        RECT 0.000 2899.025 208.565 2901.405 ;
        RECT 0.000 2898.185 208.285 2899.025 ;
        RECT 0.000 2896.265 208.565 2898.185 ;
        RECT 0.000 2895.425 208.285 2896.265 ;
        RECT 0.000 2893.045 208.565 2895.425 ;
        RECT 0.000 2892.205 208.285 2893.045 ;
        RECT 0.000 2889.825 208.565 2892.205 ;
        RECT 0.000 2888.985 208.285 2889.825 ;
        RECT 0.000 2887.065 208.565 2888.985 ;
        RECT 0.000 2886.225 208.285 2887.065 ;
        RECT 0.000 2883.845 208.565 2886.225 ;
      LAYER met2 ;
        RECT 211.300 2884.290 211.440 2923.375 ;
        RECT 209.460 2884.150 211.440 2884.290 ;
      LAYER met2 ;
        RECT 0.000 2883.005 208.285 2883.845 ;
      LAYER met2 ;
        RECT 209.460 2883.610 209.600 2884.150 ;
        RECT 208.610 2883.565 209.600 2883.610 ;
        RECT 208.565 2883.285 210.965 2883.565 ;
      LAYER met2 ;
        RECT 0.000 2880.625 208.565 2883.005 ;
        RECT 0.000 2879.785 208.285 2880.625 ;
        RECT 0.000 2877.405 208.565 2879.785 ;
      LAYER met2 ;
        RECT 208.940 2879.470 209.200 2879.790 ;
      LAYER met2 ;
        RECT 0.000 2876.565 208.285 2877.405 ;
      LAYER met2 ;
        RECT 209.000 2877.125 209.140 2879.470 ;
        RECT 208.565 2876.845 210.965 2877.125 ;
      LAYER met2 ;
        RECT 0.000 2874.645 208.565 2876.565 ;
        RECT 0.000 2873.805 208.285 2874.645 ;
        RECT 0.000 2871.425 208.565 2873.805 ;
        RECT 0.000 2870.585 208.285 2871.425 ;
        RECT 0.000 2868.205 208.565 2870.585 ;
      LAYER met2 ;
        RECT 211.760 2870.470 211.900 2924.270 ;
        RECT 212.680 2879.790 212.820 3090.610 ;
        RECT 213.140 2916.510 213.280 3127.330 ;
        RECT 213.600 3075.290 213.740 3296.310 ;
        RECT 3367.820 3181.710 3367.960 3402.050 ;
        RECT 3368.280 3368.370 3368.420 3589.050 ;
        RECT 3368.680 3415.310 3368.940 3415.630 ;
        RECT 3368.220 3368.050 3368.480 3368.370 ;
        RECT 3368.740 3215.470 3368.880 3415.310 ;
        RECT 3369.660 3402.370 3369.800 3626.110 ;
        RECT 3370.120 3589.370 3370.260 3806.310 ;
        RECT 3370.060 3589.050 3370.320 3589.370 ;
        RECT 3369.600 3402.050 3369.860 3402.370 ;
        RECT 3370.060 3368.050 3370.320 3368.370 ;
        RECT 3368.280 3215.330 3368.880 3215.470 ;
        RECT 3368.280 3194.630 3368.420 3215.330 ;
        RECT 3368.220 3194.310 3368.480 3194.630 ;
        RECT 3367.760 3181.390 3368.020 3181.710 ;
        RECT 3367.300 3147.050 3367.560 3147.370 ;
        RECT 213.540 3074.970 213.800 3075.290 ;
        RECT 3367.360 2920.930 3367.500 3147.050 ;
        RECT 3367.820 2959.690 3367.960 3181.390 ;
        RECT 3368.280 2976.010 3368.420 3194.310 ;
        RECT 3370.120 3147.370 3370.260 3368.050 ;
        RECT 3370.060 3147.050 3370.320 3147.370 ;
        RECT 3368.220 2975.690 3368.480 2976.010 ;
        RECT 3367.760 2959.370 3368.020 2959.690 ;
        RECT 3367.300 2920.610 3367.560 2920.930 ;
        RECT 213.080 2916.190 213.340 2916.510 ;
        RECT 212.620 2879.470 212.880 2879.790 ;
        RECT 211.760 2870.330 212.360 2870.470 ;
      LAYER met2 ;
        RECT 0.000 2867.365 208.285 2868.205 ;
        RECT 0.000 2865.445 208.565 2867.365 ;
        RECT 0.000 2864.605 208.285 2865.445 ;
        RECT 0.000 2862.225 208.565 2864.605 ;
        RECT 0.000 2861.385 208.285 2862.225 ;
      LAYER met2 ;
        RECT 208.565 2861.665 210.965 2861.945 ;
      LAYER met2 ;
        RECT 0.000 2859.005 208.565 2861.385 ;
      LAYER met2 ;
        RECT 209.000 2859.390 209.140 2861.665 ;
        RECT 212.220 2859.390 212.360 2870.330 ;
        RECT 208.940 2859.070 209.200 2859.390 ;
        RECT 212.160 2859.070 212.420 2859.390 ;
      LAYER met2 ;
        RECT 0.000 2858.165 208.285 2859.005 ;
        RECT 0.000 2856.245 208.565 2858.165 ;
        RECT 0.000 2855.405 208.285 2856.245 ;
        RECT 0.000 2853.025 208.565 2855.405 ;
        RECT 0.000 2852.185 208.285 2853.025 ;
        RECT 0.000 2849.805 208.565 2852.185 ;
        RECT 0.000 2848.965 208.285 2849.805 ;
        RECT 0.000 2847.045 208.565 2848.965 ;
        RECT 0.000 2846.205 208.285 2847.045 ;
        RECT 0.000 2845.210 208.565 2846.205 ;
        RECT 0.000 2707.865 208.565 2708.915 ;
        RECT 0.000 2707.025 208.285 2707.865 ;
      LAYER met2 ;
        RECT 208.565 2707.305 210.965 2707.585 ;
      LAYER met2 ;
        RECT 0.000 2704.645 208.565 2707.025 ;
      LAYER met2 ;
        RECT 209.000 2706.810 209.140 2707.305 ;
        RECT 209.000 2706.670 211.440 2706.810 ;
      LAYER met2 ;
        RECT 0.000 2703.805 208.285 2704.645 ;
        RECT 0.000 2701.425 208.565 2703.805 ;
        RECT 0.000 2700.585 208.285 2701.425 ;
      LAYER met2 ;
        RECT 208.565 2700.865 210.965 2701.145 ;
      LAYER met2 ;
        RECT 0.000 2698.665 208.565 2700.585 ;
      LAYER met2 ;
        RECT 208.940 2700.290 209.200 2700.610 ;
      LAYER met2 ;
        RECT 0.000 2697.825 208.285 2698.665 ;
      LAYER met2 ;
        RECT 209.000 2698.385 209.140 2700.290 ;
        RECT 208.565 2698.105 210.965 2698.385 ;
      LAYER met2 ;
        RECT 0.000 2695.445 208.565 2697.825 ;
        RECT 0.000 2694.605 208.285 2695.445 ;
        RECT 0.000 2692.225 208.565 2694.605 ;
        RECT 0.000 2691.385 208.285 2692.225 ;
        RECT 0.000 2689.465 208.565 2691.385 ;
        RECT 0.000 2688.625 208.285 2689.465 ;
      LAYER met2 ;
        RECT 208.565 2688.905 210.965 2689.185 ;
      LAYER met2 ;
        RECT 0.000 2686.245 208.565 2688.625 ;
        RECT 0.000 2685.405 208.285 2686.245 ;
        RECT 0.000 2683.025 208.565 2685.405 ;
        RECT 0.000 2682.185 208.285 2683.025 ;
        RECT 0.000 2680.265 208.565 2682.185 ;
        RECT 0.000 2679.425 208.285 2680.265 ;
        RECT 0.000 2677.045 208.565 2679.425 ;
        RECT 0.000 2676.205 208.285 2677.045 ;
        RECT 0.000 2673.825 208.565 2676.205 ;
        RECT 0.000 2672.985 208.285 2673.825 ;
        RECT 0.000 2671.065 208.565 2672.985 ;
        RECT 0.000 2670.225 208.285 2671.065 ;
        RECT 0.000 2667.845 208.565 2670.225 ;
      LAYER met2 ;
        RECT 211.300 2668.050 211.440 2706.670 ;
        RECT 209.460 2667.910 211.440 2668.050 ;
      LAYER met2 ;
        RECT 0.000 2667.005 208.285 2667.845 ;
      LAYER met2 ;
        RECT 209.460 2667.565 209.600 2667.910 ;
        RECT 208.565 2667.285 210.965 2667.565 ;
        RECT 208.610 2667.230 209.600 2667.285 ;
      LAYER met2 ;
        RECT 0.000 2664.625 208.565 2667.005 ;
        RECT 0.000 2663.785 208.285 2664.625 ;
        RECT 0.000 2661.405 208.565 2663.785 ;
        RECT 0.000 2660.565 208.285 2661.405 ;
      LAYER met2 ;
        RECT 208.565 2660.845 210.965 2661.125 ;
      LAYER met2 ;
        RECT 0.000 2658.645 208.565 2660.565 ;
      LAYER met2 ;
        RECT 209.000 2659.130 209.140 2660.845 ;
        RECT 208.940 2658.810 209.200 2659.130 ;
      LAYER met2 ;
        RECT 0.000 2657.805 208.285 2658.645 ;
        RECT 0.000 2655.425 208.565 2657.805 ;
        RECT 0.000 2654.585 208.285 2655.425 ;
        RECT 0.000 2652.205 208.565 2654.585 ;
        RECT 0.000 2651.365 208.285 2652.205 ;
        RECT 0.000 2649.445 208.565 2651.365 ;
        RECT 0.000 2648.605 208.285 2649.445 ;
        RECT 0.000 2646.225 208.565 2648.605 ;
        RECT 0.000 2645.385 208.285 2646.225 ;
      LAYER met2 ;
        RECT 208.565 2645.665 210.965 2645.945 ;
      LAYER met2 ;
        RECT 0.000 2643.005 208.565 2645.385 ;
      LAYER met2 ;
        RECT 209.000 2643.490 209.140 2645.665 ;
        RECT 212.220 2643.490 212.360 2859.070 ;
        RECT 212.680 2659.130 212.820 2879.470 ;
        RECT 213.140 2700.610 213.280 2916.190 ;
        RECT 3367.820 2741.410 3367.960 2959.370 ;
        RECT 3368.280 2757.050 3368.420 2975.690 ;
        RECT 3369.600 2920.610 3369.860 2920.930 ;
        RECT 3368.220 2756.730 3368.480 2757.050 ;
        RECT 3367.760 2741.090 3368.020 2741.410 ;
        RECT 3369.660 2704.690 3369.800 2920.610 ;
        RECT 3369.600 2704.370 3369.860 2704.690 ;
        RECT 213.080 2700.290 213.340 2700.610 ;
        RECT 212.620 2658.810 212.880 2659.130 ;
        RECT 208.940 2643.170 209.200 2643.490 ;
        RECT 212.160 2643.170 212.420 2643.490 ;
      LAYER met2 ;
        RECT 0.000 2642.165 208.285 2643.005 ;
        RECT 0.000 2640.245 208.565 2642.165 ;
        RECT 0.000 2639.405 208.285 2640.245 ;
        RECT 0.000 2637.025 208.565 2639.405 ;
        RECT 0.000 2636.185 208.285 2637.025 ;
        RECT 0.000 2633.805 208.565 2636.185 ;
        RECT 0.000 2632.965 208.285 2633.805 ;
        RECT 0.000 2631.045 208.565 2632.965 ;
        RECT 0.000 2630.205 208.285 2631.045 ;
        RECT 0.000 2629.210 208.565 2630.205 ;
        RECT 4.925 2467.390 200.000 2491.290 ;
        RECT 4.925 2441.395 197.965 2467.390 ;
        RECT 198.080 2442.895 200.000 2444.895 ;
        RECT 4.925 2417.495 200.000 2441.395 ;
        RECT 4.925 2417.265 197.965 2417.495 ;
        RECT 0.035 2282.200 151.405 2291.935 ;
        RECT 153.765 2281.000 158.415 2292.140 ;
        RECT 160.165 2282.200 174.575 2291.935 ;
        RECT 0.035 2280.700 197.965 2281.000 ;
        RECT 0.035 2260.095 198.000 2280.700 ;
        RECT 0.035 2259.535 197.965 2260.095 ;
        RECT 0.035 2226.925 198.000 2259.535 ;
        RECT 0.035 2226.495 197.965 2226.925 ;
        RECT 0.035 2206.500 198.000 2226.495 ;
        RECT 0.035 2206.000 197.965 2206.500 ;
        RECT 153.800 2195.025 158.450 2206.000 ;
        RECT 0.000 2068.865 208.565 2069.915 ;
        RECT 0.000 2068.025 208.285 2068.865 ;
      LAYER met2 ;
        RECT 208.565 2068.515 210.965 2068.585 ;
        RECT 208.565 2068.375 211.440 2068.515 ;
        RECT 208.565 2068.305 210.965 2068.375 ;
      LAYER met2 ;
        RECT 0.000 2065.645 208.565 2068.025 ;
        RECT 0.000 2064.805 208.285 2065.645 ;
        RECT 0.000 2062.425 208.565 2064.805 ;
        RECT 0.000 2061.585 208.285 2062.425 ;
      LAYER met2 ;
        RECT 208.565 2061.865 210.965 2062.145 ;
      LAYER met2 ;
        RECT 0.000 2059.665 208.565 2061.585 ;
        RECT 0.000 2058.825 208.285 2059.665 ;
      LAYER met2 ;
        RECT 208.610 2059.385 209.140 2059.450 ;
        RECT 208.565 2059.105 210.965 2059.385 ;
      LAYER met2 ;
        RECT 0.000 2056.445 208.565 2058.825 ;
      LAYER met2 ;
        RECT 209.000 2056.650 209.140 2059.105 ;
      LAYER met2 ;
        RECT 0.000 2055.605 208.285 2056.445 ;
      LAYER met2 ;
        RECT 208.940 2056.330 209.200 2056.650 ;
      LAYER met2 ;
        RECT 0.000 2053.225 208.565 2055.605 ;
        RECT 0.000 2052.385 208.285 2053.225 ;
        RECT 0.000 2050.465 208.565 2052.385 ;
        RECT 0.000 2049.625 208.285 2050.465 ;
      LAYER met2 ;
        RECT 208.565 2049.905 210.965 2050.185 ;
      LAYER met2 ;
        RECT 0.000 2047.245 208.565 2049.625 ;
        RECT 0.000 2046.405 208.285 2047.245 ;
        RECT 0.000 2044.025 208.565 2046.405 ;
        RECT 0.000 2043.185 208.285 2044.025 ;
        RECT 0.000 2041.265 208.565 2043.185 ;
        RECT 0.000 2040.425 208.285 2041.265 ;
        RECT 0.000 2038.045 208.565 2040.425 ;
        RECT 0.000 2037.205 208.285 2038.045 ;
        RECT 0.000 2034.825 208.565 2037.205 ;
        RECT 0.000 2033.985 208.285 2034.825 ;
        RECT 0.000 2032.065 208.565 2033.985 ;
        RECT 0.000 2031.225 208.285 2032.065 ;
        RECT 0.000 2028.845 208.565 2031.225 ;
      LAYER met2 ;
        RECT 211.300 2028.850 211.440 2068.375 ;
      LAYER met2 ;
        RECT 0.000 2028.005 208.285 2028.845 ;
      LAYER met2 ;
        RECT 209.460 2028.710 211.440 2028.850 ;
        RECT 209.460 2028.565 209.600 2028.710 ;
        RECT 208.565 2028.285 210.965 2028.565 ;
      LAYER met2 ;
        RECT 0.000 2025.625 208.565 2028.005 ;
        RECT 0.000 2024.785 208.285 2025.625 ;
        RECT 0.000 2022.405 208.565 2024.785 ;
      LAYER met2 ;
        RECT 208.940 2024.370 209.200 2024.690 ;
      LAYER met2 ;
        RECT 0.000 2021.565 208.285 2022.405 ;
      LAYER met2 ;
        RECT 209.000 2022.125 209.140 2024.370 ;
        RECT 208.565 2021.845 210.965 2022.125 ;
      LAYER met2 ;
        RECT 0.000 2019.645 208.565 2021.565 ;
        RECT 0.000 2018.805 208.285 2019.645 ;
        RECT 0.000 2016.425 208.565 2018.805 ;
        RECT 0.000 2015.585 208.285 2016.425 ;
        RECT 0.000 2013.205 208.565 2015.585 ;
        RECT 0.000 2012.365 208.285 2013.205 ;
        RECT 0.000 2010.445 208.565 2012.365 ;
        RECT 0.000 2009.605 208.285 2010.445 ;
      LAYER met2 ;
        RECT 212.220 2009.730 212.360 2643.170 ;
        RECT 213.140 2097.670 213.280 2700.290 ;
        RECT 213.540 2658.810 213.800 2659.130 ;
        RECT 212.680 2097.530 213.280 2097.670 ;
        RECT 212.680 2056.650 212.820 2097.530 ;
        RECT 212.620 2056.330 212.880 2056.650 ;
      LAYER met2 ;
        RECT 0.000 2007.225 208.565 2009.605 ;
      LAYER met2 ;
        RECT 208.940 2009.410 209.200 2009.730 ;
        RECT 212.160 2009.410 212.420 2009.730 ;
      LAYER met2 ;
        RECT 0.000 2006.385 208.285 2007.225 ;
      LAYER met2 ;
        RECT 209.000 2006.945 209.140 2009.410 ;
        RECT 208.565 2006.665 210.965 2006.945 ;
      LAYER met2 ;
        RECT 0.000 2004.005 208.565 2006.385 ;
        RECT 0.000 2003.165 208.285 2004.005 ;
        RECT 0.000 2001.245 208.565 2003.165 ;
        RECT 0.000 2000.405 208.285 2001.245 ;
        RECT 0.000 1998.025 208.565 2000.405 ;
        RECT 0.000 1997.185 208.285 1998.025 ;
        RECT 0.000 1994.805 208.565 1997.185 ;
        RECT 0.000 1993.965 208.285 1994.805 ;
        RECT 0.000 1992.045 208.565 1993.965 ;
        RECT 0.000 1991.205 208.285 1992.045 ;
        RECT 0.000 1990.210 208.565 1991.205 ;
        RECT 0.000 1852.865 208.565 1853.915 ;
        RECT 0.000 1852.025 208.285 1852.865 ;
      LAYER met2 ;
        RECT 208.565 1852.515 210.965 1852.585 ;
        RECT 208.565 1852.375 211.440 1852.515 ;
        RECT 208.565 1852.305 210.965 1852.375 ;
      LAYER met2 ;
        RECT 0.000 1849.645 208.565 1852.025 ;
        RECT 0.000 1848.805 208.285 1849.645 ;
        RECT 0.000 1846.425 208.565 1848.805 ;
        RECT 0.000 1845.585 208.285 1846.425 ;
      LAYER met2 ;
        RECT 208.565 1845.865 210.965 1846.145 ;
      LAYER met2 ;
        RECT 0.000 1843.665 208.565 1845.585 ;
      LAYER met2 ;
        RECT 208.940 1845.190 209.200 1845.510 ;
      LAYER met2 ;
        RECT 0.000 1842.825 208.285 1843.665 ;
      LAYER met2 ;
        RECT 209.000 1843.385 209.140 1845.190 ;
        RECT 208.565 1843.105 210.965 1843.385 ;
        RECT 208.610 1843.070 209.140 1843.105 ;
      LAYER met2 ;
        RECT 0.000 1840.445 208.565 1842.825 ;
        RECT 0.000 1839.605 208.285 1840.445 ;
        RECT 0.000 1837.225 208.565 1839.605 ;
        RECT 0.000 1836.385 208.285 1837.225 ;
        RECT 0.000 1834.465 208.565 1836.385 ;
        RECT 0.000 1833.625 208.285 1834.465 ;
      LAYER met2 ;
        RECT 208.565 1833.905 210.965 1834.185 ;
      LAYER met2 ;
        RECT 0.000 1831.245 208.565 1833.625 ;
        RECT 0.000 1830.405 208.285 1831.245 ;
        RECT 0.000 1828.025 208.565 1830.405 ;
        RECT 0.000 1827.185 208.285 1828.025 ;
        RECT 0.000 1825.265 208.565 1827.185 ;
        RECT 0.000 1824.425 208.285 1825.265 ;
        RECT 0.000 1822.045 208.565 1824.425 ;
        RECT 0.000 1821.205 208.285 1822.045 ;
        RECT 0.000 1818.825 208.565 1821.205 ;
        RECT 0.000 1817.985 208.285 1818.825 ;
        RECT 0.000 1816.065 208.565 1817.985 ;
        RECT 0.000 1815.225 208.285 1816.065 ;
        RECT 0.000 1812.845 208.565 1815.225 ;
      LAYER met2 ;
        RECT 211.300 1813.290 211.440 1852.375 ;
        RECT 209.000 1813.150 211.440 1813.290 ;
      LAYER met2 ;
        RECT 0.000 1812.005 208.285 1812.845 ;
      LAYER met2 ;
        RECT 209.000 1812.610 209.140 1813.150 ;
        RECT 208.610 1812.565 209.140 1812.610 ;
        RECT 208.565 1812.285 210.965 1812.565 ;
      LAYER met2 ;
        RECT 0.000 1809.625 208.565 1812.005 ;
        RECT 0.000 1808.785 208.285 1809.625 ;
        RECT 0.000 1806.405 208.565 1808.785 ;
      LAYER met2 ;
        RECT 208.940 1806.430 209.200 1806.750 ;
      LAYER met2 ;
        RECT 0.000 1805.565 208.285 1806.405 ;
      LAYER met2 ;
        RECT 209.000 1806.125 209.140 1806.430 ;
        RECT 208.565 1805.845 210.965 1806.125 ;
      LAYER met2 ;
        RECT 0.000 1803.645 208.565 1805.565 ;
        RECT 0.000 1802.805 208.285 1803.645 ;
        RECT 0.000 1800.425 208.565 1802.805 ;
        RECT 0.000 1799.585 208.285 1800.425 ;
        RECT 0.000 1797.205 208.565 1799.585 ;
        RECT 0.000 1796.365 208.285 1797.205 ;
        RECT 0.000 1794.445 208.565 1796.365 ;
        RECT 0.000 1793.605 208.285 1794.445 ;
        RECT 0.000 1791.225 208.565 1793.605 ;
        RECT 0.000 1790.385 208.285 1791.225 ;
      LAYER met2 ;
        RECT 208.565 1790.665 210.965 1790.945 ;
      LAYER met2 ;
        RECT 0.000 1788.005 208.565 1790.385 ;
      LAYER met2 ;
        RECT 209.000 1788.390 209.140 1790.665 ;
        RECT 212.220 1788.390 212.360 2009.410 ;
        RECT 212.680 1845.510 212.820 2056.330 ;
        RECT 213.600 2024.690 213.740 2658.810 ;
        RECT 3373.800 2111.390 3373.940 4982.030 ;
      LAYER met2 ;
        RECT 3390.335 4770.325 3583.075 4794.735 ;
        RECT 3388.000 4767.105 3389.920 4769.105 ;
        RECT 3390.035 4744.890 3583.075 4770.325 ;
        RECT 3413.940 4720.710 3583.075 4744.890 ;
        RECT 3429.550 4532.000 3434.200 4542.975 ;
        RECT 3390.035 4531.500 3587.965 4532.000 ;
        RECT 3390.000 4511.505 3587.965 4531.500 ;
        RECT 3390.035 4511.075 3587.965 4511.505 ;
        RECT 3390.000 4478.465 3587.965 4511.075 ;
        RECT 3390.035 4477.905 3587.965 4478.465 ;
        RECT 3390.000 4457.300 3587.965 4477.905 ;
        RECT 3390.035 4457.000 3587.965 4457.300 ;
        RECT 3413.425 4446.065 3427.835 4455.800 ;
        RECT 3429.585 4445.860 3434.235 4457.000 ;
        RECT 3436.595 4446.065 3587.965 4455.800 ;
        RECT 3379.435 4313.795 3588.000 4314.790 ;
        RECT 3379.715 4312.955 3588.000 4313.795 ;
        RECT 3379.435 4311.035 3588.000 4312.955 ;
        RECT 3379.715 4310.195 3588.000 4311.035 ;
        RECT 3379.435 4307.815 3588.000 4310.195 ;
        RECT 3379.715 4306.975 3588.000 4307.815 ;
        RECT 3379.435 4304.595 3588.000 4306.975 ;
        RECT 3379.715 4303.755 3588.000 4304.595 ;
        RECT 3379.435 4301.835 3588.000 4303.755 ;
        RECT 3379.715 4300.995 3588.000 4301.835 ;
        RECT 3379.435 4298.615 3588.000 4300.995 ;
      LAYER met2 ;
        RECT 3377.035 4298.195 3379.435 4298.335 ;
        RECT 3377.020 4298.055 3379.435 4298.195 ;
        RECT 3377.020 4295.890 3377.160 4298.055 ;
      LAYER met2 ;
        RECT 3379.715 4297.775 3588.000 4298.615 ;
      LAYER met2 ;
        RECT 3376.960 4295.570 3377.220 4295.890 ;
      LAYER met2 ;
        RECT 3379.435 4295.395 3588.000 4297.775 ;
        RECT 3379.715 4294.555 3588.000 4295.395 ;
        RECT 3379.435 4292.635 3588.000 4294.555 ;
        RECT 3379.715 4291.795 3588.000 4292.635 ;
        RECT 3379.435 4289.415 3588.000 4291.795 ;
        RECT 3379.715 4288.575 3588.000 4289.415 ;
        RECT 3379.435 4286.195 3588.000 4288.575 ;
        RECT 3379.715 4285.355 3588.000 4286.195 ;
        RECT 3379.435 4283.435 3588.000 4285.355 ;
      LAYER met2 ;
        RECT 3377.035 4282.980 3379.435 4283.155 ;
        RECT 3377.020 4282.875 3379.435 4282.980 ;
        RECT 3377.020 4280.590 3377.160 4282.875 ;
      LAYER met2 ;
        RECT 3379.715 4282.595 3588.000 4283.435 ;
      LAYER met2 ;
        RECT 3376.960 4280.270 3377.220 4280.590 ;
      LAYER met2 ;
        RECT 3379.435 4280.215 3588.000 4282.595 ;
        RECT 3379.715 4279.375 3588.000 4280.215 ;
        RECT 3379.435 4276.995 3588.000 4279.375 ;
      LAYER met2 ;
        RECT 3377.035 4276.645 3379.435 4276.715 ;
        RECT 3376.560 4276.505 3379.435 4276.645 ;
        RECT 3376.560 4236.625 3376.700 4276.505 ;
        RECT 3377.035 4276.435 3379.435 4276.505 ;
      LAYER met2 ;
        RECT 3379.715 4276.155 3588.000 4276.995 ;
        RECT 3379.435 4273.775 3588.000 4276.155 ;
        RECT 3379.715 4272.935 3588.000 4273.775 ;
        RECT 3379.435 4271.015 3588.000 4272.935 ;
        RECT 3379.715 4270.175 3588.000 4271.015 ;
        RECT 3379.435 4267.795 3588.000 4270.175 ;
        RECT 3379.715 4266.955 3588.000 4267.795 ;
        RECT 3379.435 4264.575 3588.000 4266.955 ;
        RECT 3379.715 4263.735 3588.000 4264.575 ;
        RECT 3379.435 4261.815 3588.000 4263.735 ;
        RECT 3379.715 4260.975 3588.000 4261.815 ;
        RECT 3379.435 4258.595 3588.000 4260.975 ;
        RECT 3379.715 4257.755 3588.000 4258.595 ;
        RECT 3379.435 4255.375 3588.000 4257.755 ;
      LAYER met2 ;
        RECT 3377.035 4254.815 3379.435 4255.095 ;
      LAYER met2 ;
        RECT 3379.715 4254.535 3588.000 4255.375 ;
        RECT 3379.435 4252.615 3588.000 4254.535 ;
        RECT 3379.715 4251.775 3588.000 4252.615 ;
        RECT 3379.435 4249.395 3588.000 4251.775 ;
      LAYER met2 ;
        RECT 3376.960 4248.310 3377.220 4248.630 ;
      LAYER met2 ;
        RECT 3379.715 4248.555 3588.000 4249.395 ;
      LAYER met2 ;
        RECT 3377.020 4245.895 3377.160 4248.310 ;
      LAYER met2 ;
        RECT 3379.435 4246.175 3588.000 4248.555 ;
      LAYER met2 ;
        RECT 3377.020 4245.755 3379.435 4245.895 ;
        RECT 3377.035 4245.615 3379.435 4245.755 ;
      LAYER met2 ;
        RECT 3379.715 4245.335 3588.000 4246.175 ;
        RECT 3379.435 4243.415 3588.000 4245.335 ;
      LAYER met2 ;
        RECT 3377.035 4242.855 3379.435 4243.135 ;
      LAYER met2 ;
        RECT 3379.715 4242.575 3588.000 4243.415 ;
        RECT 3379.435 4240.195 3588.000 4242.575 ;
        RECT 3379.715 4239.355 3588.000 4240.195 ;
        RECT 3379.435 4236.975 3588.000 4239.355 ;
      LAYER met2 ;
        RECT 3377.035 4236.625 3379.435 4236.695 ;
        RECT 3376.560 4236.485 3379.435 4236.625 ;
        RECT 3377.035 4236.415 3379.435 4236.485 ;
      LAYER met2 ;
        RECT 3379.715 4236.135 3588.000 4236.975 ;
        RECT 3379.435 4235.085 3588.000 4236.135 ;
        RECT 3390.035 4093.505 3583.075 4093.735 ;
        RECT 3388.000 4069.605 3583.075 4093.505 ;
        RECT 3388.000 4066.105 3389.920 4068.105 ;
        RECT 3390.035 4043.610 3583.075 4069.605 ;
        RECT 3388.000 4019.710 3583.075 4043.610 ;
      LAYER met2 ;
        RECT 3376.500 4018.810 3376.760 4019.130 ;
        RECT 3387.990 4018.955 3388.270 4019.325 ;
        RECT 3388.000 4018.810 3388.260 4018.955 ;
        RECT 3376.040 3837.930 3376.300 3838.250 ;
        RECT 3376.100 3801.190 3376.240 3837.930 ;
        RECT 3376.040 3800.870 3376.300 3801.190 ;
        RECT 3376.560 3698.470 3376.700 4018.810 ;
      LAYER met2 ;
        RECT 3379.435 3876.795 3588.000 3877.790 ;
        RECT 3379.715 3875.955 3588.000 3876.795 ;
        RECT 3379.435 3874.035 3588.000 3875.955 ;
        RECT 3379.715 3873.195 3588.000 3874.035 ;
        RECT 3379.435 3870.815 3588.000 3873.195 ;
        RECT 3379.715 3869.975 3588.000 3870.815 ;
        RECT 3379.435 3867.595 3588.000 3869.975 ;
        RECT 3379.715 3866.755 3588.000 3867.595 ;
        RECT 3379.435 3864.835 3588.000 3866.755 ;
      LAYER met2 ;
        RECT 3376.960 3863.770 3377.220 3864.090 ;
      LAYER met2 ;
        RECT 3379.715 3863.995 3588.000 3864.835 ;
      LAYER met2 ;
        RECT 3377.020 3861.335 3377.160 3863.770 ;
      LAYER met2 ;
        RECT 3379.435 3861.615 3588.000 3863.995 ;
      LAYER met2 ;
        RECT 3377.020 3861.195 3379.435 3861.335 ;
        RECT 3377.035 3861.055 3379.435 3861.195 ;
      LAYER met2 ;
        RECT 3379.715 3860.775 3588.000 3861.615 ;
        RECT 3379.435 3858.395 3588.000 3860.775 ;
        RECT 3379.715 3857.555 3588.000 3858.395 ;
        RECT 3379.435 3855.635 3588.000 3857.555 ;
        RECT 3379.715 3854.795 3588.000 3855.635 ;
        RECT 3379.435 3852.415 3588.000 3854.795 ;
        RECT 3379.715 3851.575 3588.000 3852.415 ;
        RECT 3379.435 3849.195 3588.000 3851.575 ;
      LAYER met2 ;
        RECT 3376.960 3848.130 3377.220 3848.450 ;
      LAYER met2 ;
        RECT 3379.715 3848.355 3588.000 3849.195 ;
      LAYER met2 ;
        RECT 3377.020 3846.155 3377.160 3848.130 ;
      LAYER met2 ;
        RECT 3379.435 3846.435 3588.000 3848.355 ;
      LAYER met2 ;
        RECT 3377.020 3846.015 3379.435 3846.155 ;
        RECT 3377.035 3845.875 3379.435 3846.015 ;
      LAYER met2 ;
        RECT 3379.715 3845.595 3588.000 3846.435 ;
        RECT 3379.435 3843.215 3588.000 3845.595 ;
        RECT 3379.715 3842.375 3588.000 3843.215 ;
        RECT 3379.435 3839.995 3588.000 3842.375 ;
      LAYER met2 ;
        RECT 3377.035 3839.620 3379.435 3839.715 ;
        RECT 3377.020 3839.435 3379.435 3839.620 ;
        RECT 3377.020 3838.250 3377.160 3839.435 ;
      LAYER met2 ;
        RECT 3379.715 3839.155 3588.000 3839.995 ;
      LAYER met2 ;
        RECT 3376.960 3837.930 3377.220 3838.250 ;
      LAYER met2 ;
        RECT 3379.435 3836.775 3588.000 3839.155 ;
        RECT 3379.715 3835.935 3588.000 3836.775 ;
        RECT 3379.435 3834.015 3588.000 3835.935 ;
        RECT 3379.715 3833.175 3588.000 3834.015 ;
        RECT 3379.435 3830.795 3588.000 3833.175 ;
        RECT 3379.715 3829.955 3588.000 3830.795 ;
        RECT 3379.435 3827.575 3588.000 3829.955 ;
        RECT 3379.715 3826.735 3588.000 3827.575 ;
        RECT 3379.435 3824.815 3588.000 3826.735 ;
        RECT 3379.715 3823.975 3588.000 3824.815 ;
        RECT 3379.435 3821.595 3588.000 3823.975 ;
        RECT 3379.715 3820.755 3588.000 3821.595 ;
        RECT 3379.435 3818.375 3588.000 3820.755 ;
      LAYER met2 ;
        RECT 3377.035 3817.815 3379.435 3818.095 ;
      LAYER met2 ;
        RECT 3379.715 3817.535 3588.000 3818.375 ;
        RECT 3379.435 3815.615 3588.000 3817.535 ;
        RECT 3379.715 3814.775 3588.000 3815.615 ;
        RECT 3379.435 3812.395 3588.000 3814.775 ;
        RECT 3379.715 3811.555 3588.000 3812.395 ;
        RECT 3379.435 3809.175 3588.000 3811.555 ;
      LAYER met2 ;
        RECT 3377.035 3808.755 3379.435 3808.895 ;
        RECT 3377.020 3808.615 3379.435 3808.755 ;
        RECT 3377.020 3806.630 3377.160 3808.615 ;
      LAYER met2 ;
        RECT 3379.715 3808.335 3588.000 3809.175 ;
      LAYER met2 ;
        RECT 3376.960 3806.310 3377.220 3806.630 ;
      LAYER met2 ;
        RECT 3379.435 3806.415 3588.000 3808.335 ;
      LAYER met2 ;
        RECT 3377.035 3805.855 3379.435 3806.135 ;
      LAYER met2 ;
        RECT 3379.715 3805.575 3588.000 3806.415 ;
        RECT 3379.435 3803.195 3588.000 3805.575 ;
        RECT 3379.715 3802.355 3588.000 3803.195 ;
      LAYER met2 ;
        RECT 3376.960 3800.870 3377.220 3801.190 ;
        RECT 3377.020 3799.695 3377.160 3800.870 ;
      LAYER met2 ;
        RECT 3379.435 3799.975 3588.000 3802.355 ;
      LAYER met2 ;
        RECT 3377.020 3799.500 3379.435 3799.695 ;
        RECT 3377.035 3799.415 3379.435 3799.500 ;
      LAYER met2 ;
        RECT 3379.715 3799.135 3588.000 3799.975 ;
        RECT 3379.435 3798.085 3588.000 3799.135 ;
      LAYER met2 ;
        RECT 3375.640 3698.330 3376.700 3698.470 ;
        RECT 3375.640 3546.670 3375.780 3698.330 ;
      LAYER met2 ;
        RECT 3379.435 3654.795 3588.000 3655.790 ;
        RECT 3379.715 3653.955 3588.000 3654.795 ;
        RECT 3379.435 3652.035 3588.000 3653.955 ;
        RECT 3379.715 3651.195 3588.000 3652.035 ;
        RECT 3379.435 3648.815 3588.000 3651.195 ;
        RECT 3379.715 3647.975 3588.000 3648.815 ;
        RECT 3379.435 3645.595 3588.000 3647.975 ;
        RECT 3379.715 3644.755 3588.000 3645.595 ;
        RECT 3379.435 3642.835 3588.000 3644.755 ;
      LAYER met2 ;
        RECT 3376.960 3641.750 3377.220 3642.070 ;
      LAYER met2 ;
        RECT 3379.715 3641.995 3588.000 3642.835 ;
      LAYER met2 ;
        RECT 3377.020 3639.335 3377.160 3641.750 ;
      LAYER met2 ;
        RECT 3379.435 3639.615 3588.000 3641.995 ;
      LAYER met2 ;
        RECT 3377.020 3639.195 3379.435 3639.335 ;
        RECT 3377.035 3639.055 3379.435 3639.195 ;
      LAYER met2 ;
        RECT 3379.715 3638.775 3588.000 3639.615 ;
        RECT 3379.435 3636.395 3588.000 3638.775 ;
        RECT 3379.715 3635.555 3588.000 3636.395 ;
        RECT 3379.435 3633.635 3588.000 3635.555 ;
        RECT 3379.715 3632.795 3588.000 3633.635 ;
        RECT 3379.435 3630.415 3588.000 3632.795 ;
        RECT 3379.715 3629.575 3588.000 3630.415 ;
        RECT 3379.435 3627.195 3588.000 3629.575 ;
      LAYER met2 ;
        RECT 3376.960 3626.110 3377.220 3626.430 ;
      LAYER met2 ;
        RECT 3379.715 3626.355 3588.000 3627.195 ;
      LAYER met2 ;
        RECT 3377.020 3624.155 3377.160 3626.110 ;
      LAYER met2 ;
        RECT 3379.435 3624.435 3588.000 3626.355 ;
      LAYER met2 ;
        RECT 3377.020 3624.060 3379.435 3624.155 ;
        RECT 3377.035 3623.875 3379.435 3624.060 ;
      LAYER met2 ;
        RECT 3379.715 3623.595 3588.000 3624.435 ;
        RECT 3379.435 3621.215 3588.000 3623.595 ;
        RECT 3379.715 3620.375 3588.000 3621.215 ;
        RECT 3379.435 3617.995 3588.000 3620.375 ;
      LAYER met2 ;
        RECT 3377.035 3617.645 3379.435 3617.715 ;
        RECT 3376.100 3617.505 3379.435 3617.645 ;
        RECT 3376.100 3577.625 3376.240 3617.505 ;
        RECT 3377.035 3617.435 3379.435 3617.505 ;
      LAYER met2 ;
        RECT 3379.715 3617.155 3588.000 3617.995 ;
        RECT 3379.435 3614.775 3588.000 3617.155 ;
        RECT 3379.715 3613.935 3588.000 3614.775 ;
        RECT 3379.435 3612.015 3588.000 3613.935 ;
        RECT 3379.715 3611.175 3588.000 3612.015 ;
        RECT 3379.435 3608.795 3588.000 3611.175 ;
        RECT 3379.715 3607.955 3588.000 3608.795 ;
        RECT 3379.435 3605.575 3588.000 3607.955 ;
        RECT 3379.715 3604.735 3588.000 3605.575 ;
        RECT 3379.435 3602.815 3588.000 3604.735 ;
        RECT 3379.715 3601.975 3588.000 3602.815 ;
        RECT 3379.435 3599.595 3588.000 3601.975 ;
        RECT 3379.715 3598.755 3588.000 3599.595 ;
        RECT 3379.435 3596.375 3588.000 3598.755 ;
      LAYER met2 ;
        RECT 3377.035 3595.815 3379.435 3596.095 ;
      LAYER met2 ;
        RECT 3379.715 3595.535 3588.000 3596.375 ;
        RECT 3379.435 3593.615 3588.000 3595.535 ;
        RECT 3379.715 3592.775 3588.000 3593.615 ;
        RECT 3379.435 3590.395 3588.000 3592.775 ;
        RECT 3379.715 3589.555 3588.000 3590.395 ;
      LAYER met2 ;
        RECT 3376.960 3589.050 3377.220 3589.370 ;
        RECT 3377.020 3586.895 3377.160 3589.050 ;
      LAYER met2 ;
        RECT 3379.435 3587.175 3588.000 3589.555 ;
      LAYER met2 ;
        RECT 3377.020 3586.660 3379.435 3586.895 ;
        RECT 3377.035 3586.615 3379.435 3586.660 ;
      LAYER met2 ;
        RECT 3379.715 3586.335 3588.000 3587.175 ;
        RECT 3379.435 3584.415 3588.000 3586.335 ;
      LAYER met2 ;
        RECT 3377.035 3583.855 3379.435 3584.135 ;
      LAYER met2 ;
        RECT 3379.715 3583.575 3588.000 3584.415 ;
        RECT 3379.435 3581.195 3588.000 3583.575 ;
        RECT 3379.715 3580.355 3588.000 3581.195 ;
        RECT 3379.435 3577.975 3588.000 3580.355 ;
      LAYER met2 ;
        RECT 3377.035 3577.625 3379.435 3577.695 ;
        RECT 3376.100 3577.485 3379.435 3577.625 ;
        RECT 3377.035 3577.415 3379.435 3577.485 ;
      LAYER met2 ;
        RECT 3379.715 3577.135 3588.000 3577.975 ;
        RECT 3379.435 3576.085 3588.000 3577.135 ;
      LAYER met2 ;
        RECT 3375.640 3546.530 3376.700 3546.670 ;
        RECT 3376.560 3450.070 3376.700 3546.530 ;
        RECT 3375.640 3449.930 3376.700 3450.070 ;
        RECT 3375.640 3353.470 3375.780 3449.930 ;
      LAYER met2 ;
        RECT 3379.435 3433.795 3588.000 3434.790 ;
        RECT 3379.715 3432.955 3588.000 3433.795 ;
        RECT 3379.435 3431.035 3588.000 3432.955 ;
        RECT 3379.715 3430.195 3588.000 3431.035 ;
        RECT 3379.435 3427.815 3588.000 3430.195 ;
        RECT 3379.715 3426.975 3588.000 3427.815 ;
        RECT 3379.435 3424.595 3588.000 3426.975 ;
        RECT 3379.715 3423.755 3588.000 3424.595 ;
        RECT 3379.435 3421.835 3588.000 3423.755 ;
        RECT 3379.715 3420.995 3588.000 3421.835 ;
        RECT 3379.435 3418.615 3588.000 3420.995 ;
      LAYER met2 ;
        RECT 3377.035 3418.195 3379.435 3418.335 ;
        RECT 3377.020 3418.055 3379.435 3418.195 ;
        RECT 3377.020 3415.630 3377.160 3418.055 ;
      LAYER met2 ;
        RECT 3379.715 3417.775 3588.000 3418.615 ;
      LAYER met2 ;
        RECT 3376.960 3415.310 3377.220 3415.630 ;
      LAYER met2 ;
        RECT 3379.435 3415.395 3588.000 3417.775 ;
        RECT 3379.715 3414.555 3588.000 3415.395 ;
        RECT 3379.435 3412.635 3588.000 3414.555 ;
        RECT 3379.715 3411.795 3588.000 3412.635 ;
        RECT 3379.435 3409.415 3588.000 3411.795 ;
        RECT 3379.715 3408.575 3588.000 3409.415 ;
        RECT 3379.435 3406.195 3588.000 3408.575 ;
        RECT 3379.715 3405.355 3588.000 3406.195 ;
        RECT 3379.435 3403.435 3588.000 3405.355 ;
      LAYER met2 ;
        RECT 3377.035 3403.060 3379.435 3403.155 ;
        RECT 3377.020 3402.875 3379.435 3403.060 ;
        RECT 3377.020 3402.370 3377.160 3402.875 ;
      LAYER met2 ;
        RECT 3379.715 3402.595 3588.000 3403.435 ;
      LAYER met2 ;
        RECT 3376.960 3402.050 3377.220 3402.370 ;
      LAYER met2 ;
        RECT 3379.435 3400.215 3588.000 3402.595 ;
        RECT 3379.715 3399.375 3588.000 3400.215 ;
        RECT 3379.435 3396.995 3588.000 3399.375 ;
      LAYER met2 ;
        RECT 3377.035 3396.575 3379.435 3396.715 ;
        RECT 3377.020 3396.435 3379.435 3396.575 ;
        RECT 3377.020 3394.210 3377.160 3396.435 ;
      LAYER met2 ;
        RECT 3379.715 3396.155 3588.000 3396.995 ;
      LAYER met2 ;
        RECT 3376.040 3393.890 3376.300 3394.210 ;
        RECT 3376.960 3393.890 3377.220 3394.210 ;
        RECT 3376.100 3356.625 3376.240 3393.890 ;
      LAYER met2 ;
        RECT 3379.435 3393.775 3588.000 3396.155 ;
        RECT 3379.715 3392.935 3588.000 3393.775 ;
        RECT 3379.435 3391.015 3588.000 3392.935 ;
        RECT 3379.715 3390.175 3588.000 3391.015 ;
        RECT 3379.435 3387.795 3588.000 3390.175 ;
        RECT 3379.715 3386.955 3588.000 3387.795 ;
        RECT 3379.435 3384.575 3588.000 3386.955 ;
        RECT 3379.715 3383.735 3588.000 3384.575 ;
        RECT 3379.435 3381.815 3588.000 3383.735 ;
        RECT 3379.715 3380.975 3588.000 3381.815 ;
        RECT 3379.435 3378.595 3588.000 3380.975 ;
        RECT 3379.715 3377.755 3588.000 3378.595 ;
        RECT 3379.435 3375.375 3588.000 3377.755 ;
      LAYER met2 ;
        RECT 3377.035 3374.815 3379.435 3375.095 ;
      LAYER met2 ;
        RECT 3379.715 3374.535 3588.000 3375.375 ;
        RECT 3379.435 3372.615 3588.000 3374.535 ;
        RECT 3379.715 3371.775 3588.000 3372.615 ;
        RECT 3379.435 3369.395 3588.000 3371.775 ;
        RECT 3379.715 3368.555 3588.000 3369.395 ;
      LAYER met2 ;
        RECT 3376.960 3368.050 3377.220 3368.370 ;
        RECT 3377.020 3365.895 3377.160 3368.050 ;
      LAYER met2 ;
        RECT 3379.435 3366.175 3588.000 3368.555 ;
      LAYER met2 ;
        RECT 3377.020 3365.660 3379.435 3365.895 ;
        RECT 3377.035 3365.615 3379.435 3365.660 ;
      LAYER met2 ;
        RECT 3379.715 3365.335 3588.000 3366.175 ;
        RECT 3379.435 3363.415 3588.000 3365.335 ;
      LAYER met2 ;
        RECT 3377.035 3362.855 3379.435 3363.135 ;
      LAYER met2 ;
        RECT 3379.715 3362.575 3588.000 3363.415 ;
        RECT 3379.435 3360.195 3588.000 3362.575 ;
        RECT 3379.715 3359.355 3588.000 3360.195 ;
        RECT 3379.435 3356.975 3588.000 3359.355 ;
      LAYER met2 ;
        RECT 3377.035 3356.625 3379.435 3356.695 ;
        RECT 3376.100 3356.485 3379.435 3356.625 ;
        RECT 3377.035 3356.415 3379.435 3356.485 ;
      LAYER met2 ;
        RECT 3379.715 3356.135 3588.000 3356.975 ;
        RECT 3379.435 3355.085 3588.000 3356.135 ;
      LAYER met2 ;
        RECT 3375.640 3353.330 3376.700 3353.470 ;
        RECT 3376.560 3256.870 3376.700 3353.330 ;
        RECT 3375.640 3256.730 3376.700 3256.870 ;
        RECT 3375.640 3118.870 3375.780 3256.730 ;
      LAYER met2 ;
        RECT 3379.435 3212.795 3588.000 3213.790 ;
        RECT 3379.715 3211.955 3588.000 3212.795 ;
        RECT 3379.435 3210.035 3588.000 3211.955 ;
        RECT 3379.715 3209.195 3588.000 3210.035 ;
        RECT 3379.435 3206.815 3588.000 3209.195 ;
        RECT 3379.715 3205.975 3588.000 3206.815 ;
        RECT 3379.435 3203.595 3588.000 3205.975 ;
        RECT 3379.715 3202.755 3588.000 3203.595 ;
        RECT 3379.435 3200.835 3588.000 3202.755 ;
        RECT 3379.715 3199.995 3588.000 3200.835 ;
        RECT 3379.435 3197.615 3588.000 3199.995 ;
      LAYER met2 ;
        RECT 3377.035 3197.195 3379.435 3197.335 ;
        RECT 3377.020 3197.055 3379.435 3197.195 ;
        RECT 3377.020 3194.630 3377.160 3197.055 ;
      LAYER met2 ;
        RECT 3379.715 3196.775 3588.000 3197.615 ;
      LAYER met2 ;
        RECT 3376.960 3194.310 3377.220 3194.630 ;
      LAYER met2 ;
        RECT 3379.435 3194.395 3588.000 3196.775 ;
        RECT 3379.715 3193.555 3588.000 3194.395 ;
        RECT 3379.435 3191.635 3588.000 3193.555 ;
        RECT 3379.715 3190.795 3588.000 3191.635 ;
        RECT 3379.435 3188.415 3588.000 3190.795 ;
        RECT 3379.715 3187.575 3588.000 3188.415 ;
        RECT 3379.435 3185.195 3588.000 3187.575 ;
        RECT 3379.715 3184.355 3588.000 3185.195 ;
        RECT 3379.435 3182.435 3588.000 3184.355 ;
      LAYER met2 ;
        RECT 3377.035 3182.060 3379.435 3182.155 ;
        RECT 3377.020 3181.875 3379.435 3182.060 ;
        RECT 3377.020 3181.710 3377.160 3181.875 ;
        RECT 3376.960 3181.390 3377.220 3181.710 ;
      LAYER met2 ;
        RECT 3379.715 3181.595 3588.000 3182.435 ;
        RECT 3379.435 3179.215 3588.000 3181.595 ;
        RECT 3379.715 3178.375 3588.000 3179.215 ;
        RECT 3379.435 3175.995 3588.000 3178.375 ;
      LAYER met2 ;
        RECT 3377.035 3175.575 3379.435 3175.715 ;
        RECT 3377.020 3175.435 3379.435 3175.575 ;
        RECT 3377.020 3173.210 3377.160 3175.435 ;
      LAYER met2 ;
        RECT 3379.715 3175.155 3588.000 3175.995 ;
      LAYER met2 ;
        RECT 3376.040 3172.890 3376.300 3173.210 ;
        RECT 3376.960 3172.890 3377.220 3173.210 ;
        RECT 3376.100 3135.625 3376.240 3172.890 ;
      LAYER met2 ;
        RECT 3379.435 3172.775 3588.000 3175.155 ;
        RECT 3379.715 3171.935 3588.000 3172.775 ;
        RECT 3379.435 3170.015 3588.000 3171.935 ;
        RECT 3379.715 3169.175 3588.000 3170.015 ;
        RECT 3379.435 3166.795 3588.000 3169.175 ;
        RECT 3379.715 3165.955 3588.000 3166.795 ;
        RECT 3379.435 3163.575 3588.000 3165.955 ;
        RECT 3379.715 3162.735 3588.000 3163.575 ;
        RECT 3379.435 3160.815 3588.000 3162.735 ;
        RECT 3379.715 3159.975 3588.000 3160.815 ;
        RECT 3379.435 3157.595 3588.000 3159.975 ;
        RECT 3379.715 3156.755 3588.000 3157.595 ;
        RECT 3379.435 3154.375 3588.000 3156.755 ;
      LAYER met2 ;
        RECT 3377.035 3153.815 3379.435 3154.095 ;
      LAYER met2 ;
        RECT 3379.715 3153.535 3588.000 3154.375 ;
        RECT 3379.435 3151.615 3588.000 3153.535 ;
        RECT 3379.715 3150.775 3588.000 3151.615 ;
        RECT 3379.435 3148.395 3588.000 3150.775 ;
        RECT 3379.715 3147.555 3588.000 3148.395 ;
      LAYER met2 ;
        RECT 3376.960 3147.050 3377.220 3147.370 ;
        RECT 3377.020 3144.895 3377.160 3147.050 ;
      LAYER met2 ;
        RECT 3379.435 3145.175 3588.000 3147.555 ;
      LAYER met2 ;
        RECT 3377.020 3144.660 3379.435 3144.895 ;
        RECT 3377.035 3144.615 3379.435 3144.660 ;
      LAYER met2 ;
        RECT 3379.715 3144.335 3588.000 3145.175 ;
        RECT 3379.435 3142.415 3588.000 3144.335 ;
      LAYER met2 ;
        RECT 3377.035 3141.855 3379.435 3142.135 ;
      LAYER met2 ;
        RECT 3379.715 3141.575 3588.000 3142.415 ;
        RECT 3379.435 3139.195 3588.000 3141.575 ;
        RECT 3379.715 3138.355 3588.000 3139.195 ;
        RECT 3379.435 3135.975 3588.000 3138.355 ;
      LAYER met2 ;
        RECT 3377.035 3135.625 3379.435 3135.695 ;
        RECT 3376.100 3135.485 3379.435 3135.625 ;
        RECT 3377.035 3135.415 3379.435 3135.485 ;
      LAYER met2 ;
        RECT 3379.715 3135.135 3588.000 3135.975 ;
        RECT 3379.435 3134.085 3588.000 3135.135 ;
      LAYER met2 ;
        RECT 3375.640 3118.730 3376.700 3118.870 ;
        RECT 3376.560 2951.610 3376.700 3118.730 ;
      LAYER met2 ;
        RECT 3379.435 2990.795 3588.000 2991.790 ;
        RECT 3379.715 2989.955 3588.000 2990.795 ;
        RECT 3379.435 2988.035 3588.000 2989.955 ;
        RECT 3379.715 2987.195 3588.000 2988.035 ;
        RECT 3379.435 2984.815 3588.000 2987.195 ;
        RECT 3379.715 2983.975 3588.000 2984.815 ;
        RECT 3379.435 2981.595 3588.000 2983.975 ;
        RECT 3379.715 2980.755 3588.000 2981.595 ;
        RECT 3379.435 2978.835 3588.000 2980.755 ;
        RECT 3379.715 2977.995 3588.000 2978.835 ;
      LAYER met2 ;
        RECT 3376.960 2975.690 3377.220 2976.010 ;
        RECT 3377.020 2975.335 3377.160 2975.690 ;
      LAYER met2 ;
        RECT 3379.435 2975.615 3588.000 2977.995 ;
      LAYER met2 ;
        RECT 3377.020 2975.195 3379.435 2975.335 ;
        RECT 3377.035 2975.055 3379.435 2975.195 ;
      LAYER met2 ;
        RECT 3379.715 2974.775 3588.000 2975.615 ;
        RECT 3379.435 2972.395 3588.000 2974.775 ;
        RECT 3379.715 2971.555 3588.000 2972.395 ;
        RECT 3379.435 2969.635 3588.000 2971.555 ;
        RECT 3379.715 2968.795 3588.000 2969.635 ;
        RECT 3379.435 2966.415 3588.000 2968.795 ;
        RECT 3379.715 2965.575 3588.000 2966.415 ;
        RECT 3379.435 2963.195 3588.000 2965.575 ;
        RECT 3379.715 2962.355 3588.000 2963.195 ;
        RECT 3379.435 2960.435 3588.000 2962.355 ;
      LAYER met2 ;
        RECT 3377.035 2960.015 3379.435 2960.155 ;
        RECT 3377.020 2959.875 3379.435 2960.015 ;
        RECT 3377.020 2959.690 3377.160 2959.875 ;
        RECT 3376.960 2959.370 3377.220 2959.690 ;
      LAYER met2 ;
        RECT 3379.715 2959.595 3588.000 2960.435 ;
        RECT 3379.435 2957.215 3588.000 2959.595 ;
        RECT 3379.715 2956.375 3588.000 2957.215 ;
        RECT 3379.435 2953.995 3588.000 2956.375 ;
      LAYER met2 ;
        RECT 3377.035 2953.580 3379.435 2953.715 ;
        RECT 3375.640 2951.470 3376.700 2951.610 ;
        RECT 3377.020 2953.435 3379.435 2953.580 ;
        RECT 3375.640 2677.270 3375.780 2951.470 ;
        RECT 3377.020 2950.930 3377.160 2953.435 ;
      LAYER met2 ;
        RECT 3379.715 2953.155 3588.000 2953.995 ;
      LAYER met2 ;
        RECT 3376.560 2950.790 3377.160 2950.930 ;
        RECT 3376.560 2916.250 3376.700 2950.790 ;
      LAYER met2 ;
        RECT 3379.435 2950.775 3588.000 2953.155 ;
        RECT 3379.715 2949.935 3588.000 2950.775 ;
        RECT 3379.435 2948.015 3588.000 2949.935 ;
        RECT 3379.715 2947.175 3588.000 2948.015 ;
        RECT 3379.435 2944.795 3588.000 2947.175 ;
        RECT 3379.715 2943.955 3588.000 2944.795 ;
        RECT 3379.435 2941.575 3588.000 2943.955 ;
        RECT 3379.715 2940.735 3588.000 2941.575 ;
        RECT 3379.435 2938.815 3588.000 2940.735 ;
        RECT 3379.715 2937.975 3588.000 2938.815 ;
        RECT 3379.435 2935.595 3588.000 2937.975 ;
        RECT 3379.715 2934.755 3588.000 2935.595 ;
        RECT 3379.435 2932.375 3588.000 2934.755 ;
      LAYER met2 ;
        RECT 3377.035 2931.815 3379.435 2932.095 ;
      LAYER met2 ;
        RECT 3379.715 2931.535 3588.000 2932.375 ;
        RECT 3379.435 2929.615 3588.000 2931.535 ;
        RECT 3379.715 2928.775 3588.000 2929.615 ;
        RECT 3379.435 2926.395 3588.000 2928.775 ;
        RECT 3379.715 2925.555 3588.000 2926.395 ;
        RECT 3379.435 2923.175 3588.000 2925.555 ;
      LAYER met2 ;
        RECT 3377.035 2922.755 3379.435 2922.895 ;
        RECT 3377.020 2922.615 3379.435 2922.755 ;
        RECT 3377.020 2920.930 3377.160 2922.615 ;
      LAYER met2 ;
        RECT 3379.715 2922.335 3588.000 2923.175 ;
      LAYER met2 ;
        RECT 3376.960 2920.610 3377.220 2920.930 ;
      LAYER met2 ;
        RECT 3379.435 2920.415 3588.000 2922.335 ;
      LAYER met2 ;
        RECT 3377.035 2919.855 3379.435 2920.135 ;
      LAYER met2 ;
        RECT 3379.715 2919.575 3588.000 2920.415 ;
        RECT 3379.435 2917.195 3588.000 2919.575 ;
        RECT 3379.715 2916.355 3588.000 2917.195 ;
      LAYER met2 ;
        RECT 3376.560 2916.110 3377.160 2916.250 ;
        RECT 3377.020 2913.695 3377.160 2916.110 ;
      LAYER met2 ;
        RECT 3379.435 2913.975 3588.000 2916.355 ;
      LAYER met2 ;
        RECT 3377.020 2913.460 3379.435 2913.695 ;
        RECT 3377.035 2913.415 3379.435 2913.460 ;
      LAYER met2 ;
        RECT 3379.715 2913.135 3588.000 2913.975 ;
        RECT 3379.435 2912.085 3588.000 2913.135 ;
        RECT 3379.435 2769.795 3588.000 2770.790 ;
        RECT 3379.715 2768.955 3588.000 2769.795 ;
        RECT 3379.435 2767.035 3588.000 2768.955 ;
        RECT 3379.715 2766.195 3588.000 2767.035 ;
        RECT 3379.435 2763.815 3588.000 2766.195 ;
        RECT 3379.715 2762.975 3588.000 2763.815 ;
        RECT 3379.435 2760.595 3588.000 2762.975 ;
        RECT 3379.715 2759.755 3588.000 2760.595 ;
        RECT 3379.435 2757.835 3588.000 2759.755 ;
      LAYER met2 ;
        RECT 3376.960 2756.730 3377.220 2757.050 ;
      LAYER met2 ;
        RECT 3379.715 2756.995 3588.000 2757.835 ;
      LAYER met2 ;
        RECT 3377.020 2754.335 3377.160 2756.730 ;
      LAYER met2 ;
        RECT 3379.435 2754.615 3588.000 2756.995 ;
      LAYER met2 ;
        RECT 3377.020 2754.195 3379.435 2754.335 ;
        RECT 3377.035 2754.055 3379.435 2754.195 ;
      LAYER met2 ;
        RECT 3379.715 2753.775 3588.000 2754.615 ;
        RECT 3379.435 2751.395 3588.000 2753.775 ;
        RECT 3379.715 2750.555 3588.000 2751.395 ;
        RECT 3379.435 2748.635 3588.000 2750.555 ;
        RECT 3379.715 2747.795 3588.000 2748.635 ;
        RECT 3379.435 2745.415 3588.000 2747.795 ;
        RECT 3379.715 2744.575 3588.000 2745.415 ;
        RECT 3379.435 2742.195 3588.000 2744.575 ;
      LAYER met2 ;
        RECT 3376.960 2741.090 3377.220 2741.410 ;
      LAYER met2 ;
        RECT 3379.715 2741.355 3588.000 2742.195 ;
      LAYER met2 ;
        RECT 3377.020 2739.155 3377.160 2741.090 ;
      LAYER met2 ;
        RECT 3379.435 2739.435 3588.000 2741.355 ;
      LAYER met2 ;
        RECT 3377.020 2739.015 3379.435 2739.155 ;
        RECT 3377.035 2738.875 3379.435 2739.015 ;
      LAYER met2 ;
        RECT 3379.715 2738.595 3588.000 2739.435 ;
        RECT 3379.435 2736.215 3588.000 2738.595 ;
        RECT 3379.715 2735.375 3588.000 2736.215 ;
        RECT 3379.435 2732.995 3588.000 2735.375 ;
      LAYER met2 ;
        RECT 3377.035 2732.650 3379.435 2732.715 ;
        RECT 3376.560 2732.510 3379.435 2732.650 ;
        RECT 3376.560 2695.250 3376.700 2732.510 ;
        RECT 3377.035 2732.435 3379.435 2732.510 ;
      LAYER met2 ;
        RECT 3379.715 2732.155 3588.000 2732.995 ;
        RECT 3379.435 2729.775 3588.000 2732.155 ;
        RECT 3379.715 2728.935 3588.000 2729.775 ;
        RECT 3379.435 2727.015 3588.000 2728.935 ;
        RECT 3379.715 2726.175 3588.000 2727.015 ;
        RECT 3379.435 2723.795 3588.000 2726.175 ;
        RECT 3379.715 2722.955 3588.000 2723.795 ;
        RECT 3379.435 2720.575 3588.000 2722.955 ;
        RECT 3379.715 2719.735 3588.000 2720.575 ;
        RECT 3379.435 2717.815 3588.000 2719.735 ;
        RECT 3379.715 2716.975 3588.000 2717.815 ;
        RECT 3379.435 2714.595 3588.000 2716.975 ;
        RECT 3379.715 2713.755 3588.000 2714.595 ;
        RECT 3379.435 2711.375 3588.000 2713.755 ;
      LAYER met2 ;
        RECT 3377.035 2710.815 3379.435 2711.095 ;
      LAYER met2 ;
        RECT 3379.715 2710.535 3588.000 2711.375 ;
        RECT 3379.435 2708.615 3588.000 2710.535 ;
        RECT 3379.715 2707.775 3588.000 2708.615 ;
        RECT 3379.435 2705.395 3588.000 2707.775 ;
      LAYER met2 ;
        RECT 3376.960 2704.370 3377.220 2704.690 ;
      LAYER met2 ;
        RECT 3379.715 2704.555 3588.000 2705.395 ;
      LAYER met2 ;
        RECT 3377.020 2701.895 3377.160 2704.370 ;
      LAYER met2 ;
        RECT 3379.435 2702.175 3588.000 2704.555 ;
      LAYER met2 ;
        RECT 3377.020 2701.755 3379.435 2701.895 ;
        RECT 3377.035 2701.615 3379.435 2701.755 ;
      LAYER met2 ;
        RECT 3379.715 2701.335 3588.000 2702.175 ;
        RECT 3379.435 2699.415 3588.000 2701.335 ;
      LAYER met2 ;
        RECT 3377.035 2698.855 3379.435 2699.135 ;
      LAYER met2 ;
        RECT 3379.715 2698.575 3588.000 2699.415 ;
        RECT 3379.435 2696.195 3588.000 2698.575 ;
        RECT 3379.715 2695.355 3588.000 2696.195 ;
      LAYER met2 ;
        RECT 3376.560 2695.110 3377.160 2695.250 ;
        RECT 3377.020 2692.695 3377.160 2695.110 ;
      LAYER met2 ;
        RECT 3379.435 2692.975 3588.000 2695.355 ;
      LAYER met2 ;
        RECT 3377.020 2692.460 3379.435 2692.695 ;
        RECT 3377.035 2692.415 3379.435 2692.460 ;
      LAYER met2 ;
        RECT 3379.715 2692.135 3588.000 2692.975 ;
        RECT 3379.435 2691.085 3588.000 2692.135 ;
      LAYER met2 ;
        RECT 3375.640 2677.130 3376.700 2677.270 ;
        RECT 3376.560 2497.630 3376.700 2677.130 ;
      LAYER met2 ;
        RECT 3390.035 2549.505 3583.075 2549.735 ;
        RECT 3388.000 2525.605 3583.075 2549.505 ;
        RECT 3388.000 2522.105 3389.920 2524.105 ;
        RECT 3390.035 2499.610 3583.075 2525.605 ;
      LAYER met2 ;
        RECT 3376.500 2497.310 3376.760 2497.630 ;
        RECT 3380.640 2497.310 3380.900 2497.630 ;
        RECT 3380.700 2474.510 3380.840 2497.310 ;
      LAYER met2 ;
        RECT 3388.000 2475.710 3583.075 2499.610 ;
      LAYER met2 ;
        RECT 3380.640 2474.190 3380.900 2474.510 ;
        RECT 3389.840 2474.365 3390.100 2474.510 ;
        RECT 3389.830 2473.995 3390.110 2474.365 ;
      LAYER met2 ;
        RECT 3429.550 2333.000 3434.200 2343.975 ;
        RECT 3390.035 2332.500 3587.965 2333.000 ;
        RECT 3390.000 2312.505 3587.965 2332.500 ;
        RECT 3390.035 2312.075 3587.965 2312.505 ;
        RECT 3390.000 2279.465 3587.965 2312.075 ;
        RECT 3390.035 2278.905 3587.965 2279.465 ;
        RECT 3390.000 2258.300 3587.965 2278.905 ;
        RECT 3390.035 2258.000 3587.965 2258.300 ;
        RECT 3413.425 2247.065 3427.835 2256.800 ;
        RECT 3429.585 2246.860 3434.235 2258.000 ;
        RECT 3436.595 2247.065 3587.965 2256.800 ;
        RECT 3390.035 2116.505 3583.075 2116.735 ;
      LAYER met2 ;
        RECT 3370.060 2111.070 3370.320 2111.390 ;
        RECT 3373.740 2111.070 3374.000 2111.390 ;
        RECT 3370.120 2099.685 3370.260 2111.070 ;
        RECT 3370.050 2099.315 3370.330 2099.685 ;
        RECT 3370.050 2095.915 3370.330 2096.285 ;
        RECT 3370.060 2095.770 3370.320 2095.915 ;
        RECT 3387.540 2095.770 3387.800 2096.090 ;
        RECT 3387.600 2092.205 3387.740 2095.770 ;
      LAYER met2 ;
        RECT 3388.000 2092.605 3583.075 2116.505 ;
      LAYER met2 ;
        RECT 3387.530 2091.835 3387.810 2092.205 ;
      LAYER met2 ;
        RECT 3388.000 2089.105 3389.920 2091.105 ;
        RECT 3390.035 2066.610 3583.075 2092.605 ;
        RECT 3388.000 2042.710 3583.075 2066.610 ;
      LAYER met2 ;
        RECT 213.540 2024.370 213.800 2024.690 ;
        RECT 213.600 2001.070 213.740 2024.370 ;
        RECT 213.140 2000.930 213.740 2001.070 ;
        RECT 212.620 1845.190 212.880 1845.510 ;
        RECT 208.940 1788.070 209.200 1788.390 ;
        RECT 212.160 1788.070 212.420 1788.390 ;
      LAYER met2 ;
        RECT 0.000 1787.165 208.285 1788.005 ;
        RECT 0.000 1785.245 208.565 1787.165 ;
        RECT 0.000 1784.405 208.285 1785.245 ;
        RECT 0.000 1782.025 208.565 1784.405 ;
        RECT 0.000 1781.185 208.285 1782.025 ;
        RECT 0.000 1778.805 208.565 1781.185 ;
        RECT 0.000 1777.965 208.285 1778.805 ;
        RECT 0.000 1776.045 208.565 1777.965 ;
        RECT 0.000 1775.205 208.285 1776.045 ;
        RECT 0.000 1774.210 208.565 1775.205 ;
        RECT 0.000 1635.865 208.565 1636.915 ;
        RECT 0.000 1635.025 208.285 1635.865 ;
      LAYER met2 ;
        RECT 208.565 1635.515 210.965 1635.585 ;
        RECT 208.565 1635.375 211.440 1635.515 ;
        RECT 208.565 1635.305 210.965 1635.375 ;
      LAYER met2 ;
        RECT 0.000 1632.645 208.565 1635.025 ;
        RECT 0.000 1631.805 208.285 1632.645 ;
        RECT 0.000 1629.425 208.565 1631.805 ;
        RECT 0.000 1628.585 208.285 1629.425 ;
      LAYER met2 ;
        RECT 208.565 1628.865 210.965 1629.145 ;
      LAYER met2 ;
        RECT 0.000 1626.665 208.565 1628.585 ;
      LAYER met2 ;
        RECT 208.940 1628.270 209.200 1628.590 ;
      LAYER met2 ;
        RECT 0.000 1625.825 208.285 1626.665 ;
      LAYER met2 ;
        RECT 209.000 1626.385 209.140 1628.270 ;
        RECT 208.565 1626.105 210.965 1626.385 ;
      LAYER met2 ;
        RECT 0.000 1623.445 208.565 1625.825 ;
        RECT 0.000 1622.605 208.285 1623.445 ;
        RECT 0.000 1620.225 208.565 1622.605 ;
        RECT 0.000 1619.385 208.285 1620.225 ;
        RECT 0.000 1617.465 208.565 1619.385 ;
        RECT 0.000 1616.625 208.285 1617.465 ;
      LAYER met2 ;
        RECT 208.565 1616.905 210.965 1617.185 ;
      LAYER met2 ;
        RECT 0.000 1614.245 208.565 1616.625 ;
        RECT 0.000 1613.405 208.285 1614.245 ;
        RECT 0.000 1611.025 208.565 1613.405 ;
        RECT 0.000 1610.185 208.285 1611.025 ;
        RECT 0.000 1608.265 208.565 1610.185 ;
        RECT 0.000 1607.425 208.285 1608.265 ;
        RECT 0.000 1605.045 208.565 1607.425 ;
        RECT 0.000 1604.205 208.285 1605.045 ;
        RECT 0.000 1601.825 208.565 1604.205 ;
        RECT 0.000 1600.985 208.285 1601.825 ;
        RECT 0.000 1599.065 208.565 1600.985 ;
        RECT 0.000 1598.225 208.285 1599.065 ;
        RECT 0.000 1595.845 208.565 1598.225 ;
        RECT 0.000 1595.005 208.285 1595.845 ;
      LAYER met2 ;
        RECT 208.565 1595.495 210.965 1595.565 ;
        RECT 211.300 1595.495 211.440 1635.375 ;
        RECT 212.680 1628.590 212.820 1845.190 ;
        RECT 213.140 1806.750 213.280 2000.930 ;
      LAYER met2 ;
        RECT 3379.435 1898.795 3588.000 1899.790 ;
        RECT 3379.715 1897.955 3588.000 1898.795 ;
        RECT 3379.435 1896.035 3588.000 1897.955 ;
        RECT 3379.715 1895.195 3588.000 1896.035 ;
        RECT 3379.435 1892.815 3588.000 1895.195 ;
        RECT 3379.715 1891.975 3588.000 1892.815 ;
        RECT 3379.435 1889.595 3588.000 1891.975 ;
        RECT 3379.715 1888.755 3588.000 1889.595 ;
        RECT 3379.435 1886.835 3588.000 1888.755 ;
        RECT 3379.715 1885.995 3588.000 1886.835 ;
        RECT 3379.435 1883.615 3588.000 1885.995 ;
      LAYER met2 ;
        RECT 3377.035 1883.260 3379.435 1883.335 ;
        RECT 3377.020 1883.055 3379.435 1883.260 ;
        RECT 3377.020 1880.870 3377.160 1883.055 ;
      LAYER met2 ;
        RECT 3379.715 1882.775 3588.000 1883.615 ;
      LAYER met2 ;
        RECT 3369.600 1880.550 3369.860 1880.870 ;
        RECT 3376.960 1880.550 3377.220 1880.870 ;
        RECT 3368.680 1865.250 3368.940 1865.570 ;
        RECT 213.080 1806.430 213.340 1806.750 ;
        RECT 212.620 1628.270 212.880 1628.590 ;
        RECT 212.680 1614.670 212.820 1628.270 ;
        RECT 208.565 1595.355 211.440 1595.495 ;
        RECT 212.220 1614.530 212.820 1614.670 ;
        RECT 208.565 1595.285 210.965 1595.355 ;
      LAYER met2 ;
        RECT 0.000 1592.625 208.565 1595.005 ;
        RECT 0.000 1591.785 208.285 1592.625 ;
        RECT 0.000 1589.405 208.565 1591.785 ;
        RECT 0.000 1588.565 208.285 1589.405 ;
      LAYER met2 ;
        RECT 208.565 1588.845 210.965 1589.125 ;
      LAYER met2 ;
        RECT 0.000 1586.645 208.565 1588.565 ;
      LAYER met2 ;
        RECT 209.000 1587.110 209.140 1588.845 ;
        RECT 208.940 1586.790 209.200 1587.110 ;
      LAYER met2 ;
        RECT 0.000 1585.805 208.285 1586.645 ;
        RECT 0.000 1583.425 208.565 1585.805 ;
        RECT 0.000 1582.585 208.285 1583.425 ;
        RECT 0.000 1580.205 208.565 1582.585 ;
        RECT 0.000 1579.365 208.285 1580.205 ;
        RECT 0.000 1577.445 208.565 1579.365 ;
        RECT 0.000 1576.605 208.285 1577.445 ;
        RECT 0.000 1574.225 208.565 1576.605 ;
        RECT 0.000 1573.385 208.285 1574.225 ;
      LAYER met2 ;
        RECT 208.565 1573.665 210.965 1573.945 ;
      LAYER met2 ;
        RECT 0.000 1571.005 208.565 1573.385 ;
      LAYER met2 ;
        RECT 209.000 1571.470 209.140 1573.665 ;
        RECT 208.940 1571.150 209.200 1571.470 ;
      LAYER met2 ;
        RECT 0.000 1570.165 208.285 1571.005 ;
        RECT 0.000 1568.245 208.565 1570.165 ;
        RECT 0.000 1567.405 208.285 1568.245 ;
        RECT 0.000 1565.025 208.565 1567.405 ;
      LAYER met2 ;
        RECT 212.220 1565.090 212.360 1614.530 ;
        RECT 213.140 1587.110 213.280 1806.430 ;
        RECT 213.540 1788.070 213.800 1788.390 ;
        RECT 213.080 1586.790 213.340 1587.110 ;
        RECT 212.620 1571.150 212.880 1571.470 ;
      LAYER met2 ;
        RECT 0.000 1564.185 208.285 1565.025 ;
      LAYER met2 ;
        RECT 211.300 1564.950 212.360 1565.090 ;
      LAYER met2 ;
        RECT 0.000 1561.805 208.565 1564.185 ;
        RECT 0.000 1560.965 208.285 1561.805 ;
        RECT 0.000 1559.045 208.565 1560.965 ;
        RECT 0.000 1558.205 208.285 1559.045 ;
        RECT 0.000 1557.210 208.565 1558.205 ;
        RECT 0.000 1419.865 208.565 1420.915 ;
      LAYER met2 ;
        RECT 211.300 1420.250 211.440 1564.950 ;
        RECT 211.300 1420.110 212.360 1420.250 ;
      LAYER met2 ;
        RECT 0.000 1419.025 208.285 1419.865 ;
      LAYER met2 ;
        RECT 208.565 1419.570 210.965 1419.585 ;
        RECT 208.565 1419.430 211.440 1419.570 ;
        RECT 208.565 1419.305 210.965 1419.430 ;
      LAYER met2 ;
        RECT 0.000 1416.645 208.565 1419.025 ;
        RECT 0.000 1415.805 208.285 1416.645 ;
        RECT 0.000 1413.425 208.565 1415.805 ;
        RECT 0.000 1412.585 208.285 1413.425 ;
      LAYER met2 ;
        RECT 208.565 1412.865 210.965 1413.145 ;
      LAYER met2 ;
        RECT 0.000 1410.665 208.565 1412.585 ;
        RECT 0.000 1409.825 208.285 1410.665 ;
      LAYER met2 ;
        RECT 208.565 1410.105 210.965 1410.385 ;
      LAYER met2 ;
        RECT 0.000 1407.445 208.565 1409.825 ;
      LAYER met2 ;
        RECT 209.000 1407.930 209.140 1410.105 ;
        RECT 208.940 1407.610 209.200 1407.930 ;
      LAYER met2 ;
        RECT 0.000 1406.605 208.285 1407.445 ;
        RECT 0.000 1404.225 208.565 1406.605 ;
        RECT 0.000 1403.385 208.285 1404.225 ;
        RECT 0.000 1401.465 208.565 1403.385 ;
        RECT 0.000 1400.625 208.285 1401.465 ;
      LAYER met2 ;
        RECT 208.565 1400.905 210.965 1401.185 ;
      LAYER met2 ;
        RECT 0.000 1398.245 208.565 1400.625 ;
        RECT 0.000 1397.405 208.285 1398.245 ;
        RECT 0.000 1395.025 208.565 1397.405 ;
        RECT 0.000 1394.185 208.285 1395.025 ;
        RECT 0.000 1392.265 208.565 1394.185 ;
        RECT 0.000 1391.425 208.285 1392.265 ;
        RECT 0.000 1389.045 208.565 1391.425 ;
        RECT 0.000 1388.205 208.285 1389.045 ;
        RECT 0.000 1385.825 208.565 1388.205 ;
        RECT 0.000 1384.985 208.285 1385.825 ;
        RECT 0.000 1383.065 208.565 1384.985 ;
        RECT 0.000 1382.225 208.285 1383.065 ;
        RECT 0.000 1379.845 208.565 1382.225 ;
      LAYER met2 ;
        RECT 211.300 1380.130 211.440 1419.430 ;
        RECT 212.220 1407.930 212.360 1420.110 ;
        RECT 212.160 1407.610 212.420 1407.930 ;
        RECT 209.000 1379.990 211.440 1380.130 ;
      LAYER met2 ;
        RECT 0.000 1379.005 208.285 1379.845 ;
      LAYER met2 ;
        RECT 209.000 1379.565 209.140 1379.990 ;
        RECT 208.565 1379.285 210.965 1379.565 ;
      LAYER met2 ;
        RECT 0.000 1376.625 208.565 1379.005 ;
        RECT 0.000 1375.785 208.285 1376.625 ;
        RECT 0.000 1373.405 208.565 1375.785 ;
        RECT 0.000 1372.565 208.285 1373.405 ;
      LAYER met2 ;
        RECT 208.940 1373.270 209.200 1373.590 ;
        RECT 209.000 1373.125 209.140 1373.270 ;
        RECT 208.565 1372.845 210.965 1373.125 ;
      LAYER met2 ;
        RECT 0.000 1370.645 208.565 1372.565 ;
        RECT 0.000 1369.805 208.285 1370.645 ;
        RECT 0.000 1367.425 208.565 1369.805 ;
        RECT 0.000 1366.585 208.285 1367.425 ;
        RECT 0.000 1364.205 208.565 1366.585 ;
        RECT 0.000 1363.365 208.285 1364.205 ;
        RECT 0.000 1361.445 208.565 1363.365 ;
        RECT 0.000 1360.605 208.285 1361.445 ;
      LAYER met2 ;
        RECT 212.680 1360.670 212.820 1571.150 ;
        RECT 213.140 1373.590 213.280 1586.790 ;
        RECT 213.600 1571.470 213.740 1788.070 ;
        RECT 3368.740 1670.070 3368.880 1865.250 ;
        RECT 3368.680 1669.750 3368.940 1670.070 ;
        RECT 3369.660 1659.870 3369.800 1880.550 ;
      LAYER met2 ;
        RECT 3379.435 1880.395 3588.000 1882.775 ;
        RECT 3379.715 1879.555 3588.000 1880.395 ;
        RECT 3379.435 1877.635 3588.000 1879.555 ;
        RECT 3379.715 1876.795 3588.000 1877.635 ;
        RECT 3379.435 1874.415 3588.000 1876.795 ;
        RECT 3379.715 1873.575 3588.000 1874.415 ;
        RECT 3379.435 1871.195 3588.000 1873.575 ;
        RECT 3379.715 1870.355 3588.000 1871.195 ;
        RECT 3379.435 1868.435 3588.000 1870.355 ;
      LAYER met2 ;
        RECT 3377.035 1868.015 3379.435 1868.155 ;
        RECT 3377.020 1867.875 3379.435 1868.015 ;
        RECT 3377.020 1865.570 3377.160 1867.875 ;
      LAYER met2 ;
        RECT 3379.715 1867.595 3588.000 1868.435 ;
      LAYER met2 ;
        RECT 3376.960 1865.250 3377.220 1865.570 ;
      LAYER met2 ;
        RECT 3379.435 1865.215 3588.000 1867.595 ;
        RECT 3379.715 1864.375 3588.000 1865.215 ;
        RECT 3379.435 1861.995 3588.000 1864.375 ;
      LAYER met2 ;
        RECT 3377.035 1861.570 3379.435 1861.715 ;
        RECT 3376.560 1861.435 3379.435 1861.570 ;
        RECT 3376.560 1861.430 3377.090 1861.435 ;
        RECT 3370.060 1828.530 3370.320 1828.850 ;
        RECT 3367.300 1659.550 3367.560 1659.870 ;
        RECT 3369.600 1659.550 3369.860 1659.870 ;
        RECT 213.540 1571.150 213.800 1571.470 ;
        RECT 3367.360 1443.970 3367.500 1659.550 ;
        RECT 3367.760 1644.250 3368.020 1644.570 ;
        RECT 3367.300 1443.650 3367.560 1443.970 ;
        RECT 213.540 1407.610 213.800 1407.930 ;
        RECT 213.080 1373.270 213.340 1373.590 ;
      LAYER met2 ;
        RECT 0.000 1358.225 208.565 1360.605 ;
      LAYER met2 ;
        RECT 208.940 1360.350 209.200 1360.670 ;
        RECT 212.620 1360.350 212.880 1360.670 ;
      LAYER met2 ;
        RECT 0.000 1357.385 208.285 1358.225 ;
      LAYER met2 ;
        RECT 209.000 1357.945 209.140 1360.350 ;
        RECT 208.565 1357.665 210.965 1357.945 ;
      LAYER met2 ;
        RECT 0.000 1355.005 208.565 1357.385 ;
        RECT 0.000 1354.165 208.285 1355.005 ;
        RECT 0.000 1352.245 208.565 1354.165 ;
        RECT 0.000 1351.405 208.285 1352.245 ;
        RECT 0.000 1349.025 208.565 1351.405 ;
        RECT 0.000 1348.185 208.285 1349.025 ;
        RECT 0.000 1345.805 208.565 1348.185 ;
        RECT 0.000 1344.965 208.285 1345.805 ;
        RECT 0.000 1343.045 208.565 1344.965 ;
        RECT 0.000 1342.205 208.285 1343.045 ;
        RECT 0.000 1341.210 208.565 1342.205 ;
        RECT 0.000 1203.865 208.565 1204.915 ;
        RECT 0.000 1203.025 208.285 1203.865 ;
      LAYER met2 ;
        RECT 208.565 1203.515 210.965 1203.585 ;
        RECT 208.565 1203.375 211.440 1203.515 ;
        RECT 208.565 1203.305 210.965 1203.375 ;
      LAYER met2 ;
        RECT 0.000 1200.645 208.565 1203.025 ;
        RECT 0.000 1199.805 208.285 1200.645 ;
        RECT 0.000 1197.425 208.565 1199.805 ;
        RECT 0.000 1196.585 208.285 1197.425 ;
      LAYER met2 ;
        RECT 208.565 1196.865 210.965 1197.145 ;
      LAYER met2 ;
        RECT 0.000 1194.665 208.565 1196.585 ;
        RECT 0.000 1193.825 208.285 1194.665 ;
      LAYER met2 ;
        RECT 208.565 1194.105 210.965 1194.385 ;
      LAYER met2 ;
        RECT 0.000 1191.445 208.565 1193.825 ;
      LAYER met2 ;
        RECT 209.000 1191.690 209.140 1194.105 ;
      LAYER met2 ;
        RECT 0.000 1190.605 208.285 1191.445 ;
      LAYER met2 ;
        RECT 208.940 1191.370 209.200 1191.690 ;
      LAYER met2 ;
        RECT 0.000 1188.225 208.565 1190.605 ;
        RECT 0.000 1187.385 208.285 1188.225 ;
      LAYER met2 ;
        RECT 208.565 1187.665 210.965 1187.945 ;
      LAYER met2 ;
        RECT 0.000 1185.465 208.565 1187.385 ;
        RECT 0.000 1184.625 208.285 1185.465 ;
      LAYER met2 ;
        RECT 208.565 1184.905 210.965 1185.185 ;
      LAYER met2 ;
        RECT 0.000 1182.245 208.565 1184.625 ;
        RECT 0.000 1181.405 208.285 1182.245 ;
        RECT 0.000 1179.025 208.565 1181.405 ;
        RECT 0.000 1178.185 208.285 1179.025 ;
      LAYER met2 ;
        RECT 208.565 1178.465 210.965 1178.745 ;
      LAYER met2 ;
        RECT 0.000 1176.265 208.565 1178.185 ;
        RECT 0.000 1175.425 208.285 1176.265 ;
        RECT 0.000 1173.045 208.565 1175.425 ;
        RECT 0.000 1172.205 208.285 1173.045 ;
        RECT 0.000 1169.825 208.565 1172.205 ;
        RECT 0.000 1168.985 208.285 1169.825 ;
        RECT 0.000 1167.065 208.565 1168.985 ;
        RECT 0.000 1166.225 208.285 1167.065 ;
        RECT 0.000 1163.845 208.565 1166.225 ;
      LAYER met2 ;
        RECT 211.300 1163.890 211.440 1203.375 ;
        RECT 212.160 1191.370 212.420 1191.690 ;
      LAYER met2 ;
        RECT 0.000 1163.005 208.285 1163.845 ;
      LAYER met2 ;
        RECT 209.000 1163.750 211.440 1163.890 ;
        RECT 209.000 1163.565 209.140 1163.750 ;
        RECT 208.565 1163.285 210.965 1163.565 ;
      LAYER met2 ;
        RECT 0.000 1160.625 208.565 1163.005 ;
        RECT 0.000 1159.785 208.285 1160.625 ;
        RECT 0.000 1157.405 208.565 1159.785 ;
      LAYER met2 ;
        RECT 208.940 1159.410 209.200 1159.730 ;
      LAYER met2 ;
        RECT 0.000 1156.565 208.285 1157.405 ;
      LAYER met2 ;
        RECT 209.000 1157.125 209.140 1159.410 ;
        RECT 208.565 1156.845 210.965 1157.125 ;
      LAYER met2 ;
        RECT 0.000 1154.645 208.565 1156.565 ;
        RECT 0.000 1153.805 208.285 1154.645 ;
        RECT 0.000 1151.425 208.565 1153.805 ;
        RECT 0.000 1150.585 208.285 1151.425 ;
        RECT 0.000 1148.205 208.565 1150.585 ;
        RECT 0.000 1147.365 208.285 1148.205 ;
        RECT 0.000 1145.445 208.565 1147.365 ;
        RECT 0.000 1144.605 208.285 1145.445 ;
        RECT 0.000 1142.225 208.565 1144.605 ;
      LAYER met2 ;
        RECT 208.940 1144.110 209.200 1144.430 ;
      LAYER met2 ;
        RECT 0.000 1141.385 208.285 1142.225 ;
      LAYER met2 ;
        RECT 209.000 1141.945 209.140 1144.110 ;
        RECT 208.565 1141.665 210.965 1141.945 ;
      LAYER met2 ;
        RECT 0.000 1139.005 208.565 1141.385 ;
        RECT 0.000 1138.165 208.285 1139.005 ;
        RECT 0.000 1136.245 208.565 1138.165 ;
        RECT 0.000 1135.405 208.285 1136.245 ;
        RECT 0.000 1133.025 208.565 1135.405 ;
        RECT 0.000 1132.185 208.285 1133.025 ;
        RECT 0.000 1129.805 208.565 1132.185 ;
        RECT 0.000 1128.965 208.285 1129.805 ;
        RECT 0.000 1127.045 208.565 1128.965 ;
        RECT 0.000 1126.205 208.285 1127.045 ;
        RECT 0.000 1125.210 208.565 1126.205 ;
        RECT 0.000 987.865 208.565 988.915 ;
        RECT 0.000 987.025 208.285 987.865 ;
      LAYER met2 ;
        RECT 208.565 987.515 210.965 987.585 ;
        RECT 208.565 987.375 211.440 987.515 ;
        RECT 208.565 987.305 210.965 987.375 ;
      LAYER met2 ;
        RECT 0.000 984.645 208.565 987.025 ;
        RECT 0.000 983.805 208.285 984.645 ;
        RECT 0.000 981.425 208.565 983.805 ;
        RECT 0.000 980.585 208.285 981.425 ;
      LAYER met2 ;
        RECT 208.565 980.865 210.965 981.145 ;
      LAYER met2 ;
        RECT 0.000 978.665 208.565 980.585 ;
        RECT 0.000 977.825 208.285 978.665 ;
      LAYER met2 ;
        RECT 208.565 978.105 210.965 978.385 ;
      LAYER met2 ;
        RECT 0.000 975.445 208.565 977.825 ;
      LAYER met2 ;
        RECT 209.000 975.790 209.140 978.105 ;
        RECT 208.940 975.470 209.200 975.790 ;
      LAYER met2 ;
        RECT 0.000 974.605 208.285 975.445 ;
        RECT 0.000 972.225 208.565 974.605 ;
        RECT 0.000 971.385 208.285 972.225 ;
      LAYER met2 ;
        RECT 208.565 971.665 210.965 971.945 ;
      LAYER met2 ;
        RECT 0.000 969.465 208.565 971.385 ;
        RECT 0.000 968.625 208.285 969.465 ;
      LAYER met2 ;
        RECT 208.565 968.905 210.965 969.185 ;
      LAYER met2 ;
        RECT 0.000 966.245 208.565 968.625 ;
        RECT 0.000 965.405 208.285 966.245 ;
        RECT 0.000 963.025 208.565 965.405 ;
        RECT 0.000 962.185 208.285 963.025 ;
      LAYER met2 ;
        RECT 208.565 962.465 210.965 962.745 ;
      LAYER met2 ;
        RECT 0.000 960.265 208.565 962.185 ;
        RECT 0.000 959.425 208.285 960.265 ;
        RECT 0.000 957.045 208.565 959.425 ;
        RECT 0.000 956.205 208.285 957.045 ;
        RECT 0.000 953.825 208.565 956.205 ;
        RECT 0.000 952.985 208.285 953.825 ;
        RECT 0.000 951.065 208.565 952.985 ;
        RECT 0.000 950.225 208.285 951.065 ;
        RECT 0.000 947.845 208.565 950.225 ;
        RECT 0.000 947.005 208.285 947.845 ;
      LAYER met2 ;
        RECT 211.300 947.650 211.440 987.375 ;
        RECT 212.220 975.790 212.360 1191.370 ;
        RECT 212.680 1144.430 212.820 1360.350 ;
        RECT 213.140 1159.730 213.280 1373.270 ;
        RECT 213.600 1191.690 213.740 1407.610 ;
        RECT 3367.360 1218.890 3367.500 1443.650 ;
        RECT 3367.820 1426.630 3367.960 1644.250 ;
        RECT 3370.120 1612.610 3370.260 1828.530 ;
        RECT 3376.560 1821.625 3376.700 1861.430 ;
      LAYER met2 ;
        RECT 3379.715 1861.155 3588.000 1861.995 ;
        RECT 3379.435 1858.775 3588.000 1861.155 ;
        RECT 3379.715 1857.935 3588.000 1858.775 ;
        RECT 3379.435 1856.015 3588.000 1857.935 ;
        RECT 3379.715 1855.175 3588.000 1856.015 ;
        RECT 3379.435 1852.795 3588.000 1855.175 ;
        RECT 3379.715 1851.955 3588.000 1852.795 ;
        RECT 3379.435 1849.575 3588.000 1851.955 ;
        RECT 3379.715 1848.735 3588.000 1849.575 ;
        RECT 3379.435 1846.815 3588.000 1848.735 ;
      LAYER met2 ;
        RECT 3377.035 1846.255 3379.435 1846.535 ;
      LAYER met2 ;
        RECT 3379.715 1845.975 3588.000 1846.815 ;
        RECT 3379.435 1843.595 3588.000 1845.975 ;
        RECT 3379.715 1842.755 3588.000 1843.595 ;
        RECT 3379.435 1840.375 3588.000 1842.755 ;
      LAYER met2 ;
        RECT 3377.035 1839.815 3379.435 1840.095 ;
      LAYER met2 ;
        RECT 3379.715 1839.535 3588.000 1840.375 ;
        RECT 3379.435 1837.615 3588.000 1839.535 ;
      LAYER met2 ;
        RECT 3377.035 1837.055 3379.435 1837.335 ;
      LAYER met2 ;
        RECT 3379.715 1836.775 3588.000 1837.615 ;
        RECT 3379.435 1834.395 3588.000 1836.775 ;
        RECT 3379.715 1833.555 3588.000 1834.395 ;
        RECT 3379.435 1831.175 3588.000 1833.555 ;
      LAYER met2 ;
        RECT 3377.035 1830.755 3379.435 1830.895 ;
        RECT 3377.020 1830.615 3379.435 1830.755 ;
        RECT 3377.020 1828.850 3377.160 1830.615 ;
      LAYER met2 ;
        RECT 3379.715 1830.335 3588.000 1831.175 ;
      LAYER met2 ;
        RECT 3376.960 1828.530 3377.220 1828.850 ;
      LAYER met2 ;
        RECT 3379.435 1828.415 3588.000 1830.335 ;
      LAYER met2 ;
        RECT 3377.035 1827.855 3379.435 1828.135 ;
      LAYER met2 ;
        RECT 3379.715 1827.575 3588.000 1828.415 ;
        RECT 3379.435 1825.195 3588.000 1827.575 ;
        RECT 3379.715 1824.355 3588.000 1825.195 ;
        RECT 3379.435 1821.975 3588.000 1824.355 ;
      LAYER met2 ;
        RECT 3377.035 1821.625 3379.435 1821.695 ;
        RECT 3376.560 1821.485 3379.435 1821.625 ;
        RECT 3377.035 1821.415 3379.435 1821.485 ;
      LAYER met2 ;
        RECT 3379.715 1821.135 3588.000 1821.975 ;
        RECT 3379.435 1820.085 3588.000 1821.135 ;
        RECT 3379.435 1677.795 3588.000 1678.790 ;
        RECT 3379.715 1676.955 3588.000 1677.795 ;
        RECT 3379.435 1675.035 3588.000 1676.955 ;
        RECT 3379.715 1674.195 3588.000 1675.035 ;
        RECT 3379.435 1671.815 3588.000 1674.195 ;
        RECT 3379.715 1670.975 3588.000 1671.815 ;
      LAYER met2 ;
        RECT 3376.040 1669.750 3376.300 1670.070 ;
        RECT 3376.100 1644.570 3376.240 1669.750 ;
      LAYER met2 ;
        RECT 3379.435 1668.595 3588.000 1670.975 ;
        RECT 3379.715 1667.755 3588.000 1668.595 ;
        RECT 3379.435 1665.835 3588.000 1667.755 ;
        RECT 3379.715 1664.995 3588.000 1665.835 ;
        RECT 3379.435 1662.615 3588.000 1664.995 ;
      LAYER met2 ;
        RECT 3377.035 1662.260 3379.435 1662.335 ;
        RECT 3377.020 1662.055 3379.435 1662.260 ;
        RECT 3377.020 1659.870 3377.160 1662.055 ;
      LAYER met2 ;
        RECT 3379.715 1661.775 3588.000 1662.615 ;
      LAYER met2 ;
        RECT 3376.960 1659.550 3377.220 1659.870 ;
      LAYER met2 ;
        RECT 3379.435 1659.395 3588.000 1661.775 ;
        RECT 3379.715 1658.555 3588.000 1659.395 ;
        RECT 3379.435 1656.635 3588.000 1658.555 ;
        RECT 3379.715 1655.795 3588.000 1656.635 ;
        RECT 3379.435 1653.415 3588.000 1655.795 ;
        RECT 3379.715 1652.575 3588.000 1653.415 ;
        RECT 3379.435 1650.195 3588.000 1652.575 ;
        RECT 3379.715 1649.355 3588.000 1650.195 ;
        RECT 3379.435 1647.435 3588.000 1649.355 ;
      LAYER met2 ;
        RECT 3377.035 1647.015 3379.435 1647.155 ;
        RECT 3377.020 1646.875 3379.435 1647.015 ;
        RECT 3377.020 1644.570 3377.160 1646.875 ;
      LAYER met2 ;
        RECT 3379.715 1646.595 3588.000 1647.435 ;
      LAYER met2 ;
        RECT 3376.040 1644.250 3376.300 1644.570 ;
        RECT 3376.960 1644.250 3377.220 1644.570 ;
      LAYER met2 ;
        RECT 3379.435 1644.215 3588.000 1646.595 ;
        RECT 3379.715 1643.375 3588.000 1644.215 ;
        RECT 3379.435 1640.995 3588.000 1643.375 ;
      LAYER met2 ;
        RECT 3377.035 1640.570 3379.435 1640.715 ;
        RECT 3376.560 1640.435 3379.435 1640.570 ;
        RECT 3376.560 1640.430 3377.090 1640.435 ;
        RECT 3368.220 1612.290 3368.480 1612.610 ;
        RECT 3370.060 1612.290 3370.320 1612.610 ;
        RECT 3367.760 1426.310 3368.020 1426.630 ;
        RECT 3367.300 1218.570 3367.560 1218.890 ;
        RECT 213.540 1191.370 213.800 1191.690 ;
        RECT 213.080 1159.410 213.340 1159.730 ;
        RECT 213.140 1159.130 213.280 1159.410 ;
        RECT 213.140 1158.990 214.200 1159.130 ;
        RECT 212.620 1144.110 212.880 1144.430 ;
        RECT 212.680 1131.670 212.820 1144.110 ;
        RECT 212.680 1131.530 213.740 1131.670 ;
        RECT 212.160 975.470 212.420 975.790 ;
        RECT 208.540 947.510 211.440 947.650 ;
        RECT 208.540 947.425 210.965 947.510 ;
        RECT 208.565 947.285 210.965 947.425 ;
      LAYER met2 ;
        RECT 0.000 944.625 208.565 947.005 ;
        RECT 0.000 943.785 208.285 944.625 ;
        RECT 0.000 941.405 208.565 943.785 ;
      LAYER met2 ;
        RECT 208.940 943.510 209.200 943.830 ;
      LAYER met2 ;
        RECT 0.000 940.565 208.285 941.405 ;
      LAYER met2 ;
        RECT 209.000 941.125 209.140 943.510 ;
        RECT 208.565 940.845 210.965 941.125 ;
      LAYER met2 ;
        RECT 0.000 938.645 208.565 940.565 ;
        RECT 0.000 937.805 208.285 938.645 ;
        RECT 0.000 935.425 208.565 937.805 ;
        RECT 0.000 934.585 208.285 935.425 ;
        RECT 0.000 932.205 208.565 934.585 ;
        RECT 0.000 931.365 208.285 932.205 ;
        RECT 0.000 929.445 208.565 931.365 ;
        RECT 0.000 928.605 208.285 929.445 ;
        RECT 0.000 926.225 208.565 928.605 ;
      LAYER met2 ;
        RECT 208.940 928.210 209.200 928.530 ;
      LAYER met2 ;
        RECT 0.000 925.385 208.285 926.225 ;
      LAYER met2 ;
        RECT 209.000 925.945 209.140 928.210 ;
        RECT 208.565 925.665 210.965 925.945 ;
      LAYER met2 ;
        RECT 0.000 923.005 208.565 925.385 ;
        RECT 0.000 922.165 208.285 923.005 ;
        RECT 0.000 920.245 208.565 922.165 ;
      LAYER met2 ;
        RECT 211.240 921.750 211.500 922.070 ;
      LAYER met2 ;
        RECT 0.000 919.405 208.285 920.245 ;
        RECT 0.000 917.025 208.565 919.405 ;
        RECT 0.000 916.185 208.285 917.025 ;
        RECT 0.000 913.805 208.565 916.185 ;
        RECT 0.000 912.965 208.285 913.805 ;
        RECT 0.000 911.045 208.565 912.965 ;
        RECT 0.000 910.205 208.285 911.045 ;
        RECT 0.000 909.210 208.565 910.205 ;
        RECT 4.925 601.390 200.000 625.290 ;
        RECT 4.925 575.395 197.965 601.390 ;
        RECT 198.080 576.895 200.000 578.895 ;
        RECT 4.925 551.495 200.000 575.395 ;
        RECT 4.925 551.265 197.965 551.495 ;
        RECT 153.765 415.000 158.415 426.140 ;
        RECT 159.640 415.245 163.510 426.195 ;
        RECT 3.570 414.700 197.965 415.000 ;
        RECT 3.570 394.095 198.000 414.700 ;
      LAYER met2 ;
        RECT 198.350 400.675 198.630 401.045 ;
      LAYER met2 ;
        RECT 3.570 393.535 197.965 394.095 ;
        RECT 3.570 360.925 198.000 393.535 ;
      LAYER met2 ;
        RECT 198.420 391.525 198.560 400.675 ;
        RECT 198.350 391.155 198.630 391.525 ;
      LAYER met2 ;
        RECT 3.570 360.495 197.965 360.925 ;
        RECT 3.570 340.500 198.000 360.495 ;
        RECT 3.570 340.490 197.965 340.500 ;
      LAYER met2 ;
        RECT 211.300 228.470 211.440 921.750 ;
        RECT 212.220 530.390 212.360 975.470 ;
        RECT 212.620 943.510 212.880 943.830 ;
        RECT 212.680 607.570 212.820 943.510 ;
        RECT 213.600 928.530 213.740 1131.530 ;
        RECT 214.060 943.830 214.200 1158.990 ;
        RECT 3367.360 995.850 3367.500 1218.570 ;
        RECT 3367.820 1201.550 3367.960 1426.310 ;
        RECT 3368.280 1386.850 3368.420 1612.290 ;
        RECT 3376.560 1600.625 3376.700 1640.430 ;
      LAYER met2 ;
        RECT 3379.715 1640.155 3588.000 1640.995 ;
        RECT 3379.435 1637.775 3588.000 1640.155 ;
        RECT 3379.715 1636.935 3588.000 1637.775 ;
        RECT 3379.435 1635.015 3588.000 1636.935 ;
        RECT 3379.715 1634.175 3588.000 1635.015 ;
        RECT 3379.435 1631.795 3588.000 1634.175 ;
        RECT 3379.715 1630.955 3588.000 1631.795 ;
        RECT 3379.435 1628.575 3588.000 1630.955 ;
        RECT 3379.715 1627.735 3588.000 1628.575 ;
        RECT 3379.435 1625.815 3588.000 1627.735 ;
      LAYER met2 ;
        RECT 3377.035 1625.255 3379.435 1625.535 ;
      LAYER met2 ;
        RECT 3379.715 1624.975 3588.000 1625.815 ;
        RECT 3379.435 1622.595 3588.000 1624.975 ;
        RECT 3379.715 1621.755 3588.000 1622.595 ;
        RECT 3379.435 1619.375 3588.000 1621.755 ;
      LAYER met2 ;
        RECT 3377.035 1618.815 3379.435 1619.095 ;
      LAYER met2 ;
        RECT 3379.715 1618.535 3588.000 1619.375 ;
        RECT 3379.435 1616.615 3588.000 1618.535 ;
      LAYER met2 ;
        RECT 3377.035 1616.055 3379.435 1616.335 ;
      LAYER met2 ;
        RECT 3379.715 1615.775 3588.000 1616.615 ;
        RECT 3379.435 1613.395 3588.000 1615.775 ;
      LAYER met2 ;
        RECT 3376.960 1612.290 3377.220 1612.610 ;
      LAYER met2 ;
        RECT 3379.715 1612.555 3588.000 1613.395 ;
      LAYER met2 ;
        RECT 3377.020 1609.895 3377.160 1612.290 ;
      LAYER met2 ;
        RECT 3379.435 1610.175 3588.000 1612.555 ;
      LAYER met2 ;
        RECT 3377.020 1609.755 3379.435 1609.895 ;
        RECT 3377.035 1609.615 3379.435 1609.755 ;
      LAYER met2 ;
        RECT 3379.715 1609.335 3588.000 1610.175 ;
        RECT 3379.435 1607.415 3588.000 1609.335 ;
      LAYER met2 ;
        RECT 3377.035 1606.855 3379.435 1607.135 ;
      LAYER met2 ;
        RECT 3379.715 1606.575 3588.000 1607.415 ;
        RECT 3379.435 1604.195 3588.000 1606.575 ;
        RECT 3379.715 1603.355 3588.000 1604.195 ;
        RECT 3379.435 1600.975 3588.000 1603.355 ;
      LAYER met2 ;
        RECT 3377.035 1600.625 3379.435 1600.695 ;
        RECT 3376.560 1600.485 3379.435 1600.625 ;
        RECT 3377.035 1600.415 3379.435 1600.485 ;
      LAYER met2 ;
        RECT 3379.715 1600.135 3588.000 1600.975 ;
        RECT 3379.435 1599.085 3588.000 1600.135 ;
        RECT 3379.435 1456.795 3588.000 1457.790 ;
        RECT 3379.715 1455.955 3588.000 1456.795 ;
        RECT 3379.435 1454.035 3588.000 1455.955 ;
        RECT 3379.715 1453.195 3588.000 1454.035 ;
        RECT 3379.435 1450.815 3588.000 1453.195 ;
        RECT 3379.715 1449.975 3588.000 1450.815 ;
        RECT 3379.435 1447.595 3588.000 1449.975 ;
        RECT 3379.715 1446.755 3588.000 1447.595 ;
        RECT 3379.435 1444.835 3588.000 1446.755 ;
        RECT 3379.715 1443.995 3588.000 1444.835 ;
      LAYER met2 ;
        RECT 3376.960 1443.650 3377.220 1443.970 ;
        RECT 3377.020 1441.335 3377.160 1443.650 ;
      LAYER met2 ;
        RECT 3379.435 1441.615 3588.000 1443.995 ;
      LAYER met2 ;
        RECT 3377.020 1441.260 3379.435 1441.335 ;
        RECT 3377.035 1441.055 3379.435 1441.260 ;
      LAYER met2 ;
        RECT 3379.715 1440.775 3588.000 1441.615 ;
        RECT 3379.435 1438.395 3588.000 1440.775 ;
        RECT 3379.715 1437.555 3588.000 1438.395 ;
        RECT 3379.435 1435.635 3588.000 1437.555 ;
        RECT 3379.715 1434.795 3588.000 1435.635 ;
        RECT 3379.435 1432.415 3588.000 1434.795 ;
        RECT 3379.715 1431.575 3588.000 1432.415 ;
        RECT 3379.435 1429.195 3588.000 1431.575 ;
        RECT 3379.715 1428.355 3588.000 1429.195 ;
      LAYER met2 ;
        RECT 3376.960 1426.310 3377.220 1426.630 ;
      LAYER met2 ;
        RECT 3379.435 1426.435 3588.000 1428.355 ;
      LAYER met2 ;
        RECT 3377.020 1426.155 3377.160 1426.310 ;
        RECT 3377.020 1426.015 3379.435 1426.155 ;
        RECT 3377.035 1425.875 3379.435 1426.015 ;
      LAYER met2 ;
        RECT 3379.715 1425.595 3588.000 1426.435 ;
        RECT 3379.435 1423.215 3588.000 1425.595 ;
        RECT 3379.715 1422.375 3588.000 1423.215 ;
        RECT 3379.435 1419.995 3588.000 1422.375 ;
      LAYER met2 ;
        RECT 3377.035 1419.570 3379.435 1419.715 ;
        RECT 3376.560 1419.435 3379.435 1419.570 ;
        RECT 3376.560 1419.430 3377.090 1419.435 ;
        RECT 3368.220 1386.530 3368.480 1386.850 ;
        RECT 3367.760 1201.230 3368.020 1201.550 ;
        RECT 3367.300 995.530 3367.560 995.850 ;
        RECT 214.000 943.510 214.260 943.830 ;
        RECT 213.540 928.210 213.800 928.530 ;
        RECT 213.600 922.070 213.740 928.210 ;
        RECT 213.540 921.750 213.800 922.070 ;
        RECT 3367.360 779.950 3367.500 995.530 ;
        RECT 3367.820 985.310 3367.960 1201.230 ;
        RECT 3368.280 1169.590 3368.420 1386.530 ;
        RECT 3376.560 1379.625 3376.700 1419.430 ;
      LAYER met2 ;
        RECT 3379.715 1419.155 3588.000 1419.995 ;
        RECT 3379.435 1416.775 3588.000 1419.155 ;
        RECT 3379.715 1415.935 3588.000 1416.775 ;
        RECT 3379.435 1414.015 3588.000 1415.935 ;
        RECT 3379.715 1413.175 3588.000 1414.015 ;
        RECT 3379.435 1410.795 3588.000 1413.175 ;
        RECT 3379.715 1409.955 3588.000 1410.795 ;
        RECT 3379.435 1407.575 3588.000 1409.955 ;
        RECT 3379.715 1406.735 3588.000 1407.575 ;
        RECT 3379.435 1404.815 3588.000 1406.735 ;
      LAYER met2 ;
        RECT 3377.035 1404.255 3379.435 1404.535 ;
      LAYER met2 ;
        RECT 3379.715 1403.975 3588.000 1404.815 ;
        RECT 3379.435 1401.595 3588.000 1403.975 ;
        RECT 3379.715 1400.755 3588.000 1401.595 ;
        RECT 3379.435 1398.375 3588.000 1400.755 ;
      LAYER met2 ;
        RECT 3377.035 1397.815 3379.435 1398.095 ;
      LAYER met2 ;
        RECT 3379.715 1397.535 3588.000 1398.375 ;
        RECT 3379.435 1395.615 3588.000 1397.535 ;
      LAYER met2 ;
        RECT 3377.035 1395.055 3379.435 1395.335 ;
      LAYER met2 ;
        RECT 3379.715 1394.775 3588.000 1395.615 ;
        RECT 3379.435 1392.395 3588.000 1394.775 ;
        RECT 3379.715 1391.555 3588.000 1392.395 ;
        RECT 3379.435 1389.175 3588.000 1391.555 ;
      LAYER met2 ;
        RECT 3377.035 1388.755 3379.435 1388.895 ;
        RECT 3377.020 1388.615 3379.435 1388.755 ;
        RECT 3377.020 1386.850 3377.160 1388.615 ;
      LAYER met2 ;
        RECT 3379.715 1388.335 3588.000 1389.175 ;
      LAYER met2 ;
        RECT 3376.960 1386.530 3377.220 1386.850 ;
      LAYER met2 ;
        RECT 3379.435 1386.415 3588.000 1388.335 ;
      LAYER met2 ;
        RECT 3377.035 1385.855 3379.435 1386.135 ;
      LAYER met2 ;
        RECT 3379.715 1385.575 3588.000 1386.415 ;
        RECT 3379.435 1383.195 3588.000 1385.575 ;
        RECT 3379.715 1382.355 3588.000 1383.195 ;
        RECT 3379.435 1379.975 3588.000 1382.355 ;
      LAYER met2 ;
        RECT 3377.035 1379.625 3379.435 1379.695 ;
        RECT 3376.560 1379.485 3379.435 1379.625 ;
        RECT 3377.035 1379.415 3379.435 1379.485 ;
      LAYER met2 ;
        RECT 3379.715 1379.135 3588.000 1379.975 ;
        RECT 3379.435 1378.085 3588.000 1379.135 ;
        RECT 3379.435 1234.795 3588.000 1235.790 ;
        RECT 3379.715 1233.955 3588.000 1234.795 ;
        RECT 3379.435 1232.035 3588.000 1233.955 ;
        RECT 3379.715 1231.195 3588.000 1232.035 ;
        RECT 3379.435 1228.815 3588.000 1231.195 ;
        RECT 3379.715 1227.975 3588.000 1228.815 ;
        RECT 3379.435 1225.595 3588.000 1227.975 ;
        RECT 3379.715 1224.755 3588.000 1225.595 ;
        RECT 3379.435 1222.835 3588.000 1224.755 ;
        RECT 3379.715 1221.995 3588.000 1222.835 ;
        RECT 3379.435 1219.615 3588.000 1221.995 ;
      LAYER met2 ;
        RECT 3377.035 1219.195 3379.435 1219.335 ;
        RECT 3377.020 1219.055 3379.435 1219.195 ;
        RECT 3377.020 1218.890 3377.160 1219.055 ;
        RECT 3376.960 1218.570 3377.220 1218.890 ;
      LAYER met2 ;
        RECT 3379.715 1218.775 3588.000 1219.615 ;
        RECT 3379.435 1216.395 3588.000 1218.775 ;
        RECT 3379.715 1215.555 3588.000 1216.395 ;
        RECT 3379.435 1213.635 3588.000 1215.555 ;
        RECT 3379.715 1212.795 3588.000 1213.635 ;
        RECT 3379.435 1210.415 3588.000 1212.795 ;
        RECT 3379.715 1209.575 3588.000 1210.415 ;
        RECT 3379.435 1207.195 3588.000 1209.575 ;
        RECT 3379.715 1206.355 3588.000 1207.195 ;
        RECT 3379.435 1204.435 3588.000 1206.355 ;
      LAYER met2 ;
        RECT 3377.035 1203.940 3379.435 1204.155 ;
        RECT 3377.020 1203.875 3379.435 1203.940 ;
        RECT 3377.020 1201.550 3377.160 1203.875 ;
      LAYER met2 ;
        RECT 3379.715 1203.595 3588.000 1204.435 ;
      LAYER met2 ;
        RECT 3376.960 1201.230 3377.220 1201.550 ;
      LAYER met2 ;
        RECT 3379.435 1201.215 3588.000 1203.595 ;
        RECT 3379.715 1200.375 3588.000 1201.215 ;
        RECT 3379.435 1197.995 3588.000 1200.375 ;
      LAYER met2 ;
        RECT 3377.035 1197.645 3379.435 1197.715 ;
        RECT 3376.560 1197.505 3379.435 1197.645 ;
        RECT 3368.220 1169.270 3368.480 1169.590 ;
        RECT 3367.760 984.990 3368.020 985.310 ;
        RECT 3367.300 779.630 3367.560 779.950 ;
        RECT 3367.820 764.310 3367.960 984.990 ;
        RECT 3368.280 946.550 3368.420 1169.270 ;
        RECT 3376.560 1157.625 3376.700 1197.505 ;
        RECT 3377.035 1197.435 3379.435 1197.505 ;
      LAYER met2 ;
        RECT 3379.715 1197.155 3588.000 1197.995 ;
        RECT 3379.435 1194.775 3588.000 1197.155 ;
        RECT 3379.715 1193.935 3588.000 1194.775 ;
        RECT 3379.435 1192.015 3588.000 1193.935 ;
        RECT 3379.715 1191.175 3588.000 1192.015 ;
        RECT 3379.435 1188.795 3588.000 1191.175 ;
        RECT 3379.715 1187.955 3588.000 1188.795 ;
        RECT 3379.435 1185.575 3588.000 1187.955 ;
        RECT 3379.715 1184.735 3588.000 1185.575 ;
        RECT 3379.435 1182.815 3588.000 1184.735 ;
      LAYER met2 ;
        RECT 3377.035 1182.255 3379.435 1182.535 ;
      LAYER met2 ;
        RECT 3379.715 1181.975 3588.000 1182.815 ;
        RECT 3379.435 1179.595 3588.000 1181.975 ;
        RECT 3379.715 1178.755 3588.000 1179.595 ;
        RECT 3379.435 1176.375 3588.000 1178.755 ;
      LAYER met2 ;
        RECT 3377.035 1175.815 3379.435 1176.095 ;
      LAYER met2 ;
        RECT 3379.715 1175.535 3588.000 1176.375 ;
        RECT 3379.435 1173.615 3588.000 1175.535 ;
      LAYER met2 ;
        RECT 3377.035 1173.055 3379.435 1173.335 ;
      LAYER met2 ;
        RECT 3379.715 1172.775 3588.000 1173.615 ;
        RECT 3379.435 1170.395 3588.000 1172.775 ;
      LAYER met2 ;
        RECT 3376.960 1169.270 3377.220 1169.590 ;
      LAYER met2 ;
        RECT 3379.715 1169.555 3588.000 1170.395 ;
      LAYER met2 ;
        RECT 3377.020 1166.895 3377.160 1169.270 ;
      LAYER met2 ;
        RECT 3379.435 1167.175 3588.000 1169.555 ;
      LAYER met2 ;
        RECT 3377.020 1166.755 3379.435 1166.895 ;
        RECT 3377.035 1166.615 3379.435 1166.755 ;
      LAYER met2 ;
        RECT 3379.715 1166.335 3588.000 1167.175 ;
        RECT 3379.435 1164.415 3588.000 1166.335 ;
      LAYER met2 ;
        RECT 3377.035 1163.855 3379.435 1164.135 ;
      LAYER met2 ;
        RECT 3379.715 1163.575 3588.000 1164.415 ;
        RECT 3379.435 1161.195 3588.000 1163.575 ;
        RECT 3379.715 1160.355 3588.000 1161.195 ;
        RECT 3379.435 1157.975 3588.000 1160.355 ;
      LAYER met2 ;
        RECT 3377.035 1157.625 3379.435 1157.695 ;
        RECT 3376.560 1157.485 3379.435 1157.625 ;
        RECT 3377.035 1157.415 3379.435 1157.485 ;
      LAYER met2 ;
        RECT 3379.715 1157.135 3588.000 1157.975 ;
        RECT 3379.435 1156.085 3588.000 1157.135 ;
        RECT 3379.435 1013.795 3588.000 1014.790 ;
        RECT 3379.715 1012.955 3588.000 1013.795 ;
        RECT 3379.435 1011.035 3588.000 1012.955 ;
        RECT 3379.715 1010.195 3588.000 1011.035 ;
        RECT 3379.435 1007.815 3588.000 1010.195 ;
        RECT 3379.715 1006.975 3588.000 1007.815 ;
        RECT 3379.435 1004.595 3588.000 1006.975 ;
        RECT 3379.715 1003.755 3588.000 1004.595 ;
        RECT 3379.435 1001.835 3588.000 1003.755 ;
        RECT 3379.715 1000.995 3588.000 1001.835 ;
        RECT 3379.435 998.615 3588.000 1000.995 ;
      LAYER met2 ;
        RECT 3377.035 998.195 3379.435 998.335 ;
        RECT 3377.020 998.055 3379.435 998.195 ;
        RECT 3377.020 995.850 3377.160 998.055 ;
      LAYER met2 ;
        RECT 3379.715 997.775 3588.000 998.615 ;
      LAYER met2 ;
        RECT 3376.960 995.530 3377.220 995.850 ;
      LAYER met2 ;
        RECT 3379.435 995.395 3588.000 997.775 ;
        RECT 3379.715 994.555 3588.000 995.395 ;
        RECT 3379.435 992.635 3588.000 994.555 ;
        RECT 3379.715 991.795 3588.000 992.635 ;
        RECT 3379.435 989.415 3588.000 991.795 ;
        RECT 3379.715 988.575 3588.000 989.415 ;
        RECT 3379.435 986.195 3588.000 988.575 ;
        RECT 3379.715 985.355 3588.000 986.195 ;
      LAYER met2 ;
        RECT 3376.960 984.990 3377.220 985.310 ;
        RECT 3377.020 983.155 3377.160 984.990 ;
      LAYER met2 ;
        RECT 3379.435 983.435 3588.000 985.355 ;
      LAYER met2 ;
        RECT 3377.020 982.940 3379.435 983.155 ;
        RECT 3377.035 982.875 3379.435 982.940 ;
      LAYER met2 ;
        RECT 3379.715 982.595 3588.000 983.435 ;
        RECT 3379.435 980.215 3588.000 982.595 ;
        RECT 3379.715 979.375 3588.000 980.215 ;
        RECT 3379.435 976.995 3588.000 979.375 ;
      LAYER met2 ;
        RECT 3377.035 976.645 3379.435 976.715 ;
        RECT 3376.560 976.505 3379.435 976.645 ;
        RECT 3368.220 946.230 3368.480 946.550 ;
        RECT 3367.760 763.990 3368.020 764.310 ;
        RECT 212.620 607.250 212.880 607.570 ;
        RECT 220.900 607.250 221.160 607.570 ;
        RECT 220.960 552.685 221.100 607.250 ;
        RECT 3367.300 557.610 3367.560 557.930 ;
        RECT 220.890 552.315 221.170 552.685 ;
        RECT 224.110 552.315 224.390 552.685 ;
        RECT 224.180 552.070 224.320 552.315 ;
        RECT 224.180 551.930 224.780 552.070 ;
        RECT 212.160 530.070 212.420 530.390 ;
        RECT 220.900 530.070 221.160 530.390 ;
        RECT 220.960 401.045 221.100 530.070 ;
        RECT 220.890 400.675 221.170 401.045 ;
        RECT 224.110 400.675 224.390 401.045 ;
        RECT 224.180 234.930 224.320 400.675 ;
        RECT 224.120 234.610 224.380 234.930 ;
        RECT 211.240 228.150 211.500 228.470 ;
        RECT 224.640 227.790 224.780 551.930 ;
        RECT 717.700 234.270 717.960 234.590 ;
        RECT 704.820 228.150 705.080 228.470 ;
        RECT 224.580 227.470 224.840 227.790 ;
        RECT 468.840 207.410 469.100 207.730 ;
        RECT 468.900 201.125 469.040 207.410 ;
        RECT 675.840 201.125 676.100 201.270 ;
        RECT 468.830 200.755 469.110 201.125 ;
        RECT 675.830 200.755 676.110 201.125 ;
        RECT 704.880 201.010 705.020 228.150 ;
        RECT 717.760 202.485 717.900 234.270 ;
        RECT 758.630 234.075 758.910 234.445 ;
        RECT 942.630 234.075 942.910 234.445 ;
        RECT 1004.280 234.270 1004.540 234.590 ;
        RECT 1281.200 234.270 1281.460 234.590 ;
        RECT 1488.660 234.270 1488.920 234.590 ;
        RECT 1547.080 234.270 1547.340 234.590 ;
        RECT 1762.820 234.270 1763.080 234.590 ;
        RECT 1821.240 234.270 1821.500 234.590 ;
        RECT 2036.980 234.270 2037.240 234.590 ;
        RECT 2095.400 234.270 2095.660 234.590 ;
        RECT 2310.680 234.270 2310.940 234.590 ;
        RECT 2369.100 234.270 2369.360 234.590 ;
        RECT 2584.840 234.270 2585.100 234.590 ;
        RECT 731.500 209.110 731.760 209.430 ;
        RECT 717.690 202.115 717.970 202.485 ;
        RECT 717.700 201.125 717.960 201.270 ;
        RECT 704.880 200.870 705.180 201.010 ;
        RECT 705.040 200.590 705.180 200.870 ;
        RECT 715.390 200.755 715.670 201.125 ;
        RECT 717.690 200.755 717.970 201.125 ;
        RECT 715.420 200.590 715.560 200.755 ;
        RECT 731.560 200.590 731.700 209.110 ;
        RECT 758.700 202.485 758.840 234.075 ;
        RECT 933.440 227.810 933.700 228.130 ;
        RECT 933.500 210.965 933.640 227.810 ;
        RECT 942.700 222.010 942.840 234.075 ;
        RECT 973.460 227.810 973.720 228.130 ;
        RECT 942.640 221.690 942.900 222.010 ;
        RECT 964.260 221.690 964.520 222.010 ;
        RECT 942.700 210.965 942.840 221.690 ;
        RECT 964.320 210.965 964.460 221.690 ;
        RECT 973.520 210.965 973.660 227.810 ;
        RECT 979.900 227.470 980.160 227.790 ;
        RECT 979.960 221.670 980.100 227.470 ;
        RECT 979.900 221.350 980.160 221.670 ;
        RECT 979.960 210.965 980.100 221.350 ;
        RECT 1004.340 210.965 1004.480 234.270 ;
        RECT 1007.500 221.350 1007.760 221.670 ;
        RECT 1007.560 210.965 1007.700 221.350 ;
        RECT 933.415 208.565 933.695 210.965 ;
        RECT 939.855 208.565 940.135 210.965 ;
        RECT 942.615 208.565 942.895 210.965 ;
        RECT 945.835 209.170 946.115 210.965 ;
        RECT 946.320 209.450 946.580 209.770 ;
        RECT 946.380 209.170 946.520 209.450 ;
        RECT 945.835 209.030 946.520 209.170 ;
        RECT 945.835 208.565 946.115 209.030 ;
        RECT 949.055 208.565 949.335 210.965 ;
        RECT 951.815 208.565 952.095 210.965 ;
        RECT 955.035 209.170 955.315 210.965 ;
        RECT 955.520 209.450 955.780 209.770 ;
        RECT 955.580 209.170 955.720 209.450 ;
        RECT 955.035 209.030 955.720 209.170 ;
        RECT 955.035 208.565 955.315 209.030 ;
        RECT 958.255 208.565 958.535 210.965 ;
        RECT 961.015 209.170 961.295 210.965 ;
        RECT 961.500 209.450 961.760 209.770 ;
        RECT 961.560 209.170 961.700 209.450 ;
        RECT 961.015 209.030 961.700 209.170 ;
        RECT 961.015 208.565 961.295 209.030 ;
        RECT 964.235 208.565 964.515 210.965 ;
        RECT 967.455 209.170 967.735 210.965 ;
        RECT 967.940 209.450 968.200 209.770 ;
        RECT 968.000 209.170 968.140 209.450 ;
        RECT 967.455 209.030 968.140 209.170 ;
        RECT 967.455 208.565 967.735 209.030 ;
        RECT 973.435 208.565 973.715 210.965 ;
        RECT 979.875 208.565 980.155 210.965 ;
        RECT 982.200 209.450 982.460 209.770 ;
        RECT 982.260 209.170 982.400 209.450 ;
        RECT 982.635 209.170 982.915 210.965 ;
        RECT 985.855 209.170 986.135 210.965 ;
        RECT 989.075 209.170 989.355 210.965 ;
        RECT 991.835 209.170 992.115 210.965 ;
        RECT 992.320 209.450 992.580 209.770 ;
        RECT 992.380 209.170 992.520 209.450 ;
        RECT 995.055 209.170 995.335 210.965 ;
        RECT 1000.600 209.450 1000.860 209.770 ;
        RECT 982.260 209.030 992.520 209.170 ;
        RECT 994.680 209.090 995.335 209.170 ;
        RECT 994.620 209.030 995.335 209.090 ;
        RECT 1000.660 209.170 1000.800 209.450 ;
        RECT 1001.035 209.170 1001.315 210.965 ;
        RECT 1004.255 209.170 1004.535 210.965 ;
        RECT 1000.660 209.030 1004.535 209.170 ;
        RECT 982.635 208.565 982.915 209.030 ;
        RECT 985.855 208.565 986.135 209.030 ;
        RECT 989.075 208.565 989.355 209.030 ;
        RECT 991.835 208.565 992.115 209.030 ;
        RECT 994.620 208.770 994.880 209.030 ;
        RECT 995.055 208.565 995.335 209.030 ;
        RECT 1001.035 208.565 1001.315 209.030 ;
        RECT 1004.255 208.565 1004.535 209.030 ;
        RECT 1007.475 208.565 1007.755 210.965 ;
        RECT 1010.235 208.565 1010.515 210.965 ;
      LAYER met2 ;
        RECT 932.085 208.285 933.135 208.565 ;
        RECT 933.975 208.285 936.355 208.565 ;
        RECT 937.195 208.285 939.575 208.565 ;
        RECT 940.415 208.285 942.335 208.565 ;
        RECT 943.175 208.285 945.555 208.565 ;
        RECT 946.395 208.285 948.775 208.565 ;
        RECT 949.615 208.285 951.535 208.565 ;
        RECT 952.375 208.285 954.755 208.565 ;
        RECT 955.595 208.285 957.975 208.565 ;
        RECT 958.815 208.285 960.735 208.565 ;
        RECT 961.575 208.285 963.955 208.565 ;
        RECT 964.795 208.285 967.175 208.565 ;
        RECT 968.015 208.285 969.935 208.565 ;
        RECT 970.775 208.285 973.155 208.565 ;
        RECT 973.995 208.285 976.375 208.565 ;
        RECT 977.215 208.285 979.595 208.565 ;
        RECT 980.435 208.285 982.355 208.565 ;
        RECT 983.195 208.285 985.575 208.565 ;
        RECT 986.415 208.285 988.795 208.565 ;
        RECT 989.635 208.285 991.555 208.565 ;
        RECT 992.395 208.285 994.775 208.565 ;
        RECT 995.615 208.285 997.995 208.565 ;
        RECT 998.835 208.285 1000.755 208.565 ;
        RECT 1001.595 208.285 1003.975 208.565 ;
        RECT 1004.815 208.285 1007.195 208.565 ;
        RECT 1008.035 208.285 1009.955 208.565 ;
        RECT 1010.795 208.285 1011.790 208.565 ;
      LAYER met2 ;
        RECT 758.630 202.115 758.910 202.485 ;
        RECT 704.980 200.270 705.240 200.590 ;
        RECT 715.360 200.270 715.620 200.590 ;
        RECT 722.760 200.270 723.020 200.590 ;
        RECT 731.500 200.270 731.760 200.590 ;
        RECT 705.040 200.000 705.180 200.270 ;
        RECT 715.420 200.000 715.560 200.270 ;
        RECT 722.820 200.000 722.960 200.270 ;
      LAYER met2 ;
        RECT 394.710 197.965 418.610 200.000 ;
        RECT 441.105 198.080 443.105 200.000 ;
        RECT 444.605 197.965 468.505 200.000 ;
        RECT 663.085 199.390 664.485 200.000 ;
      LAYER met2 ;
        RECT 664.765 199.670 665.785 200.000 ;
      LAYER met2 ;
        RECT 666.065 199.390 704.700 200.000 ;
        RECT 663.085 199.080 704.700 199.390 ;
      LAYER met2 ;
        RECT 704.980 199.360 705.240 200.000 ;
      LAYER met2 ;
        RECT 705.520 199.390 706.565 200.000 ;
      LAYER met2 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met2 ;
        RECT 707.775 199.390 708.055 200.000 ;
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
      LAYER met2 ;
        RECT 709.345 199.390 709.490 200.000 ;
      LAYER met2 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met2 ;
        RECT 710.700 199.390 715.060 200.000 ;
        RECT 705.520 199.080 715.060 199.390 ;
        RECT 394.710 4.925 468.735 197.965 ;
        RECT 663.085 196.020 715.060 199.080 ;
        RECT 663.085 195.735 714.775 196.020 ;
      LAYER met2 ;
        RECT 715.340 195.755 715.640 200.000 ;
      LAYER met2 ;
        RECT 715.920 198.310 716.495 200.000 ;
      LAYER met2 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met2 ;
        RECT 718.205 199.155 718.810 200.000 ;
      LAYER met2 ;
        RECT 719.090 199.435 720.755 200.000 ;
      LAYER met2 ;
        RECT 721.035 199.155 722.585 200.000 ;
      LAYER met2 ;
        RECT 722.820 199.580 723.445 200.000 ;
      LAYER met2 ;
        RECT 718.205 198.735 722.585 199.155 ;
      LAYER met2 ;
        RECT 722.865 199.015 723.445 199.580 ;
      LAYER met2 ;
        RECT 723.725 198.735 725.175 200.000 ;
        RECT 718.205 198.310 725.175 198.735 ;
        RECT 715.920 198.250 725.175 198.310 ;
        RECT 725.995 199.390 728.825 200.000 ;
      LAYER met2 ;
        RECT 729.105 199.670 729.575 200.000 ;
      LAYER met2 ;
        RECT 729.855 199.390 737.660 200.000 ;
        RECT 725.995 198.250 737.660 199.390 ;
        RECT 715.920 196.845 737.660 198.250 ;
        RECT 715.920 196.485 722.475 196.845 ;
        RECT 727.600 196.705 737.660 196.845 ;
        RECT 715.920 196.215 722.205 196.485 ;
      LAYER met2 ;
        RECT 722.755 196.425 727.320 196.565 ;
        RECT 722.755 196.355 727.650 196.425 ;
      LAYER met2 ;
        RECT 727.930 196.375 737.660 196.705 ;
      LAYER met2 ;
        RECT 722.755 196.305 727.180 196.355 ;
      LAYER met2 ;
        RECT 715.920 196.035 721.835 196.215 ;
      LAYER met2 ;
        RECT 722.755 196.205 723.115 196.305 ;
        RECT 723.125 196.205 723.225 196.305 ;
        RECT 727.070 196.235 727.305 196.305 ;
        RECT 727.320 196.235 727.650 196.355 ;
      LAYER met2 ;
        RECT 716.220 195.845 721.835 196.035 ;
      LAYER met2 ;
        RECT 722.485 196.165 722.755 196.205 ;
        RECT 722.855 196.165 723.125 196.205 ;
        RECT 722.485 196.025 723.125 196.165 ;
        RECT 727.070 196.095 727.650 196.235 ;
        RECT 727.070 196.070 727.305 196.095 ;
        RECT 722.485 195.935 722.755 196.025 ;
        RECT 722.855 195.935 723.125 196.025 ;
        RECT 715.340 195.740 715.940 195.755 ;
      LAYER met2 ;
        RECT 663.085 195.380 708.600 195.735 ;
      LAYER met2 ;
        RECT 715.055 195.455 715.940 195.740 ;
      LAYER met2 ;
        RECT 716.220 195.735 721.725 195.845 ;
      LAYER met2 ;
        RECT 722.115 195.565 722.855 195.935 ;
      LAYER met2 ;
        RECT 723.505 195.925 726.790 196.025 ;
        RECT 723.405 195.790 726.790 195.925 ;
      LAYER met2 ;
        RECT 727.305 195.955 727.625 196.070 ;
        RECT 727.650 195.955 727.995 196.095 ;
      LAYER met2 ;
        RECT 728.275 196.030 737.660 196.375 ;
      LAYER met2 ;
        RECT 727.305 195.815 727.995 195.955 ;
      LAYER met2 ;
        RECT 723.405 195.655 727.025 195.790 ;
      LAYER met2 ;
        RECT 727.305 195.750 727.625 195.815 ;
        RECT 727.650 195.750 727.995 195.815 ;
        RECT 722.005 195.455 722.485 195.565 ;
      LAYER met2 ;
        RECT 663.085 195.050 708.270 195.380 ;
      LAYER met2 ;
        RECT 708.880 195.315 722.485 195.455 ;
        RECT 708.880 195.245 709.235 195.315 ;
        RECT 715.340 195.245 715.640 195.315 ;
        RECT 722.115 195.245 722.485 195.315 ;
      LAYER met2 ;
        RECT 723.135 195.470 727.025 195.655 ;
      LAYER met2 ;
        RECT 727.625 195.675 727.955 195.750 ;
        RECT 727.995 195.675 728.265 195.750 ;
      LAYER met2 ;
        RECT 723.135 195.285 727.345 195.470 ;
      LAYER met2 ;
        RECT 727.625 195.425 728.265 195.675 ;
        RECT 727.625 195.420 727.955 195.425 ;
        RECT 708.880 195.195 722.485 195.245 ;
        RECT 708.880 195.100 709.235 195.195 ;
        RECT 709.250 195.100 709.345 195.195 ;
      LAYER met2 ;
        RECT 722.765 195.140 727.345 195.285 ;
      LAYER met2 ;
        RECT 708.550 195.055 708.880 195.100 ;
        RECT 708.920 195.055 709.250 195.100 ;
      LAYER met2 ;
        RECT 663.085 189.305 708.140 195.050 ;
      LAYER met2 ;
        RECT 708.550 194.845 709.250 195.055 ;
      LAYER met2 ;
        RECT 722.765 194.915 727.725 195.140 ;
      LAYER met2 ;
        RECT 708.550 194.770 708.880 194.845 ;
        RECT 708.920 194.770 709.250 194.845 ;
      LAYER met2 ;
        RECT 709.625 194.820 727.725 194.915 ;
      LAYER met2 ;
        RECT 708.420 194.640 708.550 194.770 ;
        RECT 708.680 194.640 708.920 194.770 ;
        RECT 708.420 194.530 708.920 194.640 ;
      LAYER met2 ;
        RECT 663.085 189.115 707.950 189.305 ;
        RECT 663.085 184.635 707.690 189.115 ;
      LAYER met2 ;
        RECT 708.420 189.025 708.680 194.530 ;
      LAYER met2 ;
        RECT 709.530 194.490 727.725 194.820 ;
        RECT 709.200 194.250 727.725 194.490 ;
      LAYER met2 ;
        RECT 708.230 188.915 708.680 189.025 ;
        RECT 708.230 188.835 708.420 188.915 ;
        RECT 708.600 188.835 708.680 188.915 ;
      LAYER met2 ;
        RECT 708.960 191.420 727.725 194.250 ;
        RECT 708.960 191.080 727.385 191.420 ;
      LAYER met2 ;
        RECT 728.005 191.140 728.265 195.425 ;
      LAYER met2 ;
        RECT 708.960 190.880 727.185 191.080 ;
      LAYER met2 ;
        RECT 727.665 190.890 728.265 191.140 ;
      LAYER met2 ;
        RECT 708.960 190.550 726.855 190.880 ;
      LAYER met2 ;
        RECT 727.665 190.800 728.005 190.890 ;
        RECT 728.035 190.800 728.265 190.890 ;
        RECT 727.465 190.750 727.665 190.800 ;
        RECT 727.835 190.750 728.035 190.800 ;
        RECT 727.465 190.680 728.035 190.750 ;
        RECT 727.465 190.600 727.665 190.680 ;
        RECT 727.835 190.600 728.035 190.680 ;
        RECT 707.970 188.465 708.600 188.835 ;
      LAYER met2 ;
        RECT 708.960 188.555 726.595 190.550 ;
      LAYER met2 ;
        RECT 727.135 190.540 727.465 190.600 ;
        RECT 727.505 190.540 727.835 190.600 ;
        RECT 727.135 190.400 727.835 190.540 ;
      LAYER met2 ;
        RECT 728.545 190.520 737.660 196.030 ;
      LAYER met2 ;
        RECT 727.135 190.270 727.465 190.400 ;
        RECT 727.505 190.270 727.835 190.400 ;
      LAYER met2 ;
        RECT 728.315 190.320 737.660 190.520 ;
        RECT 663.085 184.300 707.355 184.635 ;
      LAYER met2 ;
        RECT 707.970 184.355 708.230 188.465 ;
      LAYER met2 ;
        RECT 708.880 188.185 726.595 188.555 ;
        RECT 663.085 179.225 707.095 184.300 ;
      LAYER met2 ;
        RECT 707.635 184.105 708.230 184.355 ;
        RECT 707.635 184.020 707.970 184.105 ;
        RECT 708.005 184.020 708.230 184.105 ;
        RECT 707.375 183.650 708.005 184.020 ;
      LAYER met2 ;
        RECT 708.510 183.740 726.595 188.185 ;
      LAYER met2 ;
        RECT 707.375 179.505 707.635 183.650 ;
      LAYER met2 ;
        RECT 708.285 183.370 726.595 183.740 ;
        RECT 707.915 179.225 726.595 183.370 ;
        RECT 663.085 172.420 726.595 179.225 ;
      LAYER met2 ;
        RECT 726.875 189.900 727.505 190.270 ;
      LAYER met2 ;
        RECT 728.115 189.990 737.660 190.320 ;
      LAYER met2 ;
        RECT 726.875 173.390 727.135 189.900 ;
      LAYER met2 ;
        RECT 727.785 189.620 737.660 189.990 ;
        RECT 727.415 173.670 737.660 189.620 ;
      LAYER met2 ;
        RECT 726.875 172.700 727.350 173.390 ;
      LAYER met2 ;
        RECT 663.085 172.345 726.810 172.420 ;
        RECT 663.085 169.195 726.595 172.345 ;
      LAYER met2 ;
        RECT 727.090 172.065 727.350 172.700 ;
        RECT 726.875 171.855 727.350 172.065 ;
        RECT 726.875 171.850 727.090 171.855 ;
        RECT 726.875 171.375 727.350 171.850 ;
      LAYER met2 ;
        RECT 663.085 169.050 726.450 169.195 ;
        RECT 663.085 168.825 726.225 169.050 ;
      LAYER met2 ;
        RECT 726.875 168.915 727.135 171.375 ;
      LAYER met2 ;
        RECT 727.630 171.095 737.660 173.670 ;
        RECT 663.085 164.260 726.200 168.825 ;
      LAYER met2 ;
        RECT 726.730 168.770 727.135 168.915 ;
        RECT 726.505 168.735 726.730 168.770 ;
        RECT 726.875 168.735 727.135 168.770 ;
        RECT 726.505 168.665 727.135 168.735 ;
        RECT 726.505 168.545 726.730 168.665 ;
        RECT 726.875 168.545 727.135 168.665 ;
        RECT 726.480 168.520 726.505 168.545 ;
        RECT 726.740 168.520 726.875 168.545 ;
        RECT 726.480 168.410 726.875 168.520 ;
      LAYER met2 ;
        RECT 663.085 163.440 725.570 164.260 ;
      LAYER met2 ;
        RECT 726.480 163.980 726.740 168.410 ;
      LAYER met2 ;
        RECT 727.415 168.265 737.660 171.095 ;
        RECT 727.155 168.130 737.660 168.265 ;
      LAYER met2 ;
        RECT 725.850 163.720 726.740 163.980 ;
      LAYER met2 ;
        RECT 727.020 163.440 737.660 168.130 ;
        RECT 663.085 0.790 737.660 163.440 ;
        RECT 932.085 0.000 1011.790 208.285 ;
        RECT 1206.300 197.965 1226.905 198.000 ;
        RECT 1227.465 197.965 1260.075 198.000 ;
        RECT 1260.505 197.965 1280.500 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 158.415 1280.500 197.965 ;
      LAYER met2 ;
        RECT 1281.260 197.725 1281.400 234.270 ;
        RECT 1485.440 221.690 1485.700 222.010 ;
        RECT 1476.240 221.350 1476.500 221.670 ;
        RECT 1476.300 210.965 1476.440 221.350 ;
        RECT 1485.500 210.965 1485.640 221.690 ;
        RECT 1488.720 210.965 1488.860 234.270 ;
        RECT 1497.860 221.690 1498.120 222.010 ;
        RECT 1528.680 221.690 1528.940 222.010 ;
        RECT 1497.920 210.965 1498.060 221.690 ;
        RECT 1516.260 221.350 1516.520 221.670 ;
        RECT 1516.320 210.965 1516.460 221.350 ;
        RECT 1522.700 220.670 1522.960 220.990 ;
        RECT 1522.760 210.965 1522.900 220.670 ;
        RECT 1528.740 210.965 1528.880 221.690 ;
        RECT 1547.140 210.965 1547.280 234.270 ;
        RECT 1749.940 222.030 1750.200 222.350 ;
        RECT 1750.000 220.990 1750.140 222.030 ;
        RECT 1759.600 221.350 1759.860 221.670 ;
        RECT 1749.940 220.670 1750.200 220.990 ;
        RECT 1750.400 220.670 1750.660 220.990 ;
        RECT 1750.460 210.965 1750.600 220.670 ;
        RECT 1759.660 210.965 1759.800 221.350 ;
        RECT 1762.880 210.965 1763.020 234.270 ;
        RECT 1796.860 222.030 1797.120 222.350 ;
        RECT 1772.020 221.350 1772.280 221.670 ;
        RECT 1772.080 210.965 1772.220 221.350 ;
        RECT 1790.420 220.670 1790.680 220.990 ;
        RECT 1790.480 210.965 1790.620 220.670 ;
        RECT 1796.920 210.965 1797.060 222.030 ;
        RECT 1802.840 221.350 1803.100 221.670 ;
        RECT 1802.900 220.990 1803.040 221.350 ;
        RECT 1802.840 220.670 1803.100 220.990 ;
        RECT 1802.900 210.965 1803.040 220.670 ;
        RECT 1821.300 210.965 1821.440 234.270 ;
        RECT 2024.550 221.155 2024.830 221.525 ;
        RECT 2024.620 210.965 2024.760 221.155 ;
        RECT 2033.760 221.010 2034.020 221.330 ;
        RECT 2033.820 210.965 2033.960 221.010 ;
        RECT 2037.040 210.965 2037.180 234.270 ;
        RECT 2071.020 222.030 2071.280 222.350 ;
        RECT 2064.570 221.155 2064.850 221.525 ;
        RECT 2064.640 210.965 2064.780 221.155 ;
        RECT 2071.080 220.990 2071.220 222.030 ;
        RECT 2071.020 220.670 2071.280 220.990 ;
        RECT 2071.080 210.965 2071.220 220.670 ;
        RECT 2095.460 210.965 2095.600 234.270 ;
        RECT 2298.250 221.155 2298.530 221.525 ;
        RECT 2298.320 210.965 2298.460 221.155 ;
        RECT 2307.460 221.010 2307.720 221.330 ;
        RECT 2307.520 210.965 2307.660 221.010 ;
        RECT 2310.740 210.965 2310.880 234.270 ;
        RECT 2344.720 221.690 2344.980 222.010 ;
        RECT 2338.270 221.155 2338.550 221.525 ;
        RECT 2338.340 210.965 2338.480 221.155 ;
        RECT 2344.780 220.990 2344.920 221.690 ;
        RECT 2344.720 220.670 2344.980 220.990 ;
        RECT 2344.780 210.965 2344.920 220.670 ;
        RECT 2369.160 210.965 2369.300 234.270 ;
        RECT 2572.410 221.155 2572.690 221.525 ;
        RECT 2572.480 210.965 2572.620 221.155 ;
        RECT 2581.620 221.010 2581.880 221.330 ;
        RECT 2581.680 210.965 2581.820 221.010 ;
        RECT 2584.900 210.965 2585.040 234.270 ;
        RECT 2618.880 227.810 2619.140 228.130 ;
        RECT 2593.580 227.470 2593.840 227.790 ;
        RECT 2593.640 221.330 2593.780 227.470 ;
        RECT 2612.430 221.835 2612.710 222.205 ;
        RECT 2618.940 222.010 2619.080 227.810 ;
        RECT 2593.580 221.010 2593.840 221.330 ;
        RECT 2612.500 210.965 2612.640 221.835 ;
        RECT 2618.880 221.690 2619.140 222.010 ;
        RECT 2618.940 210.965 2619.080 221.690 ;
        RECT 3367.360 213.850 3367.500 557.610 ;
        RECT 3367.820 542.290 3367.960 763.990 ;
        RECT 3368.280 745.270 3368.420 946.230 ;
        RECT 3376.560 936.625 3376.700 976.505 ;
        RECT 3377.035 976.435 3379.435 976.505 ;
      LAYER met2 ;
        RECT 3379.715 976.155 3588.000 976.995 ;
        RECT 3379.435 973.775 3588.000 976.155 ;
        RECT 3379.715 972.935 3588.000 973.775 ;
        RECT 3379.435 971.015 3588.000 972.935 ;
        RECT 3379.715 970.175 3588.000 971.015 ;
        RECT 3379.435 967.795 3588.000 970.175 ;
        RECT 3379.715 966.955 3588.000 967.795 ;
        RECT 3379.435 964.575 3588.000 966.955 ;
        RECT 3379.715 963.735 3588.000 964.575 ;
        RECT 3379.435 961.815 3588.000 963.735 ;
      LAYER met2 ;
        RECT 3377.035 961.255 3379.435 961.535 ;
      LAYER met2 ;
        RECT 3379.715 960.975 3588.000 961.815 ;
        RECT 3379.435 958.595 3588.000 960.975 ;
        RECT 3379.715 957.755 3588.000 958.595 ;
        RECT 3379.435 955.375 3588.000 957.755 ;
      LAYER met2 ;
        RECT 3377.035 954.815 3379.435 955.095 ;
      LAYER met2 ;
        RECT 3379.715 954.535 3588.000 955.375 ;
        RECT 3379.435 952.615 3588.000 954.535 ;
      LAYER met2 ;
        RECT 3377.035 952.055 3379.435 952.335 ;
      LAYER met2 ;
        RECT 3379.715 951.775 3588.000 952.615 ;
        RECT 3379.435 949.395 3588.000 951.775 ;
        RECT 3379.715 948.555 3588.000 949.395 ;
      LAYER met2 ;
        RECT 3376.960 946.230 3377.220 946.550 ;
        RECT 3377.020 945.895 3377.160 946.230 ;
      LAYER met2 ;
        RECT 3379.435 946.175 3588.000 948.555 ;
      LAYER met2 ;
        RECT 3377.020 945.755 3379.435 945.895 ;
        RECT 3377.035 945.615 3379.435 945.755 ;
      LAYER met2 ;
        RECT 3379.715 945.335 3588.000 946.175 ;
        RECT 3379.435 943.415 3588.000 945.335 ;
      LAYER met2 ;
        RECT 3377.035 942.855 3379.435 943.135 ;
      LAYER met2 ;
        RECT 3379.715 942.575 3588.000 943.415 ;
        RECT 3379.435 940.195 3588.000 942.575 ;
        RECT 3379.715 939.355 3588.000 940.195 ;
        RECT 3379.435 936.975 3588.000 939.355 ;
      LAYER met2 ;
        RECT 3377.035 936.625 3379.435 936.695 ;
        RECT 3376.560 936.485 3379.435 936.625 ;
        RECT 3377.035 936.415 3379.435 936.485 ;
      LAYER met2 ;
        RECT 3379.715 936.135 3588.000 936.975 ;
        RECT 3379.435 935.085 3588.000 936.135 ;
        RECT 3379.435 792.795 3588.000 793.790 ;
        RECT 3379.715 791.955 3588.000 792.795 ;
        RECT 3379.435 790.035 3588.000 791.955 ;
        RECT 3379.715 789.195 3588.000 790.035 ;
        RECT 3379.435 786.815 3588.000 789.195 ;
        RECT 3379.715 785.975 3588.000 786.815 ;
        RECT 3379.435 783.595 3588.000 785.975 ;
        RECT 3379.715 782.755 3588.000 783.595 ;
        RECT 3379.435 780.835 3588.000 782.755 ;
        RECT 3379.715 779.995 3588.000 780.835 ;
      LAYER met2 ;
        RECT 3369.600 779.630 3369.860 779.950 ;
        RECT 3376.960 779.630 3377.220 779.950 ;
        RECT 3368.280 745.130 3368.880 745.270 ;
        RECT 3368.740 722.830 3368.880 745.130 ;
        RECT 3368.680 722.510 3368.940 722.830 ;
        RECT 3367.760 541.970 3368.020 542.290 ;
        RECT 3367.820 228.130 3367.960 541.970 ;
        RECT 3368.740 503.045 3368.880 722.510 ;
        RECT 3369.660 557.930 3369.800 779.630 ;
        RECT 3377.020 777.335 3377.160 779.630 ;
      LAYER met2 ;
        RECT 3379.435 777.615 3588.000 779.995 ;
      LAYER met2 ;
        RECT 3377.020 777.195 3379.435 777.335 ;
        RECT 3377.035 777.055 3379.435 777.195 ;
      LAYER met2 ;
        RECT 3379.715 776.775 3588.000 777.615 ;
        RECT 3379.435 774.395 3588.000 776.775 ;
        RECT 3379.715 773.555 3588.000 774.395 ;
        RECT 3379.435 771.635 3588.000 773.555 ;
        RECT 3379.715 770.795 3588.000 771.635 ;
        RECT 3379.435 768.415 3588.000 770.795 ;
        RECT 3379.715 767.575 3588.000 768.415 ;
        RECT 3379.435 765.195 3588.000 767.575 ;
        RECT 3379.715 764.355 3588.000 765.195 ;
      LAYER met2 ;
        RECT 3376.960 763.990 3377.220 764.310 ;
        RECT 3377.020 762.155 3377.160 763.990 ;
      LAYER met2 ;
        RECT 3379.435 762.435 3588.000 764.355 ;
      LAYER met2 ;
        RECT 3377.020 761.940 3379.435 762.155 ;
        RECT 3377.035 761.875 3379.435 761.940 ;
      LAYER met2 ;
        RECT 3379.715 761.595 3588.000 762.435 ;
        RECT 3379.435 759.215 3588.000 761.595 ;
        RECT 3379.715 758.375 3588.000 759.215 ;
        RECT 3379.435 755.995 3588.000 758.375 ;
      LAYER met2 ;
        RECT 3377.035 755.645 3379.435 755.715 ;
        RECT 3376.560 755.505 3379.435 755.645 ;
        RECT 3376.560 715.625 3376.700 755.505 ;
        RECT 3377.035 755.435 3379.435 755.505 ;
      LAYER met2 ;
        RECT 3379.715 755.155 3588.000 755.995 ;
        RECT 3379.435 752.775 3588.000 755.155 ;
        RECT 3379.715 751.935 3588.000 752.775 ;
        RECT 3379.435 750.015 3588.000 751.935 ;
        RECT 3379.715 749.175 3588.000 750.015 ;
        RECT 3379.435 746.795 3588.000 749.175 ;
        RECT 3379.715 745.955 3588.000 746.795 ;
        RECT 3379.435 743.575 3588.000 745.955 ;
        RECT 3379.715 742.735 3588.000 743.575 ;
        RECT 3379.435 740.815 3588.000 742.735 ;
      LAYER met2 ;
        RECT 3377.035 740.255 3379.435 740.535 ;
      LAYER met2 ;
        RECT 3379.715 739.975 3588.000 740.815 ;
        RECT 3379.435 737.595 3588.000 739.975 ;
        RECT 3379.715 736.755 3588.000 737.595 ;
        RECT 3379.435 734.375 3588.000 736.755 ;
      LAYER met2 ;
        RECT 3377.035 733.815 3379.435 734.095 ;
      LAYER met2 ;
        RECT 3379.715 733.535 3588.000 734.375 ;
        RECT 3379.435 731.615 3588.000 733.535 ;
      LAYER met2 ;
        RECT 3377.035 731.055 3379.435 731.335 ;
      LAYER met2 ;
        RECT 3379.715 730.775 3588.000 731.615 ;
        RECT 3379.435 728.395 3588.000 730.775 ;
        RECT 3379.715 727.555 3588.000 728.395 ;
        RECT 3379.435 725.175 3588.000 727.555 ;
      LAYER met2 ;
        RECT 3377.035 724.755 3379.435 724.895 ;
        RECT 3377.020 724.615 3379.435 724.755 ;
        RECT 3377.020 722.830 3377.160 724.615 ;
      LAYER met2 ;
        RECT 3379.715 724.335 3588.000 725.175 ;
      LAYER met2 ;
        RECT 3376.960 722.510 3377.220 722.830 ;
      LAYER met2 ;
        RECT 3379.435 722.415 3588.000 724.335 ;
      LAYER met2 ;
        RECT 3377.035 721.855 3379.435 722.135 ;
      LAYER met2 ;
        RECT 3379.715 721.575 3588.000 722.415 ;
        RECT 3379.435 719.195 3588.000 721.575 ;
        RECT 3379.715 718.355 3588.000 719.195 ;
        RECT 3379.435 715.975 3588.000 718.355 ;
      LAYER met2 ;
        RECT 3377.035 715.625 3379.435 715.695 ;
        RECT 3376.560 715.485 3379.435 715.625 ;
        RECT 3377.035 715.415 3379.435 715.485 ;
      LAYER met2 ;
        RECT 3379.715 715.135 3588.000 715.975 ;
        RECT 3379.435 714.085 3588.000 715.135 ;
        RECT 3379.435 570.795 3588.000 571.790 ;
        RECT 3379.715 569.955 3588.000 570.795 ;
        RECT 3379.435 568.035 3588.000 569.955 ;
        RECT 3379.715 567.195 3588.000 568.035 ;
        RECT 3379.435 564.815 3588.000 567.195 ;
        RECT 3379.715 563.975 3588.000 564.815 ;
        RECT 3379.435 561.595 3588.000 563.975 ;
        RECT 3379.715 560.755 3588.000 561.595 ;
        RECT 3379.435 558.835 3588.000 560.755 ;
        RECT 3379.715 557.995 3588.000 558.835 ;
      LAYER met2 ;
        RECT 3369.600 557.610 3369.860 557.930 ;
        RECT 3376.960 557.610 3377.220 557.930 ;
        RECT 3377.020 555.335 3377.160 557.610 ;
      LAYER met2 ;
        RECT 3379.435 555.615 3588.000 557.995 ;
      LAYER met2 ;
        RECT 3377.020 555.220 3379.435 555.335 ;
        RECT 3377.035 555.055 3379.435 555.220 ;
      LAYER met2 ;
        RECT 3379.715 554.775 3588.000 555.615 ;
        RECT 3379.435 552.395 3588.000 554.775 ;
        RECT 3379.715 551.555 3588.000 552.395 ;
        RECT 3379.435 549.635 3588.000 551.555 ;
        RECT 3379.715 548.795 3588.000 549.635 ;
        RECT 3379.435 546.415 3588.000 548.795 ;
        RECT 3379.715 545.575 3588.000 546.415 ;
        RECT 3379.435 543.195 3588.000 545.575 ;
        RECT 3379.715 542.355 3588.000 543.195 ;
      LAYER met2 ;
        RECT 3376.960 541.970 3377.220 542.290 ;
        RECT 3377.020 540.155 3377.160 541.970 ;
      LAYER met2 ;
        RECT 3379.435 540.435 3588.000 542.355 ;
      LAYER met2 ;
        RECT 3377.020 540.015 3379.435 540.155 ;
        RECT 3377.035 539.875 3379.435 540.015 ;
      LAYER met2 ;
        RECT 3379.715 539.595 3588.000 540.435 ;
        RECT 3379.435 537.215 3588.000 539.595 ;
        RECT 3379.715 536.375 3588.000 537.215 ;
      LAYER met2 ;
        RECT 3376.560 534.070 3377.160 534.210 ;
        RECT 3368.670 502.675 3368.950 503.045 ;
        RECT 3367.760 227.810 3368.020 228.130 ;
        RECT 3368.740 227.790 3368.880 502.675 ;
        RECT 3376.560 493.625 3376.700 534.070 ;
        RECT 3377.020 533.715 3377.160 534.070 ;
      LAYER met2 ;
        RECT 3379.435 533.995 3588.000 536.375 ;
      LAYER met2 ;
        RECT 3377.020 533.460 3379.435 533.715 ;
        RECT 3377.035 533.435 3379.435 533.460 ;
      LAYER met2 ;
        RECT 3379.715 533.155 3588.000 533.995 ;
        RECT 3379.435 530.775 3588.000 533.155 ;
        RECT 3379.715 529.935 3588.000 530.775 ;
        RECT 3379.435 528.015 3588.000 529.935 ;
        RECT 3379.715 527.175 3588.000 528.015 ;
        RECT 3379.435 524.795 3588.000 527.175 ;
        RECT 3379.715 523.955 3588.000 524.795 ;
        RECT 3379.435 521.575 3588.000 523.955 ;
        RECT 3379.715 520.735 3588.000 521.575 ;
        RECT 3379.435 518.815 3588.000 520.735 ;
      LAYER met2 ;
        RECT 3377.035 518.255 3379.435 518.535 ;
      LAYER met2 ;
        RECT 3379.715 517.975 3588.000 518.815 ;
        RECT 3379.435 515.595 3588.000 517.975 ;
        RECT 3379.715 514.755 3588.000 515.595 ;
        RECT 3379.435 512.375 3588.000 514.755 ;
      LAYER met2 ;
        RECT 3377.035 511.815 3379.435 512.095 ;
      LAYER met2 ;
        RECT 3379.715 511.535 3588.000 512.375 ;
        RECT 3379.435 509.615 3588.000 511.535 ;
      LAYER met2 ;
        RECT 3377.035 509.055 3379.435 509.335 ;
      LAYER met2 ;
        RECT 3379.715 508.775 3588.000 509.615 ;
        RECT 3379.435 506.395 3588.000 508.775 ;
        RECT 3379.715 505.555 3588.000 506.395 ;
        RECT 3379.435 503.175 3588.000 505.555 ;
      LAYER met2 ;
        RECT 3376.950 502.895 3377.230 503.045 ;
        RECT 3376.950 502.675 3379.435 502.895 ;
        RECT 3377.035 502.615 3379.435 502.675 ;
      LAYER met2 ;
        RECT 3379.715 502.335 3588.000 503.175 ;
        RECT 3379.435 500.415 3588.000 502.335 ;
      LAYER met2 ;
        RECT 3377.035 499.855 3379.435 500.135 ;
      LAYER met2 ;
        RECT 3379.715 499.575 3588.000 500.415 ;
        RECT 3379.435 497.195 3588.000 499.575 ;
        RECT 3379.715 496.355 3588.000 497.195 ;
        RECT 3379.435 493.975 3588.000 496.355 ;
      LAYER met2 ;
        RECT 3377.035 493.625 3379.435 493.695 ;
        RECT 3376.560 493.485 3379.435 493.625 ;
        RECT 3377.035 493.415 3379.435 493.485 ;
      LAYER met2 ;
        RECT 3379.715 493.135 3588.000 493.975 ;
        RECT 3379.435 492.085 3588.000 493.135 ;
      LAYER met2 ;
        RECT 3368.680 227.470 3368.940 227.790 ;
        RECT 2899.480 213.530 2899.740 213.850 ;
        RECT 3367.300 213.530 3367.560 213.850 ;
        RECT 1476.300 209.030 1476.695 210.965 ;
        RECT 1476.415 208.565 1476.695 209.030 ;
        RECT 1479.635 208.565 1479.915 210.965 ;
        RECT 1482.855 208.565 1483.135 210.965 ;
        RECT 1485.500 209.030 1485.895 210.965 ;
        RECT 1488.720 209.170 1489.115 210.965 ;
        RECT 1489.580 209.450 1489.840 209.770 ;
        RECT 1489.640 209.170 1489.780 209.450 ;
        RECT 1488.720 209.030 1489.780 209.170 ;
        RECT 1485.615 208.565 1485.895 209.030 ;
        RECT 1488.835 208.565 1489.115 209.030 ;
        RECT 1492.055 208.565 1492.335 210.965 ;
        RECT 1494.815 208.565 1495.095 210.965 ;
        RECT 1497.920 209.030 1498.315 210.965 ;
        RECT 1498.035 208.565 1498.315 209.030 ;
        RECT 1501.255 208.565 1501.535 210.965 ;
        RECT 1503.380 209.450 1503.640 209.770 ;
        RECT 1503.440 209.170 1503.580 209.450 ;
        RECT 1504.015 209.170 1504.295 210.965 ;
        RECT 1507.235 209.170 1507.515 210.965 ;
        RECT 1510.455 209.170 1510.735 210.965 ;
        RECT 1511.200 209.450 1511.460 209.770 ;
        RECT 1511.260 209.170 1511.400 209.450 ;
        RECT 1503.440 209.030 1511.400 209.170 ;
        RECT 1516.320 209.030 1516.715 210.965 ;
        RECT 1522.760 209.030 1523.155 210.965 ;
        RECT 1504.015 208.565 1504.295 209.030 ;
        RECT 1507.235 208.565 1507.515 209.030 ;
        RECT 1510.455 208.565 1510.735 209.030 ;
        RECT 1516.435 208.565 1516.715 209.030 ;
        RECT 1522.875 208.565 1523.155 209.030 ;
        RECT 1525.635 209.170 1525.915 210.965 ;
        RECT 1526.380 209.450 1526.640 209.770 ;
        RECT 1526.440 209.170 1526.580 209.450 ;
        RECT 1525.635 209.030 1526.580 209.170 ;
        RECT 1528.740 209.030 1529.135 210.965 ;
        RECT 1525.635 208.565 1525.915 209.030 ;
        RECT 1528.855 208.565 1529.135 209.030 ;
        RECT 1532.075 209.170 1532.355 210.965 ;
        RECT 1532.820 209.450 1533.080 209.770 ;
        RECT 1532.880 209.170 1533.020 209.450 ;
        RECT 1532.075 209.030 1533.020 209.170 ;
        RECT 1538.055 209.170 1538.335 210.965 ;
        RECT 1543.400 209.450 1543.660 209.770 ;
        RECT 1543.460 209.170 1543.600 209.450 ;
        RECT 1544.035 209.170 1544.315 210.965 ;
        RECT 1547.140 209.170 1547.535 210.965 ;
        RECT 1538.055 209.090 1539.000 209.170 ;
        RECT 1538.055 209.030 1539.060 209.090 ;
        RECT 1543.460 209.030 1547.535 209.170 ;
        RECT 1532.075 208.565 1532.355 209.030 ;
        RECT 1538.055 208.565 1538.335 209.030 ;
        RECT 1538.800 208.770 1539.060 209.030 ;
        RECT 1544.035 208.565 1544.315 209.030 ;
        RECT 1547.255 208.565 1547.535 209.030 ;
        RECT 1553.235 208.565 1553.515 210.965 ;
        RECT 1750.415 208.565 1750.695 210.965 ;
        RECT 1753.635 208.565 1753.915 210.965 ;
        RECT 1756.855 208.565 1757.135 210.965 ;
        RECT 1759.615 208.565 1759.895 210.965 ;
        RECT 1762.835 209.850 1763.115 210.965 ;
        RECT 1762.835 209.770 1763.480 209.850 ;
        RECT 1762.835 209.710 1763.540 209.770 ;
        RECT 1762.835 208.565 1763.115 209.710 ;
        RECT 1763.280 209.450 1763.540 209.710 ;
        RECT 1766.055 208.565 1766.335 210.965 ;
        RECT 1768.815 208.565 1769.095 210.965 ;
        RECT 1772.035 208.565 1772.315 210.965 ;
        RECT 1775.255 208.565 1775.535 210.965 ;
        RECT 1777.540 209.450 1777.800 209.770 ;
        RECT 1777.600 209.170 1777.740 209.450 ;
        RECT 1778.015 209.170 1778.295 210.965 ;
        RECT 1781.235 209.170 1781.515 210.965 ;
        RECT 1784.455 209.170 1784.735 210.965 ;
        RECT 1784.900 209.450 1785.160 209.770 ;
        RECT 1784.960 209.170 1785.100 209.450 ;
        RECT 1777.600 209.030 1785.100 209.170 ;
        RECT 1778.015 208.565 1778.295 209.030 ;
        RECT 1781.235 208.565 1781.515 209.030 ;
        RECT 1784.455 208.565 1784.735 209.030 ;
        RECT 1790.435 208.565 1790.715 210.965 ;
        RECT 1796.875 208.565 1797.155 210.965 ;
        RECT 1799.160 209.450 1799.420 209.770 ;
        RECT 1799.220 209.170 1799.360 209.450 ;
        RECT 1799.635 209.170 1799.915 210.965 ;
        RECT 1799.220 209.030 1799.915 209.170 ;
        RECT 1799.635 208.565 1799.915 209.030 ;
        RECT 1802.855 208.565 1803.135 210.965 ;
        RECT 1805.600 209.450 1805.860 209.770 ;
        RECT 1805.660 209.170 1805.800 209.450 ;
        RECT 1806.075 209.170 1806.355 210.965 ;
        RECT 1805.660 209.030 1806.355 209.170 ;
        RECT 1806.075 208.565 1806.355 209.030 ;
        RECT 1812.055 209.170 1812.335 210.965 ;
        RECT 1817.560 209.450 1817.820 209.770 ;
        RECT 1817.620 209.170 1817.760 209.450 ;
        RECT 1818.035 209.170 1818.315 210.965 ;
        RECT 1821.255 209.170 1821.535 210.965 ;
        RECT 1812.055 209.090 1812.700 209.170 ;
        RECT 1812.055 209.030 1812.760 209.090 ;
        RECT 1817.620 209.030 1821.535 209.170 ;
        RECT 1812.055 208.565 1812.335 209.030 ;
        RECT 1812.500 208.770 1812.760 209.030 ;
        RECT 1818.035 208.565 1818.315 209.030 ;
        RECT 1821.255 208.565 1821.535 209.030 ;
        RECT 1827.235 208.565 1827.515 210.965 ;
        RECT 2024.415 209.100 2024.760 210.965 ;
        RECT 2024.415 208.565 2024.695 209.100 ;
        RECT 2030.855 208.565 2031.135 210.965 ;
        RECT 2033.615 209.100 2033.960 210.965 ;
        RECT 2036.835 209.850 2037.180 210.965 ;
        RECT 2036.835 209.770 2037.640 209.850 ;
        RECT 2036.835 209.710 2037.700 209.770 ;
        RECT 2036.835 209.100 2037.180 209.710 ;
        RECT 2037.440 209.450 2037.700 209.710 ;
        RECT 2033.615 208.565 2033.895 209.100 ;
        RECT 2036.835 208.565 2037.115 209.100 ;
        RECT 2040.055 208.565 2040.335 210.965 ;
        RECT 2042.815 208.565 2043.095 210.965 ;
        RECT 2049.255 208.565 2049.535 210.965 ;
        RECT 2051.240 209.450 2051.500 209.770 ;
        RECT 2051.300 209.170 2051.440 209.450 ;
        RECT 2052.015 209.170 2052.295 210.965 ;
        RECT 2057.680 209.450 2057.940 209.770 ;
        RECT 2051.300 209.030 2052.295 209.170 ;
        RECT 2057.740 209.170 2057.880 209.450 ;
        RECT 2058.455 209.170 2058.735 210.965 ;
        RECT 2057.740 209.030 2058.735 209.170 ;
        RECT 2052.015 208.565 2052.295 209.030 ;
        RECT 2058.455 208.565 2058.735 209.030 ;
        RECT 2064.435 209.100 2064.780 210.965 ;
        RECT 2070.875 209.100 2071.220 210.965 ;
        RECT 2072.860 209.450 2073.120 209.770 ;
        RECT 2072.920 209.170 2073.060 209.450 ;
        RECT 2073.635 209.170 2073.915 210.965 ;
        RECT 2079.300 209.450 2079.560 209.770 ;
        RECT 2064.435 208.565 2064.715 209.100 ;
        RECT 2070.875 208.565 2071.155 209.100 ;
        RECT 2072.920 209.030 2073.915 209.170 ;
        RECT 2079.360 209.170 2079.500 209.450 ;
        RECT 2080.075 209.170 2080.355 210.965 ;
        RECT 2079.360 209.030 2080.355 209.170 ;
        RECT 2073.635 208.565 2073.915 209.030 ;
        RECT 2080.075 208.565 2080.355 209.030 ;
        RECT 2086.055 209.170 2086.335 210.965 ;
        RECT 2091.260 209.450 2091.520 209.770 ;
        RECT 2091.320 209.170 2091.460 209.450 ;
        RECT 2092.035 209.170 2092.315 210.965 ;
        RECT 2095.255 209.170 2095.600 210.965 ;
        RECT 2086.055 209.090 2086.860 209.170 ;
        RECT 2091.320 209.100 2095.600 209.170 ;
        RECT 2086.055 209.030 2086.920 209.090 ;
        RECT 2091.320 209.030 2095.535 209.100 ;
        RECT 2086.055 208.565 2086.335 209.030 ;
        RECT 2086.660 208.770 2086.920 209.030 ;
        RECT 2092.035 208.565 2092.315 209.030 ;
        RECT 2095.255 208.565 2095.535 209.030 ;
        RECT 2101.235 208.565 2101.515 210.965 ;
        RECT 2298.320 209.030 2298.695 210.965 ;
        RECT 2298.415 208.565 2298.695 209.030 ;
        RECT 2304.855 208.565 2305.135 210.965 ;
        RECT 2307.520 209.030 2307.895 210.965 ;
        RECT 2310.740 209.170 2311.115 210.965 ;
        RECT 2311.600 209.450 2311.860 209.770 ;
        RECT 2311.660 209.170 2311.800 209.450 ;
        RECT 2310.740 209.030 2311.800 209.170 ;
        RECT 2307.615 208.565 2307.895 209.030 ;
        RECT 2310.835 208.565 2311.115 209.030 ;
        RECT 2314.055 208.565 2314.335 210.965 ;
        RECT 2316.815 208.565 2317.095 210.965 ;
        RECT 2323.255 208.565 2323.535 210.965 ;
        RECT 2325.400 209.450 2325.660 209.770 ;
        RECT 2325.460 209.170 2325.600 209.450 ;
        RECT 2326.015 209.170 2326.295 210.965 ;
        RECT 2331.840 209.450 2332.100 209.770 ;
        RECT 2325.460 209.030 2326.295 209.170 ;
        RECT 2331.900 209.170 2332.040 209.450 ;
        RECT 2332.455 209.170 2332.735 210.965 ;
        RECT 2331.900 209.030 2332.735 209.170 ;
        RECT 2338.340 209.030 2338.715 210.965 ;
        RECT 2344.780 209.030 2345.155 210.965 ;
        RECT 2347.020 209.450 2347.280 209.770 ;
        RECT 2347.080 209.170 2347.220 209.450 ;
        RECT 2347.635 209.170 2347.915 210.965 ;
        RECT 2353.460 209.450 2353.720 209.770 ;
        RECT 2347.080 209.030 2347.915 209.170 ;
        RECT 2353.520 209.170 2353.660 209.450 ;
        RECT 2354.075 209.170 2354.355 210.965 ;
        RECT 2353.520 209.030 2354.355 209.170 ;
        RECT 2326.015 208.565 2326.295 209.030 ;
        RECT 2332.455 208.565 2332.735 209.030 ;
        RECT 2338.435 208.565 2338.715 209.030 ;
        RECT 2344.875 208.565 2345.155 209.030 ;
        RECT 2347.635 208.565 2347.915 209.030 ;
        RECT 2354.075 208.565 2354.355 209.030 ;
        RECT 2360.055 209.170 2360.335 210.965 ;
        RECT 2365.420 209.450 2365.680 209.770 ;
        RECT 2365.480 209.170 2365.620 209.450 ;
        RECT 2366.035 209.170 2366.315 210.965 ;
        RECT 2369.160 209.170 2369.535 210.965 ;
        RECT 2360.055 209.090 2361.020 209.170 ;
        RECT 2360.055 209.030 2361.080 209.090 ;
        RECT 2365.480 209.030 2369.535 209.170 ;
        RECT 2360.055 208.565 2360.335 209.030 ;
        RECT 2360.820 208.770 2361.080 209.030 ;
        RECT 2366.035 208.565 2366.315 209.030 ;
        RECT 2369.255 208.565 2369.535 209.030 ;
        RECT 2375.235 208.565 2375.515 210.965 ;
        RECT 2572.415 208.565 2572.695 210.965 ;
        RECT 2578.855 208.565 2579.135 210.965 ;
        RECT 2581.615 208.565 2581.895 210.965 ;
        RECT 2584.835 209.850 2585.115 210.965 ;
        RECT 2584.835 209.770 2585.500 209.850 ;
        RECT 2584.835 209.710 2585.560 209.770 ;
        RECT 2584.835 208.565 2585.115 209.710 ;
        RECT 2585.300 209.450 2585.560 209.710 ;
        RECT 2588.055 208.565 2588.335 210.965 ;
        RECT 2590.815 208.565 2591.095 210.965 ;
        RECT 2597.255 208.565 2597.535 210.965 ;
        RECT 2599.560 209.450 2599.820 209.770 ;
        RECT 2599.620 209.170 2599.760 209.450 ;
        RECT 2600.015 209.170 2600.295 210.965 ;
        RECT 2606.000 209.450 2606.260 209.770 ;
        RECT 2599.620 209.030 2600.295 209.170 ;
        RECT 2606.060 209.170 2606.200 209.450 ;
        RECT 2606.455 209.170 2606.735 210.965 ;
        RECT 2606.060 209.030 2606.735 209.170 ;
        RECT 2600.015 208.565 2600.295 209.030 ;
        RECT 2606.455 208.565 2606.735 209.030 ;
        RECT 2612.435 208.565 2612.715 210.965 ;
        RECT 2618.875 208.565 2619.155 210.965 ;
        RECT 2621.180 209.450 2621.440 209.770 ;
        RECT 2621.240 209.170 2621.380 209.450 ;
        RECT 2621.635 209.170 2621.915 210.965 ;
        RECT 2627.620 209.450 2627.880 209.770 ;
        RECT 2621.240 209.030 2621.915 209.170 ;
        RECT 2627.680 209.170 2627.820 209.450 ;
        RECT 2628.075 209.170 2628.355 210.965 ;
        RECT 2634.055 209.170 2634.335 210.965 ;
        RECT 2639.580 209.450 2639.840 209.770 ;
        RECT 2627.680 209.030 2628.355 209.170 ;
        RECT 2633.660 209.090 2634.335 209.170 ;
        RECT 2621.635 208.565 2621.915 209.030 ;
        RECT 2628.075 208.565 2628.355 209.030 ;
        RECT 2633.600 209.030 2634.335 209.090 ;
        RECT 2639.640 209.170 2639.780 209.450 ;
        RECT 2640.035 209.170 2640.315 210.965 ;
        RECT 2643.255 209.170 2643.535 210.965 ;
        RECT 2639.640 209.030 2643.535 209.170 ;
        RECT 2633.600 208.770 2633.860 209.030 ;
        RECT 2634.055 208.565 2634.335 209.030 ;
        RECT 2640.035 208.565 2640.315 209.030 ;
        RECT 2643.255 208.565 2643.535 209.030 ;
        RECT 2649.235 208.565 2649.515 210.965 ;
        RECT 2899.540 209.430 2899.680 213.530 ;
        RECT 2844.280 209.110 2844.540 209.430 ;
        RECT 2899.480 209.110 2899.740 209.430 ;
      LAYER met2 ;
        RECT 1475.085 208.285 1476.135 208.565 ;
        RECT 1476.975 208.285 1479.355 208.565 ;
        RECT 1480.195 208.285 1482.575 208.565 ;
        RECT 1483.415 208.285 1485.335 208.565 ;
        RECT 1486.175 208.285 1488.555 208.565 ;
        RECT 1489.395 208.285 1491.775 208.565 ;
        RECT 1492.615 208.285 1494.535 208.565 ;
        RECT 1495.375 208.285 1497.755 208.565 ;
        RECT 1498.595 208.285 1500.975 208.565 ;
        RECT 1501.815 208.285 1503.735 208.565 ;
        RECT 1504.575 208.285 1506.955 208.565 ;
        RECT 1507.795 208.285 1510.175 208.565 ;
        RECT 1511.015 208.285 1512.935 208.565 ;
        RECT 1513.775 208.285 1516.155 208.565 ;
        RECT 1516.995 208.285 1519.375 208.565 ;
        RECT 1520.215 208.285 1522.595 208.565 ;
        RECT 1523.435 208.285 1525.355 208.565 ;
        RECT 1526.195 208.285 1528.575 208.565 ;
        RECT 1529.415 208.285 1531.795 208.565 ;
        RECT 1532.635 208.285 1534.555 208.565 ;
        RECT 1535.395 208.285 1537.775 208.565 ;
        RECT 1538.615 208.285 1540.995 208.565 ;
        RECT 1541.835 208.285 1543.755 208.565 ;
        RECT 1544.595 208.285 1546.975 208.565 ;
        RECT 1547.815 208.285 1550.195 208.565 ;
        RECT 1551.035 208.285 1552.955 208.565 ;
        RECT 1553.795 208.285 1554.790 208.565 ;
      LAYER met2 ;
        RECT 1281.190 197.355 1281.470 197.725 ;
      LAYER met2 ;
        RECT 1194.860 153.765 1280.500 158.415 ;
        RECT 1206.000 3.570 1280.500 153.765 ;
        RECT 1475.085 0.000 1554.790 208.285 ;
        RECT 1749.085 208.285 1750.135 208.565 ;
        RECT 1750.975 208.285 1753.355 208.565 ;
        RECT 1754.195 208.285 1756.575 208.565 ;
        RECT 1757.415 208.285 1759.335 208.565 ;
        RECT 1760.175 208.285 1762.555 208.565 ;
        RECT 1763.395 208.285 1765.775 208.565 ;
        RECT 1766.615 208.285 1768.535 208.565 ;
        RECT 1769.375 208.285 1771.755 208.565 ;
        RECT 1772.595 208.285 1774.975 208.565 ;
        RECT 1775.815 208.285 1777.735 208.565 ;
        RECT 1778.575 208.285 1780.955 208.565 ;
        RECT 1781.795 208.285 1784.175 208.565 ;
        RECT 1785.015 208.285 1786.935 208.565 ;
        RECT 1787.775 208.285 1790.155 208.565 ;
        RECT 1790.995 208.285 1793.375 208.565 ;
        RECT 1794.215 208.285 1796.595 208.565 ;
        RECT 1797.435 208.285 1799.355 208.565 ;
        RECT 1800.195 208.285 1802.575 208.565 ;
        RECT 1803.415 208.285 1805.795 208.565 ;
        RECT 1806.635 208.285 1808.555 208.565 ;
        RECT 1809.395 208.285 1811.775 208.565 ;
        RECT 1812.615 208.285 1814.995 208.565 ;
        RECT 1815.835 208.285 1817.755 208.565 ;
        RECT 1818.595 208.285 1820.975 208.565 ;
        RECT 1821.815 208.285 1824.195 208.565 ;
        RECT 1825.035 208.285 1826.955 208.565 ;
        RECT 1827.795 208.285 1828.790 208.565 ;
        RECT 1749.085 0.000 1828.790 208.285 ;
        RECT 2023.085 208.285 2024.135 208.565 ;
        RECT 2024.975 208.285 2027.355 208.565 ;
        RECT 2028.195 208.285 2030.575 208.565 ;
        RECT 2031.415 208.285 2033.335 208.565 ;
        RECT 2034.175 208.285 2036.555 208.565 ;
        RECT 2037.395 208.285 2039.775 208.565 ;
        RECT 2040.615 208.285 2042.535 208.565 ;
        RECT 2043.375 208.285 2045.755 208.565 ;
        RECT 2046.595 208.285 2048.975 208.565 ;
        RECT 2049.815 208.285 2051.735 208.565 ;
        RECT 2052.575 208.285 2054.955 208.565 ;
        RECT 2055.795 208.285 2058.175 208.565 ;
        RECT 2059.015 208.285 2060.935 208.565 ;
        RECT 2061.775 208.285 2064.155 208.565 ;
        RECT 2064.995 208.285 2067.375 208.565 ;
        RECT 2068.215 208.285 2070.595 208.565 ;
        RECT 2071.435 208.285 2073.355 208.565 ;
        RECT 2074.195 208.285 2076.575 208.565 ;
        RECT 2077.415 208.285 2079.795 208.565 ;
        RECT 2080.635 208.285 2082.555 208.565 ;
        RECT 2083.395 208.285 2085.775 208.565 ;
        RECT 2086.615 208.285 2088.995 208.565 ;
        RECT 2089.835 208.285 2091.755 208.565 ;
        RECT 2092.595 208.285 2094.975 208.565 ;
        RECT 2095.815 208.285 2098.195 208.565 ;
        RECT 2099.035 208.285 2100.955 208.565 ;
        RECT 2101.795 208.285 2102.790 208.565 ;
        RECT 2023.085 0.000 2102.790 208.285 ;
        RECT 2297.085 208.285 2298.135 208.565 ;
        RECT 2298.975 208.285 2301.355 208.565 ;
        RECT 2302.195 208.285 2304.575 208.565 ;
        RECT 2305.415 208.285 2307.335 208.565 ;
        RECT 2308.175 208.285 2310.555 208.565 ;
        RECT 2311.395 208.285 2313.775 208.565 ;
        RECT 2314.615 208.285 2316.535 208.565 ;
        RECT 2317.375 208.285 2319.755 208.565 ;
        RECT 2320.595 208.285 2322.975 208.565 ;
        RECT 2323.815 208.285 2325.735 208.565 ;
        RECT 2326.575 208.285 2328.955 208.565 ;
        RECT 2329.795 208.285 2332.175 208.565 ;
        RECT 2333.015 208.285 2334.935 208.565 ;
        RECT 2335.775 208.285 2338.155 208.565 ;
        RECT 2338.995 208.285 2341.375 208.565 ;
        RECT 2342.215 208.285 2344.595 208.565 ;
        RECT 2345.435 208.285 2347.355 208.565 ;
        RECT 2348.195 208.285 2350.575 208.565 ;
        RECT 2351.415 208.285 2353.795 208.565 ;
        RECT 2354.635 208.285 2356.555 208.565 ;
        RECT 2357.395 208.285 2359.775 208.565 ;
        RECT 2360.615 208.285 2362.995 208.565 ;
        RECT 2363.835 208.285 2365.755 208.565 ;
        RECT 2366.595 208.285 2368.975 208.565 ;
        RECT 2369.815 208.285 2372.195 208.565 ;
        RECT 2373.035 208.285 2374.955 208.565 ;
        RECT 2375.795 208.285 2376.790 208.565 ;
        RECT 2297.085 0.000 2376.790 208.285 ;
        RECT 2571.085 208.285 2572.135 208.565 ;
        RECT 2572.975 208.285 2575.355 208.565 ;
        RECT 2576.195 208.285 2578.575 208.565 ;
        RECT 2579.415 208.285 2581.335 208.565 ;
        RECT 2582.175 208.285 2584.555 208.565 ;
        RECT 2585.395 208.285 2587.775 208.565 ;
        RECT 2588.615 208.285 2590.535 208.565 ;
        RECT 2591.375 208.285 2593.755 208.565 ;
        RECT 2594.595 208.285 2596.975 208.565 ;
        RECT 2597.815 208.285 2599.735 208.565 ;
        RECT 2600.575 208.285 2602.955 208.565 ;
        RECT 2603.795 208.285 2606.175 208.565 ;
        RECT 2607.015 208.285 2608.935 208.565 ;
        RECT 2609.775 208.285 2612.155 208.565 ;
        RECT 2612.995 208.285 2615.375 208.565 ;
        RECT 2616.215 208.285 2618.595 208.565 ;
        RECT 2619.435 208.285 2621.355 208.565 ;
        RECT 2622.195 208.285 2624.575 208.565 ;
        RECT 2625.415 208.285 2627.795 208.565 ;
        RECT 2628.635 208.285 2630.555 208.565 ;
        RECT 2631.395 208.285 2633.775 208.565 ;
        RECT 2634.615 208.285 2636.995 208.565 ;
        RECT 2637.835 208.285 2639.755 208.565 ;
        RECT 2640.595 208.285 2642.975 208.565 ;
        RECT 2643.815 208.285 2646.195 208.565 ;
        RECT 2647.035 208.285 2648.955 208.565 ;
        RECT 2649.795 208.285 2650.790 208.565 ;
        RECT 2571.085 0.000 2650.790 208.285 ;
      LAYER met2 ;
        RECT 2844.340 198.405 2844.480 209.110 ;
        RECT 2844.270 198.035 2844.550 198.405 ;
      LAYER met2 ;
        RECT 2845.710 197.965 2869.610 200.000 ;
        RECT 2892.105 198.080 2894.105 200.000 ;
        RECT 2895.605 197.965 2919.505 200.000 ;
        RECT 3114.710 197.965 3138.610 200.000 ;
        RECT 3161.105 198.080 3163.105 200.000 ;
        RECT 3164.605 197.965 3188.505 200.000 ;
        RECT 2845.710 4.925 2919.735 197.965 ;
        RECT 3114.710 4.925 3188.735 197.965 ;
      LAYER via2 ;
        RECT 2928.910 4987.320 2929.190 4987.600 ;
        RECT 1697.490 4985.280 1697.770 4985.560 ;
        RECT 220.890 4429.040 221.170 4429.320 ;
        RECT 224.110 4429.040 224.390 4429.320 ;
        RECT 220.890 4354.920 221.170 4355.200 ;
        RECT 3387.990 4019.000 3388.270 4019.280 ;
        RECT 3389.830 2474.040 3390.110 2474.320 ;
        RECT 3370.050 2099.360 3370.330 2099.640 ;
        RECT 3370.050 2095.960 3370.330 2096.240 ;
        RECT 3387.530 2091.880 3387.810 2092.160 ;
        RECT 198.350 400.720 198.630 401.000 ;
        RECT 198.350 391.200 198.630 391.480 ;
        RECT 220.890 552.360 221.170 552.640 ;
        RECT 224.110 552.360 224.390 552.640 ;
        RECT 220.890 400.720 221.170 401.000 ;
        RECT 224.110 400.720 224.390 401.000 ;
        RECT 468.830 200.800 469.110 201.080 ;
        RECT 675.830 200.800 676.110 201.080 ;
        RECT 758.630 234.120 758.910 234.400 ;
        RECT 942.630 234.120 942.910 234.400 ;
        RECT 717.690 202.160 717.970 202.440 ;
        RECT 715.390 200.800 715.670 201.080 ;
        RECT 717.690 200.800 717.970 201.080 ;
        RECT 758.630 202.160 758.910 202.440 ;
        RECT 2024.550 221.200 2024.830 221.480 ;
        RECT 2064.570 221.200 2064.850 221.480 ;
        RECT 2298.250 221.200 2298.530 221.480 ;
        RECT 2338.270 221.200 2338.550 221.480 ;
        RECT 2572.410 221.200 2572.690 221.480 ;
        RECT 2612.430 221.880 2612.710 222.160 ;
        RECT 3368.670 502.720 3368.950 503.000 ;
        RECT 3376.950 502.720 3377.230 503.000 ;
        RECT 1281.190 197.400 1281.470 197.680 ;
        RECT 2844.270 198.080 2844.550 198.360 ;
      LAYER met3 ;
        RECT 375.455 5070.750 449.250 5161.315 ;
        RECT 375.455 5002.905 399.320 5070.750 ;
        RECT 425.120 5002.905 449.250 5070.750 ;
        RECT 615.455 5070.750 689.250 5161.315 ;
        RECT 615.455 5002.905 639.320 5070.750 ;
        RECT 665.120 5002.905 689.250 5070.750 ;
        RECT 855.455 5070.750 929.250 5161.315 ;
        RECT 855.455 5002.905 879.320 5070.750 ;
        RECT 905.120 5002.905 929.250 5070.750 ;
        RECT 1100.000 5004.085 1269.000 5188.000 ;
        RECT 1357.000 5004.085 1526.000 5188.000 ;
        RECT 1697.240 5014.250 1771.290 5188.000 ;
        RECT 2124.455 5070.750 2198.250 5161.315 ;
      LAYER met3 ;
        RECT 1100.000 4988.000 1171.395 5003.685 ;
      LAYER met3 ;
        RECT 1171.795 4999.730 1196.990 5004.085 ;
        RECT 1171.795 4991.125 1184.490 4999.730 ;
        RECT 1171.795 4990.725 1172.495 4991.125 ;
        RECT 1184.295 4990.725 1184.490 4991.125 ;
      LAYER met3 ;
        RECT 1172.895 4988.000 1183.895 4990.725 ;
        RECT 1184.890 4988.000 1195.890 4999.330 ;
      LAYER met3 ;
        RECT 1196.290 4990.725 1196.990 4999.730 ;
      LAYER met3 ;
        RECT 1357.000 4988.000 1428.395 5003.685 ;
      LAYER met3 ;
        RECT 1428.795 4999.730 1453.990 5004.085 ;
        RECT 1428.795 4991.125 1441.490 4999.730 ;
        RECT 1428.795 4990.725 1429.495 4991.125 ;
        RECT 1441.295 4990.725 1441.490 4991.125 ;
      LAYER met3 ;
        RECT 1429.895 4988.000 1440.895 4990.725 ;
        RECT 1441.890 4988.000 1452.890 4999.330 ;
      LAYER met3 ;
        RECT 1453.290 4990.725 1453.990 4999.730 ;
      LAYER met3 ;
        RECT 1697.495 4988.000 1721.395 5013.850 ;
      LAYER met3 ;
        RECT 1721.795 4990.035 1746.990 5014.250 ;
        RECT 1722.895 4988.000 1733.895 4990.035 ;
        RECT 1734.890 4988.000 1745.890 4990.035 ;
      LAYER met3 ;
        RECT 1747.390 4988.000 1771.290 5013.850 ;
      LAYER met3 ;
        RECT 2124.455 5002.905 2148.320 5070.750 ;
        RECT 2174.120 5002.905 2198.250 5070.750 ;
        RECT 2371.455 5070.750 2445.250 5161.315 ;
        RECT 2371.455 5002.905 2395.320 5070.750 ;
        RECT 2421.120 5002.905 2445.250 5070.750 ;
        RECT 2629.455 5070.750 2703.250 5161.315 ;
        RECT 2629.455 5002.905 2653.320 5070.750 ;
        RECT 2679.120 5002.905 2703.250 5070.750 ;
        RECT 2878.240 5025.160 2952.290 5183.100 ;
        RECT 3135.455 5070.750 3209.250 5161.315 ;
        RECT 2878.240 5020.915 2927.990 5025.160 ;
      LAYER met3 ;
        RECT 2878.495 4988.000 2902.395 5020.515 ;
      LAYER met3 ;
        RECT 2902.795 4990.035 2927.990 5020.915 ;
        RECT 2903.895 4988.000 2914.895 4990.035 ;
        RECT 2915.890 4988.000 2926.890 4990.035 ;
      LAYER met3 ;
        RECT 2928.390 4988.000 2952.290 5024.760 ;
      LAYER met3 ;
        RECT 3135.455 5002.905 3159.320 5070.750 ;
        RECT 3185.120 5002.905 3209.250 5070.750 ;
      LAYER met3 ;
        RECT 1697.710 4985.585 1698.010 4988.000 ;
        RECT 2928.670 4987.625 2928.970 4988.000 ;
        RECT 2928.670 4987.310 2929.215 4987.625 ;
        RECT 2928.885 4987.295 2929.215 4987.310 ;
        RECT 1697.465 4985.270 1698.010 4985.585 ;
        RECT 1697.465 4985.255 1697.795 4985.270 ;
      LAYER met3 ;
        RECT 26.685 4826.120 185.095 4850.250 ;
        RECT 26.685 4800.320 117.250 4826.120 ;
        RECT 26.685 4776.455 185.095 4800.320 ;
      LAYER met3 ;
        RECT 3388.000 4770.605 3403.685 4842.000 ;
      LAYER met3 ;
        RECT 3404.085 4770.205 3588.000 4842.000 ;
        RECT 3390.725 4769.505 3588.000 4770.205 ;
      LAYER met3 ;
        RECT 3388.000 4758.105 3390.725 4769.105 ;
      LAYER met3 ;
        RECT 3391.125 4757.705 3588.000 4769.505 ;
        RECT 3390.725 4757.510 3588.000 4757.705 ;
      LAYER met3 ;
        RECT 3388.000 4746.110 3399.330 4757.110 ;
      LAYER met3 ;
        RECT 3399.730 4745.710 3588.000 4757.510 ;
        RECT 3390.725 4745.010 3588.000 4745.710 ;
        RECT 3404.085 4673.000 3588.000 4745.010 ;
        RECT 0.035 4641.200 24.250 4650.935 ;
        RECT 153.765 4640.605 158.415 4651.140 ;
        RECT 169.550 4641.200 174.200 4650.935 ;
        RECT 0.035 4615.355 190.700 4640.000 ;
      LAYER met3 ;
        RECT 191.100 4615.755 198.000 4639.700 ;
      LAYER met3 ;
        RECT 0.035 4614.255 197.965 4615.355 ;
        RECT 0.035 4603.380 198.000 4614.255 ;
        RECT 0.035 4601.880 197.965 4603.380 ;
        RECT 0.035 4591.000 198.000 4601.880 ;
        RECT 0.035 4589.900 197.965 4591.000 ;
        RECT 0.035 4565.100 190.700 4589.900 ;
      LAYER met3 ;
        RECT 191.100 4565.500 198.000 4589.500 ;
      LAYER met3 ;
        RECT 0.035 4565.000 197.965 4565.100 ;
        RECT 153.800 4554.025 158.450 4564.105 ;
        RECT 3429.550 4532.895 3434.200 4542.975 ;
        RECT 3390.035 4531.900 3587.965 4532.000 ;
      LAYER met3 ;
        RECT 3390.000 4507.500 3396.900 4531.500 ;
      LAYER met3 ;
        RECT 3397.300 4507.100 3587.965 4531.900 ;
        RECT 3390.035 4506.000 3587.965 4507.100 ;
        RECT 3390.000 4495.120 3587.965 4506.000 ;
        RECT 3390.035 4493.620 3587.965 4495.120 ;
        RECT 3390.000 4482.745 3587.965 4493.620 ;
        RECT 3390.035 4481.645 3587.965 4482.745 ;
      LAYER met3 ;
        RECT 3390.000 4457.300 3396.900 4481.245 ;
      LAYER met3 ;
        RECT 3397.300 4457.000 3587.965 4481.645 ;
        RECT 3413.800 4446.065 3418.450 4455.800 ;
        RECT 3429.585 4445.860 3434.235 4456.395 ;
        RECT 3563.750 4446.065 3587.965 4455.800 ;
      LAYER met3 ;
        RECT 220.865 4429.330 221.195 4429.345 ;
        RECT 224.085 4429.330 224.415 4429.345 ;
        RECT 220.865 4429.030 224.415 4429.330 ;
        RECT 220.865 4429.015 221.195 4429.030 ;
        RECT 224.085 4429.015 224.415 4429.030 ;
      LAYER met3 ;
        RECT 0.000 4403.990 179.800 4428.290 ;
      LAYER met3 ;
        RECT 180.200 4404.390 200.000 4428.290 ;
      LAYER met3 ;
        RECT 0.000 4402.890 197.965 4403.990 ;
        RECT 0.000 4391.890 200.000 4402.890 ;
        RECT 0.000 4390.895 197.965 4391.890 ;
        RECT 0.000 4379.895 200.000 4390.895 ;
        RECT 0.000 4378.795 197.965 4379.895 ;
        RECT 0.000 4354.240 179.800 4378.795 ;
      LAYER met3 ;
        RECT 180.200 4355.210 200.000 4378.395 ;
        RECT 220.865 4355.210 221.195 4355.225 ;
        RECT 180.200 4354.910 221.195 4355.210 ;
        RECT 180.200 4354.495 200.000 4354.910 ;
        RECT 220.865 4354.895 221.195 4354.910 ;
      LAYER met3 ;
        RECT 3386.690 4235.430 3588.000 4314.690 ;
        RECT 4.900 4191.990 162.840 4216.290 ;
      LAYER met3 ;
        RECT 163.240 4192.390 200.000 4216.290 ;
      LAYER met3 ;
        RECT 4.900 4190.890 197.965 4191.990 ;
        RECT 4.900 4179.890 200.000 4190.890 ;
        RECT 4.900 4178.895 197.965 4179.890 ;
        RECT 4.900 4167.895 200.000 4178.895 ;
        RECT 4.900 4166.795 197.965 4167.895 ;
        RECT 4.900 4142.240 167.085 4166.795 ;
      LAYER met3 ;
        RECT 167.485 4142.495 200.000 4166.395 ;
        RECT 3388.000 4069.605 3402.960 4093.505 ;
      LAYER met3 ;
        RECT 3403.360 4069.205 3588.000 4093.760 ;
        RECT 3390.035 4068.105 3588.000 4069.205 ;
        RECT 3388.000 4057.105 3588.000 4068.105 ;
        RECT 3390.035 4056.110 3588.000 4057.105 ;
        RECT 3388.000 4045.110 3588.000 4056.110 ;
        RECT 3390.035 4044.010 3588.000 4045.110 ;
      LAYER met3 ;
        RECT 3388.000 4019.710 3402.960 4043.610 ;
      LAYER met3 ;
        RECT 3403.360 4019.710 3588.000 4044.010 ;
      LAYER met3 ;
        RECT 3387.965 4019.290 3388.295 4019.305 ;
        RECT 3388.670 4019.290 3388.970 4019.710 ;
        RECT 3387.965 4018.990 3388.970 4019.290 ;
        RECT 3387.965 4018.975 3388.295 4018.990 ;
      LAYER met3 ;
        RECT 0.000 3926.310 201.310 4005.570 ;
        RECT 3386.690 3798.430 3588.000 3877.690 ;
        RECT 0.000 3710.310 201.310 3789.570 ;
        RECT 3386.690 3576.430 3588.000 3655.690 ;
        RECT 0.000 3494.310 201.310 3573.570 ;
        RECT 0.000 3277.310 201.310 3356.570 ;
        RECT 3386.690 3355.430 3588.000 3434.690 ;
        RECT 0.000 3061.310 201.310 3140.570 ;
        RECT 3386.690 3134.430 3588.000 3213.690 ;
        RECT 0.000 2845.310 201.310 2924.570 ;
        RECT 3386.690 2912.430 3588.000 2991.690 ;
        RECT 0.000 2629.310 201.310 2708.570 ;
        RECT 3386.690 2691.430 3588.000 2770.690 ;
      LAYER met3 ;
        RECT 3388.000 2525.605 3402.960 2549.505 ;
      LAYER met3 ;
        RECT 3403.360 2525.205 3588.000 2549.760 ;
        RECT 3390.035 2524.105 3588.000 2525.205 ;
        RECT 3388.000 2513.105 3588.000 2524.105 ;
        RECT 3390.035 2512.110 3588.000 2513.105 ;
        RECT 3388.000 2501.110 3588.000 2512.110 ;
        RECT 3390.035 2500.010 3588.000 2501.110 ;
        RECT 0.000 2466.990 184.640 2491.290 ;
      LAYER met3 ;
        RECT 185.040 2467.390 200.000 2491.290 ;
        RECT 3388.000 2475.710 3402.960 2499.610 ;
      LAYER met3 ;
        RECT 3403.360 2475.710 3588.000 2500.010 ;
      LAYER met3 ;
        RECT 3389.590 2474.345 3389.890 2475.710 ;
        RECT 3389.590 2474.030 3390.135 2474.345 ;
        RECT 3389.805 2474.015 3390.135 2474.030 ;
      LAYER met3 ;
        RECT 0.000 2465.890 197.965 2466.990 ;
        RECT 0.000 2454.890 200.000 2465.890 ;
        RECT 0.000 2453.895 197.965 2454.890 ;
        RECT 0.000 2442.895 200.000 2453.895 ;
        RECT 0.000 2441.795 197.965 2442.895 ;
        RECT 0.000 2417.240 184.640 2441.795 ;
      LAYER met3 ;
        RECT 185.040 2417.495 200.000 2441.395 ;
      LAYER met3 ;
        RECT 3429.550 2333.895 3434.200 2343.975 ;
        RECT 3390.035 2332.900 3587.965 2333.000 ;
        RECT 3430.000 2308.100 3587.965 2332.900 ;
        RECT 3390.035 2307.000 3587.965 2308.100 ;
        RECT 3390.000 2296.120 3587.965 2307.000 ;
        RECT 3390.035 2294.620 3587.965 2296.120 ;
        RECT 0.035 2282.200 24.250 2291.935 ;
        RECT 153.765 2281.605 158.415 2292.140 ;
        RECT 169.550 2282.200 174.200 2291.935 ;
        RECT 3390.000 2283.745 3587.965 2294.620 ;
        RECT 3390.035 2282.645 3587.965 2283.745 ;
        RECT 0.035 2256.355 158.000 2281.000 ;
      LAYER met3 ;
        RECT 158.400 2256.755 198.000 2280.700 ;
        RECT 3390.000 2258.300 3429.600 2282.245 ;
      LAYER met3 ;
        RECT 3430.000 2258.000 3587.965 2282.645 ;
        RECT 0.035 2255.255 197.965 2256.355 ;
        RECT 0.035 2244.380 198.000 2255.255 ;
        RECT 3413.800 2247.065 3418.450 2256.800 ;
        RECT 3429.585 2246.860 3434.235 2257.395 ;
        RECT 3563.750 2247.065 3587.965 2256.800 ;
        RECT 0.035 2242.880 197.965 2244.380 ;
        RECT 0.035 2232.000 198.000 2242.880 ;
        RECT 0.035 2230.900 197.965 2232.000 ;
        RECT 0.035 2206.100 158.000 2230.900 ;
        RECT 0.035 2206.000 197.965 2206.100 ;
        RECT 153.800 2195.025 158.450 2205.105 ;
      LAYER met3 ;
        RECT 3369.310 2099.650 3369.690 2099.660 ;
        RECT 3370.025 2099.650 3370.355 2099.665 ;
        RECT 3369.310 2099.350 3370.355 2099.650 ;
        RECT 3369.310 2099.340 3369.690 2099.350 ;
        RECT 3370.025 2099.335 3370.355 2099.350 ;
        RECT 3369.310 2096.250 3369.690 2096.260 ;
        RECT 3370.025 2096.250 3370.355 2096.265 ;
        RECT 3369.310 2095.950 3370.355 2096.250 ;
        RECT 3369.310 2095.940 3369.690 2095.950 ;
        RECT 3370.025 2095.935 3370.355 2095.950 ;
        RECT 3388.000 2092.605 3420.515 2116.505 ;
        RECT 3387.505 2092.170 3387.835 2092.185 ;
        RECT 3388.670 2092.170 3388.970 2092.605 ;
      LAYER met3 ;
        RECT 3420.915 2092.205 3583.100 2116.760 ;
      LAYER met3 ;
        RECT 3387.505 2091.870 3388.970 2092.170 ;
        RECT 3387.505 2091.855 3387.835 2091.870 ;
      LAYER met3 ;
        RECT 3390.035 2091.105 3583.100 2092.205 ;
        RECT 3388.000 2080.105 3583.100 2091.105 ;
        RECT 3390.035 2079.110 3583.100 2080.105 ;
        RECT 0.000 1990.310 201.310 2069.570 ;
        RECT 3388.000 2068.110 3583.100 2079.110 ;
        RECT 3390.035 2067.010 3583.100 2068.110 ;
      LAYER met3 ;
        RECT 3388.000 2042.710 3424.760 2066.610 ;
      LAYER met3 ;
        RECT 3425.160 2042.710 3583.100 2067.010 ;
        RECT 0.000 1774.310 201.310 1853.570 ;
        RECT 3386.690 1820.430 3588.000 1899.690 ;
        RECT 0.000 1557.310 201.310 1636.570 ;
        RECT 3386.690 1599.430 3588.000 1678.690 ;
        RECT 0.000 1341.310 201.310 1420.570 ;
        RECT 3386.690 1378.430 3588.000 1457.690 ;
        RECT 0.000 1125.310 201.310 1204.570 ;
        RECT 3386.690 1156.430 3588.000 1235.690 ;
        RECT 0.000 909.310 201.310 988.570 ;
        RECT 3386.690 935.430 3588.000 1014.690 ;
        RECT 3386.690 714.430 3588.000 793.690 ;
        RECT 0.000 600.990 179.800 625.290 ;
      LAYER met3 ;
        RECT 180.200 601.390 200.000 625.290 ;
      LAYER met3 ;
        RECT 0.000 599.890 197.965 600.990 ;
        RECT 0.000 588.890 200.000 599.890 ;
        RECT 0.000 587.895 197.965 588.890 ;
        RECT 0.000 576.895 200.000 587.895 ;
        RECT 0.000 575.795 197.965 576.895 ;
        RECT 0.000 551.240 179.800 575.795 ;
      LAYER met3 ;
        RECT 180.200 552.650 200.000 575.395 ;
        RECT 220.865 552.650 221.195 552.665 ;
        RECT 224.085 552.650 224.415 552.665 ;
        RECT 180.200 552.350 224.415 552.650 ;
        RECT 180.200 551.495 200.000 552.350 ;
        RECT 220.865 552.335 221.195 552.350 ;
        RECT 224.085 552.335 224.415 552.350 ;
        RECT 3368.645 503.010 3368.975 503.025 ;
        RECT 3376.925 503.010 3377.255 503.025 ;
        RECT 3368.645 502.710 3377.255 503.010 ;
        RECT 3368.645 502.695 3368.975 502.710 ;
        RECT 3376.925 502.695 3377.255 502.710 ;
      LAYER met3 ;
        RECT 3386.690 492.430 3588.000 571.690 ;
        RECT 153.765 415.605 158.415 426.140 ;
        RECT 159.805 415.440 163.270 426.140 ;
        RECT 4.395 390.355 190.700 415.000 ;
      LAYER met3 ;
        RECT 191.100 391.490 198.000 414.700 ;
        RECT 198.325 401.010 198.655 401.025 ;
        RECT 220.865 401.010 221.195 401.025 ;
        RECT 224.085 401.010 224.415 401.025 ;
        RECT 198.325 400.710 224.415 401.010 ;
        RECT 198.325 400.695 198.655 400.710 ;
        RECT 220.865 400.695 221.195 400.710 ;
        RECT 224.085 400.695 224.415 400.710 ;
        RECT 198.325 391.490 198.655 391.505 ;
        RECT 191.100 391.190 198.655 391.490 ;
        RECT 191.100 390.755 198.000 391.190 ;
        RECT 198.325 391.175 198.655 391.190 ;
      LAYER met3 ;
        RECT 4.395 389.255 197.965 390.355 ;
        RECT 4.395 378.380 198.000 389.255 ;
        RECT 4.395 376.880 197.965 378.380 ;
        RECT 4.395 366.000 198.000 376.880 ;
        RECT 4.395 364.900 197.965 366.000 ;
        RECT 4.395 340.490 190.700 364.900 ;
      LAYER met3 ;
        RECT 191.100 340.500 198.000 364.500 ;
        RECT 758.605 234.410 758.935 234.425 ;
        RECT 942.605 234.410 942.935 234.425 ;
        RECT 758.605 234.110 942.935 234.410 ;
        RECT 758.605 234.095 758.935 234.110 ;
        RECT 942.605 234.095 942.935 234.110 ;
        RECT 2612.405 222.170 2612.735 222.185 ;
        RECT 2580.450 221.870 2612.735 222.170 ;
        RECT 2024.525 221.490 2024.855 221.505 ;
        RECT 2064.545 221.490 2064.875 221.505 ;
        RECT 2024.525 221.190 2064.875 221.490 ;
        RECT 2024.525 221.175 2024.855 221.190 ;
        RECT 2064.545 221.175 2064.875 221.190 ;
        RECT 2298.225 221.490 2298.555 221.505 ;
        RECT 2338.245 221.490 2338.575 221.505 ;
        RECT 2298.225 221.190 2338.575 221.490 ;
        RECT 2298.225 221.175 2298.555 221.190 ;
        RECT 2338.245 221.175 2338.575 221.190 ;
        RECT 2572.385 221.490 2572.715 221.505 ;
        RECT 2580.450 221.490 2580.750 221.870 ;
        RECT 2612.405 221.855 2612.735 221.870 ;
        RECT 2572.385 221.190 2580.750 221.490 ;
        RECT 2572.385 221.175 2572.715 221.190 ;
        RECT 717.665 202.450 717.995 202.465 ;
        RECT 758.605 202.450 758.935 202.465 ;
        RECT 717.665 202.150 758.935 202.450 ;
        RECT 717.665 202.135 717.995 202.150 ;
        RECT 728.950 201.770 729.250 202.150 ;
        RECT 758.605 202.135 758.935 202.150 ;
        RECT 728.950 201.470 729.490 201.770 ;
        RECT 468.805 201.090 469.135 201.105 ;
        RECT 675.805 201.090 676.135 201.105 ;
        RECT 455.710 200.790 469.135 201.090 ;
        RECT 455.710 200.000 456.010 200.790 ;
        RECT 468.805 200.775 469.135 200.790 ;
        RECT 665.470 200.790 676.135 201.090 ;
        RECT 665.470 200.000 665.770 200.790 ;
        RECT 675.805 200.775 676.135 200.790 ;
        RECT 715.365 201.090 715.695 201.105 ;
        RECT 717.665 201.090 717.995 201.105 ;
        RECT 715.365 200.790 717.290 201.090 ;
        RECT 715.365 200.775 715.695 200.790 ;
        RECT 716.990 200.000 717.290 200.790 ;
        RECT 717.665 200.790 720.050 201.090 ;
        RECT 717.665 200.775 717.995 200.790 ;
        RECT 719.750 200.000 720.050 200.790 ;
        RECT 729.190 200.070 729.490 201.470 ;
        RECT 729.100 200.000 729.490 200.070 ;
        RECT 238.000 164.765 256.010 180.085 ;
        RECT 258.000 164.765 276.010 180.085 ;
        RECT 278.000 164.765 296.010 180.085 ;
        RECT 298.000 164.765 316.010 180.085 ;
        RECT 318.000 164.765 336.010 180.085 ;
        RECT 338.000 164.765 356.010 180.085 ;
        RECT 394.710 163.240 418.610 200.000 ;
      LAYER met3 ;
        RECT 420.110 197.965 431.110 200.000 ;
        RECT 432.105 197.965 443.105 200.000 ;
        RECT 419.010 167.085 444.205 197.965 ;
      LAYER met3 ;
        RECT 444.605 167.485 468.505 200.000 ;
      LAYER met3 ;
        RECT 419.010 162.840 468.760 167.085 ;
      LAYER met3 ;
        RECT 507.000 164.765 525.010 180.085 ;
        RECT 527.000 164.765 545.010 180.085 ;
        RECT 547.000 164.765 565.010 180.085 ;
        RECT 567.000 164.765 585.010 180.085 ;
        RECT 587.000 164.765 605.010 180.085 ;
        RECT 607.000 164.765 625.010 180.085 ;
      LAYER met3 ;
        RECT 394.710 4.900 468.760 162.840 ;
        RECT 663.300 151.080 664.340 199.375 ;
        RECT 663.300 133.400 663.675 151.080 ;
      LAYER met3 ;
        RECT 664.740 150.680 665.810 200.000 ;
        RECT 664.075 135.400 665.810 150.680 ;
      LAYER met3 ;
        RECT 666.210 188.690 707.935 199.375 ;
        RECT 709.465 193.730 716.375 199.375 ;
        RECT 709.465 192.265 714.910 193.730 ;
      LAYER met3 ;
        RECT 716.775 193.330 717.925 200.000 ;
      LAYER met3 ;
        RECT 709.465 191.985 714.630 192.265 ;
        RECT 709.465 190.555 713.550 191.985 ;
      LAYER met3 ;
        RECT 715.310 191.950 717.925 193.330 ;
        RECT 715.310 191.865 716.875 191.950 ;
        RECT 716.940 191.865 717.925 191.950 ;
      LAYER met3 ;
        RECT 718.325 196.465 718.690 199.375 ;
      LAYER met3 ;
        RECT 719.090 196.865 720.755 200.000 ;
      LAYER met3 ;
        RECT 721.155 196.465 728.680 199.375 ;
      LAYER met3 ;
        RECT 715.030 191.800 715.310 191.865 ;
        RECT 715.395 191.800 716.940 191.865 ;
        RECT 715.030 191.650 716.940 191.800 ;
        RECT 715.030 191.585 716.575 191.650 ;
        RECT 716.660 191.585 716.940 191.650 ;
      LAYER met3 ;
        RECT 709.765 190.255 713.550 190.555 ;
        RECT 666.210 184.830 708.700 188.690 ;
        RECT 710.230 187.335 713.550 190.255 ;
      LAYER met3 ;
        RECT 713.950 191.500 715.030 191.585 ;
        RECT 715.095 191.500 716.660 191.585 ;
        RECT 713.950 190.020 716.660 191.500 ;
      LAYER met3 ;
        RECT 718.325 191.465 728.680 196.465 ;
        RECT 717.340 191.185 728.680 191.465 ;
      LAYER met3 ;
        RECT 713.950 187.735 715.095 190.020 ;
      LAYER met3 ;
        RECT 717.060 189.620 728.680 191.185 ;
        RECT 715.495 187.335 728.680 189.620 ;
        RECT 710.230 184.830 728.680 187.335 ;
        RECT 666.210 183.015 728.680 184.830 ;
      LAYER met3 ;
        RECT 729.080 184.215 729.600 200.000 ;
      LAYER met3 ;
        RECT 730.000 184.615 737.035 199.375 ;
        RECT 730.210 184.405 737.035 184.615 ;
      LAYER met3 ;
        RECT 729.080 184.005 729.810 184.215 ;
        RECT 729.080 183.555 730.260 184.005 ;
      LAYER met3 ;
        RECT 730.660 183.955 737.035 184.405 ;
      LAYER met3 ;
        RECT 729.080 183.415 729.670 183.555 ;
        RECT 729.680 183.415 730.710 183.555 ;
      LAYER met3 ;
        RECT 731.110 183.505 737.035 183.955 ;
      LAYER met3 ;
        RECT 729.670 183.105 730.710 183.415 ;
      LAYER met3 ;
        RECT 666.210 182.555 729.270 183.015 ;
      LAYER met3 ;
        RECT 729.670 182.955 731.225 183.105 ;
      LAYER met3 ;
        RECT 666.210 181.980 729.730 182.555 ;
      LAYER met3 ;
        RECT 730.130 182.380 731.225 182.955 ;
      LAYER met3 ;
        RECT 666.210 169.105 730.305 181.980 ;
        RECT 666.210 168.520 729.720 169.105 ;
      LAYER met3 ;
        RECT 730.705 168.705 731.225 182.380 ;
      LAYER met3 ;
        RECT 666.210 167.805 729.005 168.520 ;
      LAYER met3 ;
        RECT 730.120 168.195 731.225 168.705 ;
        RECT 730.120 168.120 730.775 168.195 ;
        RECT 730.850 168.120 731.225 168.195 ;
        RECT 729.405 168.045 730.120 168.120 ;
        RECT 730.135 168.045 730.850 168.120 ;
      LAYER met3 ;
        RECT 666.210 167.220 728.420 167.805 ;
      LAYER met3 ;
        RECT 729.405 167.445 730.850 168.045 ;
      LAYER met3 ;
        RECT 731.625 167.720 737.035 183.505 ;
      LAYER met3 ;
        RECT 729.405 167.405 730.120 167.445 ;
        RECT 730.135 167.405 730.850 167.445 ;
        RECT 728.820 167.295 729.405 167.405 ;
        RECT 729.445 167.295 730.135 167.405 ;
      LAYER met3 ;
        RECT 666.210 167.005 728.205 167.220 ;
        RECT 666.210 165.475 715.325 167.005 ;
      LAYER met3 ;
        RECT 728.820 166.845 730.135 167.295 ;
      LAYER met3 ;
        RECT 731.250 167.005 737.035 167.720 ;
      LAYER met3 ;
        RECT 728.820 166.820 729.425 166.845 ;
        RECT 729.550 166.820 730.135 166.845 ;
        RECT 728.605 166.695 728.820 166.820 ;
        RECT 728.845 166.695 729.550 166.820 ;
        RECT 728.605 166.605 729.550 166.695 ;
        RECT 715.725 166.305 729.550 166.605 ;
      LAYER met3 ;
        RECT 730.535 166.420 737.035 167.005 ;
      LAYER met3 ;
        RECT 715.725 166.300 728.885 166.305 ;
        RECT 729.030 166.300 729.550 166.305 ;
        RECT 715.725 165.875 729.030 166.300 ;
      LAYER met3 ;
        RECT 729.950 165.900 737.035 166.420 ;
        RECT 729.430 165.475 737.035 165.900 ;
        RECT 666.210 135.800 737.035 165.475 ;
      LAYER met3 ;
        RECT 776.000 164.765 794.010 180.085 ;
        RECT 796.000 164.765 814.010 180.085 ;
        RECT 816.000 164.765 834.010 180.085 ;
        RECT 836.000 164.765 854.010 180.085 ;
        RECT 856.000 164.765 874.010 180.085 ;
        RECT 876.000 164.765 894.010 180.085 ;
        RECT 664.075 133.800 667.410 135.400 ;
      LAYER met3 ;
        RECT 667.810 134.200 737.035 135.800 ;
        RECT 663.300 131.800 665.410 133.400 ;
      LAYER met3 ;
        RECT 665.810 132.400 668.810 133.800 ;
      LAYER met3 ;
        RECT 669.210 132.800 737.035 134.200 ;
      LAYER met3 ;
        RECT 665.810 132.250 669.745 132.400 ;
        RECT 665.810 132.200 667.410 132.250 ;
        RECT 667.510 132.200 669.745 132.250 ;
      LAYER met3 ;
        RECT 663.300 130.515 667.010 131.800 ;
      LAYER met3 ;
        RECT 667.410 131.465 669.745 132.200 ;
      LAYER met3 ;
        RECT 670.145 131.865 737.035 132.800 ;
      LAYER met3 ;
        RECT 667.410 131.350 669.710 131.465 ;
        RECT 669.745 131.350 670.610 131.465 ;
        RECT 667.410 131.050 670.610 131.350 ;
        RECT 667.410 130.915 668.695 131.050 ;
        RECT 668.710 130.915 670.610 131.050 ;
      LAYER met3 ;
        RECT 671.010 131.000 737.035 131.865 ;
      LAYER met3 ;
        RECT 668.695 130.600 670.610 130.915 ;
      LAYER met3 ;
        RECT 663.300 129.565 668.295 130.515 ;
      LAYER met3 ;
        RECT 668.695 130.000 671.960 130.600 ;
        RECT 668.695 129.965 669.645 130.000 ;
        RECT 669.760 129.965 671.960 130.000 ;
      LAYER met3 ;
        RECT 663.300 128.600 669.245 129.565 ;
      LAYER met3 ;
        RECT 669.645 129.250 671.960 129.965 ;
      LAYER met3 ;
        RECT 672.360 129.650 737.035 131.000 ;
      LAYER met3 ;
        RECT 669.645 129.100 673.140 129.250 ;
        RECT 669.645 129.000 670.610 129.100 ;
        RECT 670.660 129.000 673.140 129.100 ;
      LAYER met3 ;
        RECT 663.300 127.390 670.210 128.600 ;
      LAYER met3 ;
        RECT 670.610 127.920 673.140 129.000 ;
        RECT 670.610 127.790 671.820 127.920 ;
        RECT 671.840 127.790 673.140 127.920 ;
        RECT 671.820 127.600 673.140 127.790 ;
      LAYER met3 ;
        RECT 663.300 127.200 671.420 127.390 ;
        RECT 663.300 104.955 671.610 127.200 ;
      LAYER met3 ;
        RECT 672.010 105.355 673.140 127.600 ;
      LAYER met3 ;
        RECT 673.540 104.955 737.035 129.650 ;
        RECT 663.300 0.000 737.035 104.955 ;
        RECT 932.430 0.000 1011.690 201.310 ;
      LAYER met3 ;
        RECT 1050.000 164.765 1068.010 180.085 ;
        RECT 1070.000 164.765 1088.010 180.085 ;
        RECT 1090.000 164.765 1108.010 180.085 ;
        RECT 1110.000 164.765 1128.010 180.085 ;
        RECT 1130.000 164.765 1148.010 180.085 ;
        RECT 1150.000 164.765 1168.010 180.085 ;
      LAYER met3 ;
        RECT 1194.860 159.805 1205.560 163.270 ;
        RECT 1194.860 153.765 1205.395 158.415 ;
      LAYER met3 ;
        RECT 1206.300 158.400 1230.245 198.000 ;
      LAYER met3 ;
        RECT 1231.745 197.965 1242.620 198.000 ;
        RECT 1244.120 197.965 1255.000 198.000 ;
        RECT 1230.645 158.000 1256.100 197.965 ;
      LAYER met3 ;
        RECT 1256.500 197.690 1280.500 198.000 ;
        RECT 1281.165 197.690 1281.495 197.705 ;
        RECT 1256.500 197.390 1281.495 197.690 ;
        RECT 1256.500 158.400 1280.500 197.390 ;
        RECT 1281.165 197.375 1281.495 197.390 ;
        RECT 1319.000 164.765 1337.010 180.085 ;
        RECT 1339.000 164.765 1357.010 180.085 ;
        RECT 1359.000 164.765 1377.010 180.085 ;
        RECT 1379.000 164.765 1397.010 180.085 ;
        RECT 1399.000 164.765 1417.010 180.085 ;
        RECT 1419.000 164.765 1437.010 180.085 ;
      LAYER met3 ;
        RECT 1206.000 4.395 1280.500 158.000 ;
        RECT 1475.430 0.000 1554.690 201.310 ;
      LAYER met3 ;
        RECT 1593.000 164.765 1611.010 180.085 ;
        RECT 1613.000 164.765 1631.010 180.085 ;
        RECT 1633.000 164.765 1651.010 180.085 ;
        RECT 1653.000 164.765 1671.010 180.085 ;
        RECT 1673.000 164.765 1691.010 180.085 ;
        RECT 1693.000 164.765 1711.010 180.085 ;
      LAYER met3 ;
        RECT 1749.430 0.000 1828.690 201.310 ;
      LAYER met3 ;
        RECT 1867.000 164.765 1885.010 180.085 ;
        RECT 1887.000 164.765 1905.010 180.085 ;
        RECT 1907.000 164.765 1925.010 180.085 ;
        RECT 1927.000 164.765 1945.010 180.085 ;
        RECT 1947.000 164.765 1965.010 180.085 ;
        RECT 1967.000 164.765 1985.010 180.085 ;
      LAYER met3 ;
        RECT 2023.430 0.000 2102.690 201.310 ;
      LAYER met3 ;
        RECT 2141.000 164.765 2159.010 180.085 ;
        RECT 2161.000 164.765 2179.010 180.085 ;
        RECT 2181.000 164.765 2199.010 180.085 ;
        RECT 2201.000 164.765 2219.010 180.085 ;
        RECT 2221.000 164.765 2239.010 180.085 ;
        RECT 2241.000 164.765 2259.010 180.085 ;
      LAYER met3 ;
        RECT 2297.430 0.000 2376.690 201.310 ;
      LAYER met3 ;
        RECT 2415.000 164.765 2433.010 180.085 ;
        RECT 2435.000 164.765 2453.010 180.085 ;
        RECT 2455.000 164.765 2473.010 180.085 ;
        RECT 2475.000 164.765 2493.010 180.085 ;
        RECT 2495.000 164.765 2513.010 180.085 ;
        RECT 2515.000 164.765 2533.010 180.085 ;
      LAYER met3 ;
        RECT 2571.430 0.000 2650.690 201.310 ;
      LAYER met3 ;
        RECT 2844.245 198.370 2844.575 198.385 ;
        RECT 2845.710 198.370 2869.610 200.000 ;
        RECT 2844.245 198.070 2869.610 198.370 ;
        RECT 2844.245 198.055 2844.575 198.070 ;
        RECT 2689.000 164.765 2707.010 180.085 ;
        RECT 2709.000 164.765 2727.010 180.085 ;
        RECT 2729.000 164.765 2747.010 180.085 ;
        RECT 2749.000 164.765 2767.010 180.085 ;
        RECT 2769.000 164.765 2787.010 180.085 ;
        RECT 2789.000 164.765 2807.010 180.085 ;
        RECT 2845.710 174.150 2869.610 198.070 ;
      LAYER met3 ;
        RECT 2871.110 197.965 2882.110 200.000 ;
        RECT 2883.105 197.965 2894.105 200.000 ;
        RECT 2870.010 173.750 2895.205 197.965 ;
      LAYER met3 ;
        RECT 2895.605 174.150 2919.505 200.000 ;
        RECT 3114.710 185.040 3138.610 200.000 ;
      LAYER met3 ;
        RECT 3140.110 197.965 3151.110 200.000 ;
        RECT 3152.105 197.965 3163.105 200.000 ;
        RECT 3139.010 184.640 3164.205 197.965 ;
      LAYER met3 ;
        RECT 3164.605 185.040 3188.505 200.000 ;
      LAYER met3 ;
        RECT 2845.710 0.000 2919.760 173.750 ;
      LAYER met3 ;
        RECT 2958.000 164.765 2976.010 180.085 ;
        RECT 2978.000 164.765 2996.010 180.085 ;
        RECT 2998.000 164.765 3016.010 180.085 ;
        RECT 3018.000 164.765 3036.010 180.085 ;
        RECT 3038.000 164.765 3056.010 180.085 ;
        RECT 3058.000 164.765 3076.010 180.085 ;
      LAYER met3 ;
        RECT 3114.710 0.000 3188.760 184.640 ;
      LAYER met3 ;
        RECT 3227.000 164.765 3245.010 180.085 ;
        RECT 3247.000 164.765 3265.010 180.085 ;
        RECT 3267.000 164.765 3285.010 180.085 ;
        RECT 3287.000 164.765 3305.010 180.085 ;
        RECT 3307.000 164.765 3325.010 180.085 ;
        RECT 3327.000 164.765 3345.010 180.085 ;
      LAYER via3 ;
        RECT 3369.340 2099.340 3369.660 2099.660 ;
        RECT 3369.340 2095.940 3369.660 2096.260 ;
        RECT 238.230 175.875 255.720 179.885 ;
        RECT 238.260 164.935 255.910 167.885 ;
        RECT 258.230 175.875 275.720 179.885 ;
        RECT 258.260 164.935 275.910 167.885 ;
        RECT 278.230 175.875 295.720 179.885 ;
        RECT 278.260 164.935 295.910 167.885 ;
        RECT 298.230 175.875 315.720 179.885 ;
        RECT 298.260 164.935 315.910 167.885 ;
        RECT 318.230 175.875 335.720 179.885 ;
        RECT 318.260 164.935 335.910 167.885 ;
        RECT 338.230 175.875 355.720 179.885 ;
        RECT 338.260 164.935 355.910 167.885 ;
        RECT 507.230 175.875 524.720 179.885 ;
        RECT 507.260 164.935 524.910 167.885 ;
        RECT 527.230 175.875 544.720 179.885 ;
        RECT 527.260 164.935 544.910 167.885 ;
        RECT 547.230 175.875 564.720 179.885 ;
        RECT 547.260 164.935 564.910 167.885 ;
        RECT 567.230 175.875 584.720 179.885 ;
        RECT 567.260 164.935 584.910 167.885 ;
        RECT 587.230 175.875 604.720 179.885 ;
        RECT 587.260 164.935 604.910 167.885 ;
        RECT 607.230 175.875 624.720 179.885 ;
        RECT 607.260 164.935 624.910 167.885 ;
        RECT 776.230 175.875 793.720 179.885 ;
        RECT 776.260 164.935 793.910 167.885 ;
        RECT 796.230 175.875 813.720 179.885 ;
        RECT 796.260 164.935 813.910 167.885 ;
        RECT 816.230 175.875 833.720 179.885 ;
        RECT 816.260 164.935 833.910 167.885 ;
        RECT 836.230 175.875 853.720 179.885 ;
        RECT 836.260 164.935 853.910 167.885 ;
        RECT 856.230 175.875 873.720 179.885 ;
        RECT 856.260 164.935 873.910 167.885 ;
        RECT 876.230 175.875 893.720 179.885 ;
        RECT 876.260 164.935 893.910 167.885 ;
        RECT 1050.230 175.875 1067.720 179.885 ;
        RECT 1050.260 164.935 1067.910 167.885 ;
        RECT 1070.230 175.875 1087.720 179.885 ;
        RECT 1070.260 164.935 1087.910 167.885 ;
        RECT 1090.230 175.875 1107.720 179.885 ;
        RECT 1090.260 164.935 1107.910 167.885 ;
        RECT 1110.230 175.875 1127.720 179.885 ;
        RECT 1110.260 164.935 1127.910 167.885 ;
        RECT 1130.230 175.875 1147.720 179.885 ;
        RECT 1130.260 164.935 1147.910 167.885 ;
        RECT 1150.230 175.875 1167.720 179.885 ;
        RECT 1150.260 164.935 1167.910 167.885 ;
        RECT 1319.230 175.875 1336.720 179.885 ;
        RECT 1319.260 164.935 1336.910 167.885 ;
        RECT 1339.230 175.875 1356.720 179.885 ;
        RECT 1339.260 164.935 1356.910 167.885 ;
        RECT 1359.230 175.875 1376.720 179.885 ;
        RECT 1359.260 164.935 1376.910 167.885 ;
        RECT 1379.230 175.875 1396.720 179.885 ;
        RECT 1379.260 164.935 1396.910 167.885 ;
        RECT 1399.230 175.875 1416.720 179.885 ;
        RECT 1399.260 164.935 1416.910 167.885 ;
        RECT 1419.230 175.875 1436.720 179.885 ;
        RECT 1419.260 164.935 1436.910 167.885 ;
        RECT 1593.230 175.875 1610.720 179.885 ;
        RECT 1593.260 164.935 1610.910 167.885 ;
        RECT 1613.230 175.875 1630.720 179.885 ;
        RECT 1613.260 164.935 1630.910 167.885 ;
        RECT 1633.230 175.875 1650.720 179.885 ;
        RECT 1633.260 164.935 1650.910 167.885 ;
        RECT 1653.230 175.875 1670.720 179.885 ;
        RECT 1653.260 164.935 1670.910 167.885 ;
        RECT 1673.230 175.875 1690.720 179.885 ;
        RECT 1673.260 164.935 1690.910 167.885 ;
        RECT 1693.230 175.875 1710.720 179.885 ;
        RECT 1693.260 164.935 1710.910 167.885 ;
        RECT 1867.230 175.875 1884.720 179.885 ;
        RECT 1867.260 164.935 1884.910 167.885 ;
        RECT 1887.230 175.875 1904.720 179.885 ;
        RECT 1887.260 164.935 1904.910 167.885 ;
        RECT 1907.230 175.875 1924.720 179.885 ;
        RECT 1907.260 164.935 1924.910 167.885 ;
        RECT 1927.230 175.875 1944.720 179.885 ;
        RECT 1927.260 164.935 1944.910 167.885 ;
        RECT 1947.230 175.875 1964.720 179.885 ;
        RECT 1947.260 164.935 1964.910 167.885 ;
        RECT 1967.230 175.875 1984.720 179.885 ;
        RECT 1967.260 164.935 1984.910 167.885 ;
        RECT 2141.230 175.875 2158.720 179.885 ;
        RECT 2141.260 164.935 2158.910 167.885 ;
        RECT 2161.230 175.875 2178.720 179.885 ;
        RECT 2161.260 164.935 2178.910 167.885 ;
        RECT 2181.230 175.875 2198.720 179.885 ;
        RECT 2181.260 164.935 2198.910 167.885 ;
        RECT 2201.230 175.875 2218.720 179.885 ;
        RECT 2201.260 164.935 2218.910 167.885 ;
        RECT 2221.230 175.875 2238.720 179.885 ;
        RECT 2221.260 164.935 2238.910 167.885 ;
        RECT 2241.230 175.875 2258.720 179.885 ;
        RECT 2241.260 164.935 2258.910 167.885 ;
        RECT 2415.230 175.875 2432.720 179.885 ;
        RECT 2415.260 164.935 2432.910 167.885 ;
        RECT 2435.230 175.875 2452.720 179.885 ;
        RECT 2435.260 164.935 2452.910 167.885 ;
        RECT 2455.230 175.875 2472.720 179.885 ;
        RECT 2455.260 164.935 2472.910 167.885 ;
        RECT 2475.230 175.875 2492.720 179.885 ;
        RECT 2475.260 164.935 2492.910 167.885 ;
        RECT 2495.230 175.875 2512.720 179.885 ;
        RECT 2495.260 164.935 2512.910 167.885 ;
        RECT 2515.230 175.875 2532.720 179.885 ;
        RECT 2515.260 164.935 2532.910 167.885 ;
        RECT 2689.230 175.875 2706.720 179.885 ;
        RECT 2689.260 164.935 2706.910 167.885 ;
        RECT 2709.230 175.875 2726.720 179.885 ;
        RECT 2709.260 164.935 2726.910 167.885 ;
        RECT 2729.230 175.875 2746.720 179.885 ;
        RECT 2729.260 164.935 2746.910 167.885 ;
        RECT 2749.230 175.875 2766.720 179.885 ;
        RECT 2749.260 164.935 2766.910 167.885 ;
        RECT 2769.230 175.875 2786.720 179.885 ;
        RECT 2769.260 164.935 2786.910 167.885 ;
        RECT 2789.230 175.875 2806.720 179.885 ;
        RECT 2958.230 175.875 2975.720 179.885 ;
        RECT 2789.260 164.935 2806.910 167.885 ;
        RECT 2958.260 164.935 2975.910 167.885 ;
        RECT 2978.230 175.875 2995.720 179.885 ;
        RECT 2978.260 164.935 2995.910 167.885 ;
        RECT 2998.230 175.875 3015.720 179.885 ;
        RECT 2998.260 164.935 3015.910 167.885 ;
        RECT 3018.230 175.875 3035.720 179.885 ;
        RECT 3018.260 164.935 3035.910 167.885 ;
        RECT 3038.230 175.875 3055.720 179.885 ;
        RECT 3038.260 164.935 3055.910 167.885 ;
        RECT 3058.230 175.875 3075.720 179.885 ;
        RECT 3058.260 164.935 3075.910 167.885 ;
        RECT 3227.230 175.875 3244.720 179.885 ;
        RECT 3227.260 164.935 3244.910 167.885 ;
        RECT 3247.230 175.875 3264.720 179.885 ;
        RECT 3247.260 164.935 3264.910 167.885 ;
        RECT 3267.230 175.875 3284.720 179.885 ;
        RECT 3267.260 164.935 3284.910 167.885 ;
        RECT 3287.230 175.875 3304.720 179.885 ;
        RECT 3287.260 164.935 3304.910 167.885 ;
        RECT 3307.230 175.875 3324.720 179.885 ;
        RECT 3307.260 164.935 3324.910 167.885 ;
        RECT 3327.230 175.875 3344.720 179.885 ;
        RECT 3327.260 164.935 3344.910 167.885 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 204.000 5083.400 375.000 5188.000 ;
      LAYER met4 ;
        RECT 375.000 5163.785 376.270 5188.000 ;
      LAYER met4 ;
        RECT 376.670 5163.385 448.330 5188.000 ;
      LAYER met4 ;
        RECT 448.730 5163.785 450.000 5188.000 ;
      LAYER met4 ;
        RECT 375.965 5083.400 449.035 5163.385 ;
        RECT 450.000 5083.400 615.000 5188.000 ;
      LAYER met4 ;
        RECT 615.000 5163.785 616.270 5188.000 ;
      LAYER met4 ;
        RECT 616.670 5163.385 688.330 5188.000 ;
      LAYER met4 ;
        RECT 688.730 5163.785 690.000 5188.000 ;
      LAYER met4 ;
        RECT 615.965 5083.400 689.035 5163.385 ;
        RECT 690.000 5083.400 855.000 5188.000 ;
      LAYER met4 ;
        RECT 855.000 5163.785 856.270 5188.000 ;
      LAYER met4 ;
        RECT 856.670 5163.385 928.330 5188.000 ;
      LAYER met4 ;
        RECT 928.730 5163.785 930.000 5188.000 ;
      LAYER met4 ;
        RECT 855.965 5083.400 929.035 5163.385 ;
        RECT 930.000 5083.400 1100.000 5188.000 ;
      LAYER met4 ;
        RECT 1100.000 5163.785 1148.205 5188.000 ;
      LAYER met4 ;
        RECT 1148.605 5163.385 1225.485 5188.000 ;
      LAYER met4 ;
        RECT 1225.885 5163.785 1269.000 5188.000 ;
      LAYER met4 ;
        RECT 1147.240 5083.400 1225.885 5163.385 ;
        RECT 1269.000 5083.400 1357.000 5188.000 ;
      LAYER met4 ;
        RECT 1357.000 5163.785 1405.205 5188.000 ;
      LAYER met4 ;
        RECT 1405.605 5163.385 1482.485 5188.000 ;
      LAYER met4 ;
        RECT 1482.885 5163.785 1526.000 5188.000 ;
      LAYER met4 ;
        RECT 1404.240 5083.400 1482.885 5163.385 ;
        RECT 1526.000 5083.400 1697.000 5188.000 ;
      LAYER met4 ;
        RECT 1697.000 5163.785 1698.270 5188.000 ;
      LAYER met4 ;
        RECT 1698.670 5163.385 1770.330 5188.000 ;
      LAYER met4 ;
        RECT 1770.730 5163.785 1772.000 5188.000 ;
      LAYER met4 ;
        RECT 1772.000 5163.785 2124.000 5188.000 ;
      LAYER met4 ;
        RECT 2124.000 5163.785 2125.270 5188.000 ;
      LAYER met4 ;
        RECT 1697.965 5083.400 1771.035 5163.385 ;
        RECT 1772.000 5083.400 1943.000 5163.785 ;
        RECT 1948.000 5083.400 2124.000 5163.785 ;
        RECT 2125.670 5163.385 2197.330 5188.000 ;
      LAYER met4 ;
        RECT 2197.730 5163.785 2199.000 5188.000 ;
      LAYER met4 ;
        RECT 2124.965 5083.400 2198.035 5163.385 ;
        RECT 2199.000 5083.400 2371.000 5188.000 ;
      LAYER met4 ;
        RECT 2371.000 5163.785 2372.270 5188.000 ;
      LAYER met4 ;
        RECT 2372.670 5163.385 2444.330 5188.000 ;
      LAYER met4 ;
        RECT 2444.730 5163.785 2446.000 5188.000 ;
      LAYER met4 ;
        RECT 2371.965 5083.400 2445.035 5163.385 ;
        RECT 2446.000 5083.400 2629.000 5188.000 ;
      LAYER met4 ;
        RECT 2629.000 5163.785 2630.270 5188.000 ;
      LAYER met4 ;
        RECT 2630.670 5163.385 2702.330 5188.000 ;
      LAYER met4 ;
        RECT 2702.730 5163.785 2704.000 5188.000 ;
      LAYER met4 ;
        RECT 2629.965 5083.400 2703.035 5163.385 ;
        RECT 2704.000 5083.400 2878.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.000 5163.785 2879.270 5188.000 ;
      LAYER met4 ;
        RECT 2879.670 5163.385 2951.330 5188.000 ;
      LAYER met4 ;
        RECT 2951.730 5163.785 2953.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.965 5083.400 2952.035 5163.385 ;
        RECT 2953.000 5083.400 3135.000 5188.000 ;
      LAYER met4 ;
        RECT 3135.000 5163.785 3136.270 5188.000 ;
      LAYER met4 ;
        RECT 3136.670 5163.385 3208.330 5188.000 ;
      LAYER met4 ;
        RECT 3208.730 5163.785 3210.000 5188.000 ;
      LAYER met4 ;
        RECT 3210.000 5163.385 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
        RECT 3135.965 5083.400 3209.035 5163.385 ;
        RECT 3210.000 5083.400 3588.000 5163.385 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
      LAYER met4 ;
        RECT 202.145 5058.035 376.270 5083.000 ;
      LAYER met4 ;
        RECT 376.670 5057.635 448.330 5083.400 ;
      LAYER met4 ;
        RECT 448.730 5058.035 616.270 5083.000 ;
      LAYER met4 ;
        RECT 616.670 5057.635 688.330 5083.400 ;
      LAYER met4 ;
        RECT 688.730 5058.035 856.270 5083.000 ;
      LAYER met4 ;
        RECT 856.670 5057.635 928.330 5083.400 ;
      LAYER met4 ;
        RECT 928.730 5058.035 1147.715 5083.000 ;
      LAYER met4 ;
        RECT 1148.115 5057.635 1225.485 5083.400 ;
      LAYER met4 ;
        RECT 1225.885 5058.035 1404.715 5083.000 ;
      LAYER met4 ;
        RECT 1405.115 5057.635 1482.485 5083.400 ;
      LAYER met4 ;
        RECT 1482.885 5058.035 1698.270 5083.000 ;
      LAYER met4 ;
        RECT 1698.670 5057.635 1770.330 5083.400 ;
      LAYER met4 ;
        RECT 1770.730 5058.035 2125.270 5083.000 ;
      LAYER met4 ;
        RECT 2125.670 5057.635 2197.330 5083.400 ;
      LAYER met4 ;
        RECT 2197.730 5058.035 2372.270 5083.000 ;
      LAYER met4 ;
        RECT 2372.670 5057.635 2444.330 5083.400 ;
      LAYER met4 ;
        RECT 2444.730 5058.035 2630.270 5083.000 ;
      LAYER met4 ;
        RECT 2630.670 5057.635 2702.330 5083.400 ;
      LAYER met4 ;
        RECT 2702.730 5058.035 2879.270 5083.000 ;
      LAYER met4 ;
        RECT 2879.670 5057.635 2951.330 5083.400 ;
      LAYER met4 ;
        RECT 2951.730 5058.035 3136.270 5083.000 ;
      LAYER met4 ;
        RECT 3136.670 5057.635 3208.330 5083.400 ;
      LAYER met4 ;
        RECT 3208.730 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 375.000 5057.635 ;
        RECT 375.965 5056.935 449.035 5057.635 ;
        RECT 450.000 5056.935 615.000 5057.635 ;
        RECT 615.965 5056.935 689.035 5057.635 ;
        RECT 690.000 5056.935 855.000 5057.635 ;
        RECT 855.965 5056.935 929.035 5057.635 ;
        RECT 930.000 5056.935 1100.000 5057.635 ;
        RECT 1147.240 5056.935 1225.885 5057.635 ;
        RECT 1269.000 5056.935 1357.000 5057.635 ;
        RECT 1404.240 5056.935 1482.885 5057.635 ;
        RECT 1526.000 5056.935 1697.000 5057.635 ;
        RECT 1697.965 5056.935 1771.035 5057.635 ;
        RECT 1772.000 5056.935 1943.000 5057.635 ;
        RECT 1948.000 5056.935 2124.000 5057.635 ;
        RECT 2124.965 5056.935 2198.035 5057.635 ;
        RECT 2199.000 5056.935 2371.000 5057.635 ;
        RECT 2371.965 5056.935 2445.035 5057.635 ;
        RECT 2446.000 5056.935 2629.000 5057.635 ;
        RECT 2629.965 5056.935 2703.035 5057.635 ;
        RECT 2704.000 5056.935 2878.000 5057.635 ;
        RECT 2878.965 5056.935 2952.035 5057.635 ;
        RECT 2953.000 5056.935 3135.000 5057.635 ;
        RECT 3135.965 5056.935 3209.035 5057.635 ;
        RECT 3210.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 376.270 5056.535 ;
      LAYER met4 ;
        RECT 376.670 5051.685 448.330 5056.935 ;
      LAYER met4 ;
        RECT 448.730 5052.085 616.270 5056.535 ;
      LAYER met4 ;
        RECT 616.670 5051.685 688.330 5056.935 ;
      LAYER met4 ;
        RECT 688.730 5052.085 856.270 5056.535 ;
      LAYER met4 ;
        RECT 856.670 5051.685 928.330 5056.935 ;
      LAYER met4 ;
        RECT 928.730 5052.085 1147.715 5056.535 ;
      LAYER met4 ;
        RECT 1148.115 5051.685 1225.485 5056.935 ;
      LAYER met4 ;
        RECT 1225.885 5052.085 1404.715 5056.535 ;
      LAYER met4 ;
        RECT 1405.115 5051.685 1482.485 5056.935 ;
      LAYER met4 ;
        RECT 1482.885 5052.085 1698.270 5056.535 ;
      LAYER met4 ;
        RECT 1698.670 5051.685 1770.330 5056.935 ;
      LAYER met4 ;
        RECT 1770.730 5052.085 2125.270 5056.535 ;
      LAYER met4 ;
        RECT 2125.670 5051.685 2197.330 5056.935 ;
      LAYER met4 ;
        RECT 2197.730 5052.085 2372.270 5056.535 ;
      LAYER met4 ;
        RECT 2372.670 5051.685 2444.330 5056.935 ;
      LAYER met4 ;
        RECT 2444.730 5052.085 2630.270 5056.535 ;
      LAYER met4 ;
        RECT 2630.670 5051.685 2702.330 5056.935 ;
      LAYER met4 ;
        RECT 2702.730 5052.085 2879.270 5056.535 ;
      LAYER met4 ;
        RECT 2879.670 5051.685 2951.330 5056.935 ;
      LAYER met4 ;
        RECT 2951.730 5052.085 3136.270 5056.535 ;
      LAYER met4 ;
        RECT 3136.670 5051.685 3208.330 5056.935 ;
      LAYER met4 ;
        RECT 3208.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 375.000 5051.685 ;
        RECT 375.965 5051.085 449.035 5051.685 ;
        RECT 450.000 5051.085 615.000 5051.685 ;
        RECT 615.965 5051.085 689.035 5051.685 ;
        RECT 690.000 5051.085 855.000 5051.685 ;
        RECT 855.965 5051.085 929.035 5051.685 ;
        RECT 930.000 5051.085 1100.000 5051.685 ;
        RECT 1147.240 5051.085 1225.885 5051.685 ;
        RECT 1269.000 5051.085 1357.000 5051.685 ;
        RECT 1404.240 5051.085 1482.885 5051.685 ;
        RECT 1526.000 5051.085 1697.000 5051.685 ;
        RECT 1697.965 5051.085 1771.035 5051.685 ;
        RECT 1772.000 5051.085 1943.000 5051.685 ;
        RECT 1948.000 5051.085 2124.000 5051.685 ;
        RECT 2124.965 5051.085 2198.035 5051.685 ;
        RECT 2199.000 5051.085 2371.000 5051.685 ;
        RECT 2371.965 5051.085 2445.035 5051.685 ;
        RECT 2446.000 5051.085 2629.000 5051.685 ;
        RECT 2629.965 5051.085 2703.035 5051.685 ;
        RECT 2704.000 5051.085 2878.000 5051.685 ;
        RECT 2878.965 5051.085 2952.035 5051.685 ;
        RECT 2953.000 5051.085 3135.000 5051.685 ;
        RECT 3135.965 5051.085 3209.035 5051.685 ;
        RECT 3210.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 376.270 5050.685 ;
      LAYER met4 ;
        RECT 376.670 5045.835 448.330 5051.085 ;
      LAYER met4 ;
        RECT 448.730 5046.235 616.270 5050.685 ;
      LAYER met4 ;
        RECT 616.670 5045.835 688.330 5051.085 ;
      LAYER met4 ;
        RECT 688.730 5046.235 856.270 5050.685 ;
      LAYER met4 ;
        RECT 856.670 5045.835 928.330 5051.085 ;
      LAYER met4 ;
        RECT 928.730 5046.235 1147.715 5050.685 ;
      LAYER met4 ;
        RECT 1148.115 5045.835 1225.485 5051.085 ;
      LAYER met4 ;
        RECT 1225.885 5046.235 1404.715 5050.685 ;
      LAYER met4 ;
        RECT 1405.115 5045.835 1482.485 5051.085 ;
      LAYER met4 ;
        RECT 1482.885 5046.235 1698.270 5050.685 ;
      LAYER met4 ;
        RECT 1698.670 5045.835 1770.330 5051.085 ;
      LAYER met4 ;
        RECT 1770.730 5046.235 2125.270 5050.685 ;
      LAYER met4 ;
        RECT 2125.670 5045.835 2197.330 5051.085 ;
      LAYER met4 ;
        RECT 2197.730 5046.235 2372.270 5050.685 ;
      LAYER met4 ;
        RECT 2372.670 5045.835 2444.330 5051.085 ;
      LAYER met4 ;
        RECT 2444.730 5046.235 2630.270 5050.685 ;
      LAYER met4 ;
        RECT 2630.670 5045.835 2702.330 5051.085 ;
      LAYER met4 ;
        RECT 2702.730 5046.235 2879.270 5050.685 ;
      LAYER met4 ;
        RECT 2879.670 5045.835 2951.330 5051.085 ;
      LAYER met4 ;
        RECT 2951.730 5046.235 3136.270 5050.685 ;
      LAYER met4 ;
        RECT 3136.670 5045.835 3208.330 5051.085 ;
      LAYER met4 ;
        RECT 3208.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 375.000 5045.835 ;
        RECT 375.965 5045.135 449.035 5045.835 ;
        RECT 450.000 5045.135 615.000 5045.835 ;
        RECT 615.965 5045.135 689.035 5045.835 ;
        RECT 690.000 5045.135 855.000 5045.835 ;
        RECT 855.965 5045.135 929.035 5045.835 ;
        RECT 930.000 5045.135 1100.000 5045.835 ;
        RECT 1147.240 5045.135 1225.885 5045.835 ;
        RECT 1269.000 5045.135 1357.000 5045.835 ;
        RECT 1404.240 5045.135 1482.885 5045.835 ;
        RECT 1526.000 5045.135 1697.000 5045.835 ;
        RECT 1697.965 5045.135 1771.035 5045.835 ;
        RECT 1772.000 5045.135 1943.000 5045.835 ;
        RECT 1948.000 5045.135 2124.000 5045.835 ;
        RECT 2124.965 5045.135 2198.035 5045.835 ;
        RECT 2199.000 5045.135 2371.000 5045.835 ;
        RECT 2371.965 5045.135 2445.035 5045.835 ;
        RECT 2446.000 5045.135 2629.000 5045.835 ;
        RECT 2629.965 5045.135 2703.035 5045.835 ;
        RECT 2704.000 5045.135 2878.000 5045.835 ;
        RECT 2878.965 5045.135 2952.035 5045.835 ;
        RECT 2953.000 5045.135 3135.000 5045.835 ;
        RECT 3135.965 5045.135 3209.035 5045.835 ;
        RECT 3210.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 1943.000 5044.735 ;
        RECT 1948.000 5044.405 2879.270 5044.735 ;
      LAYER met4 ;
        RECT 2879.670 5044.505 2951.330 5045.135 ;
      LAYER met4 ;
        RECT 2951.730 5044.405 3411.175 5044.735 ;
      LAYER met4 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.645 375.000 5040.825 ;
      LAYER met4 ;
        RECT 375.000 5039.645 376.270 5040.825 ;
      LAYER met4 ;
        RECT 376.670 5039.745 448.330 5040.725 ;
      LAYER met4 ;
        RECT 448.730 5039.645 450.000 5040.825 ;
      LAYER met4 ;
        RECT 450.000 5039.645 615.000 5040.825 ;
      LAYER met4 ;
        RECT 615.000 5039.645 616.270 5040.825 ;
      LAYER met4 ;
        RECT 616.670 5039.745 688.330 5040.725 ;
      LAYER met4 ;
        RECT 688.730 5039.645 690.000 5040.825 ;
      LAYER met4 ;
        RECT 690.000 5039.645 855.000 5040.825 ;
      LAYER met4 ;
        RECT 855.000 5039.645 856.270 5040.825 ;
      LAYER met4 ;
        RECT 856.670 5039.745 928.330 5040.725 ;
      LAYER met4 ;
        RECT 928.730 5039.645 930.000 5040.825 ;
      LAYER met4 ;
        RECT 930.000 5039.645 1100.000 5040.825 ;
      LAYER met4 ;
        RECT 1100.000 5039.645 1147.240 5040.825 ;
      LAYER met4 ;
        RECT 1147.640 5039.745 1225.485 5040.725 ;
      LAYER met4 ;
        RECT 1225.885 5039.645 1269.000 5040.825 ;
      LAYER met4 ;
        RECT 1269.000 5039.645 1357.000 5040.825 ;
      LAYER met4 ;
        RECT 1357.000 5039.645 1404.240 5040.825 ;
      LAYER met4 ;
        RECT 1404.640 5039.745 1482.485 5040.725 ;
      LAYER met4 ;
        RECT 1482.885 5039.645 1526.000 5040.825 ;
      LAYER met4 ;
        RECT 1526.000 5039.645 1697.000 5040.825 ;
      LAYER met4 ;
        RECT 1697.000 5039.645 1698.270 5040.825 ;
      LAYER met4 ;
        RECT 1698.670 5039.745 1770.330 5040.725 ;
      LAYER met4 ;
        RECT 1770.730 5039.645 1772.000 5040.825 ;
      LAYER met4 ;
        RECT 1772.000 5039.645 1943.000 5040.825 ;
        RECT 1948.000 5039.645 2124.000 5040.825 ;
      LAYER met4 ;
        RECT 2124.000 5039.645 2125.270 5040.825 ;
      LAYER met4 ;
        RECT 2125.670 5039.745 2197.330 5040.725 ;
      LAYER met4 ;
        RECT 2197.730 5039.645 2199.000 5040.825 ;
      LAYER met4 ;
        RECT 2199.000 5039.645 2371.000 5040.825 ;
      LAYER met4 ;
        RECT 2371.000 5039.645 2372.270 5040.825 ;
      LAYER met4 ;
        RECT 2372.670 5039.745 2444.330 5040.725 ;
      LAYER met4 ;
        RECT 2444.730 5039.645 2446.000 5040.825 ;
      LAYER met4 ;
        RECT 2446.000 5039.645 2629.000 5040.825 ;
      LAYER met4 ;
        RECT 2629.000 5039.645 2630.270 5040.825 ;
      LAYER met4 ;
        RECT 2630.670 5039.745 2702.330 5040.725 ;
      LAYER met4 ;
        RECT 2702.730 5039.645 2704.000 5040.825 ;
      LAYER met4 ;
        RECT 2704.000 5039.645 2878.000 5040.825 ;
      LAYER met4 ;
        RECT 2878.000 5039.645 2879.270 5040.825 ;
      LAYER met4 ;
        RECT 2879.670 5039.745 2951.330 5040.725 ;
      LAYER met4 ;
        RECT 2951.730 5039.645 2953.000 5040.825 ;
      LAYER met4 ;
        RECT 2953.000 5039.645 3135.000 5040.825 ;
      LAYER met4 ;
        RECT 3135.000 5039.645 3136.270 5040.825 ;
      LAYER met4 ;
        RECT 3136.670 5039.745 3208.330 5040.725 ;
      LAYER met4 ;
        RECT 3208.730 5039.645 3210.000 5040.825 ;
      LAYER met4 ;
        RECT 3210.000 5039.645 3388.000 5040.825 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 1943.000 5036.065 ;
        RECT 1948.000 5035.735 2879.270 5036.065 ;
      LAYER met4 ;
        RECT 2879.670 5035.335 2951.330 5035.965 ;
      LAYER met4 ;
        RECT 2951.730 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 375.965 5034.635 449.035 5035.335 ;
        RECT 615.965 5034.635 689.035 5035.335 ;
        RECT 855.965 5034.635 929.035 5035.335 ;
        RECT 1147.240 5034.635 1225.885 5035.335 ;
        RECT 1404.240 5034.635 1482.885 5035.335 ;
        RECT 1697.965 5034.635 1771.035 5035.335 ;
        RECT 2124.965 5034.635 2198.035 5035.335 ;
        RECT 2371.965 5034.635 2445.035 5035.335 ;
        RECT 2629.965 5034.635 2703.035 5035.335 ;
        RECT 2878.965 5034.635 2952.035 5035.335 ;
        RECT 3135.965 5034.635 3209.035 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 376.270 5034.235 ;
      LAYER met4 ;
        RECT 376.670 5029.185 448.330 5034.635 ;
      LAYER met4 ;
        RECT 448.730 5029.585 616.270 5034.235 ;
      LAYER met4 ;
        RECT 616.670 5029.185 688.330 5034.635 ;
      LAYER met4 ;
        RECT 688.730 5029.585 856.270 5034.235 ;
      LAYER met4 ;
        RECT 856.670 5029.185 928.330 5034.635 ;
      LAYER met4 ;
        RECT 928.730 5029.585 1147.250 5034.235 ;
      LAYER met4 ;
        RECT 1147.650 5029.185 1225.485 5034.635 ;
      LAYER met4 ;
        RECT 1225.885 5029.585 1404.250 5034.235 ;
      LAYER met4 ;
        RECT 1404.650 5029.185 1482.485 5034.635 ;
      LAYER met4 ;
        RECT 1482.885 5029.585 1698.270 5034.235 ;
      LAYER met4 ;
        RECT 1698.670 5029.185 1770.330 5034.635 ;
      LAYER met4 ;
        RECT 1770.730 5029.585 1948.000 5034.235 ;
        RECT 1953.000 5029.585 2125.270 5034.235 ;
      LAYER met4 ;
        RECT 2125.670 5029.185 2197.330 5034.635 ;
      LAYER met4 ;
        RECT 2197.730 5029.585 2372.270 5034.235 ;
      LAYER met4 ;
        RECT 2372.670 5029.185 2444.330 5034.635 ;
      LAYER met4 ;
        RECT 2444.730 5029.585 2630.270 5034.235 ;
      LAYER met4 ;
        RECT 2630.670 5029.185 2702.330 5034.635 ;
      LAYER met4 ;
        RECT 2702.730 5029.585 2879.270 5034.235 ;
      LAYER met4 ;
        RECT 2879.670 5029.185 2951.330 5034.635 ;
      LAYER met4 ;
        RECT 2951.730 5029.585 3136.270 5034.235 ;
      LAYER met4 ;
        RECT 3136.670 5029.185 3208.330 5034.635 ;
      LAYER met4 ;
        RECT 3208.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 375.965 5028.585 449.035 5029.185 ;
        RECT 615.965 5028.585 689.035 5029.185 ;
        RECT 855.965 5028.585 929.035 5029.185 ;
        RECT 1147.240 5028.585 1225.885 5029.185 ;
        RECT 1404.240 5028.585 1482.885 5029.185 ;
        RECT 1697.965 5028.585 1771.035 5029.185 ;
        RECT 2124.965 5028.585 2198.035 5029.185 ;
        RECT 2371.965 5028.585 2445.035 5029.185 ;
        RECT 2629.965 5028.585 2703.035 5029.185 ;
        RECT 2878.965 5028.585 2952.035 5029.185 ;
        RECT 3135.965 5028.585 3209.035 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 376.270 5028.185 ;
      LAYER met4 ;
        RECT 376.670 5024.335 448.330 5028.585 ;
      LAYER met4 ;
        RECT 448.730 5024.735 616.270 5028.185 ;
      LAYER met4 ;
        RECT 616.670 5024.335 688.330 5028.585 ;
      LAYER met4 ;
        RECT 688.730 5024.735 856.270 5028.185 ;
      LAYER met4 ;
        RECT 856.670 5024.335 928.330 5028.585 ;
      LAYER met4 ;
        RECT 928.730 5024.735 1147.715 5028.185 ;
      LAYER met4 ;
        RECT 1148.115 5024.335 1225.485 5028.585 ;
      LAYER met4 ;
        RECT 1225.885 5024.735 1404.715 5028.185 ;
      LAYER met4 ;
        RECT 1405.115 5024.335 1482.485 5028.585 ;
      LAYER met4 ;
        RECT 1482.885 5024.735 1698.270 5028.185 ;
      LAYER met4 ;
        RECT 1698.670 5024.335 1770.330 5028.585 ;
      LAYER met4 ;
        RECT 1770.730 5024.735 1943.000 5028.185 ;
        RECT 1948.000 5024.735 2125.270 5028.185 ;
      LAYER met4 ;
        RECT 2125.670 5024.335 2197.330 5028.585 ;
      LAYER met4 ;
        RECT 2197.730 5024.735 2372.270 5028.185 ;
      LAYER met4 ;
        RECT 2372.670 5024.335 2444.330 5028.585 ;
      LAYER met4 ;
        RECT 2444.730 5024.735 2630.270 5028.185 ;
      LAYER met4 ;
        RECT 2630.670 5024.335 2702.330 5028.585 ;
      LAYER met4 ;
        RECT 2702.730 5024.735 2879.270 5028.185 ;
      LAYER met4 ;
        RECT 2879.670 5024.335 2951.330 5028.585 ;
      LAYER met4 ;
        RECT 2951.730 5024.735 3136.270 5028.185 ;
      LAYER met4 ;
        RECT 3136.670 5024.335 3208.330 5028.585 ;
      LAYER met4 ;
        RECT 3208.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 375.965 5023.735 449.035 5024.335 ;
        RECT 615.965 5023.735 689.035 5024.335 ;
        RECT 855.965 5023.735 929.035 5024.335 ;
        RECT 1147.240 5023.735 1225.885 5024.335 ;
        RECT 1404.240 5023.735 1482.885 5024.335 ;
        RECT 1697.965 5023.735 1771.035 5024.335 ;
        RECT 2124.965 5023.735 2198.035 5024.335 ;
        RECT 2371.965 5023.735 2445.035 5024.335 ;
        RECT 2629.965 5023.735 2703.035 5024.335 ;
        RECT 2878.965 5023.735 2952.035 5024.335 ;
        RECT 3135.965 5023.735 3209.035 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 376.270 5023.335 ;
      LAYER met4 ;
        RECT 376.670 5019.485 448.330 5023.735 ;
      LAYER met4 ;
        RECT 448.730 5019.885 616.270 5023.335 ;
      LAYER met4 ;
        RECT 616.670 5019.485 688.330 5023.735 ;
      LAYER met4 ;
        RECT 688.730 5019.885 856.270 5023.335 ;
      LAYER met4 ;
        RECT 856.670 5019.485 928.330 5023.735 ;
      LAYER met4 ;
        RECT 928.730 5019.885 1147.715 5023.335 ;
      LAYER met4 ;
        RECT 1148.115 5019.485 1225.485 5023.735 ;
      LAYER met4 ;
        RECT 1225.885 5019.885 1404.715 5023.335 ;
      LAYER met4 ;
        RECT 1405.115 5019.485 1482.485 5023.735 ;
      LAYER met4 ;
        RECT 1482.885 5019.885 1698.270 5023.335 ;
      LAYER met4 ;
        RECT 1698.670 5019.485 1770.330 5023.735 ;
      LAYER met4 ;
        RECT 1770.730 5019.885 2125.270 5023.335 ;
      LAYER met4 ;
        RECT 2125.670 5019.485 2197.330 5023.735 ;
      LAYER met4 ;
        RECT 2197.730 5019.885 2372.270 5023.335 ;
      LAYER met4 ;
        RECT 2372.670 5019.485 2444.330 5023.735 ;
      LAYER met4 ;
        RECT 2444.730 5019.885 2630.270 5023.335 ;
      LAYER met4 ;
        RECT 2630.670 5019.485 2702.330 5023.735 ;
      LAYER met4 ;
        RECT 2702.730 5019.885 2879.270 5023.335 ;
      LAYER met4 ;
        RECT 2879.670 5019.485 2951.330 5023.735 ;
      LAYER met4 ;
        RECT 2951.730 5019.885 3136.270 5023.335 ;
      LAYER met4 ;
        RECT 3136.670 5019.485 3208.330 5023.735 ;
      LAYER met4 ;
        RECT 3208.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 375.965 5018.885 449.035 5019.485 ;
        RECT 615.965 5018.885 689.035 5019.485 ;
        RECT 855.965 5018.885 929.035 5019.485 ;
        RECT 1147.240 5018.885 1225.885 5019.485 ;
        RECT 1404.240 5018.885 1482.885 5019.485 ;
        RECT 1697.965 5018.885 1771.035 5019.485 ;
        RECT 2124.965 5018.885 2198.035 5019.485 ;
        RECT 2371.965 5018.885 2445.035 5019.485 ;
        RECT 2629.965 5018.885 2703.035 5019.485 ;
        RECT 2878.965 5018.885 2952.035 5019.485 ;
        RECT 3135.965 5018.885 3209.035 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 376.270 5018.485 ;
      LAYER met4 ;
        RECT 376.670 5013.435 448.330 5018.885 ;
      LAYER met4 ;
        RECT 448.730 5013.835 616.270 5018.485 ;
      LAYER met4 ;
        RECT 616.670 5013.435 688.330 5018.885 ;
      LAYER met4 ;
        RECT 688.730 5013.835 856.270 5018.485 ;
      LAYER met4 ;
        RECT 856.670 5013.435 928.330 5018.885 ;
      LAYER met4 ;
        RECT 928.730 5013.835 1147.715 5018.485 ;
      LAYER met4 ;
        RECT 1148.115 5013.435 1225.485 5018.885 ;
      LAYER met4 ;
        RECT 1225.885 5013.835 1404.715 5018.485 ;
      LAYER met4 ;
        RECT 1405.115 5013.435 1482.485 5018.885 ;
      LAYER met4 ;
        RECT 1482.885 5013.835 1698.270 5018.485 ;
      LAYER met4 ;
        RECT 1698.670 5013.435 1770.330 5018.885 ;
      LAYER met4 ;
        RECT 1770.730 5013.835 2125.270 5018.485 ;
      LAYER met4 ;
        RECT 2125.670 5013.435 2197.330 5018.885 ;
      LAYER met4 ;
        RECT 2197.730 5013.835 2372.270 5018.485 ;
      LAYER met4 ;
        RECT 2372.670 5013.435 2444.330 5018.885 ;
      LAYER met4 ;
        RECT 2444.730 5013.835 2630.270 5018.485 ;
      LAYER met4 ;
        RECT 2630.670 5013.435 2702.330 5018.885 ;
      LAYER met4 ;
        RECT 2702.730 5013.835 2879.270 5018.485 ;
      LAYER met4 ;
        RECT 2879.670 5013.435 2951.330 5018.885 ;
      LAYER met4 ;
        RECT 2951.730 5013.835 3136.270 5018.485 ;
      LAYER met4 ;
        RECT 3136.670 5013.435 3208.330 5018.885 ;
      LAYER met4 ;
        RECT 3208.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 375.965 5012.835 449.035 5013.435 ;
        RECT 615.965 5012.835 689.035 5013.435 ;
        RECT 855.965 5012.835 929.035 5013.435 ;
        RECT 1147.240 5012.835 1225.885 5013.435 ;
        RECT 1404.240 5012.835 1482.885 5013.435 ;
        RECT 1697.965 5012.835 1771.035 5013.435 ;
        RECT 2124.965 5012.835 2198.035 5013.435 ;
        RECT 2371.965 5012.835 2445.035 5013.435 ;
        RECT 2629.965 5012.835 2703.035 5013.435 ;
        RECT 2878.965 5012.835 2952.035 5013.435 ;
        RECT 3135.965 5012.835 3209.035 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4851.000 104.600 4988.000 ;
      LAYER met4 ;
        RECT 0.000 4849.730 24.215 4851.000 ;
      LAYER met4 ;
        RECT 24.615 4849.330 104.600 4850.035 ;
      LAYER met4 ;
        RECT 105.000 4849.730 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4851.000 131.065 4989.880 ;
        RECT 130.365 4849.330 131.065 4850.035 ;
      LAYER met4 ;
        RECT 131.465 4849.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4851.000 136.915 4989.880 ;
        RECT 136.315 4849.330 136.915 4850.035 ;
      LAYER met4 ;
        RECT 137.315 4849.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4851.000 142.865 4990.025 ;
        RECT 142.165 4849.330 142.865 4850.035 ;
        RECT 0.000 4777.670 142.865 4849.330 ;
      LAYER met4 ;
        RECT 0.000 4776.000 24.215 4777.270 ;
      LAYER met4 ;
        RECT 24.615 4776.965 104.600 4777.670 ;
        RECT 0.000 4640.000 104.600 4776.000 ;
      LAYER met4 ;
        RECT 0.000 4638.730 24.215 4640.000 ;
      LAYER met4 ;
        RECT 24.215 4639.785 24.250 4640.000 ;
        RECT 24.615 4638.330 104.600 4640.000 ;
      LAYER met4 ;
        RECT 105.000 4638.730 129.965 4777.270 ;
      LAYER met4 ;
        RECT 130.365 4776.965 131.065 4777.670 ;
        RECT 130.365 4638.330 131.065 4776.000 ;
      LAYER met4 ;
        RECT 131.465 4638.730 135.915 4777.270 ;
      LAYER met4 ;
        RECT 136.315 4776.965 136.915 4777.670 ;
        RECT 136.315 4638.330 136.915 4776.000 ;
      LAYER met4 ;
        RECT 137.315 4638.730 141.765 4777.270 ;
      LAYER met4 ;
        RECT 142.165 4776.965 142.865 4777.670 ;
        RECT 142.165 4638.330 142.865 4776.000 ;
        RECT 0.000 4566.670 142.865 4638.330 ;
      LAYER met4 ;
        RECT 0.000 4565.000 24.215 4566.270 ;
      LAYER met4 ;
        RECT 24.615 4565.000 104.600 4566.670 ;
        RECT 0.000 4429.000 104.600 4565.000 ;
      LAYER met4 ;
        RECT 0.000 4427.730 24.215 4429.000 ;
      LAYER met4 ;
        RECT 24.615 4427.330 104.600 4428.035 ;
      LAYER met4 ;
        RECT 105.000 4427.730 129.965 4566.270 ;
      LAYER met4 ;
        RECT 130.365 4429.000 131.065 4566.670 ;
        RECT 130.365 4427.330 131.065 4428.035 ;
      LAYER met4 ;
        RECT 131.465 4427.730 135.915 4566.270 ;
      LAYER met4 ;
        RECT 136.315 4429.000 136.915 4566.670 ;
        RECT 136.315 4427.330 136.915 4428.035 ;
      LAYER met4 ;
        RECT 137.315 4427.730 141.765 4566.270 ;
      LAYER met4 ;
        RECT 142.165 4429.000 142.865 4566.670 ;
        RECT 142.165 4427.330 142.865 4428.035 ;
        RECT 0.000 4355.670 142.865 4427.330 ;
      LAYER met4 ;
        RECT 0.000 4354.000 24.215 4355.270 ;
      LAYER met4 ;
        RECT 24.615 4354.965 104.600 4355.670 ;
        RECT 0.000 4217.000 104.600 4354.000 ;
      LAYER met4 ;
        RECT 0.000 4215.730 24.215 4217.000 ;
      LAYER met4 ;
        RECT 24.615 4215.330 104.600 4216.035 ;
      LAYER met4 ;
        RECT 105.000 4215.730 129.965 4355.270 ;
      LAYER met4 ;
        RECT 130.365 4354.965 131.065 4355.670 ;
        RECT 130.365 4217.000 131.065 4354.000 ;
        RECT 130.365 4215.330 131.065 4216.035 ;
      LAYER met4 ;
        RECT 131.465 4215.730 135.915 4355.270 ;
      LAYER met4 ;
        RECT 136.315 4354.965 136.915 4355.670 ;
        RECT 136.315 4217.000 136.915 4354.000 ;
        RECT 136.315 4215.330 136.915 4216.035 ;
      LAYER met4 ;
        RECT 137.315 4215.730 141.765 4355.270 ;
      LAYER met4 ;
        RECT 142.165 4354.965 142.865 4355.670 ;
        RECT 142.165 4217.000 142.865 4354.000 ;
        RECT 142.165 4215.330 142.865 4216.035 ;
      LAYER met4 ;
        RECT 143.265 4215.730 143.595 5011.175 ;
      LAYER met4 ;
        RECT 0.000 4143.670 143.495 4215.330 ;
      LAYER met4 ;
        RECT 0.000 4142.000 24.215 4143.270 ;
      LAYER met4 ;
        RECT 24.615 4142.965 104.600 4143.670 ;
        RECT 0.000 4006.000 104.600 4142.000 ;
      LAYER met4 ;
        RECT 0.000 4004.730 24.215 4006.000 ;
      LAYER met4 ;
        RECT 24.615 4004.330 104.600 4004.970 ;
      LAYER met4 ;
        RECT 105.000 4004.730 129.965 4143.270 ;
      LAYER met4 ;
        RECT 130.365 4142.965 131.065 4143.670 ;
        RECT 130.365 4006.000 131.065 4142.000 ;
        RECT 130.365 4004.330 131.065 4004.970 ;
      LAYER met4 ;
        RECT 131.465 4004.730 135.915 4143.270 ;
      LAYER met4 ;
        RECT 136.315 4142.965 136.915 4143.670 ;
        RECT 136.315 4006.000 136.915 4142.000 ;
        RECT 136.315 4004.330 136.915 4004.970 ;
      LAYER met4 ;
        RECT 137.315 4004.730 141.765 4143.270 ;
      LAYER met4 ;
        RECT 142.165 4142.965 142.865 4143.670 ;
        RECT 142.165 4006.000 142.865 4142.000 ;
        RECT 142.165 4004.330 142.865 4004.970 ;
        RECT 0.000 3972.690 142.865 4004.330 ;
      LAYER met4 ;
        RECT 143.265 3973.090 143.595 4143.270 ;
      LAYER met4 ;
        RECT 0.000 3964.360 143.495 3972.690 ;
      LAYER met4 ;
        RECT 143.895 3964.760 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.175 4851.000 148.355 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4849.730 148.355 4851.000 ;
      LAYER met4 ;
        RECT 147.275 4777.670 148.255 4849.330 ;
      LAYER met4 ;
        RECT 147.175 4776.000 148.355 4777.270 ;
      LAYER met4 ;
        RECT 147.175 4640.000 148.355 4776.000 ;
      LAYER met4 ;
        RECT 147.175 4638.730 148.355 4640.000 ;
      LAYER met4 ;
        RECT 147.275 4566.670 148.255 4638.330 ;
      LAYER met4 ;
        RECT 147.175 4565.000 148.355 4566.270 ;
      LAYER met4 ;
        RECT 147.175 4429.000 148.355 4565.000 ;
      LAYER met4 ;
        RECT 147.175 4427.730 148.355 4429.000 ;
      LAYER met4 ;
        RECT 147.275 4355.670 148.255 4427.330 ;
      LAYER met4 ;
        RECT 147.175 4354.000 148.355 4355.270 ;
      LAYER met4 ;
        RECT 147.175 4217.000 148.355 4354.000 ;
      LAYER met4 ;
        RECT 147.175 4215.730 148.355 4217.000 ;
      LAYER met4 ;
        RECT 147.275 4143.670 148.255 4215.330 ;
      LAYER met4 ;
        RECT 147.175 4142.000 148.355 4143.270 ;
      LAYER met4 ;
        RECT 147.175 4006.000 148.355 4142.000 ;
      LAYER met4 ;
        RECT 147.175 4004.730 148.355 4006.000 ;
      LAYER met4 ;
        RECT 147.275 3980.065 148.255 4004.330 ;
      LAYER met4 ;
        RECT 148.655 3980.465 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
      LAYER met4 ;
        RECT 151.935 4215.730 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 376.270 5012.435 ;
      LAYER met4 ;
        RECT 376.670 5007.385 448.330 5012.835 ;
      LAYER met4 ;
        RECT 448.730 5007.785 616.270 5012.435 ;
      LAYER met4 ;
        RECT 616.670 5007.385 688.330 5012.835 ;
      LAYER met4 ;
        RECT 688.730 5007.785 856.270 5012.435 ;
      LAYER met4 ;
        RECT 856.670 5007.385 928.330 5012.835 ;
      LAYER met4 ;
        RECT 928.730 5007.785 1147.715 5012.435 ;
      LAYER met4 ;
        RECT 1148.115 5007.385 1220.805 5012.835 ;
      LAYER met4 ;
        RECT 1221.205 5007.785 1404.715 5012.435 ;
      LAYER met4 ;
        RECT 1405.115 5007.385 1477.805 5012.835 ;
      LAYER met4 ;
        RECT 1478.205 5007.785 1698.270 5012.435 ;
      LAYER met4 ;
        RECT 1698.670 5007.385 1770.330 5012.835 ;
      LAYER met4 ;
        RECT 1770.730 5007.785 2125.270 5012.435 ;
      LAYER met4 ;
        RECT 2125.670 5007.385 2197.330 5012.835 ;
      LAYER met4 ;
        RECT 2197.730 5007.785 2372.270 5012.435 ;
      LAYER met4 ;
        RECT 2372.670 5007.385 2444.330 5012.835 ;
      LAYER met4 ;
        RECT 2444.730 5007.785 2630.270 5012.435 ;
      LAYER met4 ;
        RECT 2630.670 5007.385 2702.330 5012.835 ;
      LAYER met4 ;
        RECT 2702.730 5007.785 2879.270 5012.435 ;
      LAYER met4 ;
        RECT 2879.670 5007.385 2951.330 5012.835 ;
      LAYER met4 ;
        RECT 2951.730 5007.785 3136.270 5012.435 ;
      LAYER met4 ;
        RECT 3136.670 5007.385 3208.330 5012.835 ;
      LAYER met4 ;
        RECT 3208.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 375.965 5006.785 449.035 5007.385 ;
        RECT 615.965 5006.785 689.035 5007.385 ;
        RECT 855.965 5006.785 929.035 5007.385 ;
        RECT 1147.240 5006.785 1225.885 5007.385 ;
        RECT 1404.240 5006.785 1482.885 5007.385 ;
        RECT 1697.965 5006.785 1771.035 5007.385 ;
        RECT 2124.965 5006.785 2198.035 5007.385 ;
        RECT 2371.965 5006.785 2445.035 5007.385 ;
        RECT 2629.965 5006.785 2703.035 5007.385 ;
        RECT 2878.965 5006.785 2952.035 5007.385 ;
        RECT 3135.965 5006.785 3209.035 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 375.965 5006.385 ;
      LAYER met4 ;
        RECT 376.365 5002.535 448.635 5006.785 ;
      LAYER met4 ;
        RECT 449.035 5002.935 615.965 5006.385 ;
      LAYER met4 ;
        RECT 616.365 5002.535 688.635 5006.785 ;
      LAYER met4 ;
        RECT 689.035 5002.935 855.965 5006.385 ;
      LAYER met4 ;
        RECT 856.365 5002.535 928.635 5006.785 ;
      LAYER met4 ;
        RECT 929.035 5002.935 1147.715 5006.385 ;
      LAYER met4 ;
        RECT 1148.115 5002.535 1220.805 5006.785 ;
      LAYER met4 ;
        RECT 1221.205 5002.935 1404.715 5006.385 ;
      LAYER met4 ;
        RECT 1405.115 5002.535 1477.805 5006.785 ;
      LAYER met4 ;
        RECT 1478.205 5002.935 1697.965 5006.385 ;
      LAYER met4 ;
        RECT 1698.365 5002.535 1770.635 5006.785 ;
      LAYER met4 ;
        RECT 1771.035 5002.935 1943.000 5006.385 ;
        RECT 1948.000 5002.935 2124.965 5006.385 ;
      LAYER met4 ;
        RECT 2125.365 5002.535 2197.635 5006.785 ;
      LAYER met4 ;
        RECT 2198.035 5002.935 2371.965 5006.385 ;
      LAYER met4 ;
        RECT 2372.365 5002.535 2444.635 5006.785 ;
      LAYER met4 ;
        RECT 2445.035 5002.935 2629.965 5006.385 ;
      LAYER met4 ;
        RECT 2630.365 5002.535 2702.635 5006.785 ;
      LAYER met4 ;
        RECT 2703.035 5002.935 2878.965 5006.385 ;
      LAYER met4 ;
        RECT 2879.365 5002.535 2951.635 5006.785 ;
      LAYER met4 ;
        RECT 2952.035 5002.935 3135.965 5006.385 ;
      LAYER met4 ;
        RECT 3136.365 5002.535 3208.635 5006.785 ;
      LAYER met4 ;
        RECT 3209.035 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 375.965 5001.935 449.035 5002.535 ;
        RECT 615.965 5001.935 689.035 5002.535 ;
        RECT 855.965 5001.935 929.035 5002.535 ;
        RECT 1147.240 5001.935 1225.885 5002.535 ;
        RECT 1404.240 5001.935 1482.885 5002.535 ;
        RECT 1697.965 5001.935 1771.035 5002.535 ;
        RECT 2124.965 5001.935 2198.035 5002.535 ;
        RECT 2371.965 5001.935 2445.035 5002.535 ;
        RECT 2629.965 5001.935 2703.035 5002.535 ;
        RECT 2878.965 5001.935 2952.035 5002.535 ;
        RECT 3135.965 5001.935 3209.035 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 376.270 5001.535 ;
      LAYER met4 ;
        RECT 376.670 4996.485 448.330 5001.935 ;
      LAYER met4 ;
        RECT 448.730 4996.885 616.270 5001.535 ;
      LAYER met4 ;
        RECT 616.670 4996.485 688.330 5001.935 ;
      LAYER met4 ;
        RECT 688.730 4996.885 856.270 5001.535 ;
      LAYER met4 ;
        RECT 856.670 4996.485 928.330 5001.935 ;
      LAYER met4 ;
        RECT 928.730 4996.885 1147.715 5001.535 ;
      LAYER met4 ;
        RECT 1148.115 4996.485 1225.485 5001.935 ;
      LAYER met4 ;
        RECT 1225.885 4996.885 1404.715 5001.535 ;
      LAYER met4 ;
        RECT 1405.115 4996.485 1482.485 5001.935 ;
      LAYER met4 ;
        RECT 1482.885 4996.885 1698.270 5001.535 ;
      LAYER met4 ;
        RECT 1698.670 4996.485 1770.330 5001.935 ;
      LAYER met4 ;
        RECT 1770.730 4996.885 1948.000 5001.535 ;
        RECT 1953.000 4996.885 2125.270 5001.535 ;
      LAYER met4 ;
        RECT 2125.670 4996.485 2197.330 5001.935 ;
      LAYER met4 ;
        RECT 2197.730 4996.885 2372.270 5001.535 ;
      LAYER met4 ;
        RECT 2372.670 4996.485 2444.330 5001.935 ;
      LAYER met4 ;
        RECT 2444.730 4996.885 2630.270 5001.535 ;
      LAYER met4 ;
        RECT 2630.670 4996.485 2702.330 5001.935 ;
      LAYER met4 ;
        RECT 2702.730 4996.885 2879.270 5001.535 ;
      LAYER met4 ;
        RECT 2879.670 4996.485 2951.330 5001.935 ;
      LAYER met4 ;
        RECT 2951.730 4996.885 3136.270 5001.535 ;
      LAYER met4 ;
        RECT 3136.670 4996.485 3208.330 5001.935 ;
      LAYER met4 ;
        RECT 3208.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 375.965 4995.885 449.035 4996.485 ;
        RECT 615.965 4995.885 689.035 4996.485 ;
        RECT 855.965 4995.885 929.035 4996.485 ;
        RECT 1147.240 4995.885 1225.885 4996.485 ;
        RECT 1404.240 4995.885 1482.885 4996.485 ;
        RECT 1697.965 4995.885 1771.035 4996.485 ;
        RECT 2124.965 4995.885 2198.035 4996.485 ;
        RECT 2371.965 4995.885 2445.035 4996.485 ;
        RECT 2629.965 4995.885 2703.035 4996.485 ;
        RECT 2878.965 4995.885 2952.035 4996.485 ;
        RECT 3135.965 4995.885 3209.035 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4849.330 153.365 4850.035 ;
      LAYER met4 ;
        RECT 153.765 4849.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4849.330 159.415 4850.035 ;
      LAYER met4 ;
        RECT 159.815 4849.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4849.330 164.265 4850.035 ;
      LAYER met4 ;
        RECT 164.665 4849.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4849.330 169.115 4850.035 ;
      LAYER met4 ;
        RECT 169.515 4849.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4849.330 175.165 4850.035 ;
      LAYER met4 ;
        RECT 175.565 4849.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4850.035 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4849.635 181.215 4850.035 ;
        RECT 185.465 4849.635 186.065 4850.035 ;
      LAYER met4 ;
        RECT 186.465 4849.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4849.330 186.065 4849.635 ;
        RECT 191.515 4849.330 192.115 4850.035 ;
      LAYER met4 ;
        RECT 192.515 4849.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4989.635 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 376.270 4995.485 ;
      LAYER met4 ;
        RECT 376.670 4990.035 448.330 4995.885 ;
      LAYER met4 ;
        RECT 448.730 4990.035 616.270 4995.485 ;
      LAYER met4 ;
        RECT 616.670 4990.035 688.330 4995.885 ;
      LAYER met4 ;
        RECT 688.730 4990.035 856.270 4995.485 ;
      LAYER met4 ;
        RECT 856.670 4990.035 928.330 4995.885 ;
      LAYER met4 ;
        RECT 928.730 4990.035 1147.715 4995.485 ;
      LAYER met4 ;
        RECT 1148.115 4990.035 1225.485 4995.885 ;
      LAYER met4 ;
        RECT 1225.885 4990.035 1404.715 4995.485 ;
      LAYER met4 ;
        RECT 1405.115 4990.035 1482.485 4995.885 ;
      LAYER met4 ;
        RECT 1482.885 4990.035 1698.270 4995.485 ;
      LAYER met4 ;
        RECT 1698.670 4990.035 1770.330 4995.885 ;
      LAYER met4 ;
        RECT 1770.730 4990.035 2125.270 4995.485 ;
      LAYER met4 ;
        RECT 2125.670 4990.035 2197.330 4995.885 ;
      LAYER met4 ;
        RECT 2197.730 4990.035 2372.270 4995.485 ;
      LAYER met4 ;
        RECT 2372.670 4990.035 2444.330 4995.885 ;
      LAYER met4 ;
        RECT 2444.730 4990.035 2630.270 4995.485 ;
      LAYER met4 ;
        RECT 2630.670 4990.035 2702.330 4995.885 ;
      LAYER met4 ;
        RECT 2702.730 4990.035 2879.270 4995.485 ;
      LAYER met4 ;
        RECT 2879.670 4990.035 2951.330 4995.885 ;
      LAYER met4 ;
        RECT 2951.730 4990.035 3136.270 4995.485 ;
      LAYER met4 ;
        RECT 3136.670 4990.035 3208.330 4995.885 ;
      LAYER met4 ;
        RECT 3208.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 198.365 4988.000 202.745 4989.635 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 152.665 4777.670 197.965 4849.330 ;
      LAYER met4 ;
        RECT 3390.035 4794.285 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4793.885 3396.485 4794.760 ;
      LAYER met4 ;
        RECT 3396.885 4794.285 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
        RECT 3401.935 4793.885 3402.535 4794.760 ;
      LAYER met4 ;
        RECT 3402.935 4794.285 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3406.785 4793.885 3407.385 4794.760 ;
      LAYER met4 ;
        RECT 3407.785 4794.285 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3412.835 4793.885 3413.435 4794.760 ;
      LAYER met4 ;
        RECT 3413.835 4794.285 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4793.885 3419.485 4794.760 ;
      LAYER met4 ;
        RECT 3419.885 4794.285 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4793.885 3424.335 4794.760 ;
      LAYER met4 ;
        RECT 3424.735 4794.285 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4794.350 3429.185 4794.760 ;
      LAYER met4 ;
        RECT 3429.585 4794.750 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4794.350 3435.335 4794.760 ;
        RECT 3428.585 4793.885 3435.335 4794.350 ;
        RECT 152.665 4776.965 153.365 4777.670 ;
        RECT 152.665 4638.330 153.365 4640.000 ;
      LAYER met4 ;
        RECT 153.765 4638.730 158.415 4777.270 ;
      LAYER met4 ;
        RECT 158.815 4776.965 159.415 4777.670 ;
        RECT 158.815 4638.330 159.415 4640.000 ;
      LAYER met4 ;
        RECT 159.815 4638.730 163.265 4777.270 ;
      LAYER met4 ;
        RECT 163.665 4776.965 164.265 4777.670 ;
        RECT 163.665 4638.330 164.265 4640.000 ;
      LAYER met4 ;
        RECT 164.665 4638.730 168.115 4777.270 ;
      LAYER met4 ;
        RECT 168.515 4776.965 169.115 4777.670 ;
        RECT 168.515 4638.330 169.115 4640.000 ;
      LAYER met4 ;
        RECT 169.515 4638.730 174.165 4777.270 ;
      LAYER met4 ;
        RECT 174.565 4776.965 175.165 4777.670 ;
        RECT 180.615 4777.365 186.065 4777.670 ;
        RECT 174.165 4639.935 174.200 4650.935 ;
        RECT 174.565 4638.330 175.165 4640.000 ;
      LAYER met4 ;
        RECT 175.565 4638.730 180.215 4777.270 ;
      LAYER met4 ;
        RECT 180.615 4776.965 181.215 4777.365 ;
        RECT 185.465 4776.965 186.065 4777.365 ;
        RECT 180.615 4638.635 181.215 4640.000 ;
      LAYER met4 ;
        RECT 181.615 4639.035 185.065 4776.965 ;
      LAYER met4 ;
        RECT 185.465 4638.635 186.065 4640.000 ;
      LAYER met4 ;
        RECT 186.465 4638.730 191.115 4777.270 ;
      LAYER met4 ;
        RECT 191.515 4776.965 192.115 4777.670 ;
        RECT 180.615 4638.330 186.065 4638.635 ;
        RECT 191.515 4638.330 192.115 4640.000 ;
      LAYER met4 ;
        RECT 192.515 4638.730 197.965 4777.270 ;
      LAYER met4 ;
        RECT 3390.035 4721.195 3435.335 4793.885 ;
        RECT 3390.035 4716.515 3402.535 4721.195 ;
        RECT 3395.885 4716.115 3396.485 4716.515 ;
        RECT 3401.935 4716.115 3402.535 4716.515 ;
        RECT 152.665 4566.670 197.965 4638.330 ;
        RECT 152.665 4565.000 153.365 4566.670 ;
        RECT 152.665 4427.330 153.365 4428.035 ;
      LAYER met4 ;
        RECT 153.765 4427.730 158.415 4566.270 ;
      LAYER met4 ;
        RECT 158.415 4554.025 158.450 4565.070 ;
        RECT 158.815 4565.000 159.415 4566.670 ;
        RECT 158.815 4427.330 159.415 4428.035 ;
      LAYER met4 ;
        RECT 159.815 4427.730 163.265 4566.270 ;
      LAYER met4 ;
        RECT 163.665 4565.000 164.265 4566.670 ;
        RECT 163.665 4427.330 164.265 4428.035 ;
      LAYER met4 ;
        RECT 164.665 4427.730 168.115 4566.270 ;
      LAYER met4 ;
        RECT 168.515 4565.000 169.115 4566.670 ;
        RECT 168.515 4427.330 169.115 4428.035 ;
      LAYER met4 ;
        RECT 169.515 4427.730 174.165 4566.270 ;
      LAYER met4 ;
        RECT 174.565 4565.000 175.165 4566.670 ;
        RECT 180.615 4566.365 186.065 4566.670 ;
        RECT 174.565 4427.330 175.165 4428.035 ;
      LAYER met4 ;
        RECT 175.565 4427.730 180.215 4566.270 ;
      LAYER met4 ;
        RECT 180.615 4565.000 181.215 4566.365 ;
      LAYER met4 ;
        RECT 181.615 4428.035 185.065 4565.965 ;
      LAYER met4 ;
        RECT 185.465 4565.000 186.065 4566.365 ;
        RECT 180.615 4427.635 181.215 4428.035 ;
        RECT 185.465 4427.635 186.065 4428.035 ;
      LAYER met4 ;
        RECT 186.465 4427.730 191.115 4566.270 ;
      LAYER met4 ;
        RECT 191.515 4565.000 192.115 4566.670 ;
        RECT 180.615 4427.330 186.065 4427.635 ;
        RECT 191.515 4427.330 192.115 4428.035 ;
      LAYER met4 ;
        RECT 192.515 4427.730 197.965 4566.270 ;
        RECT 3390.035 4530.730 3395.485 4716.115 ;
      LAYER met4 ;
        RECT 3395.885 4530.330 3396.485 4532.000 ;
      LAYER met4 ;
        RECT 3396.885 4530.730 3401.535 4716.115 ;
      LAYER met4 ;
        RECT 3401.935 4530.635 3402.535 4532.000 ;
      LAYER met4 ;
        RECT 3402.935 4531.035 3406.385 4720.795 ;
      LAYER met4 ;
        RECT 3406.785 4716.115 3407.385 4721.195 ;
        RECT 3406.785 4530.635 3407.385 4532.000 ;
      LAYER met4 ;
        RECT 3407.785 4530.730 3412.435 4720.795 ;
      LAYER met4 ;
        RECT 3412.835 4716.515 3435.335 4721.195 ;
        RECT 3412.835 4716.115 3413.435 4716.515 ;
        RECT 3418.885 4716.115 3419.485 4716.515 ;
        RECT 3423.735 4716.115 3424.335 4716.515 ;
        RECT 3428.585 4716.115 3429.185 4716.515 ;
        RECT 3434.635 4716.115 3435.335 4716.515 ;
        RECT 3401.935 4530.330 3407.385 4530.635 ;
        RECT 3412.835 4530.330 3413.435 4532.000 ;
      LAYER met4 ;
        RECT 3413.835 4530.730 3418.485 4716.115 ;
      LAYER met4 ;
        RECT 3418.885 4530.330 3419.485 4532.000 ;
      LAYER met4 ;
        RECT 3419.885 4530.730 3423.335 4716.115 ;
      LAYER met4 ;
        RECT 3423.735 4530.330 3424.335 4532.000 ;
      LAYER met4 ;
        RECT 3424.735 4530.730 3428.185 4716.115 ;
      LAYER met4 ;
        RECT 3428.585 4530.330 3429.185 4532.000 ;
        RECT 3429.550 4531.930 3429.585 4542.975 ;
      LAYER met4 ;
        RECT 3429.585 4530.730 3434.235 4716.115 ;
      LAYER met4 ;
        RECT 3434.635 4530.330 3435.335 4532.000 ;
        RECT 3390.035 4458.670 3435.335 4530.330 ;
        RECT 152.665 4355.670 197.965 4427.330 ;
        RECT 152.665 4354.965 153.365 4355.670 ;
        RECT 152.665 4215.330 153.365 4216.035 ;
      LAYER met4 ;
        RECT 153.765 4215.730 158.415 4355.270 ;
      LAYER met4 ;
        RECT 158.815 4354.965 159.415 4355.670 ;
        RECT 158.815 4215.330 159.415 4216.035 ;
      LAYER met4 ;
        RECT 159.815 4215.730 163.265 4355.270 ;
      LAYER met4 ;
        RECT 163.665 4354.965 164.265 4355.670 ;
        RECT 163.665 4215.330 164.265 4216.035 ;
      LAYER met4 ;
        RECT 164.665 4215.730 168.115 4355.270 ;
      LAYER met4 ;
        RECT 168.515 4354.965 169.115 4355.670 ;
        RECT 168.515 4215.330 169.115 4216.035 ;
      LAYER met4 ;
        RECT 169.515 4215.730 174.165 4355.270 ;
      LAYER met4 ;
        RECT 174.565 4354.965 175.165 4355.670 ;
        RECT 180.615 4355.365 186.065 4355.670 ;
        RECT 174.565 4215.330 175.165 4216.035 ;
      LAYER met4 ;
        RECT 175.565 4215.730 180.215 4355.270 ;
      LAYER met4 ;
        RECT 180.615 4354.965 181.215 4355.365 ;
        RECT 185.465 4354.965 186.065 4355.365 ;
      LAYER met4 ;
        RECT 181.615 4216.035 185.065 4354.965 ;
      LAYER met4 ;
        RECT 180.615 4215.635 181.215 4216.035 ;
        RECT 185.465 4215.635 186.065 4216.035 ;
      LAYER met4 ;
        RECT 186.465 4215.730 191.115 4355.270 ;
      LAYER met4 ;
        RECT 191.515 4354.965 192.115 4355.670 ;
        RECT 180.615 4215.330 186.065 4215.635 ;
        RECT 191.515 4215.330 192.115 4216.035 ;
      LAYER met4 ;
        RECT 192.515 4215.730 197.965 4355.270 ;
      LAYER met4 ;
        RECT 3388.535 4313.330 3389.635 4314.035 ;
      LAYER met4 ;
        RECT 3390.035 4313.730 3395.485 4458.270 ;
      LAYER met4 ;
        RECT 3395.885 4457.000 3396.485 4458.670 ;
        RECT 3401.935 4458.365 3407.385 4458.670 ;
        RECT 3395.885 4313.330 3396.485 4314.035 ;
      LAYER met4 ;
        RECT 3396.885 4313.730 3401.535 4458.270 ;
      LAYER met4 ;
        RECT 3401.935 4457.000 3402.535 4458.365 ;
      LAYER met4 ;
        RECT 3402.935 4314.035 3406.385 4457.965 ;
      LAYER met4 ;
        RECT 3406.785 4457.000 3407.385 4458.365 ;
        RECT 3401.935 4313.635 3402.535 4314.035 ;
        RECT 3406.785 4313.635 3407.385 4314.035 ;
      LAYER met4 ;
        RECT 3407.785 4313.730 3412.435 4458.270 ;
      LAYER met4 ;
        RECT 3412.835 4457.000 3413.435 4458.670 ;
        RECT 3413.800 4446.065 3413.835 4457.065 ;
        RECT 3401.935 4313.330 3407.385 4313.635 ;
        RECT 3412.835 4313.330 3413.435 4314.035 ;
      LAYER met4 ;
        RECT 3413.835 4313.730 3418.485 4458.270 ;
      LAYER met4 ;
        RECT 3418.885 4457.000 3419.485 4458.670 ;
        RECT 3418.885 4313.330 3419.485 4314.035 ;
      LAYER met4 ;
        RECT 3419.885 4313.730 3423.335 4458.270 ;
      LAYER met4 ;
        RECT 3423.735 4457.000 3424.335 4458.670 ;
        RECT 3423.735 4313.330 3424.335 4314.035 ;
      LAYER met4 ;
        RECT 3424.735 4313.730 3428.185 4458.270 ;
      LAYER met4 ;
        RECT 3428.585 4457.000 3429.185 4458.670 ;
        RECT 3428.585 4313.330 3429.185 4314.035 ;
      LAYER met4 ;
        RECT 3429.585 4313.730 3434.235 4458.270 ;
      LAYER met4 ;
        RECT 3434.635 4457.000 3435.335 4458.670 ;
        RECT 3434.635 4313.330 3435.335 4314.035 ;
        RECT 3388.535 4311.990 3435.335 4313.330 ;
      LAYER met4 ;
        RECT 3435.735 4312.390 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
        RECT 3388.535 4268.310 3435.965 4311.990 ;
        RECT 3388.535 4236.670 3435.335 4268.310 ;
        RECT 3388.535 4236.030 3389.635 4236.670 ;
        RECT 152.035 4143.670 197.965 4215.330 ;
        RECT 147.275 3978.545 151.535 3980.065 ;
        RECT 147.275 3964.360 148.255 3978.545 ;
        RECT 0.000 3962.840 148.255 3964.360 ;
        RECT 0.000 3929.010 143.495 3962.840 ;
        RECT 0.000 3927.670 142.865 3929.010 ;
      LAYER met4 ;
        RECT 0.000 3926.000 24.215 3927.270 ;
      LAYER met4 ;
        RECT 24.615 3926.965 104.600 3927.670 ;
        RECT 0.000 3790.000 104.600 3926.000 ;
      LAYER met4 ;
        RECT 0.000 3788.730 24.215 3790.000 ;
      LAYER met4 ;
        RECT 24.615 3788.330 104.600 3788.970 ;
      LAYER met4 ;
        RECT 105.000 3788.730 129.965 3927.270 ;
      LAYER met4 ;
        RECT 130.365 3926.965 131.065 3927.670 ;
        RECT 130.365 3790.000 131.065 3926.000 ;
        RECT 130.365 3788.330 131.065 3788.970 ;
      LAYER met4 ;
        RECT 131.465 3788.730 135.915 3927.270 ;
      LAYER met4 ;
        RECT 136.315 3926.965 136.915 3927.670 ;
        RECT 136.315 3790.000 136.915 3926.000 ;
        RECT 136.315 3788.330 136.915 3788.970 ;
      LAYER met4 ;
        RECT 137.315 3788.730 141.765 3927.270 ;
      LAYER met4 ;
        RECT 142.165 3926.965 142.865 3927.670 ;
        RECT 142.165 3790.000 142.865 3926.000 ;
        RECT 142.165 3788.330 142.865 3788.970 ;
        RECT 0.000 3756.690 142.865 3788.330 ;
      LAYER met4 ;
        RECT 143.265 3757.090 143.595 3928.610 ;
      LAYER met4 ;
        RECT 0.000 3748.360 143.495 3756.690 ;
      LAYER met4 ;
        RECT 143.895 3748.760 146.875 3962.440 ;
      LAYER met4 ;
        RECT 147.275 3927.670 148.255 3962.840 ;
      LAYER met4 ;
        RECT 147.175 3926.000 148.355 3927.270 ;
      LAYER met4 ;
        RECT 147.175 3790.000 148.355 3926.000 ;
      LAYER met4 ;
        RECT 147.175 3788.730 148.355 3790.000 ;
      LAYER met4 ;
        RECT 147.275 3764.065 148.255 3788.330 ;
      LAYER met4 ;
        RECT 148.655 3764.465 151.635 3978.145 ;
        RECT 151.935 3973.090 152.265 4143.270 ;
      LAYER met4 ;
        RECT 152.665 4142.965 153.365 4143.670 ;
        RECT 152.665 4004.330 153.365 4004.970 ;
      LAYER met4 ;
        RECT 153.765 4004.730 158.415 4143.270 ;
      LAYER met4 ;
        RECT 158.815 4142.965 159.415 4143.670 ;
        RECT 158.815 4004.330 159.415 4004.970 ;
      LAYER met4 ;
        RECT 159.815 4004.730 163.265 4143.270 ;
      LAYER met4 ;
        RECT 163.665 4142.965 164.265 4143.670 ;
        RECT 163.665 4004.330 164.265 4004.970 ;
      LAYER met4 ;
        RECT 164.665 4004.730 168.115 4143.270 ;
      LAYER met4 ;
        RECT 168.515 4142.965 169.115 4143.670 ;
        RECT 168.515 4004.330 169.115 4004.970 ;
      LAYER met4 ;
        RECT 169.515 4004.730 174.165 4143.270 ;
      LAYER met4 ;
        RECT 174.565 4142.965 175.165 4143.670 ;
        RECT 180.615 4143.365 186.065 4143.670 ;
        RECT 174.565 4004.330 175.165 4004.970 ;
      LAYER met4 ;
        RECT 175.565 4004.730 180.215 4143.270 ;
      LAYER met4 ;
        RECT 180.615 4142.965 181.215 4143.365 ;
        RECT 185.465 4142.965 186.065 4143.365 ;
      LAYER met4 ;
        RECT 181.615 4004.970 185.065 4142.965 ;
      LAYER met4 ;
        RECT 180.615 4004.570 181.215 4004.970 ;
        RECT 185.465 4004.570 186.065 4004.970 ;
      LAYER met4 ;
        RECT 186.465 4004.730 191.115 4143.270 ;
      LAYER met4 ;
        RECT 191.515 4142.965 192.115 4143.670 ;
        RECT 180.615 4004.330 186.065 4004.570 ;
        RECT 191.515 4004.330 192.115 4004.970 ;
      LAYER met4 ;
        RECT 192.515 4004.730 197.965 4143.270 ;
        RECT 3390.035 4092.730 3395.485 4236.270 ;
      LAYER met4 ;
        RECT 3395.885 4236.030 3396.485 4236.670 ;
        RECT 3401.935 4236.430 3407.385 4236.670 ;
        RECT 3395.885 4092.330 3396.485 4093.035 ;
      LAYER met4 ;
        RECT 3396.885 4092.730 3401.535 4236.270 ;
      LAYER met4 ;
        RECT 3401.935 4236.030 3402.535 4236.430 ;
        RECT 3406.785 4236.030 3407.385 4236.430 ;
      LAYER met4 ;
        RECT 3402.935 4093.035 3406.385 4236.030 ;
      LAYER met4 ;
        RECT 3401.935 4092.635 3402.535 4093.035 ;
        RECT 3406.785 4092.635 3407.385 4093.035 ;
      LAYER met4 ;
        RECT 3407.785 4092.730 3412.435 4236.270 ;
      LAYER met4 ;
        RECT 3412.835 4236.030 3413.435 4236.670 ;
        RECT 3401.935 4092.330 3407.385 4092.635 ;
        RECT 3412.835 4092.330 3413.435 4093.035 ;
      LAYER met4 ;
        RECT 3413.835 4092.730 3418.485 4236.270 ;
      LAYER met4 ;
        RECT 3418.885 4236.030 3419.485 4236.670 ;
        RECT 3418.885 4092.330 3419.485 4093.035 ;
      LAYER met4 ;
        RECT 3419.885 4092.730 3423.335 4236.270 ;
      LAYER met4 ;
        RECT 3423.735 4236.030 3424.335 4236.670 ;
        RECT 3423.735 4092.330 3424.335 4093.035 ;
      LAYER met4 ;
        RECT 3424.735 4092.730 3428.185 4236.270 ;
      LAYER met4 ;
        RECT 3428.585 4236.030 3429.185 4236.670 ;
        RECT 3428.585 4092.330 3429.185 4093.035 ;
      LAYER met4 ;
        RECT 3429.585 4092.730 3434.235 4236.270 ;
      LAYER met4 ;
        RECT 3434.635 4236.030 3435.335 4236.670 ;
        RECT 3434.635 4092.330 3435.335 4093.035 ;
        RECT 3390.035 4020.670 3435.335 4092.330 ;
        RECT 198.365 4004.330 199.465 4004.970 ;
        RECT 152.665 3972.690 199.465 4004.330 ;
        RECT 152.035 3929.010 199.465 3972.690 ;
        RECT 147.275 3762.545 151.535 3764.065 ;
        RECT 147.275 3748.360 148.255 3762.545 ;
        RECT 0.000 3746.840 148.255 3748.360 ;
        RECT 0.000 3713.010 143.495 3746.840 ;
        RECT 0.000 3711.670 142.865 3713.010 ;
      LAYER met4 ;
        RECT 0.000 3710.000 24.215 3711.270 ;
      LAYER met4 ;
        RECT 24.615 3710.965 104.600 3711.670 ;
        RECT 0.000 3574.000 104.600 3710.000 ;
      LAYER met4 ;
        RECT 0.000 3572.730 24.215 3574.000 ;
      LAYER met4 ;
        RECT 24.615 3572.330 104.600 3572.970 ;
      LAYER met4 ;
        RECT 105.000 3572.730 129.965 3711.270 ;
      LAYER met4 ;
        RECT 130.365 3710.965 131.065 3711.670 ;
        RECT 130.365 3574.000 131.065 3710.000 ;
        RECT 130.365 3572.330 131.065 3572.970 ;
      LAYER met4 ;
        RECT 131.465 3572.730 135.915 3711.270 ;
      LAYER met4 ;
        RECT 136.315 3710.965 136.915 3711.670 ;
        RECT 136.315 3574.000 136.915 3710.000 ;
        RECT 136.315 3572.330 136.915 3572.970 ;
      LAYER met4 ;
        RECT 137.315 3572.730 141.765 3711.270 ;
      LAYER met4 ;
        RECT 142.165 3710.965 142.865 3711.670 ;
        RECT 142.165 3574.000 142.865 3710.000 ;
        RECT 142.165 3572.330 142.865 3572.970 ;
        RECT 0.000 3540.690 142.865 3572.330 ;
      LAYER met4 ;
        RECT 143.265 3541.090 143.595 3712.610 ;
      LAYER met4 ;
        RECT 0.000 3532.360 143.495 3540.690 ;
      LAYER met4 ;
        RECT 143.895 3532.760 146.875 3746.440 ;
      LAYER met4 ;
        RECT 147.275 3711.670 148.255 3746.840 ;
      LAYER met4 ;
        RECT 147.175 3710.000 148.355 3711.270 ;
      LAYER met4 ;
        RECT 147.175 3574.000 148.355 3710.000 ;
      LAYER met4 ;
        RECT 147.175 3572.730 148.355 3574.000 ;
      LAYER met4 ;
        RECT 147.275 3548.065 148.255 3572.330 ;
      LAYER met4 ;
        RECT 148.655 3548.465 151.635 3762.145 ;
        RECT 151.935 3757.090 152.265 3928.610 ;
      LAYER met4 ;
        RECT 152.665 3927.670 199.465 3929.010 ;
        RECT 152.665 3926.965 153.365 3927.670 ;
        RECT 152.665 3788.330 153.365 3788.970 ;
      LAYER met4 ;
        RECT 153.765 3788.730 158.415 3927.270 ;
      LAYER met4 ;
        RECT 158.815 3926.965 159.415 3927.670 ;
        RECT 158.815 3788.330 159.415 3788.970 ;
      LAYER met4 ;
        RECT 159.815 3788.730 163.265 3927.270 ;
      LAYER met4 ;
        RECT 163.665 3926.965 164.265 3927.670 ;
        RECT 163.665 3788.330 164.265 3788.970 ;
      LAYER met4 ;
        RECT 164.665 3788.730 168.115 3927.270 ;
      LAYER met4 ;
        RECT 168.515 3926.965 169.115 3927.670 ;
        RECT 168.515 3788.330 169.115 3788.970 ;
      LAYER met4 ;
        RECT 169.515 3788.730 174.165 3927.270 ;
      LAYER met4 ;
        RECT 174.565 3926.965 175.165 3927.670 ;
        RECT 180.615 3927.365 186.065 3927.670 ;
        RECT 174.565 3788.330 175.165 3788.970 ;
      LAYER met4 ;
        RECT 175.565 3788.730 180.215 3927.270 ;
      LAYER met4 ;
        RECT 180.615 3926.965 181.215 3927.365 ;
        RECT 185.465 3926.965 186.065 3927.365 ;
      LAYER met4 ;
        RECT 181.615 3788.970 185.065 3926.965 ;
      LAYER met4 ;
        RECT 180.615 3788.570 181.215 3788.970 ;
        RECT 185.465 3788.570 186.065 3788.970 ;
      LAYER met4 ;
        RECT 186.465 3788.730 191.115 3927.270 ;
      LAYER met4 ;
        RECT 191.515 3926.965 192.115 3927.670 ;
        RECT 180.615 3788.330 186.065 3788.570 ;
        RECT 191.515 3788.330 192.115 3788.970 ;
      LAYER met4 ;
        RECT 192.515 3788.730 197.965 3927.270 ;
      LAYER met4 ;
        RECT 198.365 3926.965 199.465 3927.670 ;
        RECT 3388.535 3876.330 3389.635 3877.035 ;
      LAYER met4 ;
        RECT 3390.035 3876.730 3395.485 4020.270 ;
      LAYER met4 ;
        RECT 3395.885 4019.965 3396.485 4020.670 ;
        RECT 3401.935 4020.365 3407.385 4020.670 ;
        RECT 3395.885 3876.330 3396.485 3877.035 ;
      LAYER met4 ;
        RECT 3396.885 3876.730 3401.535 4020.270 ;
      LAYER met4 ;
        RECT 3401.935 4019.965 3402.535 4020.365 ;
        RECT 3406.785 4019.965 3407.385 4020.365 ;
      LAYER met4 ;
        RECT 3402.935 3877.035 3406.385 4019.965 ;
      LAYER met4 ;
        RECT 3401.935 3876.635 3402.535 3877.035 ;
        RECT 3406.785 3876.635 3407.385 3877.035 ;
      LAYER met4 ;
        RECT 3407.785 3876.730 3412.435 4020.270 ;
      LAYER met4 ;
        RECT 3412.835 4019.965 3413.435 4020.670 ;
        RECT 3401.935 3876.330 3407.385 3876.635 ;
        RECT 3412.835 3876.330 3413.435 3877.035 ;
      LAYER met4 ;
        RECT 3413.835 3876.730 3418.485 4020.270 ;
      LAYER met4 ;
        RECT 3418.885 4019.965 3419.485 4020.670 ;
        RECT 3418.885 3876.330 3419.485 3877.035 ;
      LAYER met4 ;
        RECT 3419.885 3876.730 3423.335 4020.270 ;
      LAYER met4 ;
        RECT 3423.735 4019.965 3424.335 4020.670 ;
        RECT 3423.735 3876.330 3424.335 3877.035 ;
      LAYER met4 ;
        RECT 3424.735 3876.730 3428.185 4020.270 ;
      LAYER met4 ;
        RECT 3428.585 4019.965 3429.185 4020.670 ;
        RECT 3428.585 3876.330 3429.185 3877.035 ;
      LAYER met4 ;
        RECT 3429.585 3876.730 3434.235 4020.270 ;
      LAYER met4 ;
        RECT 3434.635 4019.965 3435.335 4020.670 ;
        RECT 3434.635 3876.330 3435.335 3877.035 ;
        RECT 3388.535 3874.990 3435.335 3876.330 ;
      LAYER met4 ;
        RECT 3435.735 3875.390 3436.065 4267.910 ;
        RECT 3436.365 4262.855 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.645 4842.000 3440.825 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4794.760 3440.825 4842.000 ;
      LAYER met4 ;
        RECT 3439.745 4716.515 3440.725 4794.360 ;
      LAYER met4 ;
        RECT 3439.645 4673.000 3440.825 4716.115 ;
      LAYER met4 ;
        RECT 3439.645 4532.000 3440.825 4673.000 ;
      LAYER met4 ;
        RECT 3439.645 4530.730 3440.825 4532.000 ;
      LAYER met4 ;
        RECT 3439.745 4458.670 3440.725 4530.330 ;
      LAYER met4 ;
        RECT 3439.645 4457.000 3440.825 4458.270 ;
      LAYER met4 ;
        RECT 3439.645 4315.000 3440.825 4457.000 ;
      LAYER met4 ;
        RECT 3439.645 4313.730 3440.825 4315.000 ;
      LAYER met4 ;
        RECT 3439.745 4278.160 3440.725 4313.330 ;
      LAYER met4 ;
        RECT 3441.125 4278.560 3444.105 5010.910 ;
        RECT 3444.405 4312.390 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4842.000 3445.835 4984.000 ;
        RECT 3445.135 4793.885 3445.835 4794.760 ;
      LAYER met4 ;
        RECT 3446.235 4794.285 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4842.000 3451.685 4984.000 ;
        RECT 3451.085 4793.885 3451.685 4794.760 ;
      LAYER met4 ;
        RECT 3452.085 4794.285 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4842.000 3457.635 4984.000 ;
        RECT 3456.935 4793.885 3457.635 4794.760 ;
      LAYER met4 ;
        RECT 3458.035 4794.285 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3483.400 4842.000 3588.000 4984.000 ;
        RECT 3483.400 4793.885 3563.385 4794.760 ;
        RECT 3445.135 4793.395 3563.385 4793.885 ;
      LAYER met4 ;
        RECT 3563.785 4793.795 3588.000 4842.000 ;
      LAYER met4 ;
        RECT 3445.135 4716.515 3588.000 4793.395 ;
        RECT 3445.135 4716.115 3445.835 4716.515 ;
        RECT 3451.085 4716.115 3451.685 4716.515 ;
        RECT 3456.935 4716.115 3457.635 4716.515 ;
        RECT 3483.400 4716.115 3563.385 4716.515 ;
        RECT 3445.135 4530.330 3445.835 4673.000 ;
      LAYER met4 ;
        RECT 3446.235 4530.730 3450.685 4716.115 ;
      LAYER met4 ;
        RECT 3451.085 4530.330 3451.685 4673.000 ;
      LAYER met4 ;
        RECT 3452.085 4530.730 3456.535 4716.115 ;
      LAYER met4 ;
        RECT 3456.935 4530.330 3457.635 4673.000 ;
      LAYER met4 ;
        RECT 3458.035 4530.730 3483.000 4716.115 ;
        RECT 3563.785 4673.000 3588.000 4716.115 ;
      LAYER met4 ;
        RECT 3483.400 4532.000 3588.000 4673.000 ;
        RECT 3483.400 4530.330 3563.385 4532.000 ;
      LAYER met4 ;
        RECT 3563.785 4530.730 3588.000 4532.000 ;
      LAYER met4 ;
        RECT 3445.135 4458.670 3588.000 4530.330 ;
        RECT 3445.135 4315.000 3445.835 4458.670 ;
        RECT 3445.135 4313.330 3445.835 4314.035 ;
      LAYER met4 ;
        RECT 3446.235 4313.730 3450.685 4458.270 ;
      LAYER met4 ;
        RECT 3451.085 4315.000 3451.685 4458.670 ;
        RECT 3451.085 4313.330 3451.685 4314.035 ;
      LAYER met4 ;
        RECT 3452.085 4313.730 3456.535 4458.270 ;
      LAYER met4 ;
        RECT 3456.935 4315.000 3457.635 4458.670 ;
        RECT 3456.935 4313.330 3457.635 4314.035 ;
      LAYER met4 ;
        RECT 3458.035 4313.730 3483.000 4458.270 ;
      LAYER met4 ;
        RECT 3483.400 4457.000 3563.385 4458.670 ;
        RECT 3563.750 4457.000 3563.785 4457.215 ;
      LAYER met4 ;
        RECT 3563.785 4457.000 3588.000 4458.270 ;
      LAYER met4 ;
        RECT 3483.400 4315.000 3588.000 4457.000 ;
        RECT 3483.400 4313.330 3563.385 4314.035 ;
      LAYER met4 ;
        RECT 3563.785 4313.730 3588.000 4315.000 ;
      LAYER met4 ;
        RECT 3445.135 4311.990 3588.000 4313.330 ;
        RECT 3444.505 4278.160 3588.000 4311.990 ;
        RECT 3439.745 4276.640 3588.000 4278.160 ;
        RECT 3439.745 4262.455 3440.725 4276.640 ;
        RECT 3436.465 4260.935 3440.725 4262.455 ;
        RECT 3388.535 3831.310 3435.965 3874.990 ;
        RECT 3388.535 3799.670 3435.335 3831.310 ;
        RECT 3388.535 3799.030 3389.635 3799.670 ;
        RECT 198.365 3788.330 199.465 3788.970 ;
        RECT 152.665 3756.690 199.465 3788.330 ;
        RECT 152.035 3713.010 199.465 3756.690 ;
        RECT 147.275 3546.545 151.535 3548.065 ;
        RECT 147.275 3532.360 148.255 3546.545 ;
        RECT 0.000 3530.840 148.255 3532.360 ;
        RECT 0.000 3497.010 143.495 3530.840 ;
        RECT 0.000 3495.670 142.865 3497.010 ;
      LAYER met4 ;
        RECT 0.000 3494.000 24.215 3495.270 ;
      LAYER met4 ;
        RECT 24.615 3494.965 104.600 3495.670 ;
        RECT 0.000 3357.000 104.600 3494.000 ;
      LAYER met4 ;
        RECT 0.000 3355.730 24.215 3357.000 ;
      LAYER met4 ;
        RECT 24.615 3355.330 104.600 3355.970 ;
      LAYER met4 ;
        RECT 105.000 3355.730 129.965 3495.270 ;
      LAYER met4 ;
        RECT 130.365 3494.965 131.065 3495.670 ;
        RECT 130.365 3357.000 131.065 3494.000 ;
        RECT 130.365 3355.330 131.065 3355.970 ;
      LAYER met4 ;
        RECT 131.465 3355.730 135.915 3495.270 ;
      LAYER met4 ;
        RECT 136.315 3494.965 136.915 3495.670 ;
        RECT 136.315 3357.000 136.915 3494.000 ;
        RECT 136.315 3355.330 136.915 3355.970 ;
      LAYER met4 ;
        RECT 137.315 3355.730 141.765 3495.270 ;
      LAYER met4 ;
        RECT 142.165 3494.965 142.865 3495.670 ;
        RECT 142.165 3357.000 142.865 3494.000 ;
        RECT 142.165 3355.330 142.865 3355.970 ;
        RECT 0.000 3323.690 142.865 3355.330 ;
      LAYER met4 ;
        RECT 143.265 3324.090 143.595 3496.610 ;
      LAYER met4 ;
        RECT 0.000 3315.360 143.495 3323.690 ;
      LAYER met4 ;
        RECT 143.895 3315.760 146.875 3530.440 ;
      LAYER met4 ;
        RECT 147.275 3495.670 148.255 3530.840 ;
      LAYER met4 ;
        RECT 147.175 3494.000 148.355 3495.270 ;
      LAYER met4 ;
        RECT 147.175 3357.000 148.355 3494.000 ;
      LAYER met4 ;
        RECT 147.175 3355.730 148.355 3357.000 ;
      LAYER met4 ;
        RECT 147.275 3331.065 148.255 3355.330 ;
      LAYER met4 ;
        RECT 148.655 3331.465 151.635 3546.145 ;
        RECT 151.935 3541.090 152.265 3712.610 ;
      LAYER met4 ;
        RECT 152.665 3711.670 199.465 3713.010 ;
        RECT 152.665 3710.965 153.365 3711.670 ;
        RECT 152.665 3572.330 153.365 3572.970 ;
      LAYER met4 ;
        RECT 153.765 3572.730 158.415 3711.270 ;
      LAYER met4 ;
        RECT 158.815 3710.965 159.415 3711.670 ;
        RECT 158.815 3572.330 159.415 3572.970 ;
      LAYER met4 ;
        RECT 159.815 3572.730 163.265 3711.270 ;
      LAYER met4 ;
        RECT 163.665 3710.965 164.265 3711.670 ;
        RECT 163.665 3572.330 164.265 3572.970 ;
      LAYER met4 ;
        RECT 164.665 3572.730 168.115 3711.270 ;
      LAYER met4 ;
        RECT 168.515 3710.965 169.115 3711.670 ;
        RECT 168.515 3572.330 169.115 3572.970 ;
      LAYER met4 ;
        RECT 169.515 3572.730 174.165 3711.270 ;
      LAYER met4 ;
        RECT 174.565 3710.965 175.165 3711.670 ;
        RECT 180.615 3711.365 186.065 3711.670 ;
        RECT 174.565 3572.330 175.165 3572.970 ;
      LAYER met4 ;
        RECT 175.565 3572.730 180.215 3711.270 ;
      LAYER met4 ;
        RECT 180.615 3710.965 181.215 3711.365 ;
        RECT 185.465 3710.965 186.065 3711.365 ;
      LAYER met4 ;
        RECT 181.615 3572.970 185.065 3710.965 ;
      LAYER met4 ;
        RECT 180.615 3572.570 181.215 3572.970 ;
        RECT 185.465 3572.570 186.065 3572.970 ;
      LAYER met4 ;
        RECT 186.465 3572.730 191.115 3711.270 ;
      LAYER met4 ;
        RECT 191.515 3710.965 192.115 3711.670 ;
        RECT 180.615 3572.330 186.065 3572.570 ;
        RECT 191.515 3572.330 192.115 3572.970 ;
      LAYER met4 ;
        RECT 192.515 3572.730 197.965 3711.270 ;
      LAYER met4 ;
        RECT 198.365 3710.965 199.465 3711.670 ;
        RECT 3388.535 3654.330 3389.635 3655.035 ;
      LAYER met4 ;
        RECT 3390.035 3654.730 3395.485 3799.270 ;
      LAYER met4 ;
        RECT 3395.885 3799.030 3396.485 3799.670 ;
        RECT 3401.935 3799.430 3407.385 3799.670 ;
        RECT 3395.885 3654.330 3396.485 3655.035 ;
      LAYER met4 ;
        RECT 3396.885 3654.730 3401.535 3799.270 ;
      LAYER met4 ;
        RECT 3401.935 3799.030 3402.535 3799.430 ;
        RECT 3406.785 3799.030 3407.385 3799.430 ;
      LAYER met4 ;
        RECT 3402.935 3655.035 3406.385 3799.030 ;
      LAYER met4 ;
        RECT 3401.935 3654.635 3402.535 3655.035 ;
        RECT 3406.785 3654.635 3407.385 3655.035 ;
      LAYER met4 ;
        RECT 3407.785 3654.730 3412.435 3799.270 ;
      LAYER met4 ;
        RECT 3412.835 3799.030 3413.435 3799.670 ;
        RECT 3401.935 3654.330 3407.385 3654.635 ;
        RECT 3412.835 3654.330 3413.435 3655.035 ;
      LAYER met4 ;
        RECT 3413.835 3654.730 3418.485 3799.270 ;
      LAYER met4 ;
        RECT 3418.885 3799.030 3419.485 3799.670 ;
        RECT 3418.885 3654.330 3419.485 3655.035 ;
      LAYER met4 ;
        RECT 3419.885 3654.730 3423.335 3799.270 ;
      LAYER met4 ;
        RECT 3423.735 3799.030 3424.335 3799.670 ;
        RECT 3423.735 3654.330 3424.335 3655.035 ;
      LAYER met4 ;
        RECT 3424.735 3654.730 3428.185 3799.270 ;
      LAYER met4 ;
        RECT 3428.585 3799.030 3429.185 3799.670 ;
        RECT 3428.585 3654.330 3429.185 3655.035 ;
      LAYER met4 ;
        RECT 3429.585 3654.730 3434.235 3799.270 ;
      LAYER met4 ;
        RECT 3434.635 3799.030 3435.335 3799.670 ;
        RECT 3434.635 3654.330 3435.335 3655.035 ;
        RECT 3388.535 3652.990 3435.335 3654.330 ;
      LAYER met4 ;
        RECT 3435.735 3653.390 3436.065 3830.910 ;
        RECT 3436.365 3825.855 3439.345 4260.535 ;
      LAYER met4 ;
        RECT 3439.745 4236.670 3440.725 4260.935 ;
      LAYER met4 ;
        RECT 3439.645 4235.000 3440.825 4236.270 ;
      LAYER met4 ;
        RECT 3439.645 4094.000 3440.825 4235.000 ;
      LAYER met4 ;
        RECT 3439.645 4092.730 3440.825 4094.000 ;
      LAYER met4 ;
        RECT 3439.745 4020.670 3440.725 4092.330 ;
      LAYER met4 ;
        RECT 3439.645 4019.000 3440.825 4020.270 ;
      LAYER met4 ;
        RECT 3439.645 3878.000 3440.825 4019.000 ;
      LAYER met4 ;
        RECT 3439.645 3876.730 3440.825 3878.000 ;
      LAYER met4 ;
        RECT 3439.745 3841.160 3440.725 3876.330 ;
      LAYER met4 ;
        RECT 3441.125 3841.560 3444.105 4276.240 ;
      LAYER met4 ;
        RECT 3444.505 4268.310 3588.000 4276.640 ;
      LAYER met4 ;
        RECT 3444.405 3875.390 3444.735 4267.910 ;
      LAYER met4 ;
        RECT 3445.135 4236.670 3588.000 4268.310 ;
        RECT 3445.135 4236.030 3445.835 4236.670 ;
        RECT 3445.135 4094.000 3445.835 4235.000 ;
        RECT 3445.135 4092.330 3445.835 4093.035 ;
      LAYER met4 ;
        RECT 3446.235 4092.730 3450.685 4236.270 ;
      LAYER met4 ;
        RECT 3451.085 4236.030 3451.685 4236.670 ;
        RECT 3451.085 4094.000 3451.685 4235.000 ;
        RECT 3451.085 4092.330 3451.685 4093.035 ;
      LAYER met4 ;
        RECT 3452.085 4092.730 3456.535 4236.270 ;
      LAYER met4 ;
        RECT 3456.935 4236.030 3457.635 4236.670 ;
        RECT 3456.935 4094.000 3457.635 4235.000 ;
        RECT 3456.935 4092.330 3457.635 4093.035 ;
      LAYER met4 ;
        RECT 3458.035 4092.730 3483.000 4236.270 ;
      LAYER met4 ;
        RECT 3483.400 4236.030 3563.385 4236.670 ;
      LAYER met4 ;
        RECT 3563.785 4235.000 3588.000 4236.270 ;
      LAYER met4 ;
        RECT 3483.400 4094.000 3588.000 4235.000 ;
        RECT 3483.400 4092.330 3563.385 4093.035 ;
      LAYER met4 ;
        RECT 3563.785 4092.730 3588.000 4094.000 ;
      LAYER met4 ;
        RECT 3445.135 4020.670 3588.000 4092.330 ;
        RECT 3445.135 4019.965 3445.835 4020.670 ;
        RECT 3445.135 3878.000 3445.835 4019.000 ;
        RECT 3445.135 3876.330 3445.835 3877.035 ;
      LAYER met4 ;
        RECT 3446.235 3876.730 3450.685 4020.270 ;
      LAYER met4 ;
        RECT 3451.085 4019.965 3451.685 4020.670 ;
        RECT 3451.085 3878.000 3451.685 4019.000 ;
        RECT 3451.085 3876.330 3451.685 3877.035 ;
      LAYER met4 ;
        RECT 3452.085 3876.730 3456.535 4020.270 ;
      LAYER met4 ;
        RECT 3456.935 4019.965 3457.635 4020.670 ;
        RECT 3456.935 3878.000 3457.635 4019.000 ;
        RECT 3456.935 3876.330 3457.635 3877.035 ;
      LAYER met4 ;
        RECT 3458.035 3876.730 3483.000 4020.270 ;
      LAYER met4 ;
        RECT 3483.400 4019.965 3563.385 4020.670 ;
      LAYER met4 ;
        RECT 3563.785 4019.000 3588.000 4020.270 ;
      LAYER met4 ;
        RECT 3483.400 3878.000 3588.000 4019.000 ;
        RECT 3483.400 3876.330 3563.385 3877.035 ;
      LAYER met4 ;
        RECT 3563.785 3876.730 3588.000 3878.000 ;
      LAYER met4 ;
        RECT 3445.135 3874.990 3588.000 3876.330 ;
        RECT 3444.505 3841.160 3588.000 3874.990 ;
        RECT 3439.745 3839.640 3588.000 3841.160 ;
        RECT 3439.745 3825.455 3440.725 3839.640 ;
        RECT 3436.465 3823.935 3440.725 3825.455 ;
        RECT 3388.535 3609.310 3435.965 3652.990 ;
        RECT 3388.535 3577.670 3435.335 3609.310 ;
        RECT 3388.535 3577.030 3389.635 3577.670 ;
        RECT 198.365 3572.330 199.465 3572.970 ;
        RECT 152.665 3540.690 199.465 3572.330 ;
        RECT 152.035 3497.010 199.465 3540.690 ;
        RECT 147.275 3329.545 151.535 3331.065 ;
        RECT 147.275 3315.360 148.255 3329.545 ;
        RECT 0.000 3313.840 148.255 3315.360 ;
        RECT 0.000 3280.010 143.495 3313.840 ;
        RECT 0.000 3278.670 142.865 3280.010 ;
      LAYER met4 ;
        RECT 0.000 3277.000 24.215 3278.270 ;
      LAYER met4 ;
        RECT 24.615 3277.965 104.600 3278.670 ;
        RECT 0.000 3141.000 104.600 3277.000 ;
      LAYER met4 ;
        RECT 0.000 3139.730 24.215 3141.000 ;
      LAYER met4 ;
        RECT 24.615 3139.330 104.600 3139.970 ;
      LAYER met4 ;
        RECT 105.000 3139.730 129.965 3278.270 ;
      LAYER met4 ;
        RECT 130.365 3277.965 131.065 3278.670 ;
        RECT 130.365 3141.000 131.065 3277.000 ;
        RECT 130.365 3139.330 131.065 3139.970 ;
      LAYER met4 ;
        RECT 131.465 3139.730 135.915 3278.270 ;
      LAYER met4 ;
        RECT 136.315 3277.965 136.915 3278.670 ;
        RECT 136.315 3141.000 136.915 3277.000 ;
        RECT 136.315 3139.330 136.915 3139.970 ;
      LAYER met4 ;
        RECT 137.315 3139.730 141.765 3278.270 ;
      LAYER met4 ;
        RECT 142.165 3277.965 142.865 3278.670 ;
        RECT 142.165 3141.000 142.865 3277.000 ;
        RECT 142.165 3139.330 142.865 3139.970 ;
        RECT 0.000 3107.690 142.865 3139.330 ;
      LAYER met4 ;
        RECT 143.265 3108.090 143.595 3279.610 ;
      LAYER met4 ;
        RECT 0.000 3099.360 143.495 3107.690 ;
      LAYER met4 ;
        RECT 143.895 3099.760 146.875 3313.440 ;
      LAYER met4 ;
        RECT 147.275 3278.670 148.255 3313.840 ;
      LAYER met4 ;
        RECT 147.175 3277.000 148.355 3278.270 ;
      LAYER met4 ;
        RECT 147.175 3141.000 148.355 3277.000 ;
      LAYER met4 ;
        RECT 147.175 3139.730 148.355 3141.000 ;
      LAYER met4 ;
        RECT 147.275 3115.065 148.255 3139.330 ;
      LAYER met4 ;
        RECT 148.655 3115.465 151.635 3329.145 ;
        RECT 151.935 3324.090 152.265 3496.610 ;
      LAYER met4 ;
        RECT 152.665 3495.670 199.465 3497.010 ;
        RECT 152.665 3494.965 153.365 3495.670 ;
        RECT 152.665 3355.330 153.365 3355.970 ;
      LAYER met4 ;
        RECT 153.765 3355.730 158.415 3495.270 ;
      LAYER met4 ;
        RECT 158.815 3494.965 159.415 3495.670 ;
        RECT 158.815 3355.330 159.415 3355.970 ;
      LAYER met4 ;
        RECT 159.815 3355.730 163.265 3495.270 ;
      LAYER met4 ;
        RECT 163.665 3494.965 164.265 3495.670 ;
        RECT 163.665 3355.330 164.265 3355.970 ;
      LAYER met4 ;
        RECT 164.665 3355.730 168.115 3495.270 ;
      LAYER met4 ;
        RECT 168.515 3494.965 169.115 3495.670 ;
        RECT 168.515 3355.330 169.115 3355.970 ;
      LAYER met4 ;
        RECT 169.515 3355.730 174.165 3495.270 ;
      LAYER met4 ;
        RECT 174.565 3494.965 175.165 3495.670 ;
        RECT 180.615 3495.365 186.065 3495.670 ;
        RECT 174.565 3355.330 175.165 3355.970 ;
      LAYER met4 ;
        RECT 175.565 3355.730 180.215 3495.270 ;
      LAYER met4 ;
        RECT 180.615 3494.965 181.215 3495.365 ;
        RECT 185.465 3494.965 186.065 3495.365 ;
      LAYER met4 ;
        RECT 181.615 3355.970 185.065 3494.965 ;
      LAYER met4 ;
        RECT 180.615 3355.570 181.215 3355.970 ;
        RECT 185.465 3355.570 186.065 3355.970 ;
      LAYER met4 ;
        RECT 186.465 3355.730 191.115 3495.270 ;
      LAYER met4 ;
        RECT 191.515 3494.965 192.115 3495.670 ;
        RECT 180.615 3355.330 186.065 3355.570 ;
        RECT 191.515 3355.330 192.115 3355.970 ;
      LAYER met4 ;
        RECT 192.515 3355.730 197.965 3495.270 ;
      LAYER met4 ;
        RECT 198.365 3494.965 199.465 3495.670 ;
        RECT 3388.535 3433.330 3389.635 3434.035 ;
      LAYER met4 ;
        RECT 3390.035 3433.730 3395.485 3577.270 ;
      LAYER met4 ;
        RECT 3395.885 3577.030 3396.485 3577.670 ;
        RECT 3401.935 3577.430 3407.385 3577.670 ;
        RECT 3395.885 3433.330 3396.485 3434.035 ;
      LAYER met4 ;
        RECT 3396.885 3433.730 3401.535 3577.270 ;
      LAYER met4 ;
        RECT 3401.935 3577.030 3402.535 3577.430 ;
        RECT 3406.785 3577.030 3407.385 3577.430 ;
      LAYER met4 ;
        RECT 3402.935 3434.035 3406.385 3577.030 ;
      LAYER met4 ;
        RECT 3401.935 3433.635 3402.535 3434.035 ;
        RECT 3406.785 3433.635 3407.385 3434.035 ;
      LAYER met4 ;
        RECT 3407.785 3433.730 3412.435 3577.270 ;
      LAYER met4 ;
        RECT 3412.835 3577.030 3413.435 3577.670 ;
        RECT 3401.935 3433.330 3407.385 3433.635 ;
        RECT 3412.835 3433.330 3413.435 3434.035 ;
      LAYER met4 ;
        RECT 3413.835 3433.730 3418.485 3577.270 ;
      LAYER met4 ;
        RECT 3418.885 3577.030 3419.485 3577.670 ;
        RECT 3418.885 3433.330 3419.485 3434.035 ;
      LAYER met4 ;
        RECT 3419.885 3433.730 3423.335 3577.270 ;
      LAYER met4 ;
        RECT 3423.735 3577.030 3424.335 3577.670 ;
        RECT 3423.735 3433.330 3424.335 3434.035 ;
      LAYER met4 ;
        RECT 3424.735 3433.730 3428.185 3577.270 ;
      LAYER met4 ;
        RECT 3428.585 3577.030 3429.185 3577.670 ;
        RECT 3428.585 3433.330 3429.185 3434.035 ;
      LAYER met4 ;
        RECT 3429.585 3433.730 3434.235 3577.270 ;
      LAYER met4 ;
        RECT 3434.635 3577.030 3435.335 3577.670 ;
        RECT 3434.635 3433.330 3435.335 3434.035 ;
        RECT 3388.535 3431.990 3435.335 3433.330 ;
      LAYER met4 ;
        RECT 3435.735 3432.390 3436.065 3608.910 ;
        RECT 3436.365 3603.855 3439.345 3823.535 ;
      LAYER met4 ;
        RECT 3439.745 3799.670 3440.725 3823.935 ;
      LAYER met4 ;
        RECT 3439.645 3798.000 3440.825 3799.270 ;
      LAYER met4 ;
        RECT 3439.645 3656.000 3440.825 3798.000 ;
      LAYER met4 ;
        RECT 3439.645 3654.730 3440.825 3656.000 ;
      LAYER met4 ;
        RECT 3439.745 3619.160 3440.725 3654.330 ;
      LAYER met4 ;
        RECT 3441.125 3619.560 3444.105 3839.240 ;
      LAYER met4 ;
        RECT 3444.505 3831.310 3588.000 3839.640 ;
      LAYER met4 ;
        RECT 3444.405 3653.390 3444.735 3830.910 ;
      LAYER met4 ;
        RECT 3445.135 3799.670 3588.000 3831.310 ;
        RECT 3445.135 3799.030 3445.835 3799.670 ;
        RECT 3445.135 3656.000 3445.835 3798.000 ;
        RECT 3445.135 3654.330 3445.835 3655.035 ;
      LAYER met4 ;
        RECT 3446.235 3654.730 3450.685 3799.270 ;
      LAYER met4 ;
        RECT 3451.085 3799.030 3451.685 3799.670 ;
        RECT 3451.085 3656.000 3451.685 3798.000 ;
        RECT 3451.085 3654.330 3451.685 3655.035 ;
      LAYER met4 ;
        RECT 3452.085 3654.730 3456.535 3799.270 ;
      LAYER met4 ;
        RECT 3456.935 3799.030 3457.635 3799.670 ;
        RECT 3456.935 3656.000 3457.635 3798.000 ;
        RECT 3456.935 3654.330 3457.635 3655.035 ;
      LAYER met4 ;
        RECT 3458.035 3654.730 3483.000 3799.270 ;
      LAYER met4 ;
        RECT 3483.400 3799.030 3563.385 3799.670 ;
      LAYER met4 ;
        RECT 3563.785 3798.000 3588.000 3799.270 ;
      LAYER met4 ;
        RECT 3483.400 3656.000 3588.000 3798.000 ;
        RECT 3483.400 3654.330 3563.385 3655.035 ;
      LAYER met4 ;
        RECT 3563.785 3654.730 3588.000 3656.000 ;
      LAYER met4 ;
        RECT 3445.135 3652.990 3588.000 3654.330 ;
        RECT 3444.505 3619.160 3588.000 3652.990 ;
        RECT 3439.745 3617.640 3588.000 3619.160 ;
        RECT 3439.745 3603.455 3440.725 3617.640 ;
        RECT 3436.465 3601.935 3440.725 3603.455 ;
        RECT 3388.535 3388.310 3435.965 3431.990 ;
        RECT 3388.535 3356.670 3435.335 3388.310 ;
        RECT 3388.535 3356.030 3389.635 3356.670 ;
        RECT 198.365 3355.330 199.465 3355.970 ;
        RECT 152.665 3323.690 199.465 3355.330 ;
        RECT 152.035 3280.010 199.465 3323.690 ;
        RECT 147.275 3113.545 151.535 3115.065 ;
        RECT 147.275 3099.360 148.255 3113.545 ;
        RECT 0.000 3097.840 148.255 3099.360 ;
        RECT 0.000 3064.010 143.495 3097.840 ;
        RECT 0.000 3062.670 142.865 3064.010 ;
      LAYER met4 ;
        RECT 0.000 3061.000 24.215 3062.270 ;
      LAYER met4 ;
        RECT 24.615 3061.965 104.600 3062.670 ;
        RECT 0.000 2925.000 104.600 3061.000 ;
      LAYER met4 ;
        RECT 0.000 2923.730 24.215 2925.000 ;
      LAYER met4 ;
        RECT 24.615 2923.330 104.600 2923.970 ;
      LAYER met4 ;
        RECT 105.000 2923.730 129.965 3062.270 ;
      LAYER met4 ;
        RECT 130.365 3061.965 131.065 3062.670 ;
        RECT 130.365 2925.000 131.065 3061.000 ;
        RECT 130.365 2923.330 131.065 2923.970 ;
      LAYER met4 ;
        RECT 131.465 2923.730 135.915 3062.270 ;
      LAYER met4 ;
        RECT 136.315 3061.965 136.915 3062.670 ;
        RECT 136.315 2925.000 136.915 3061.000 ;
        RECT 136.315 2923.330 136.915 2923.970 ;
      LAYER met4 ;
        RECT 137.315 2923.730 141.765 3062.270 ;
      LAYER met4 ;
        RECT 142.165 3061.965 142.865 3062.670 ;
        RECT 142.165 2925.000 142.865 3061.000 ;
        RECT 142.165 2923.330 142.865 2923.970 ;
        RECT 0.000 2891.690 142.865 2923.330 ;
      LAYER met4 ;
        RECT 143.265 2892.090 143.595 3063.610 ;
      LAYER met4 ;
        RECT 0.000 2883.360 143.495 2891.690 ;
      LAYER met4 ;
        RECT 143.895 2883.760 146.875 3097.440 ;
      LAYER met4 ;
        RECT 147.275 3062.670 148.255 3097.840 ;
      LAYER met4 ;
        RECT 147.175 3061.000 148.355 3062.270 ;
      LAYER met4 ;
        RECT 147.175 2925.000 148.355 3061.000 ;
      LAYER met4 ;
        RECT 147.175 2923.730 148.355 2925.000 ;
      LAYER met4 ;
        RECT 147.275 2899.065 148.255 2923.330 ;
      LAYER met4 ;
        RECT 148.655 2899.465 151.635 3113.145 ;
        RECT 151.935 3108.090 152.265 3279.610 ;
      LAYER met4 ;
        RECT 152.665 3278.670 199.465 3280.010 ;
        RECT 152.665 3277.965 153.365 3278.670 ;
        RECT 152.665 3139.330 153.365 3139.970 ;
      LAYER met4 ;
        RECT 153.765 3139.730 158.415 3278.270 ;
      LAYER met4 ;
        RECT 158.815 3277.965 159.415 3278.670 ;
        RECT 158.815 3139.330 159.415 3139.970 ;
      LAYER met4 ;
        RECT 159.815 3139.730 163.265 3278.270 ;
      LAYER met4 ;
        RECT 163.665 3277.965 164.265 3278.670 ;
        RECT 163.665 3139.330 164.265 3139.970 ;
      LAYER met4 ;
        RECT 164.665 3139.730 168.115 3278.270 ;
      LAYER met4 ;
        RECT 168.515 3277.965 169.115 3278.670 ;
        RECT 168.515 3139.330 169.115 3139.970 ;
      LAYER met4 ;
        RECT 169.515 3139.730 174.165 3278.270 ;
      LAYER met4 ;
        RECT 174.565 3277.965 175.165 3278.670 ;
        RECT 180.615 3278.365 186.065 3278.670 ;
        RECT 174.565 3139.330 175.165 3139.970 ;
      LAYER met4 ;
        RECT 175.565 3139.730 180.215 3278.270 ;
      LAYER met4 ;
        RECT 180.615 3277.965 181.215 3278.365 ;
        RECT 185.465 3277.965 186.065 3278.365 ;
      LAYER met4 ;
        RECT 181.615 3139.970 185.065 3277.965 ;
      LAYER met4 ;
        RECT 180.615 3139.570 181.215 3139.970 ;
        RECT 185.465 3139.570 186.065 3139.970 ;
      LAYER met4 ;
        RECT 186.465 3139.730 191.115 3278.270 ;
      LAYER met4 ;
        RECT 191.515 3277.965 192.115 3278.670 ;
        RECT 180.615 3139.330 186.065 3139.570 ;
        RECT 191.515 3139.330 192.115 3139.970 ;
      LAYER met4 ;
        RECT 192.515 3139.730 197.965 3278.270 ;
      LAYER met4 ;
        RECT 198.365 3277.965 199.465 3278.670 ;
        RECT 3388.535 3212.330 3389.635 3213.035 ;
      LAYER met4 ;
        RECT 3390.035 3212.730 3395.485 3356.270 ;
      LAYER met4 ;
        RECT 3395.885 3356.030 3396.485 3356.670 ;
        RECT 3401.935 3356.430 3407.385 3356.670 ;
        RECT 3395.885 3212.330 3396.485 3213.035 ;
      LAYER met4 ;
        RECT 3396.885 3212.730 3401.535 3356.270 ;
      LAYER met4 ;
        RECT 3401.935 3356.030 3402.535 3356.430 ;
        RECT 3406.785 3356.030 3407.385 3356.430 ;
      LAYER met4 ;
        RECT 3402.935 3213.035 3406.385 3356.030 ;
      LAYER met4 ;
        RECT 3401.935 3212.635 3402.535 3213.035 ;
        RECT 3406.785 3212.635 3407.385 3213.035 ;
      LAYER met4 ;
        RECT 3407.785 3212.730 3412.435 3356.270 ;
      LAYER met4 ;
        RECT 3412.835 3356.030 3413.435 3356.670 ;
        RECT 3401.935 3212.330 3407.385 3212.635 ;
        RECT 3412.835 3212.330 3413.435 3213.035 ;
      LAYER met4 ;
        RECT 3413.835 3212.730 3418.485 3356.270 ;
      LAYER met4 ;
        RECT 3418.885 3356.030 3419.485 3356.670 ;
        RECT 3418.885 3212.330 3419.485 3213.035 ;
      LAYER met4 ;
        RECT 3419.885 3212.730 3423.335 3356.270 ;
      LAYER met4 ;
        RECT 3423.735 3356.030 3424.335 3356.670 ;
        RECT 3423.735 3212.330 3424.335 3213.035 ;
      LAYER met4 ;
        RECT 3424.735 3212.730 3428.185 3356.270 ;
      LAYER met4 ;
        RECT 3428.585 3356.030 3429.185 3356.670 ;
        RECT 3428.585 3212.330 3429.185 3213.035 ;
      LAYER met4 ;
        RECT 3429.585 3212.730 3434.235 3356.270 ;
      LAYER met4 ;
        RECT 3434.635 3356.030 3435.335 3356.670 ;
        RECT 3434.635 3212.330 3435.335 3213.035 ;
        RECT 3388.535 3210.990 3435.335 3212.330 ;
      LAYER met4 ;
        RECT 3435.735 3211.390 3436.065 3387.910 ;
        RECT 3436.365 3382.855 3439.345 3601.535 ;
      LAYER met4 ;
        RECT 3439.745 3577.670 3440.725 3601.935 ;
      LAYER met4 ;
        RECT 3439.645 3576.000 3440.825 3577.270 ;
      LAYER met4 ;
        RECT 3439.645 3435.000 3440.825 3576.000 ;
      LAYER met4 ;
        RECT 3439.645 3433.730 3440.825 3435.000 ;
      LAYER met4 ;
        RECT 3439.745 3398.160 3440.725 3433.330 ;
      LAYER met4 ;
        RECT 3441.125 3398.560 3444.105 3617.240 ;
      LAYER met4 ;
        RECT 3444.505 3609.310 3588.000 3617.640 ;
      LAYER met4 ;
        RECT 3444.405 3432.390 3444.735 3608.910 ;
      LAYER met4 ;
        RECT 3445.135 3577.670 3588.000 3609.310 ;
        RECT 3445.135 3577.030 3445.835 3577.670 ;
        RECT 3445.135 3435.000 3445.835 3576.000 ;
        RECT 3445.135 3433.330 3445.835 3434.035 ;
      LAYER met4 ;
        RECT 3446.235 3433.730 3450.685 3577.270 ;
      LAYER met4 ;
        RECT 3451.085 3577.030 3451.685 3577.670 ;
        RECT 3451.085 3435.000 3451.685 3576.000 ;
        RECT 3451.085 3433.330 3451.685 3434.035 ;
      LAYER met4 ;
        RECT 3452.085 3433.730 3456.535 3577.270 ;
      LAYER met4 ;
        RECT 3456.935 3577.030 3457.635 3577.670 ;
        RECT 3456.935 3435.000 3457.635 3576.000 ;
        RECT 3456.935 3433.330 3457.635 3434.035 ;
      LAYER met4 ;
        RECT 3458.035 3433.730 3483.000 3577.270 ;
      LAYER met4 ;
        RECT 3483.400 3577.030 3563.385 3577.670 ;
      LAYER met4 ;
        RECT 3563.785 3576.000 3588.000 3577.270 ;
      LAYER met4 ;
        RECT 3483.400 3435.000 3588.000 3576.000 ;
        RECT 3483.400 3433.330 3563.385 3434.035 ;
      LAYER met4 ;
        RECT 3563.785 3433.730 3588.000 3435.000 ;
      LAYER met4 ;
        RECT 3445.135 3431.990 3588.000 3433.330 ;
        RECT 3444.505 3398.160 3588.000 3431.990 ;
        RECT 3439.745 3396.640 3588.000 3398.160 ;
        RECT 3439.745 3382.455 3440.725 3396.640 ;
        RECT 3436.465 3380.935 3440.725 3382.455 ;
        RECT 3388.535 3167.310 3435.965 3210.990 ;
        RECT 198.365 3139.330 199.465 3139.970 ;
        RECT 152.665 3107.690 199.465 3139.330 ;
        RECT 3388.535 3135.670 3435.335 3167.310 ;
        RECT 3388.535 3135.030 3389.635 3135.670 ;
        RECT 152.035 3064.010 199.465 3107.690 ;
        RECT 147.275 2897.545 151.535 2899.065 ;
        RECT 147.275 2883.360 148.255 2897.545 ;
        RECT 0.000 2881.840 148.255 2883.360 ;
        RECT 0.000 2848.010 143.495 2881.840 ;
        RECT 0.000 2846.670 142.865 2848.010 ;
      LAYER met4 ;
        RECT 0.000 2845.000 24.215 2846.270 ;
      LAYER met4 ;
        RECT 24.615 2845.965 104.600 2846.670 ;
        RECT 0.000 2709.000 104.600 2845.000 ;
      LAYER met4 ;
        RECT 0.000 2707.730 24.215 2709.000 ;
      LAYER met4 ;
        RECT 24.615 2707.330 104.600 2707.970 ;
      LAYER met4 ;
        RECT 105.000 2707.730 129.965 2846.270 ;
      LAYER met4 ;
        RECT 130.365 2845.965 131.065 2846.670 ;
        RECT 130.365 2709.000 131.065 2845.000 ;
        RECT 130.365 2707.330 131.065 2707.970 ;
      LAYER met4 ;
        RECT 131.465 2707.730 135.915 2846.270 ;
      LAYER met4 ;
        RECT 136.315 2845.965 136.915 2846.670 ;
        RECT 136.315 2709.000 136.915 2845.000 ;
        RECT 136.315 2707.330 136.915 2707.970 ;
      LAYER met4 ;
        RECT 137.315 2707.730 141.765 2846.270 ;
      LAYER met4 ;
        RECT 142.165 2845.965 142.865 2846.670 ;
        RECT 142.165 2709.000 142.865 2845.000 ;
        RECT 142.165 2707.330 142.865 2707.970 ;
        RECT 0.000 2675.690 142.865 2707.330 ;
      LAYER met4 ;
        RECT 143.265 2676.090 143.595 2847.610 ;
      LAYER met4 ;
        RECT 0.000 2667.360 143.495 2675.690 ;
      LAYER met4 ;
        RECT 143.895 2667.760 146.875 2881.440 ;
      LAYER met4 ;
        RECT 147.275 2846.670 148.255 2881.840 ;
      LAYER met4 ;
        RECT 147.175 2845.000 148.355 2846.270 ;
      LAYER met4 ;
        RECT 147.175 2709.000 148.355 2845.000 ;
      LAYER met4 ;
        RECT 147.175 2707.730 148.355 2709.000 ;
      LAYER met4 ;
        RECT 147.275 2683.065 148.255 2707.330 ;
      LAYER met4 ;
        RECT 148.655 2683.465 151.635 2897.145 ;
        RECT 151.935 2892.090 152.265 3063.610 ;
      LAYER met4 ;
        RECT 152.665 3062.670 199.465 3064.010 ;
        RECT 152.665 3061.965 153.365 3062.670 ;
        RECT 152.665 2923.330 153.365 2923.970 ;
      LAYER met4 ;
        RECT 153.765 2923.730 158.415 3062.270 ;
      LAYER met4 ;
        RECT 158.815 3061.965 159.415 3062.670 ;
        RECT 158.815 2923.330 159.415 2923.970 ;
      LAYER met4 ;
        RECT 159.815 2923.730 163.265 3062.270 ;
      LAYER met4 ;
        RECT 163.665 3061.965 164.265 3062.670 ;
        RECT 163.665 2923.330 164.265 2923.970 ;
      LAYER met4 ;
        RECT 164.665 2923.730 168.115 3062.270 ;
      LAYER met4 ;
        RECT 168.515 3061.965 169.115 3062.670 ;
        RECT 168.515 2923.330 169.115 2923.970 ;
      LAYER met4 ;
        RECT 169.515 2923.730 174.165 3062.270 ;
      LAYER met4 ;
        RECT 174.565 3061.965 175.165 3062.670 ;
        RECT 180.615 3062.365 186.065 3062.670 ;
        RECT 174.565 2923.330 175.165 2923.970 ;
      LAYER met4 ;
        RECT 175.565 2923.730 180.215 3062.270 ;
      LAYER met4 ;
        RECT 180.615 3061.965 181.215 3062.365 ;
        RECT 185.465 3061.965 186.065 3062.365 ;
      LAYER met4 ;
        RECT 181.615 2923.970 185.065 3061.965 ;
      LAYER met4 ;
        RECT 180.615 2923.570 181.215 2923.970 ;
        RECT 185.465 2923.570 186.065 2923.970 ;
      LAYER met4 ;
        RECT 186.465 2923.730 191.115 3062.270 ;
      LAYER met4 ;
        RECT 191.515 3061.965 192.115 3062.670 ;
        RECT 180.615 2923.330 186.065 2923.570 ;
        RECT 191.515 2923.330 192.115 2923.970 ;
      LAYER met4 ;
        RECT 192.515 2923.730 197.965 3062.270 ;
      LAYER met4 ;
        RECT 198.365 3061.965 199.465 3062.670 ;
        RECT 3388.535 2990.330 3389.635 2991.035 ;
      LAYER met4 ;
        RECT 3390.035 2990.730 3395.485 3135.270 ;
      LAYER met4 ;
        RECT 3395.885 3135.030 3396.485 3135.670 ;
        RECT 3401.935 3135.430 3407.385 3135.670 ;
        RECT 3395.885 2990.330 3396.485 2991.035 ;
      LAYER met4 ;
        RECT 3396.885 2990.730 3401.535 3135.270 ;
      LAYER met4 ;
        RECT 3401.935 3135.030 3402.535 3135.430 ;
        RECT 3406.785 3135.030 3407.385 3135.430 ;
      LAYER met4 ;
        RECT 3402.935 2991.035 3406.385 3135.030 ;
      LAYER met4 ;
        RECT 3401.935 2990.635 3402.535 2991.035 ;
        RECT 3406.785 2990.635 3407.385 2991.035 ;
      LAYER met4 ;
        RECT 3407.785 2990.730 3412.435 3135.270 ;
      LAYER met4 ;
        RECT 3412.835 3135.030 3413.435 3135.670 ;
        RECT 3401.935 2990.330 3407.385 2990.635 ;
        RECT 3412.835 2990.330 3413.435 2991.035 ;
      LAYER met4 ;
        RECT 3413.835 2990.730 3418.485 3135.270 ;
      LAYER met4 ;
        RECT 3418.885 3135.030 3419.485 3135.670 ;
        RECT 3418.885 2990.330 3419.485 2991.035 ;
      LAYER met4 ;
        RECT 3419.885 2990.730 3423.335 3135.270 ;
      LAYER met4 ;
        RECT 3423.735 3135.030 3424.335 3135.670 ;
        RECT 3423.735 2990.330 3424.335 2991.035 ;
      LAYER met4 ;
        RECT 3424.735 2990.730 3428.185 3135.270 ;
      LAYER met4 ;
        RECT 3428.585 3135.030 3429.185 3135.670 ;
        RECT 3428.585 2990.330 3429.185 2991.035 ;
      LAYER met4 ;
        RECT 3429.585 2990.730 3434.235 3135.270 ;
      LAYER met4 ;
        RECT 3434.635 3135.030 3435.335 3135.670 ;
        RECT 3434.635 2990.330 3435.335 2991.035 ;
        RECT 3388.535 2988.990 3435.335 2990.330 ;
      LAYER met4 ;
        RECT 3435.735 2989.390 3436.065 3166.910 ;
        RECT 3436.365 3161.855 3439.345 3380.535 ;
      LAYER met4 ;
        RECT 3439.745 3356.670 3440.725 3380.935 ;
      LAYER met4 ;
        RECT 3439.645 3355.000 3440.825 3356.270 ;
      LAYER met4 ;
        RECT 3439.645 3214.000 3440.825 3355.000 ;
      LAYER met4 ;
        RECT 3439.645 3212.730 3440.825 3214.000 ;
      LAYER met4 ;
        RECT 3439.745 3177.160 3440.725 3212.330 ;
      LAYER met4 ;
        RECT 3441.125 3177.560 3444.105 3396.240 ;
      LAYER met4 ;
        RECT 3444.505 3388.310 3588.000 3396.640 ;
      LAYER met4 ;
        RECT 3444.405 3211.390 3444.735 3387.910 ;
      LAYER met4 ;
        RECT 3445.135 3356.670 3588.000 3388.310 ;
        RECT 3445.135 3356.030 3445.835 3356.670 ;
        RECT 3445.135 3214.000 3445.835 3355.000 ;
        RECT 3445.135 3212.330 3445.835 3213.035 ;
      LAYER met4 ;
        RECT 3446.235 3212.730 3450.685 3356.270 ;
      LAYER met4 ;
        RECT 3451.085 3356.030 3451.685 3356.670 ;
        RECT 3451.085 3214.000 3451.685 3355.000 ;
        RECT 3451.085 3212.330 3451.685 3213.035 ;
      LAYER met4 ;
        RECT 3452.085 3212.730 3456.535 3356.270 ;
      LAYER met4 ;
        RECT 3456.935 3356.030 3457.635 3356.670 ;
        RECT 3456.935 3214.000 3457.635 3355.000 ;
        RECT 3456.935 3212.330 3457.635 3213.035 ;
      LAYER met4 ;
        RECT 3458.035 3212.730 3483.000 3356.270 ;
      LAYER met4 ;
        RECT 3483.400 3356.030 3563.385 3356.670 ;
      LAYER met4 ;
        RECT 3563.785 3355.000 3588.000 3356.270 ;
      LAYER met4 ;
        RECT 3483.400 3214.000 3588.000 3355.000 ;
        RECT 3483.400 3212.330 3563.385 3213.035 ;
      LAYER met4 ;
        RECT 3563.785 3212.730 3588.000 3214.000 ;
      LAYER met4 ;
        RECT 3445.135 3210.990 3588.000 3212.330 ;
        RECT 3444.505 3177.160 3588.000 3210.990 ;
        RECT 3439.745 3175.640 3588.000 3177.160 ;
        RECT 3439.745 3161.455 3440.725 3175.640 ;
        RECT 3436.465 3159.935 3440.725 3161.455 ;
        RECT 3388.535 2945.310 3435.965 2988.990 ;
        RECT 198.365 2923.330 199.465 2923.970 ;
        RECT 152.665 2891.690 199.465 2923.330 ;
        RECT 3388.535 2913.670 3435.335 2945.310 ;
        RECT 3388.535 2913.030 3389.635 2913.670 ;
        RECT 152.035 2848.010 199.465 2891.690 ;
        RECT 147.275 2681.545 151.535 2683.065 ;
        RECT 147.275 2667.360 148.255 2681.545 ;
        RECT 0.000 2665.840 148.255 2667.360 ;
        RECT 0.000 2632.010 143.495 2665.840 ;
        RECT 0.000 2630.670 142.865 2632.010 ;
      LAYER met4 ;
        RECT 0.000 2629.000 24.215 2630.270 ;
      LAYER met4 ;
        RECT 24.615 2629.965 104.600 2630.670 ;
        RECT 0.000 2492.000 104.600 2629.000 ;
      LAYER met4 ;
        RECT 0.000 2490.730 24.215 2492.000 ;
      LAYER met4 ;
        RECT 24.615 2490.330 104.600 2491.035 ;
      LAYER met4 ;
        RECT 105.000 2490.730 129.965 2630.270 ;
      LAYER met4 ;
        RECT 130.365 2629.965 131.065 2630.670 ;
        RECT 130.365 2492.000 131.065 2629.000 ;
        RECT 130.365 2490.330 131.065 2491.035 ;
      LAYER met4 ;
        RECT 131.465 2490.730 135.915 2630.270 ;
      LAYER met4 ;
        RECT 136.315 2629.965 136.915 2630.670 ;
        RECT 136.315 2492.000 136.915 2629.000 ;
        RECT 136.315 2490.330 136.915 2491.035 ;
      LAYER met4 ;
        RECT 137.315 2490.730 141.765 2630.270 ;
      LAYER met4 ;
        RECT 142.165 2629.965 142.865 2630.670 ;
        RECT 142.165 2492.000 142.865 2629.000 ;
        RECT 142.165 2490.330 142.865 2491.035 ;
        RECT 0.000 2418.670 142.865 2490.330 ;
      LAYER met4 ;
        RECT 0.000 2417.000 24.215 2418.270 ;
      LAYER met4 ;
        RECT 24.615 2417.965 104.600 2418.670 ;
        RECT 0.000 2282.465 104.600 2417.000 ;
        RECT 0.000 2281.000 0.035 2282.465 ;
        RECT 24.215 2281.000 104.600 2282.465 ;
        RECT 24.215 2280.785 24.250 2281.000 ;
        RECT 24.615 2279.330 104.600 2281.000 ;
      LAYER met4 ;
        RECT 105.000 2279.730 129.965 2418.270 ;
      LAYER met4 ;
        RECT 130.365 2417.965 131.065 2418.670 ;
        RECT 130.365 2279.330 131.065 2417.000 ;
      LAYER met4 ;
        RECT 131.465 2279.730 135.915 2418.270 ;
      LAYER met4 ;
        RECT 136.315 2417.965 136.915 2418.670 ;
        RECT 136.315 2279.330 136.915 2417.000 ;
      LAYER met4 ;
        RECT 137.315 2279.730 141.765 2418.270 ;
      LAYER met4 ;
        RECT 142.165 2417.965 142.865 2418.670 ;
        RECT 142.165 2279.330 142.865 2417.000 ;
        RECT 0.000 2207.670 142.865 2279.330 ;
      LAYER met4 ;
        RECT 0.000 2206.000 24.215 2207.270 ;
      LAYER met4 ;
        RECT 24.615 2206.000 104.600 2207.670 ;
        RECT 0.000 2070.000 104.600 2206.000 ;
      LAYER met4 ;
        RECT 0.000 2068.730 24.215 2070.000 ;
      LAYER met4 ;
        RECT 24.615 2068.330 104.600 2068.970 ;
      LAYER met4 ;
        RECT 105.000 2068.730 129.965 2207.270 ;
      LAYER met4 ;
        RECT 130.365 2070.000 131.065 2207.670 ;
        RECT 130.365 2068.330 131.065 2068.970 ;
      LAYER met4 ;
        RECT 131.465 2068.730 135.915 2207.270 ;
      LAYER met4 ;
        RECT 136.315 2070.000 136.915 2207.670 ;
        RECT 136.315 2068.330 136.915 2068.970 ;
      LAYER met4 ;
        RECT 137.315 2068.730 141.765 2207.270 ;
      LAYER met4 ;
        RECT 142.165 2070.000 142.865 2207.670 ;
        RECT 142.165 2068.330 142.865 2068.970 ;
        RECT 0.000 2036.690 142.865 2068.330 ;
        RECT 0.000 2028.360 143.495 2036.690 ;
      LAYER met4 ;
        RECT 143.895 2028.760 146.875 2665.440 ;
      LAYER met4 ;
        RECT 147.275 2630.670 148.255 2665.840 ;
      LAYER met4 ;
        RECT 147.175 2629.000 148.355 2630.270 ;
      LAYER met4 ;
        RECT 147.175 2492.000 148.355 2629.000 ;
      LAYER met4 ;
        RECT 147.175 2490.730 148.355 2492.000 ;
      LAYER met4 ;
        RECT 147.275 2418.670 148.255 2490.330 ;
      LAYER met4 ;
        RECT 147.175 2417.000 148.355 2418.270 ;
      LAYER met4 ;
        RECT 147.175 2281.000 148.355 2417.000 ;
      LAYER met4 ;
        RECT 147.175 2279.730 148.355 2281.000 ;
      LAYER met4 ;
        RECT 147.275 2207.670 148.255 2279.330 ;
      LAYER met4 ;
        RECT 147.175 2206.000 148.355 2207.270 ;
      LAYER met4 ;
        RECT 147.175 2070.000 148.355 2206.000 ;
      LAYER met4 ;
        RECT 147.175 2068.730 148.355 2070.000 ;
      LAYER met4 ;
        RECT 147.275 2044.065 148.255 2068.330 ;
      LAYER met4 ;
        RECT 148.655 2044.465 151.635 2681.145 ;
        RECT 151.935 2676.090 152.265 2847.610 ;
      LAYER met4 ;
        RECT 152.665 2846.670 199.465 2848.010 ;
        RECT 152.665 2845.965 153.365 2846.670 ;
        RECT 152.665 2707.330 153.365 2707.970 ;
      LAYER met4 ;
        RECT 153.765 2707.730 158.415 2846.270 ;
      LAYER met4 ;
        RECT 158.815 2845.965 159.415 2846.670 ;
        RECT 158.815 2707.330 159.415 2707.970 ;
      LAYER met4 ;
        RECT 159.815 2707.730 163.265 2846.270 ;
      LAYER met4 ;
        RECT 163.665 2845.965 164.265 2846.670 ;
        RECT 163.665 2707.330 164.265 2707.970 ;
      LAYER met4 ;
        RECT 164.665 2707.730 168.115 2846.270 ;
      LAYER met4 ;
        RECT 168.515 2845.965 169.115 2846.670 ;
        RECT 168.515 2707.330 169.115 2707.970 ;
      LAYER met4 ;
        RECT 169.515 2707.730 174.165 2846.270 ;
      LAYER met4 ;
        RECT 174.565 2845.965 175.165 2846.670 ;
        RECT 180.615 2846.365 186.065 2846.670 ;
        RECT 174.565 2707.330 175.165 2707.970 ;
      LAYER met4 ;
        RECT 175.565 2707.730 180.215 2846.270 ;
      LAYER met4 ;
        RECT 180.615 2845.965 181.215 2846.365 ;
        RECT 185.465 2845.965 186.065 2846.365 ;
      LAYER met4 ;
        RECT 181.615 2707.970 185.065 2845.965 ;
      LAYER met4 ;
        RECT 180.615 2707.570 181.215 2707.970 ;
        RECT 185.465 2707.570 186.065 2707.970 ;
      LAYER met4 ;
        RECT 186.465 2707.730 191.115 2846.270 ;
      LAYER met4 ;
        RECT 191.515 2845.965 192.115 2846.670 ;
        RECT 180.615 2707.330 186.065 2707.570 ;
        RECT 191.515 2707.330 192.115 2707.970 ;
      LAYER met4 ;
        RECT 192.515 2707.730 197.965 2846.270 ;
      LAYER met4 ;
        RECT 198.365 2845.965 199.465 2846.670 ;
        RECT 3388.535 2769.330 3389.635 2770.035 ;
      LAYER met4 ;
        RECT 3390.035 2769.730 3395.485 2913.270 ;
      LAYER met4 ;
        RECT 3395.885 2913.030 3396.485 2913.670 ;
        RECT 3401.935 2913.430 3407.385 2913.670 ;
        RECT 3395.885 2769.330 3396.485 2770.035 ;
      LAYER met4 ;
        RECT 3396.885 2769.730 3401.535 2913.270 ;
      LAYER met4 ;
        RECT 3401.935 2913.030 3402.535 2913.430 ;
        RECT 3406.785 2913.030 3407.385 2913.430 ;
      LAYER met4 ;
        RECT 3402.935 2770.035 3406.385 2913.030 ;
      LAYER met4 ;
        RECT 3401.935 2769.635 3402.535 2770.035 ;
        RECT 3406.785 2769.635 3407.385 2770.035 ;
      LAYER met4 ;
        RECT 3407.785 2769.730 3412.435 2913.270 ;
      LAYER met4 ;
        RECT 3412.835 2913.030 3413.435 2913.670 ;
        RECT 3401.935 2769.330 3407.385 2769.635 ;
        RECT 3412.835 2769.330 3413.435 2770.035 ;
      LAYER met4 ;
        RECT 3413.835 2769.730 3418.485 2913.270 ;
      LAYER met4 ;
        RECT 3418.885 2913.030 3419.485 2913.670 ;
        RECT 3418.885 2769.330 3419.485 2770.035 ;
      LAYER met4 ;
        RECT 3419.885 2769.730 3423.335 2913.270 ;
      LAYER met4 ;
        RECT 3423.735 2913.030 3424.335 2913.670 ;
        RECT 3423.735 2769.330 3424.335 2770.035 ;
      LAYER met4 ;
        RECT 3424.735 2769.730 3428.185 2913.270 ;
      LAYER met4 ;
        RECT 3428.585 2913.030 3429.185 2913.670 ;
        RECT 3428.585 2769.330 3429.185 2770.035 ;
      LAYER met4 ;
        RECT 3429.585 2769.730 3434.235 2913.270 ;
      LAYER met4 ;
        RECT 3434.635 2913.030 3435.335 2913.670 ;
        RECT 3434.635 2769.330 3435.335 2770.035 ;
        RECT 3388.535 2767.990 3435.335 2769.330 ;
      LAYER met4 ;
        RECT 3435.735 2768.390 3436.065 2944.910 ;
        RECT 3436.365 2939.855 3439.345 3159.535 ;
      LAYER met4 ;
        RECT 3439.745 3135.670 3440.725 3159.935 ;
      LAYER met4 ;
        RECT 3439.645 3134.000 3440.825 3135.270 ;
      LAYER met4 ;
        RECT 3439.645 2992.000 3440.825 3134.000 ;
      LAYER met4 ;
        RECT 3439.645 2990.730 3440.825 2992.000 ;
      LAYER met4 ;
        RECT 3439.745 2955.160 3440.725 2990.330 ;
      LAYER met4 ;
        RECT 3441.125 2955.560 3444.105 3175.240 ;
      LAYER met4 ;
        RECT 3444.505 3167.310 3588.000 3175.640 ;
      LAYER met4 ;
        RECT 3444.405 2989.390 3444.735 3166.910 ;
      LAYER met4 ;
        RECT 3445.135 3135.670 3588.000 3167.310 ;
        RECT 3445.135 3135.030 3445.835 3135.670 ;
        RECT 3445.135 2992.000 3445.835 3134.000 ;
        RECT 3445.135 2990.330 3445.835 2991.035 ;
      LAYER met4 ;
        RECT 3446.235 2990.730 3450.685 3135.270 ;
      LAYER met4 ;
        RECT 3451.085 3135.030 3451.685 3135.670 ;
        RECT 3451.085 2992.000 3451.685 3134.000 ;
        RECT 3451.085 2990.330 3451.685 2991.035 ;
      LAYER met4 ;
        RECT 3452.085 2990.730 3456.535 3135.270 ;
      LAYER met4 ;
        RECT 3456.935 3135.030 3457.635 3135.670 ;
        RECT 3456.935 2992.000 3457.635 3134.000 ;
        RECT 3456.935 2990.330 3457.635 2991.035 ;
      LAYER met4 ;
        RECT 3458.035 2990.730 3483.000 3135.270 ;
      LAYER met4 ;
        RECT 3483.400 3135.030 3563.385 3135.670 ;
      LAYER met4 ;
        RECT 3563.785 3134.000 3588.000 3135.270 ;
      LAYER met4 ;
        RECT 3483.400 2992.000 3588.000 3134.000 ;
        RECT 3483.400 2990.330 3563.385 2991.035 ;
      LAYER met4 ;
        RECT 3563.785 2990.730 3588.000 2992.000 ;
      LAYER met4 ;
        RECT 3445.135 2988.990 3588.000 2990.330 ;
        RECT 3444.505 2955.160 3588.000 2988.990 ;
        RECT 3439.745 2953.640 3588.000 2955.160 ;
        RECT 3439.745 2939.455 3440.725 2953.640 ;
        RECT 3436.465 2937.935 3440.725 2939.455 ;
        RECT 3388.535 2724.310 3435.965 2767.990 ;
        RECT 198.365 2707.330 199.465 2707.970 ;
        RECT 152.665 2675.690 199.465 2707.330 ;
        RECT 3388.535 2692.670 3435.335 2724.310 ;
        RECT 3388.535 2692.030 3389.635 2692.670 ;
        RECT 152.035 2632.010 199.465 2675.690 ;
        RECT 147.275 2042.545 151.535 2044.065 ;
        RECT 147.275 2028.360 148.255 2042.545 ;
        RECT 0.000 2026.840 148.255 2028.360 ;
        RECT 0.000 1993.010 143.495 2026.840 ;
        RECT 0.000 1991.670 142.865 1993.010 ;
      LAYER met4 ;
        RECT 0.000 1990.000 24.215 1991.270 ;
      LAYER met4 ;
        RECT 24.615 1990.965 104.600 1991.670 ;
        RECT 0.000 1854.000 104.600 1990.000 ;
      LAYER met4 ;
        RECT 0.000 1852.730 24.215 1854.000 ;
      LAYER met4 ;
        RECT 24.615 1852.330 104.600 1852.970 ;
      LAYER met4 ;
        RECT 105.000 1852.730 129.965 1991.270 ;
      LAYER met4 ;
        RECT 130.365 1990.965 131.065 1991.670 ;
        RECT 130.365 1854.000 131.065 1990.000 ;
        RECT 130.365 1852.330 131.065 1852.970 ;
      LAYER met4 ;
        RECT 131.465 1852.730 135.915 1991.270 ;
      LAYER met4 ;
        RECT 136.315 1990.965 136.915 1991.670 ;
        RECT 136.315 1854.000 136.915 1990.000 ;
        RECT 136.315 1852.330 136.915 1852.970 ;
      LAYER met4 ;
        RECT 137.315 1852.730 141.765 1991.270 ;
      LAYER met4 ;
        RECT 142.165 1990.965 142.865 1991.670 ;
        RECT 142.165 1854.000 142.865 1990.000 ;
        RECT 142.165 1852.330 142.865 1852.970 ;
        RECT 0.000 1820.690 142.865 1852.330 ;
      LAYER met4 ;
        RECT 143.265 1821.090 143.595 1992.610 ;
      LAYER met4 ;
        RECT 0.000 1812.360 143.495 1820.690 ;
      LAYER met4 ;
        RECT 143.895 1812.760 146.875 2026.440 ;
      LAYER met4 ;
        RECT 147.275 1991.670 148.255 2026.840 ;
      LAYER met4 ;
        RECT 147.175 1990.000 148.355 1991.270 ;
      LAYER met4 ;
        RECT 147.175 1854.000 148.355 1990.000 ;
      LAYER met4 ;
        RECT 147.175 1852.730 148.355 1854.000 ;
      LAYER met4 ;
        RECT 147.275 1828.065 148.255 1852.330 ;
      LAYER met4 ;
        RECT 148.655 1828.465 151.635 2042.145 ;
        RECT 151.935 2037.090 152.265 2631.610 ;
      LAYER met4 ;
        RECT 152.665 2630.670 199.465 2632.010 ;
        RECT 152.665 2629.965 153.365 2630.670 ;
        RECT 152.665 2490.330 153.365 2491.035 ;
      LAYER met4 ;
        RECT 153.765 2490.730 158.415 2630.270 ;
      LAYER met4 ;
        RECT 158.815 2629.965 159.415 2630.670 ;
        RECT 158.815 2490.330 159.415 2491.035 ;
      LAYER met4 ;
        RECT 159.815 2490.730 163.265 2630.270 ;
      LAYER met4 ;
        RECT 163.665 2629.965 164.265 2630.670 ;
        RECT 163.665 2490.330 164.265 2491.035 ;
      LAYER met4 ;
        RECT 164.665 2490.730 168.115 2630.270 ;
      LAYER met4 ;
        RECT 168.515 2629.965 169.115 2630.670 ;
        RECT 168.515 2490.330 169.115 2491.035 ;
      LAYER met4 ;
        RECT 169.515 2490.730 174.165 2630.270 ;
      LAYER met4 ;
        RECT 174.565 2629.965 175.165 2630.670 ;
        RECT 180.615 2630.365 186.065 2630.670 ;
        RECT 174.565 2490.330 175.165 2491.035 ;
      LAYER met4 ;
        RECT 175.565 2490.730 180.215 2630.270 ;
      LAYER met4 ;
        RECT 180.615 2629.965 181.215 2630.365 ;
        RECT 185.465 2629.965 186.065 2630.365 ;
      LAYER met4 ;
        RECT 181.615 2491.035 185.065 2629.965 ;
      LAYER met4 ;
        RECT 180.615 2490.635 181.215 2491.035 ;
        RECT 185.465 2490.635 186.065 2491.035 ;
      LAYER met4 ;
        RECT 186.465 2490.730 191.115 2630.270 ;
      LAYER met4 ;
        RECT 191.515 2629.965 192.115 2630.670 ;
        RECT 180.615 2490.330 186.065 2490.635 ;
        RECT 191.515 2490.330 192.115 2491.035 ;
      LAYER met4 ;
        RECT 192.515 2490.730 197.965 2630.270 ;
      LAYER met4 ;
        RECT 198.365 2629.965 199.465 2630.670 ;
      LAYER met4 ;
        RECT 3390.035 2548.730 3395.485 2692.270 ;
      LAYER met4 ;
        RECT 3395.885 2692.030 3396.485 2692.670 ;
        RECT 3401.935 2692.430 3407.385 2692.670 ;
        RECT 3395.885 2548.330 3396.485 2549.035 ;
      LAYER met4 ;
        RECT 3396.885 2548.730 3401.535 2692.270 ;
      LAYER met4 ;
        RECT 3401.935 2692.030 3402.535 2692.430 ;
        RECT 3406.785 2692.030 3407.385 2692.430 ;
      LAYER met4 ;
        RECT 3402.935 2549.035 3406.385 2692.030 ;
      LAYER met4 ;
        RECT 3401.935 2548.635 3402.535 2549.035 ;
        RECT 3406.785 2548.635 3407.385 2549.035 ;
      LAYER met4 ;
        RECT 3407.785 2548.730 3412.435 2692.270 ;
      LAYER met4 ;
        RECT 3412.835 2692.030 3413.435 2692.670 ;
        RECT 3401.935 2548.330 3407.385 2548.635 ;
        RECT 3412.835 2548.330 3413.435 2549.035 ;
      LAYER met4 ;
        RECT 3413.835 2548.730 3418.485 2692.270 ;
      LAYER met4 ;
        RECT 3418.885 2692.030 3419.485 2692.670 ;
        RECT 3418.885 2548.330 3419.485 2549.035 ;
      LAYER met4 ;
        RECT 3419.885 2548.730 3423.335 2692.270 ;
      LAYER met4 ;
        RECT 3423.735 2692.030 3424.335 2692.670 ;
        RECT 3423.735 2548.330 3424.335 2549.035 ;
      LAYER met4 ;
        RECT 3424.735 2548.730 3428.185 2692.270 ;
      LAYER met4 ;
        RECT 3428.585 2692.030 3429.185 2692.670 ;
        RECT 3428.585 2548.330 3429.185 2549.035 ;
      LAYER met4 ;
        RECT 3429.585 2548.730 3434.235 2692.270 ;
      LAYER met4 ;
        RECT 3434.635 2692.030 3435.335 2692.670 ;
        RECT 3434.635 2548.330 3435.335 2549.035 ;
        RECT 152.665 2418.670 197.965 2490.330 ;
        RECT 3390.035 2476.670 3435.335 2548.330 ;
        RECT 152.665 2417.965 153.365 2418.670 ;
        RECT 152.665 2279.330 153.365 2281.000 ;
      LAYER met4 ;
        RECT 153.765 2279.730 158.415 2418.270 ;
      LAYER met4 ;
        RECT 158.815 2417.965 159.415 2418.670 ;
        RECT 158.815 2279.330 159.415 2281.000 ;
      LAYER met4 ;
        RECT 159.815 2279.730 163.265 2418.270 ;
      LAYER met4 ;
        RECT 163.665 2417.965 164.265 2418.670 ;
        RECT 168.515 2417.965 169.115 2418.670 ;
        RECT 163.665 2279.330 164.265 2281.000 ;
        RECT 168.515 2279.330 169.115 2281.000 ;
      LAYER met4 ;
        RECT 169.515 2279.730 174.165 2418.270 ;
      LAYER met4 ;
        RECT 174.565 2417.965 175.165 2418.670 ;
        RECT 180.615 2418.365 186.065 2418.670 ;
        RECT 174.165 2280.935 174.200 2291.935 ;
        RECT 174.565 2279.330 175.165 2281.000 ;
      LAYER met4 ;
        RECT 175.565 2279.730 180.215 2418.270 ;
      LAYER met4 ;
        RECT 180.615 2417.965 181.215 2418.365 ;
        RECT 185.465 2417.965 186.065 2418.365 ;
        RECT 191.515 2417.965 192.115 2418.670 ;
      LAYER met4 ;
        RECT 3390.035 2331.730 3395.485 2476.270 ;
      LAYER met4 ;
        RECT 3395.885 2475.965 3396.485 2476.670 ;
        RECT 3401.935 2476.365 3407.385 2476.670 ;
        RECT 3395.885 2331.330 3396.485 2333.000 ;
      LAYER met4 ;
        RECT 3396.885 2331.730 3401.535 2476.270 ;
      LAYER met4 ;
        RECT 3401.935 2475.965 3402.535 2476.365 ;
        RECT 3406.785 2475.965 3407.385 2476.365 ;
        RECT 3401.935 2331.635 3402.535 2333.000 ;
      LAYER met4 ;
        RECT 3402.935 2332.035 3406.385 2475.965 ;
      LAYER met4 ;
        RECT 3406.785 2331.635 3407.385 2333.000 ;
      LAYER met4 ;
        RECT 3407.785 2331.730 3412.435 2476.270 ;
      LAYER met4 ;
        RECT 3412.835 2475.965 3413.435 2476.670 ;
        RECT 3401.935 2331.330 3407.385 2331.635 ;
        RECT 3412.835 2331.330 3413.435 2333.000 ;
      LAYER met4 ;
        RECT 3413.835 2331.730 3418.485 2476.270 ;
      LAYER met4 ;
        RECT 3418.885 2475.965 3419.485 2476.670 ;
        RECT 3418.885 2331.330 3419.485 2333.000 ;
      LAYER met4 ;
        RECT 3419.885 2331.730 3423.335 2476.270 ;
      LAYER met4 ;
        RECT 3423.735 2475.965 3424.335 2476.670 ;
        RECT 3423.735 2331.330 3424.335 2333.000 ;
      LAYER met4 ;
        RECT 3424.735 2331.730 3428.185 2476.270 ;
      LAYER met4 ;
        RECT 3428.585 2475.965 3429.185 2476.670 ;
        RECT 3428.585 2331.330 3429.185 2333.000 ;
        RECT 3429.550 2332.930 3429.585 2343.975 ;
      LAYER met4 ;
        RECT 3429.585 2331.730 3434.235 2476.270 ;
      LAYER met4 ;
        RECT 3434.635 2475.965 3435.335 2476.670 ;
        RECT 3434.635 2331.330 3435.335 2333.000 ;
        RECT 180.615 2279.635 181.215 2281.000 ;
        RECT 185.465 2279.635 186.065 2281.000 ;
        RECT 180.615 2279.330 186.065 2279.635 ;
        RECT 191.515 2279.330 192.115 2281.000 ;
        RECT 152.665 2207.670 197.965 2279.330 ;
        RECT 3390.035 2259.670 3435.335 2331.330 ;
        RECT 152.665 2206.000 153.365 2207.670 ;
        RECT 152.665 2068.330 153.365 2068.970 ;
      LAYER met4 ;
        RECT 153.765 2068.730 158.415 2207.270 ;
      LAYER met4 ;
        RECT 158.415 2195.025 158.450 2206.070 ;
        RECT 158.815 2206.000 159.415 2207.670 ;
        RECT 158.815 2068.330 159.415 2068.970 ;
      LAYER met4 ;
        RECT 159.815 2068.730 163.265 2207.270 ;
      LAYER met4 ;
        RECT 163.665 2206.000 164.265 2207.670 ;
        RECT 163.665 2068.330 164.265 2068.970 ;
      LAYER met4 ;
        RECT 164.665 2068.730 168.115 2207.270 ;
      LAYER met4 ;
        RECT 168.515 2206.000 169.115 2207.670 ;
        RECT 168.515 2068.330 169.115 2068.970 ;
      LAYER met4 ;
        RECT 169.515 2068.730 174.165 2207.270 ;
      LAYER met4 ;
        RECT 174.565 2206.000 175.165 2207.670 ;
        RECT 180.615 2207.365 186.065 2207.670 ;
        RECT 174.565 2068.330 175.165 2068.970 ;
      LAYER met4 ;
        RECT 175.565 2068.730 180.215 2207.270 ;
      LAYER met4 ;
        RECT 180.615 2206.000 181.215 2207.365 ;
      LAYER met4 ;
        RECT 181.615 2068.970 185.065 2206.965 ;
      LAYER met4 ;
        RECT 185.465 2206.000 186.065 2207.365 ;
        RECT 180.615 2068.570 181.215 2068.970 ;
        RECT 185.465 2068.570 186.065 2068.970 ;
      LAYER met4 ;
        RECT 186.465 2068.730 191.115 2207.270 ;
      LAYER met4 ;
        RECT 191.515 2206.000 192.115 2207.670 ;
        RECT 180.615 2068.330 186.065 2068.570 ;
        RECT 191.515 2068.330 192.115 2068.970 ;
      LAYER met4 ;
        RECT 192.515 2068.730 197.965 2207.270 ;
        RECT 3390.035 2115.730 3395.485 2259.270 ;
      LAYER met4 ;
        RECT 3395.885 2258.000 3396.485 2259.670 ;
        RECT 3401.935 2259.365 3407.385 2259.670 ;
        RECT 3401.935 2258.000 3402.535 2259.365 ;
        RECT 3406.785 2258.000 3407.385 2259.365 ;
        RECT 3395.885 2115.330 3396.485 2116.035 ;
        RECT 3401.935 2115.635 3402.535 2116.035 ;
        RECT 3406.785 2115.635 3407.385 2116.035 ;
      LAYER met4 ;
        RECT 3407.785 2115.730 3412.435 2259.270 ;
      LAYER met4 ;
        RECT 3412.835 2258.000 3413.435 2259.670 ;
        RECT 3413.800 2247.065 3413.835 2258.065 ;
        RECT 3401.935 2115.330 3407.385 2115.635 ;
        RECT 3412.835 2115.330 3413.435 2116.035 ;
      LAYER met4 ;
        RECT 3413.835 2115.730 3418.485 2259.270 ;
      LAYER met4 ;
        RECT 3418.885 2258.000 3419.485 2259.670 ;
        RECT 3418.885 2115.330 3419.485 2116.035 ;
      LAYER met4 ;
        RECT 3419.885 2115.730 3423.335 2259.270 ;
      LAYER met4 ;
        RECT 3423.735 2258.000 3424.335 2259.670 ;
        RECT 3423.735 2115.330 3424.335 2116.035 ;
      LAYER met4 ;
        RECT 3424.735 2115.730 3428.185 2259.270 ;
      LAYER met4 ;
        RECT 3428.585 2258.000 3429.185 2259.670 ;
        RECT 3428.585 2115.330 3429.185 2116.035 ;
      LAYER met4 ;
        RECT 3429.585 2115.730 3434.235 2259.270 ;
      LAYER met4 ;
        RECT 3434.635 2258.000 3435.335 2259.670 ;
        RECT 3434.635 2115.330 3435.335 2116.035 ;
      LAYER met4 ;
        RECT 3435.735 2115.730 3436.065 2723.910 ;
        RECT 3436.365 2718.855 3439.345 2937.535 ;
      LAYER met4 ;
        RECT 3439.745 2913.670 3440.725 2937.935 ;
      LAYER met4 ;
        RECT 3439.645 2912.000 3440.825 2913.270 ;
      LAYER met4 ;
        RECT 3439.645 2771.000 3440.825 2912.000 ;
      LAYER met4 ;
        RECT 3439.645 2769.730 3440.825 2771.000 ;
      LAYER met4 ;
        RECT 3439.745 2734.160 3440.725 2769.330 ;
      LAYER met4 ;
        RECT 3441.125 2734.560 3444.105 2953.240 ;
      LAYER met4 ;
        RECT 3444.505 2945.310 3588.000 2953.640 ;
      LAYER met4 ;
        RECT 3444.405 2768.390 3444.735 2944.910 ;
      LAYER met4 ;
        RECT 3445.135 2913.670 3588.000 2945.310 ;
        RECT 3445.135 2913.030 3445.835 2913.670 ;
        RECT 3445.135 2771.000 3445.835 2912.000 ;
        RECT 3445.135 2769.330 3445.835 2770.035 ;
      LAYER met4 ;
        RECT 3446.235 2769.730 3450.685 2913.270 ;
      LAYER met4 ;
        RECT 3451.085 2913.030 3451.685 2913.670 ;
        RECT 3451.085 2771.000 3451.685 2912.000 ;
        RECT 3451.085 2769.330 3451.685 2770.035 ;
      LAYER met4 ;
        RECT 3452.085 2769.730 3456.535 2913.270 ;
      LAYER met4 ;
        RECT 3456.935 2913.030 3457.635 2913.670 ;
        RECT 3456.935 2771.000 3457.635 2912.000 ;
        RECT 3456.935 2769.330 3457.635 2770.035 ;
      LAYER met4 ;
        RECT 3458.035 2769.730 3483.000 2913.270 ;
      LAYER met4 ;
        RECT 3483.400 2913.030 3563.385 2913.670 ;
      LAYER met4 ;
        RECT 3563.785 2912.000 3588.000 2913.270 ;
      LAYER met4 ;
        RECT 3483.400 2771.000 3588.000 2912.000 ;
        RECT 3483.400 2769.330 3563.385 2770.035 ;
      LAYER met4 ;
        RECT 3563.785 2769.730 3588.000 2771.000 ;
      LAYER met4 ;
        RECT 3445.135 2767.990 3588.000 2769.330 ;
        RECT 3444.505 2734.160 3588.000 2767.990 ;
        RECT 3439.745 2732.640 3588.000 2734.160 ;
        RECT 3439.745 2718.455 3440.725 2732.640 ;
        RECT 3436.465 2716.935 3440.725 2718.455 ;
      LAYER met4 ;
        RECT 3369.335 2099.650 3369.665 2099.665 ;
        RECT 3369.335 2099.350 3370.570 2099.650 ;
        RECT 3369.335 2099.335 3369.665 2099.350 ;
        RECT 3369.335 2096.250 3369.665 2096.265 ;
        RECT 3370.270 2096.250 3370.570 2099.350 ;
        RECT 3369.335 2095.950 3370.570 2096.250 ;
        RECT 3369.335 2095.935 3369.665 2095.950 ;
      LAYER met4 ;
        RECT 198.365 2068.330 199.465 2068.970 ;
        RECT 152.665 2036.690 199.465 2068.330 ;
        RECT 3390.035 2043.670 3435.965 2115.330 ;
        RECT 152.035 1993.010 199.465 2036.690 ;
        RECT 147.275 1826.545 151.535 1828.065 ;
        RECT 147.275 1812.360 148.255 1826.545 ;
        RECT 0.000 1810.840 148.255 1812.360 ;
        RECT 0.000 1777.010 143.495 1810.840 ;
        RECT 0.000 1775.670 142.865 1777.010 ;
      LAYER met4 ;
        RECT 0.000 1774.000 24.215 1775.270 ;
      LAYER met4 ;
        RECT 24.615 1774.965 104.600 1775.670 ;
        RECT 0.000 1637.000 104.600 1774.000 ;
      LAYER met4 ;
        RECT 0.000 1635.730 24.215 1637.000 ;
      LAYER met4 ;
        RECT 24.615 1635.330 104.600 1635.970 ;
      LAYER met4 ;
        RECT 105.000 1635.730 129.965 1775.270 ;
      LAYER met4 ;
        RECT 130.365 1774.965 131.065 1775.670 ;
        RECT 130.365 1637.000 131.065 1774.000 ;
        RECT 130.365 1635.330 131.065 1635.970 ;
      LAYER met4 ;
        RECT 131.465 1635.730 135.915 1775.270 ;
      LAYER met4 ;
        RECT 136.315 1774.965 136.915 1775.670 ;
        RECT 136.315 1637.000 136.915 1774.000 ;
        RECT 136.315 1635.330 136.915 1635.970 ;
      LAYER met4 ;
        RECT 137.315 1635.730 141.765 1775.270 ;
      LAYER met4 ;
        RECT 142.165 1774.965 142.865 1775.670 ;
        RECT 142.165 1637.000 142.865 1774.000 ;
        RECT 142.165 1635.330 142.865 1635.970 ;
        RECT 0.000 1603.690 142.865 1635.330 ;
      LAYER met4 ;
        RECT 143.265 1604.090 143.595 1776.610 ;
      LAYER met4 ;
        RECT 0.000 1595.360 143.495 1603.690 ;
      LAYER met4 ;
        RECT 143.895 1595.760 146.875 1810.440 ;
      LAYER met4 ;
        RECT 147.275 1775.670 148.255 1810.840 ;
      LAYER met4 ;
        RECT 147.175 1774.000 148.355 1775.270 ;
      LAYER met4 ;
        RECT 147.175 1637.000 148.355 1774.000 ;
      LAYER met4 ;
        RECT 147.175 1635.730 148.355 1637.000 ;
      LAYER met4 ;
        RECT 147.275 1611.065 148.255 1635.330 ;
      LAYER met4 ;
        RECT 148.655 1611.465 151.635 1826.145 ;
        RECT 151.935 1821.090 152.265 1992.610 ;
      LAYER met4 ;
        RECT 152.665 1991.670 199.465 1993.010 ;
        RECT 152.665 1990.965 153.365 1991.670 ;
        RECT 152.665 1852.330 153.365 1852.970 ;
      LAYER met4 ;
        RECT 153.765 1852.730 158.415 1991.270 ;
      LAYER met4 ;
        RECT 158.815 1990.965 159.415 1991.670 ;
        RECT 158.815 1852.330 159.415 1852.970 ;
      LAYER met4 ;
        RECT 159.815 1852.730 163.265 1991.270 ;
      LAYER met4 ;
        RECT 163.665 1990.965 164.265 1991.670 ;
        RECT 163.665 1852.330 164.265 1852.970 ;
      LAYER met4 ;
        RECT 164.665 1852.730 168.115 1991.270 ;
      LAYER met4 ;
        RECT 168.515 1990.965 169.115 1991.670 ;
        RECT 168.515 1852.330 169.115 1852.970 ;
      LAYER met4 ;
        RECT 169.515 1852.730 174.165 1991.270 ;
      LAYER met4 ;
        RECT 174.565 1990.965 175.165 1991.670 ;
        RECT 180.615 1991.365 186.065 1991.670 ;
        RECT 174.565 1852.330 175.165 1852.970 ;
      LAYER met4 ;
        RECT 175.565 1852.730 180.215 1991.270 ;
      LAYER met4 ;
        RECT 180.615 1990.965 181.215 1991.365 ;
        RECT 185.465 1990.965 186.065 1991.365 ;
      LAYER met4 ;
        RECT 181.615 1852.970 185.065 1990.965 ;
      LAYER met4 ;
        RECT 180.615 1852.570 181.215 1852.970 ;
        RECT 185.465 1852.570 186.065 1852.970 ;
      LAYER met4 ;
        RECT 186.465 1852.730 191.115 1991.270 ;
      LAYER met4 ;
        RECT 191.515 1990.965 192.115 1991.670 ;
        RECT 180.615 1852.330 186.065 1852.570 ;
        RECT 191.515 1852.330 192.115 1852.970 ;
      LAYER met4 ;
        RECT 192.515 1852.730 197.965 1991.270 ;
      LAYER met4 ;
        RECT 198.365 1990.965 199.465 1991.670 ;
        RECT 3388.535 1898.330 3389.635 1899.035 ;
      LAYER met4 ;
        RECT 3390.035 1898.730 3395.485 2043.270 ;
      LAYER met4 ;
        RECT 3395.885 2042.965 3396.485 2043.670 ;
        RECT 3401.935 2043.365 3407.385 2043.670 ;
        RECT 3395.885 1898.330 3396.485 1899.035 ;
      LAYER met4 ;
        RECT 3396.885 1898.730 3401.535 2043.270 ;
      LAYER met4 ;
        RECT 3401.935 2042.965 3402.535 2043.365 ;
        RECT 3406.785 2042.965 3407.385 2043.365 ;
      LAYER met4 ;
        RECT 3402.935 1899.035 3406.385 2042.965 ;
      LAYER met4 ;
        RECT 3401.935 1898.635 3402.535 1899.035 ;
        RECT 3406.785 1898.635 3407.385 1899.035 ;
      LAYER met4 ;
        RECT 3407.785 1898.730 3412.435 2043.270 ;
      LAYER met4 ;
        RECT 3412.835 2042.965 3413.435 2043.670 ;
        RECT 3401.935 1898.330 3407.385 1898.635 ;
        RECT 3412.835 1898.330 3413.435 1899.035 ;
      LAYER met4 ;
        RECT 3413.835 1898.730 3418.485 2043.270 ;
      LAYER met4 ;
        RECT 3418.885 2042.965 3419.485 2043.670 ;
        RECT 3418.885 1898.330 3419.485 1899.035 ;
      LAYER met4 ;
        RECT 3419.885 1898.730 3423.335 2043.270 ;
      LAYER met4 ;
        RECT 3423.735 2042.965 3424.335 2043.670 ;
        RECT 3423.735 1898.330 3424.335 1899.035 ;
      LAYER met4 ;
        RECT 3424.735 1898.730 3428.185 2043.270 ;
      LAYER met4 ;
        RECT 3428.585 2042.965 3429.185 2043.670 ;
        RECT 3428.585 1898.330 3429.185 1899.035 ;
      LAYER met4 ;
        RECT 3429.585 1898.730 3434.235 2043.270 ;
      LAYER met4 ;
        RECT 3434.635 2042.965 3435.335 2043.670 ;
        RECT 3434.635 1898.330 3435.335 1899.035 ;
        RECT 3388.535 1896.990 3435.335 1898.330 ;
      LAYER met4 ;
        RECT 3435.735 1897.390 3436.065 2043.270 ;
      LAYER met4 ;
        RECT 3388.535 1853.310 3435.965 1896.990 ;
        RECT 198.365 1852.330 199.465 1852.970 ;
        RECT 152.665 1820.690 199.465 1852.330 ;
        RECT 3388.535 1821.670 3435.335 1853.310 ;
        RECT 3388.535 1821.030 3389.635 1821.670 ;
        RECT 152.035 1777.010 199.465 1820.690 ;
        RECT 147.275 1609.545 151.535 1611.065 ;
        RECT 147.275 1595.360 148.255 1609.545 ;
        RECT 0.000 1593.840 148.255 1595.360 ;
        RECT 0.000 1560.010 143.495 1593.840 ;
        RECT 0.000 1558.670 142.865 1560.010 ;
      LAYER met4 ;
        RECT 0.000 1557.000 24.215 1558.270 ;
      LAYER met4 ;
        RECT 24.615 1557.965 104.600 1558.670 ;
        RECT 0.000 1421.000 104.600 1557.000 ;
      LAYER met4 ;
        RECT 0.000 1419.730 24.215 1421.000 ;
      LAYER met4 ;
        RECT 24.615 1419.330 104.600 1419.970 ;
      LAYER met4 ;
        RECT 105.000 1419.730 129.965 1558.270 ;
      LAYER met4 ;
        RECT 130.365 1557.965 131.065 1558.670 ;
        RECT 130.365 1421.000 131.065 1557.000 ;
        RECT 130.365 1419.330 131.065 1419.970 ;
      LAYER met4 ;
        RECT 131.465 1419.730 135.915 1558.270 ;
      LAYER met4 ;
        RECT 136.315 1557.965 136.915 1558.670 ;
        RECT 136.315 1421.000 136.915 1557.000 ;
        RECT 136.315 1419.330 136.915 1419.970 ;
      LAYER met4 ;
        RECT 137.315 1419.730 141.765 1558.270 ;
      LAYER met4 ;
        RECT 142.165 1557.965 142.865 1558.670 ;
        RECT 142.165 1421.000 142.865 1557.000 ;
        RECT 142.165 1419.330 142.865 1419.970 ;
        RECT 0.000 1387.690 142.865 1419.330 ;
      LAYER met4 ;
        RECT 143.265 1388.090 143.595 1559.610 ;
      LAYER met4 ;
        RECT 0.000 1379.360 143.495 1387.690 ;
      LAYER met4 ;
        RECT 143.895 1379.760 146.875 1593.440 ;
      LAYER met4 ;
        RECT 147.275 1558.670 148.255 1593.840 ;
      LAYER met4 ;
        RECT 147.175 1557.000 148.355 1558.270 ;
      LAYER met4 ;
        RECT 147.175 1421.000 148.355 1557.000 ;
      LAYER met4 ;
        RECT 147.175 1419.730 148.355 1421.000 ;
      LAYER met4 ;
        RECT 147.275 1395.065 148.255 1419.330 ;
      LAYER met4 ;
        RECT 148.655 1395.465 151.635 1609.145 ;
        RECT 151.935 1604.090 152.265 1776.610 ;
      LAYER met4 ;
        RECT 152.665 1775.670 199.465 1777.010 ;
        RECT 152.665 1774.965 153.365 1775.670 ;
        RECT 152.665 1635.330 153.365 1635.970 ;
      LAYER met4 ;
        RECT 153.765 1635.730 158.415 1775.270 ;
      LAYER met4 ;
        RECT 158.815 1774.965 159.415 1775.670 ;
        RECT 158.815 1635.330 159.415 1635.970 ;
      LAYER met4 ;
        RECT 159.815 1635.730 163.265 1775.270 ;
      LAYER met4 ;
        RECT 163.665 1774.965 164.265 1775.670 ;
        RECT 163.665 1635.330 164.265 1635.970 ;
      LAYER met4 ;
        RECT 164.665 1635.730 168.115 1775.270 ;
      LAYER met4 ;
        RECT 168.515 1774.965 169.115 1775.670 ;
        RECT 168.515 1635.330 169.115 1635.970 ;
      LAYER met4 ;
        RECT 169.515 1635.730 174.165 1775.270 ;
      LAYER met4 ;
        RECT 174.565 1774.965 175.165 1775.670 ;
        RECT 180.615 1775.365 186.065 1775.670 ;
        RECT 174.565 1635.330 175.165 1635.970 ;
      LAYER met4 ;
        RECT 175.565 1635.730 180.215 1775.270 ;
      LAYER met4 ;
        RECT 180.615 1774.965 181.215 1775.365 ;
        RECT 185.465 1774.965 186.065 1775.365 ;
      LAYER met4 ;
        RECT 181.615 1635.970 185.065 1774.965 ;
      LAYER met4 ;
        RECT 180.615 1635.570 181.215 1635.970 ;
        RECT 185.465 1635.570 186.065 1635.970 ;
      LAYER met4 ;
        RECT 186.465 1635.730 191.115 1775.270 ;
      LAYER met4 ;
        RECT 191.515 1774.965 192.115 1775.670 ;
        RECT 180.615 1635.330 186.065 1635.570 ;
        RECT 191.515 1635.330 192.115 1635.970 ;
      LAYER met4 ;
        RECT 192.515 1635.730 197.965 1775.270 ;
      LAYER met4 ;
        RECT 198.365 1774.965 199.465 1775.670 ;
        RECT 3388.535 1677.330 3389.635 1678.035 ;
      LAYER met4 ;
        RECT 3390.035 1677.730 3395.485 1821.270 ;
      LAYER met4 ;
        RECT 3395.885 1821.030 3396.485 1821.670 ;
        RECT 3401.935 1821.430 3407.385 1821.670 ;
        RECT 3395.885 1677.330 3396.485 1678.035 ;
      LAYER met4 ;
        RECT 3396.885 1677.730 3401.535 1821.270 ;
      LAYER met4 ;
        RECT 3401.935 1821.030 3402.535 1821.430 ;
        RECT 3406.785 1821.030 3407.385 1821.430 ;
      LAYER met4 ;
        RECT 3402.935 1678.035 3406.385 1821.030 ;
      LAYER met4 ;
        RECT 3401.935 1677.635 3402.535 1678.035 ;
        RECT 3406.785 1677.635 3407.385 1678.035 ;
      LAYER met4 ;
        RECT 3407.785 1677.730 3412.435 1821.270 ;
      LAYER met4 ;
        RECT 3412.835 1821.030 3413.435 1821.670 ;
        RECT 3401.935 1677.330 3407.385 1677.635 ;
        RECT 3412.835 1677.330 3413.435 1678.035 ;
      LAYER met4 ;
        RECT 3413.835 1677.730 3418.485 1821.270 ;
      LAYER met4 ;
        RECT 3418.885 1821.030 3419.485 1821.670 ;
        RECT 3418.885 1677.330 3419.485 1678.035 ;
      LAYER met4 ;
        RECT 3419.885 1677.730 3423.335 1821.270 ;
      LAYER met4 ;
        RECT 3423.735 1821.030 3424.335 1821.670 ;
        RECT 3423.735 1677.330 3424.335 1678.035 ;
      LAYER met4 ;
        RECT 3424.735 1677.730 3428.185 1821.270 ;
      LAYER met4 ;
        RECT 3428.585 1821.030 3429.185 1821.670 ;
        RECT 3428.585 1677.330 3429.185 1678.035 ;
      LAYER met4 ;
        RECT 3429.585 1677.730 3434.235 1821.270 ;
      LAYER met4 ;
        RECT 3434.635 1821.030 3435.335 1821.670 ;
        RECT 3434.635 1677.330 3435.335 1678.035 ;
        RECT 3388.535 1675.990 3435.335 1677.330 ;
      LAYER met4 ;
        RECT 3435.735 1676.390 3436.065 1852.910 ;
        RECT 3436.365 1847.855 3439.345 2716.535 ;
      LAYER met4 ;
        RECT 3439.745 2692.670 3440.725 2716.935 ;
      LAYER met4 ;
        RECT 3439.645 2691.000 3440.825 2692.270 ;
      LAYER met4 ;
        RECT 3439.645 2550.000 3440.825 2691.000 ;
      LAYER met4 ;
        RECT 3439.645 2548.730 3440.825 2550.000 ;
      LAYER met4 ;
        RECT 3439.745 2476.670 3440.725 2548.330 ;
      LAYER met4 ;
        RECT 3439.645 2475.000 3440.825 2476.270 ;
      LAYER met4 ;
        RECT 3439.645 2333.000 3440.825 2475.000 ;
      LAYER met4 ;
        RECT 3439.645 2331.730 3440.825 2333.000 ;
      LAYER met4 ;
        RECT 3439.745 2259.670 3440.725 2331.330 ;
      LAYER met4 ;
        RECT 3439.645 2258.000 3440.825 2259.270 ;
      LAYER met4 ;
        RECT 3439.645 2117.000 3440.825 2258.000 ;
      LAYER met4 ;
        RECT 3439.645 2115.730 3440.825 2117.000 ;
      LAYER met4 ;
        RECT 3439.745 2043.670 3440.725 2115.330 ;
      LAYER met4 ;
        RECT 3439.645 2042.000 3440.825 2043.270 ;
      LAYER met4 ;
        RECT 3439.645 1900.000 3440.825 2042.000 ;
      LAYER met4 ;
        RECT 3439.645 1898.730 3440.825 1900.000 ;
      LAYER met4 ;
        RECT 3439.745 1863.160 3440.725 1898.330 ;
      LAYER met4 ;
        RECT 3441.125 1863.560 3444.105 2732.240 ;
      LAYER met4 ;
        RECT 3444.505 2724.310 3588.000 2732.640 ;
        RECT 3445.135 2692.670 3588.000 2724.310 ;
        RECT 3445.135 2692.030 3445.835 2692.670 ;
        RECT 3445.135 2550.000 3445.835 2691.000 ;
        RECT 3445.135 2548.330 3445.835 2549.035 ;
      LAYER met4 ;
        RECT 3446.235 2548.730 3450.685 2692.270 ;
      LAYER met4 ;
        RECT 3451.085 2692.030 3451.685 2692.670 ;
        RECT 3451.085 2550.000 3451.685 2691.000 ;
        RECT 3451.085 2548.330 3451.685 2549.035 ;
      LAYER met4 ;
        RECT 3452.085 2548.730 3456.535 2692.270 ;
      LAYER met4 ;
        RECT 3456.935 2692.030 3457.635 2692.670 ;
        RECT 3456.935 2550.000 3457.635 2691.000 ;
        RECT 3456.935 2548.330 3457.635 2549.035 ;
      LAYER met4 ;
        RECT 3458.035 2548.730 3483.000 2692.270 ;
      LAYER met4 ;
        RECT 3483.400 2692.030 3563.385 2692.670 ;
      LAYER met4 ;
        RECT 3563.785 2691.000 3588.000 2692.270 ;
      LAYER met4 ;
        RECT 3483.400 2550.000 3588.000 2691.000 ;
        RECT 3483.400 2548.330 3563.385 2549.035 ;
      LAYER met4 ;
        RECT 3563.785 2548.730 3588.000 2550.000 ;
      LAYER met4 ;
        RECT 3445.135 2476.670 3588.000 2548.330 ;
        RECT 3445.135 2475.965 3445.835 2476.670 ;
        RECT 3445.135 2331.330 3445.835 2475.000 ;
      LAYER met4 ;
        RECT 3446.235 2331.730 3450.685 2476.270 ;
      LAYER met4 ;
        RECT 3451.085 2475.965 3451.685 2476.670 ;
        RECT 3451.085 2331.330 3451.685 2475.000 ;
      LAYER met4 ;
        RECT 3452.085 2331.730 3456.535 2476.270 ;
      LAYER met4 ;
        RECT 3456.935 2475.965 3457.635 2476.670 ;
        RECT 3456.935 2331.330 3457.635 2475.000 ;
      LAYER met4 ;
        RECT 3458.035 2331.730 3483.000 2476.270 ;
      LAYER met4 ;
        RECT 3483.400 2475.965 3563.385 2476.670 ;
      LAYER met4 ;
        RECT 3563.785 2475.000 3588.000 2476.270 ;
      LAYER met4 ;
        RECT 3483.400 2333.000 3588.000 2475.000 ;
        RECT 3483.400 2331.330 3563.385 2333.000 ;
      LAYER met4 ;
        RECT 3563.785 2331.730 3588.000 2333.000 ;
      LAYER met4 ;
        RECT 3445.135 2259.670 3588.000 2331.330 ;
        RECT 3445.135 2117.000 3445.835 2259.670 ;
        RECT 3445.135 2115.330 3445.835 2116.035 ;
      LAYER met4 ;
        RECT 3446.235 2115.730 3450.685 2259.270 ;
      LAYER met4 ;
        RECT 3451.085 2117.000 3451.685 2259.670 ;
        RECT 3451.085 2115.330 3451.685 2116.035 ;
      LAYER met4 ;
        RECT 3452.085 2115.730 3456.535 2259.270 ;
      LAYER met4 ;
        RECT 3456.935 2117.000 3457.635 2259.670 ;
        RECT 3456.935 2115.330 3457.635 2116.035 ;
      LAYER met4 ;
        RECT 3458.035 2115.730 3483.000 2259.270 ;
      LAYER met4 ;
        RECT 3483.400 2258.000 3563.385 2259.670 ;
        RECT 3563.750 2258.000 3563.785 2258.215 ;
      LAYER met4 ;
        RECT 3563.785 2258.000 3588.000 2259.270 ;
      LAYER met4 ;
        RECT 3483.400 2117.000 3588.000 2258.000 ;
        RECT 3483.400 2115.330 3563.385 2116.035 ;
      LAYER met4 ;
        RECT 3563.785 2115.730 3588.000 2117.000 ;
      LAYER met4 ;
        RECT 3444.505 2043.670 3588.000 2115.330 ;
      LAYER met4 ;
        RECT 3444.405 1897.390 3444.735 2043.270 ;
      LAYER met4 ;
        RECT 3445.135 2042.965 3445.835 2043.670 ;
        RECT 3445.135 1900.000 3445.835 2042.000 ;
        RECT 3445.135 1898.330 3445.835 1899.035 ;
      LAYER met4 ;
        RECT 3446.235 1898.730 3450.685 2043.270 ;
      LAYER met4 ;
        RECT 3451.085 2042.965 3451.685 2043.670 ;
        RECT 3451.085 1900.000 3451.685 2042.000 ;
        RECT 3451.085 1898.330 3451.685 1899.035 ;
      LAYER met4 ;
        RECT 3452.085 1898.730 3456.535 2043.270 ;
      LAYER met4 ;
        RECT 3456.935 2042.965 3457.635 2043.670 ;
        RECT 3456.935 1900.000 3457.635 2042.000 ;
        RECT 3456.935 1898.330 3457.635 1899.035 ;
      LAYER met4 ;
        RECT 3458.035 1898.730 3483.000 2043.270 ;
      LAYER met4 ;
        RECT 3483.400 2042.965 3563.385 2043.670 ;
      LAYER met4 ;
        RECT 3563.785 2042.000 3588.000 2043.270 ;
      LAYER met4 ;
        RECT 3483.400 1900.000 3588.000 2042.000 ;
        RECT 3483.400 1898.330 3563.385 1899.035 ;
      LAYER met4 ;
        RECT 3563.785 1898.730 3588.000 1900.000 ;
      LAYER met4 ;
        RECT 3445.135 1896.990 3588.000 1898.330 ;
        RECT 3444.505 1863.160 3588.000 1896.990 ;
        RECT 3439.745 1861.640 3588.000 1863.160 ;
        RECT 3439.745 1847.455 3440.725 1861.640 ;
        RECT 3436.465 1845.935 3440.725 1847.455 ;
        RECT 198.365 1635.330 199.465 1635.970 ;
        RECT 152.665 1603.690 199.465 1635.330 ;
        RECT 152.035 1560.010 199.465 1603.690 ;
        RECT 3388.535 1632.310 3435.965 1675.990 ;
        RECT 3388.535 1600.670 3435.335 1632.310 ;
        RECT 3388.535 1600.030 3389.635 1600.670 ;
        RECT 147.275 1393.545 151.535 1395.065 ;
        RECT 147.275 1379.360 148.255 1393.545 ;
        RECT 0.000 1377.840 148.255 1379.360 ;
        RECT 0.000 1344.010 143.495 1377.840 ;
        RECT 0.000 1342.670 142.865 1344.010 ;
      LAYER met4 ;
        RECT 0.000 1341.000 24.215 1342.270 ;
      LAYER met4 ;
        RECT 24.615 1341.965 104.600 1342.670 ;
        RECT 0.000 1205.000 104.600 1341.000 ;
      LAYER met4 ;
        RECT 0.000 1203.730 24.215 1205.000 ;
      LAYER met4 ;
        RECT 24.615 1203.330 104.600 1203.970 ;
      LAYER met4 ;
        RECT 105.000 1203.730 129.965 1342.270 ;
      LAYER met4 ;
        RECT 130.365 1341.965 131.065 1342.670 ;
        RECT 130.365 1205.000 131.065 1341.000 ;
        RECT 130.365 1203.330 131.065 1203.970 ;
      LAYER met4 ;
        RECT 131.465 1203.730 135.915 1342.270 ;
      LAYER met4 ;
        RECT 136.315 1341.965 136.915 1342.670 ;
        RECT 136.315 1205.000 136.915 1341.000 ;
        RECT 136.315 1203.330 136.915 1203.970 ;
      LAYER met4 ;
        RECT 137.315 1203.730 141.765 1342.270 ;
      LAYER met4 ;
        RECT 142.165 1341.965 142.865 1342.670 ;
        RECT 142.165 1205.000 142.865 1341.000 ;
        RECT 142.165 1203.330 142.865 1203.970 ;
        RECT 0.000 1171.690 142.865 1203.330 ;
      LAYER met4 ;
        RECT 143.265 1172.090 143.595 1343.610 ;
      LAYER met4 ;
        RECT 0.000 1163.360 143.495 1171.690 ;
      LAYER met4 ;
        RECT 143.895 1163.760 146.875 1377.440 ;
      LAYER met4 ;
        RECT 147.275 1342.670 148.255 1377.840 ;
      LAYER met4 ;
        RECT 147.175 1341.000 148.355 1342.270 ;
      LAYER met4 ;
        RECT 147.175 1205.000 148.355 1341.000 ;
      LAYER met4 ;
        RECT 147.175 1203.730 148.355 1205.000 ;
      LAYER met4 ;
        RECT 147.275 1179.065 148.255 1203.330 ;
      LAYER met4 ;
        RECT 148.655 1179.465 151.635 1393.145 ;
        RECT 151.935 1388.090 152.265 1559.610 ;
      LAYER met4 ;
        RECT 152.665 1558.670 199.465 1560.010 ;
        RECT 152.665 1557.965 153.365 1558.670 ;
        RECT 152.665 1419.330 153.365 1419.970 ;
      LAYER met4 ;
        RECT 153.765 1419.730 158.415 1558.270 ;
      LAYER met4 ;
        RECT 158.815 1557.965 159.415 1558.670 ;
        RECT 158.815 1419.330 159.415 1419.970 ;
      LAYER met4 ;
        RECT 159.815 1419.730 163.265 1558.270 ;
      LAYER met4 ;
        RECT 163.665 1557.965 164.265 1558.670 ;
        RECT 163.665 1419.330 164.265 1419.970 ;
      LAYER met4 ;
        RECT 164.665 1419.730 168.115 1558.270 ;
      LAYER met4 ;
        RECT 168.515 1557.965 169.115 1558.670 ;
        RECT 168.515 1419.330 169.115 1419.970 ;
      LAYER met4 ;
        RECT 169.515 1419.730 174.165 1558.270 ;
      LAYER met4 ;
        RECT 174.565 1557.965 175.165 1558.670 ;
        RECT 180.615 1558.365 186.065 1558.670 ;
        RECT 174.565 1419.330 175.165 1419.970 ;
      LAYER met4 ;
        RECT 175.565 1419.730 180.215 1558.270 ;
      LAYER met4 ;
        RECT 180.615 1557.965 181.215 1558.365 ;
        RECT 185.465 1557.965 186.065 1558.365 ;
      LAYER met4 ;
        RECT 181.615 1419.970 185.065 1557.965 ;
      LAYER met4 ;
        RECT 180.615 1419.570 181.215 1419.970 ;
        RECT 185.465 1419.570 186.065 1419.970 ;
      LAYER met4 ;
        RECT 186.465 1419.730 191.115 1558.270 ;
      LAYER met4 ;
        RECT 191.515 1557.965 192.115 1558.670 ;
        RECT 180.615 1419.330 186.065 1419.570 ;
        RECT 191.515 1419.330 192.115 1419.970 ;
      LAYER met4 ;
        RECT 192.515 1419.730 197.965 1558.270 ;
      LAYER met4 ;
        RECT 198.365 1557.965 199.465 1558.670 ;
        RECT 3388.535 1456.330 3389.635 1457.035 ;
      LAYER met4 ;
        RECT 3390.035 1456.730 3395.485 1600.270 ;
      LAYER met4 ;
        RECT 3395.885 1600.030 3396.485 1600.670 ;
        RECT 3401.935 1600.430 3407.385 1600.670 ;
        RECT 3395.885 1456.330 3396.485 1457.035 ;
      LAYER met4 ;
        RECT 3396.885 1456.730 3401.535 1600.270 ;
      LAYER met4 ;
        RECT 3401.935 1600.030 3402.535 1600.430 ;
        RECT 3406.785 1600.030 3407.385 1600.430 ;
      LAYER met4 ;
        RECT 3402.935 1457.035 3406.385 1600.030 ;
      LAYER met4 ;
        RECT 3401.935 1456.635 3402.535 1457.035 ;
        RECT 3406.785 1456.635 3407.385 1457.035 ;
      LAYER met4 ;
        RECT 3407.785 1456.730 3412.435 1600.270 ;
      LAYER met4 ;
        RECT 3412.835 1600.030 3413.435 1600.670 ;
        RECT 3401.935 1456.330 3407.385 1456.635 ;
        RECT 3412.835 1456.330 3413.435 1457.035 ;
      LAYER met4 ;
        RECT 3413.835 1456.730 3418.485 1600.270 ;
      LAYER met4 ;
        RECT 3418.885 1600.030 3419.485 1600.670 ;
        RECT 3418.885 1456.330 3419.485 1457.035 ;
      LAYER met4 ;
        RECT 3419.885 1456.730 3423.335 1600.270 ;
      LAYER met4 ;
        RECT 3423.735 1600.030 3424.335 1600.670 ;
        RECT 3423.735 1456.330 3424.335 1457.035 ;
      LAYER met4 ;
        RECT 3424.735 1456.730 3428.185 1600.270 ;
      LAYER met4 ;
        RECT 3428.585 1600.030 3429.185 1600.670 ;
        RECT 3428.585 1456.330 3429.185 1457.035 ;
      LAYER met4 ;
        RECT 3429.585 1456.730 3434.235 1600.270 ;
      LAYER met4 ;
        RECT 3434.635 1600.030 3435.335 1600.670 ;
        RECT 3434.635 1456.330 3435.335 1457.035 ;
        RECT 3388.535 1454.990 3435.335 1456.330 ;
      LAYER met4 ;
        RECT 3435.735 1455.390 3436.065 1631.910 ;
        RECT 3436.365 1626.855 3439.345 1845.535 ;
      LAYER met4 ;
        RECT 3439.745 1821.670 3440.725 1845.935 ;
      LAYER met4 ;
        RECT 3439.645 1820.000 3440.825 1821.270 ;
      LAYER met4 ;
        RECT 3439.645 1679.000 3440.825 1820.000 ;
      LAYER met4 ;
        RECT 3439.645 1677.730 3440.825 1679.000 ;
      LAYER met4 ;
        RECT 3439.745 1642.160 3440.725 1677.330 ;
      LAYER met4 ;
        RECT 3441.125 1642.560 3444.105 1861.240 ;
      LAYER met4 ;
        RECT 3444.505 1853.310 3588.000 1861.640 ;
      LAYER met4 ;
        RECT 3444.405 1676.390 3444.735 1852.910 ;
      LAYER met4 ;
        RECT 3445.135 1821.670 3588.000 1853.310 ;
        RECT 3445.135 1821.030 3445.835 1821.670 ;
        RECT 3445.135 1679.000 3445.835 1820.000 ;
        RECT 3445.135 1677.330 3445.835 1678.035 ;
      LAYER met4 ;
        RECT 3446.235 1677.730 3450.685 1821.270 ;
      LAYER met4 ;
        RECT 3451.085 1821.030 3451.685 1821.670 ;
        RECT 3451.085 1679.000 3451.685 1820.000 ;
        RECT 3451.085 1677.330 3451.685 1678.035 ;
      LAYER met4 ;
        RECT 3452.085 1677.730 3456.535 1821.270 ;
      LAYER met4 ;
        RECT 3456.935 1821.030 3457.635 1821.670 ;
        RECT 3456.935 1679.000 3457.635 1820.000 ;
        RECT 3456.935 1677.330 3457.635 1678.035 ;
      LAYER met4 ;
        RECT 3458.035 1677.730 3483.000 1821.270 ;
      LAYER met4 ;
        RECT 3483.400 1821.030 3563.385 1821.670 ;
      LAYER met4 ;
        RECT 3563.785 1820.000 3588.000 1821.270 ;
      LAYER met4 ;
        RECT 3483.400 1679.000 3588.000 1820.000 ;
        RECT 3483.400 1677.330 3563.385 1678.035 ;
      LAYER met4 ;
        RECT 3563.785 1677.730 3588.000 1679.000 ;
      LAYER met4 ;
        RECT 3445.135 1675.990 3588.000 1677.330 ;
        RECT 3444.505 1642.160 3588.000 1675.990 ;
        RECT 3439.745 1640.640 3588.000 1642.160 ;
        RECT 3439.745 1626.455 3440.725 1640.640 ;
        RECT 3436.465 1624.935 3440.725 1626.455 ;
        RECT 198.365 1419.330 199.465 1419.970 ;
        RECT 152.665 1387.690 199.465 1419.330 ;
        RECT 152.035 1344.010 199.465 1387.690 ;
        RECT 3388.535 1411.310 3435.965 1454.990 ;
        RECT 3388.535 1379.670 3435.335 1411.310 ;
        RECT 3388.535 1379.030 3389.635 1379.670 ;
        RECT 147.275 1177.545 151.535 1179.065 ;
        RECT 147.275 1163.360 148.255 1177.545 ;
        RECT 0.000 1161.840 148.255 1163.360 ;
        RECT 0.000 1128.010 143.495 1161.840 ;
        RECT 0.000 1126.670 142.865 1128.010 ;
      LAYER met4 ;
        RECT 0.000 1125.000 24.215 1126.270 ;
      LAYER met4 ;
        RECT 24.615 1125.965 104.600 1126.670 ;
        RECT 0.000 989.000 104.600 1125.000 ;
      LAYER met4 ;
        RECT 0.000 987.730 24.215 989.000 ;
      LAYER met4 ;
        RECT 24.615 987.330 104.600 987.970 ;
      LAYER met4 ;
        RECT 105.000 987.730 129.965 1126.270 ;
      LAYER met4 ;
        RECT 130.365 1125.965 131.065 1126.670 ;
        RECT 130.365 989.000 131.065 1125.000 ;
        RECT 130.365 987.330 131.065 987.970 ;
      LAYER met4 ;
        RECT 131.465 987.730 135.915 1126.270 ;
      LAYER met4 ;
        RECT 136.315 1125.965 136.915 1126.670 ;
        RECT 136.315 989.000 136.915 1125.000 ;
        RECT 136.315 987.330 136.915 987.970 ;
      LAYER met4 ;
        RECT 137.315 987.730 141.765 1126.270 ;
      LAYER met4 ;
        RECT 142.165 1125.965 142.865 1126.670 ;
        RECT 142.165 989.000 142.865 1125.000 ;
        RECT 142.165 987.330 142.865 987.970 ;
        RECT 0.000 955.690 142.865 987.330 ;
      LAYER met4 ;
        RECT 143.265 956.090 143.595 1127.610 ;
      LAYER met4 ;
        RECT 0.000 947.360 143.495 955.690 ;
      LAYER met4 ;
        RECT 143.895 947.760 146.875 1161.440 ;
      LAYER met4 ;
        RECT 147.275 1126.670 148.255 1161.840 ;
      LAYER met4 ;
        RECT 147.175 1125.000 148.355 1126.270 ;
      LAYER met4 ;
        RECT 147.175 989.000 148.355 1125.000 ;
      LAYER met4 ;
        RECT 147.175 987.730 148.355 989.000 ;
      LAYER met4 ;
        RECT 147.275 963.065 148.255 987.330 ;
      LAYER met4 ;
        RECT 148.655 963.465 151.635 1177.145 ;
        RECT 151.935 1172.090 152.265 1343.610 ;
      LAYER met4 ;
        RECT 152.665 1342.670 199.465 1344.010 ;
        RECT 152.665 1341.965 153.365 1342.670 ;
        RECT 152.665 1203.330 153.365 1203.970 ;
      LAYER met4 ;
        RECT 153.765 1203.730 158.415 1342.270 ;
      LAYER met4 ;
        RECT 158.815 1341.965 159.415 1342.670 ;
        RECT 158.815 1203.330 159.415 1203.970 ;
      LAYER met4 ;
        RECT 159.815 1203.730 163.265 1342.270 ;
      LAYER met4 ;
        RECT 163.665 1341.965 164.265 1342.670 ;
        RECT 163.665 1203.330 164.265 1203.970 ;
      LAYER met4 ;
        RECT 164.665 1203.730 168.115 1342.270 ;
      LAYER met4 ;
        RECT 168.515 1341.965 169.115 1342.670 ;
        RECT 168.515 1203.330 169.115 1203.970 ;
      LAYER met4 ;
        RECT 169.515 1203.730 174.165 1342.270 ;
      LAYER met4 ;
        RECT 174.565 1341.965 175.165 1342.670 ;
        RECT 180.615 1342.365 186.065 1342.670 ;
        RECT 174.565 1203.330 175.165 1203.970 ;
      LAYER met4 ;
        RECT 175.565 1203.730 180.215 1342.270 ;
      LAYER met4 ;
        RECT 180.615 1341.965 181.215 1342.365 ;
        RECT 185.465 1341.965 186.065 1342.365 ;
      LAYER met4 ;
        RECT 181.615 1203.970 185.065 1341.965 ;
      LAYER met4 ;
        RECT 180.615 1203.570 181.215 1203.970 ;
        RECT 185.465 1203.570 186.065 1203.970 ;
      LAYER met4 ;
        RECT 186.465 1203.730 191.115 1342.270 ;
      LAYER met4 ;
        RECT 191.515 1341.965 192.115 1342.670 ;
        RECT 180.615 1203.330 186.065 1203.570 ;
        RECT 191.515 1203.330 192.115 1203.970 ;
      LAYER met4 ;
        RECT 192.515 1203.730 197.965 1342.270 ;
      LAYER met4 ;
        RECT 198.365 1341.965 199.465 1342.670 ;
        RECT 3388.535 1234.330 3389.635 1235.035 ;
      LAYER met4 ;
        RECT 3390.035 1234.730 3395.485 1379.270 ;
      LAYER met4 ;
        RECT 3395.885 1379.030 3396.485 1379.670 ;
        RECT 3401.935 1379.430 3407.385 1379.670 ;
        RECT 3395.885 1234.330 3396.485 1235.035 ;
      LAYER met4 ;
        RECT 3396.885 1234.730 3401.535 1379.270 ;
      LAYER met4 ;
        RECT 3401.935 1379.030 3402.535 1379.430 ;
        RECT 3406.785 1379.030 3407.385 1379.430 ;
      LAYER met4 ;
        RECT 3402.935 1235.035 3406.385 1379.030 ;
      LAYER met4 ;
        RECT 3401.935 1234.635 3402.535 1235.035 ;
        RECT 3406.785 1234.635 3407.385 1235.035 ;
      LAYER met4 ;
        RECT 3407.785 1234.730 3412.435 1379.270 ;
      LAYER met4 ;
        RECT 3412.835 1379.030 3413.435 1379.670 ;
        RECT 3401.935 1234.330 3407.385 1234.635 ;
        RECT 3412.835 1234.330 3413.435 1235.035 ;
      LAYER met4 ;
        RECT 3413.835 1234.730 3418.485 1379.270 ;
      LAYER met4 ;
        RECT 3418.885 1379.030 3419.485 1379.670 ;
        RECT 3418.885 1234.330 3419.485 1235.035 ;
      LAYER met4 ;
        RECT 3419.885 1234.730 3423.335 1379.270 ;
      LAYER met4 ;
        RECT 3423.735 1379.030 3424.335 1379.670 ;
        RECT 3423.735 1234.330 3424.335 1235.035 ;
      LAYER met4 ;
        RECT 3424.735 1234.730 3428.185 1379.270 ;
      LAYER met4 ;
        RECT 3428.585 1379.030 3429.185 1379.670 ;
        RECT 3428.585 1234.330 3429.185 1235.035 ;
      LAYER met4 ;
        RECT 3429.585 1234.730 3434.235 1379.270 ;
      LAYER met4 ;
        RECT 3434.635 1379.030 3435.335 1379.670 ;
        RECT 3434.635 1234.330 3435.335 1235.035 ;
        RECT 3388.535 1232.990 3435.335 1234.330 ;
      LAYER met4 ;
        RECT 3435.735 1233.390 3436.065 1410.910 ;
        RECT 3436.365 1405.855 3439.345 1624.535 ;
      LAYER met4 ;
        RECT 3439.745 1600.670 3440.725 1624.935 ;
      LAYER met4 ;
        RECT 3439.645 1599.000 3440.825 1600.270 ;
      LAYER met4 ;
        RECT 3439.645 1458.000 3440.825 1599.000 ;
      LAYER met4 ;
        RECT 3439.645 1456.730 3440.825 1458.000 ;
      LAYER met4 ;
        RECT 3439.745 1421.160 3440.725 1456.330 ;
      LAYER met4 ;
        RECT 3441.125 1421.560 3444.105 1640.240 ;
      LAYER met4 ;
        RECT 3444.505 1632.310 3588.000 1640.640 ;
      LAYER met4 ;
        RECT 3444.405 1455.390 3444.735 1631.910 ;
      LAYER met4 ;
        RECT 3445.135 1600.670 3588.000 1632.310 ;
        RECT 3445.135 1600.030 3445.835 1600.670 ;
        RECT 3445.135 1458.000 3445.835 1599.000 ;
        RECT 3445.135 1456.330 3445.835 1457.035 ;
      LAYER met4 ;
        RECT 3446.235 1456.730 3450.685 1600.270 ;
      LAYER met4 ;
        RECT 3451.085 1600.030 3451.685 1600.670 ;
        RECT 3451.085 1458.000 3451.685 1599.000 ;
        RECT 3451.085 1456.330 3451.685 1457.035 ;
      LAYER met4 ;
        RECT 3452.085 1456.730 3456.535 1600.270 ;
      LAYER met4 ;
        RECT 3456.935 1600.030 3457.635 1600.670 ;
        RECT 3456.935 1458.000 3457.635 1599.000 ;
        RECT 3456.935 1456.330 3457.635 1457.035 ;
      LAYER met4 ;
        RECT 3458.035 1456.730 3483.000 1600.270 ;
      LAYER met4 ;
        RECT 3483.400 1600.030 3563.385 1600.670 ;
      LAYER met4 ;
        RECT 3563.785 1599.000 3588.000 1600.270 ;
      LAYER met4 ;
        RECT 3483.400 1458.000 3588.000 1599.000 ;
        RECT 3483.400 1456.330 3563.385 1457.035 ;
      LAYER met4 ;
        RECT 3563.785 1456.730 3588.000 1458.000 ;
      LAYER met4 ;
        RECT 3445.135 1454.990 3588.000 1456.330 ;
        RECT 3444.505 1421.160 3588.000 1454.990 ;
        RECT 3439.745 1419.640 3588.000 1421.160 ;
        RECT 3439.745 1405.455 3440.725 1419.640 ;
        RECT 3436.465 1403.935 3440.725 1405.455 ;
        RECT 198.365 1203.330 199.465 1203.970 ;
        RECT 152.665 1171.690 199.465 1203.330 ;
        RECT 152.035 1128.010 199.465 1171.690 ;
        RECT 3388.535 1189.310 3435.965 1232.990 ;
        RECT 3388.535 1157.670 3435.335 1189.310 ;
        RECT 3388.535 1157.030 3389.635 1157.670 ;
        RECT 147.275 961.545 151.535 963.065 ;
        RECT 147.275 947.360 148.255 961.545 ;
        RECT 0.000 945.840 148.255 947.360 ;
        RECT 0.000 912.010 143.495 945.840 ;
        RECT 0.000 910.670 142.865 912.010 ;
      LAYER met4 ;
        RECT 0.000 909.000 24.215 910.270 ;
      LAYER met4 ;
        RECT 24.615 909.965 104.600 910.670 ;
        RECT 0.000 767.000 104.600 909.000 ;
        RECT 0.000 762.000 24.215 767.000 ;
        RECT 0.000 626.000 104.600 762.000 ;
      LAYER met4 ;
        RECT 0.000 624.730 24.215 626.000 ;
      LAYER met4 ;
        RECT 24.615 624.330 104.600 625.035 ;
      LAYER met4 ;
        RECT 105.000 624.730 129.965 910.270 ;
      LAYER met4 ;
        RECT 130.365 909.965 131.065 910.670 ;
        RECT 130.365 767.000 131.065 909.000 ;
        RECT 130.365 626.000 131.065 762.000 ;
        RECT 130.365 624.330 131.065 625.035 ;
      LAYER met4 ;
        RECT 131.465 624.730 135.915 910.270 ;
      LAYER met4 ;
        RECT 136.315 909.965 136.915 910.670 ;
        RECT 136.315 767.000 136.915 909.000 ;
        RECT 136.315 626.000 136.915 762.000 ;
        RECT 136.315 624.330 136.915 625.035 ;
      LAYER met4 ;
        RECT 137.315 624.730 141.765 910.270 ;
      LAYER met4 ;
        RECT 142.165 909.965 142.865 910.670 ;
        RECT 142.165 767.000 142.865 909.000 ;
      LAYER met4 ;
        RECT 143.265 767.000 143.595 911.610 ;
      LAYER met4 ;
        RECT 142.165 626.000 142.865 762.000 ;
        RECT 142.165 624.330 142.865 625.035 ;
        RECT 0.000 552.670 142.865 624.330 ;
      LAYER met4 ;
        RECT 0.000 551.000 24.215 552.270 ;
      LAYER met4 ;
        RECT 24.615 551.965 104.600 552.670 ;
        RECT 0.000 415.000 104.600 551.000 ;
      LAYER met4 ;
        RECT 0.000 413.730 24.215 415.000 ;
      LAYER met4 ;
        RECT 24.615 413.330 104.600 415.000 ;
      LAYER met4 ;
        RECT 105.000 413.730 129.965 552.270 ;
      LAYER met4 ;
        RECT 130.365 551.965 131.065 552.670 ;
        RECT 130.365 413.330 131.065 551.000 ;
      LAYER met4 ;
        RECT 131.465 413.730 135.915 552.270 ;
      LAYER met4 ;
        RECT 136.315 551.965 136.915 552.670 ;
        RECT 136.315 413.330 136.915 551.000 ;
      LAYER met4 ;
        RECT 137.315 413.730 141.765 552.270 ;
      LAYER met4 ;
        RECT 142.165 551.965 142.865 552.670 ;
        RECT 142.165 413.330 142.865 551.000 ;
        RECT 0.000 341.670 142.865 413.330 ;
      LAYER met4 ;
        RECT 0.000 340.000 24.215 341.270 ;
      LAYER met4 ;
        RECT 24.615 340.965 104.600 341.670 ;
        RECT 0.000 204.000 104.600 340.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 341.270 ;
      LAYER met4 ;
        RECT 130.365 340.965 131.065 341.670 ;
        RECT 130.365 204.000 131.065 340.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 341.270 ;
      LAYER met4 ;
        RECT 136.315 340.965 136.915 341.670 ;
        RECT 136.315 204.000 136.915 340.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 341.270 ;
      LAYER met4 ;
        RECT 142.165 340.965 142.865 341.670 ;
        RECT 142.165 204.000 142.865 340.000 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 762.000 ;
        RECT 143.895 177.090 146.875 945.440 ;
      LAYER met4 ;
        RECT 147.275 910.670 148.255 945.840 ;
      LAYER met4 ;
        RECT 147.175 909.000 148.355 910.270 ;
      LAYER met4 ;
        RECT 147.175 767.000 148.355 909.000 ;
        RECT 147.175 626.000 148.355 762.000 ;
      LAYER met4 ;
        RECT 147.175 624.730 148.355 626.000 ;
      LAYER met4 ;
        RECT 147.275 552.670 148.255 624.330 ;
      LAYER met4 ;
        RECT 147.175 551.000 148.355 552.270 ;
      LAYER met4 ;
        RECT 147.175 415.000 148.355 551.000 ;
      LAYER met4 ;
        RECT 147.175 413.730 148.355 415.000 ;
      LAYER met4 ;
        RECT 147.275 341.670 148.255 413.330 ;
      LAYER met4 ;
        RECT 147.175 340.000 148.355 341.270 ;
      LAYER met4 ;
        RECT 147.175 204.000 148.355 340.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 961.145 ;
        RECT 151.935 956.090 152.265 1127.610 ;
      LAYER met4 ;
        RECT 152.665 1126.670 199.465 1128.010 ;
        RECT 152.665 1125.965 153.365 1126.670 ;
        RECT 152.665 987.330 153.365 987.970 ;
      LAYER met4 ;
        RECT 153.765 987.730 158.415 1126.270 ;
      LAYER met4 ;
        RECT 158.815 1125.965 159.415 1126.670 ;
        RECT 158.815 987.330 159.415 987.970 ;
      LAYER met4 ;
        RECT 159.815 987.730 163.265 1126.270 ;
      LAYER met4 ;
        RECT 163.665 1125.965 164.265 1126.670 ;
        RECT 163.665 987.330 164.265 987.970 ;
      LAYER met4 ;
        RECT 164.665 987.730 168.115 1126.270 ;
      LAYER met4 ;
        RECT 168.515 1125.965 169.115 1126.670 ;
        RECT 168.515 987.330 169.115 987.970 ;
      LAYER met4 ;
        RECT 169.515 987.730 174.165 1126.270 ;
      LAYER met4 ;
        RECT 174.565 1125.965 175.165 1126.670 ;
        RECT 180.615 1126.365 186.065 1126.670 ;
        RECT 174.565 987.330 175.165 987.970 ;
      LAYER met4 ;
        RECT 175.565 987.730 180.215 1126.270 ;
      LAYER met4 ;
        RECT 180.615 1125.965 181.215 1126.365 ;
        RECT 185.465 1125.965 186.065 1126.365 ;
      LAYER met4 ;
        RECT 181.615 987.970 185.065 1125.965 ;
      LAYER met4 ;
        RECT 180.615 987.570 181.215 987.970 ;
        RECT 185.465 987.570 186.065 987.970 ;
      LAYER met4 ;
        RECT 186.465 987.730 191.115 1126.270 ;
      LAYER met4 ;
        RECT 191.515 1125.965 192.115 1126.670 ;
        RECT 180.615 987.330 186.065 987.570 ;
        RECT 191.515 987.330 192.115 987.970 ;
      LAYER met4 ;
        RECT 192.515 987.730 197.965 1126.270 ;
      LAYER met4 ;
        RECT 198.365 1125.965 199.465 1126.670 ;
        RECT 3388.535 1013.330 3389.635 1014.035 ;
      LAYER met4 ;
        RECT 3390.035 1013.730 3395.485 1157.270 ;
      LAYER met4 ;
        RECT 3395.885 1157.030 3396.485 1157.670 ;
        RECT 3401.935 1157.430 3407.385 1157.670 ;
        RECT 3395.885 1013.330 3396.485 1014.035 ;
      LAYER met4 ;
        RECT 3396.885 1013.730 3401.535 1157.270 ;
      LAYER met4 ;
        RECT 3401.935 1157.030 3402.535 1157.430 ;
        RECT 3406.785 1157.030 3407.385 1157.430 ;
      LAYER met4 ;
        RECT 3402.935 1014.035 3406.385 1157.030 ;
      LAYER met4 ;
        RECT 3401.935 1013.635 3402.535 1014.035 ;
        RECT 3406.785 1013.635 3407.385 1014.035 ;
      LAYER met4 ;
        RECT 3407.785 1013.730 3412.435 1157.270 ;
      LAYER met4 ;
        RECT 3412.835 1157.030 3413.435 1157.670 ;
        RECT 3401.935 1013.330 3407.385 1013.635 ;
        RECT 3412.835 1013.330 3413.435 1014.035 ;
      LAYER met4 ;
        RECT 3413.835 1013.730 3418.485 1157.270 ;
      LAYER met4 ;
        RECT 3418.885 1157.030 3419.485 1157.670 ;
        RECT 3418.885 1013.330 3419.485 1014.035 ;
      LAYER met4 ;
        RECT 3419.885 1013.730 3423.335 1157.270 ;
      LAYER met4 ;
        RECT 3423.735 1157.030 3424.335 1157.670 ;
        RECT 3423.735 1013.330 3424.335 1014.035 ;
      LAYER met4 ;
        RECT 3424.735 1013.730 3428.185 1157.270 ;
      LAYER met4 ;
        RECT 3428.585 1157.030 3429.185 1157.670 ;
        RECT 3428.585 1013.330 3429.185 1014.035 ;
      LAYER met4 ;
        RECT 3429.585 1013.730 3434.235 1157.270 ;
      LAYER met4 ;
        RECT 3434.635 1157.030 3435.335 1157.670 ;
        RECT 3434.635 1013.330 3435.335 1014.035 ;
        RECT 3388.535 1011.990 3435.335 1013.330 ;
      LAYER met4 ;
        RECT 3435.735 1012.390 3436.065 1188.910 ;
        RECT 3436.365 1183.855 3439.345 1403.535 ;
      LAYER met4 ;
        RECT 3439.745 1379.670 3440.725 1403.935 ;
      LAYER met4 ;
        RECT 3439.645 1378.000 3440.825 1379.270 ;
      LAYER met4 ;
        RECT 3439.645 1236.000 3440.825 1378.000 ;
      LAYER met4 ;
        RECT 3439.645 1234.730 3440.825 1236.000 ;
      LAYER met4 ;
        RECT 3439.745 1199.160 3440.725 1234.330 ;
      LAYER met4 ;
        RECT 3441.125 1199.560 3444.105 1419.240 ;
      LAYER met4 ;
        RECT 3444.505 1411.310 3588.000 1419.640 ;
      LAYER met4 ;
        RECT 3444.405 1233.390 3444.735 1410.910 ;
      LAYER met4 ;
        RECT 3445.135 1379.670 3588.000 1411.310 ;
        RECT 3445.135 1379.030 3445.835 1379.670 ;
        RECT 3445.135 1236.000 3445.835 1378.000 ;
        RECT 3445.135 1234.330 3445.835 1235.035 ;
      LAYER met4 ;
        RECT 3446.235 1234.730 3450.685 1379.270 ;
      LAYER met4 ;
        RECT 3451.085 1379.030 3451.685 1379.670 ;
        RECT 3451.085 1236.000 3451.685 1378.000 ;
        RECT 3451.085 1234.330 3451.685 1235.035 ;
      LAYER met4 ;
        RECT 3452.085 1234.730 3456.535 1379.270 ;
      LAYER met4 ;
        RECT 3456.935 1379.030 3457.635 1379.670 ;
        RECT 3456.935 1236.000 3457.635 1378.000 ;
        RECT 3456.935 1234.330 3457.635 1235.035 ;
      LAYER met4 ;
        RECT 3458.035 1234.730 3483.000 1379.270 ;
      LAYER met4 ;
        RECT 3483.400 1379.030 3563.385 1379.670 ;
      LAYER met4 ;
        RECT 3563.785 1378.000 3588.000 1379.270 ;
      LAYER met4 ;
        RECT 3483.400 1236.000 3588.000 1378.000 ;
        RECT 3483.400 1234.330 3563.385 1235.035 ;
      LAYER met4 ;
        RECT 3563.785 1234.730 3588.000 1236.000 ;
      LAYER met4 ;
        RECT 3445.135 1232.990 3588.000 1234.330 ;
        RECT 3444.505 1199.160 3588.000 1232.990 ;
        RECT 3439.745 1197.640 3588.000 1199.160 ;
        RECT 3439.745 1183.455 3440.725 1197.640 ;
        RECT 3436.465 1181.935 3440.725 1183.455 ;
        RECT 198.365 987.330 199.465 987.970 ;
        RECT 152.665 955.690 199.465 987.330 ;
        RECT 152.035 912.010 199.465 955.690 ;
        RECT 3388.535 968.310 3435.965 1011.990 ;
        RECT 3388.535 936.670 3435.335 968.310 ;
        RECT 3388.535 936.030 3389.635 936.670 ;
      LAYER met4 ;
        RECT 151.935 767.000 152.265 911.610 ;
      LAYER met4 ;
        RECT 152.665 910.670 199.465 912.010 ;
        RECT 152.665 909.965 153.365 910.670 ;
      LAYER met4 ;
        RECT 153.765 772.000 158.415 910.270 ;
      LAYER met4 ;
        RECT 158.815 909.965 159.415 910.670 ;
      LAYER met4 ;
        RECT 159.815 767.000 163.265 910.270 ;
      LAYER met4 ;
        RECT 163.665 909.965 164.265 910.670 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 762.000 ;
      LAYER met4 ;
        RECT 152.665 624.330 153.365 625.035 ;
      LAYER met4 ;
        RECT 153.765 624.730 158.415 767.000 ;
      LAYER met4 ;
        RECT 158.815 624.330 159.415 625.035 ;
      LAYER met4 ;
        RECT 159.815 624.730 163.265 762.000 ;
      LAYER met4 ;
        RECT 163.665 624.330 164.265 625.035 ;
      LAYER met4 ;
        RECT 164.665 624.730 168.115 910.270 ;
      LAYER met4 ;
        RECT 168.515 909.965 169.115 910.670 ;
        RECT 168.515 624.330 169.115 625.035 ;
      LAYER met4 ;
        RECT 169.515 624.730 174.165 910.270 ;
      LAYER met4 ;
        RECT 174.565 909.965 175.165 910.670 ;
        RECT 180.615 910.365 186.065 910.670 ;
        RECT 174.565 624.330 175.165 625.035 ;
      LAYER met4 ;
        RECT 175.565 624.730 180.215 910.270 ;
      LAYER met4 ;
        RECT 180.615 909.965 181.215 910.365 ;
        RECT 185.465 909.965 186.065 910.365 ;
      LAYER met4 ;
        RECT 181.615 767.000 185.065 909.965 ;
        RECT 186.465 772.000 191.115 910.270 ;
      LAYER met4 ;
        RECT 191.515 909.965 192.115 910.670 ;
      LAYER met4 ;
        RECT 181.615 625.035 185.065 762.000 ;
      LAYER met4 ;
        RECT 180.615 624.635 181.215 625.035 ;
        RECT 185.465 624.635 186.065 625.035 ;
      LAYER met4 ;
        RECT 186.465 624.730 191.115 767.000 ;
      LAYER met4 ;
        RECT 180.615 624.330 186.065 624.635 ;
        RECT 191.515 624.330 192.115 625.035 ;
      LAYER met4 ;
        RECT 192.515 624.730 197.965 910.270 ;
      LAYER met4 ;
        RECT 198.365 909.965 199.465 910.670 ;
        RECT 3388.535 792.330 3389.635 793.035 ;
      LAYER met4 ;
        RECT 3390.035 792.730 3395.485 936.270 ;
      LAYER met4 ;
        RECT 3395.885 936.030 3396.485 936.670 ;
        RECT 3401.935 936.430 3407.385 936.670 ;
        RECT 3395.885 792.330 3396.485 793.035 ;
      LAYER met4 ;
        RECT 3396.885 792.730 3401.535 936.270 ;
      LAYER met4 ;
        RECT 3401.935 936.030 3402.535 936.430 ;
        RECT 3406.785 936.030 3407.385 936.430 ;
      LAYER met4 ;
        RECT 3402.935 793.035 3406.385 936.030 ;
      LAYER met4 ;
        RECT 3401.935 792.635 3402.535 793.035 ;
        RECT 3406.785 792.635 3407.385 793.035 ;
      LAYER met4 ;
        RECT 3407.785 792.730 3412.435 936.270 ;
      LAYER met4 ;
        RECT 3412.835 936.030 3413.435 936.670 ;
        RECT 3401.935 792.330 3407.385 792.635 ;
        RECT 3412.835 792.330 3413.435 793.035 ;
      LAYER met4 ;
        RECT 3413.835 792.730 3418.485 936.270 ;
      LAYER met4 ;
        RECT 3418.885 936.030 3419.485 936.670 ;
        RECT 3418.885 792.330 3419.485 793.035 ;
      LAYER met4 ;
        RECT 3419.885 792.730 3423.335 936.270 ;
      LAYER met4 ;
        RECT 3423.735 936.030 3424.335 936.670 ;
        RECT 3423.735 792.330 3424.335 793.035 ;
      LAYER met4 ;
        RECT 3424.735 792.730 3428.185 936.270 ;
      LAYER met4 ;
        RECT 3428.585 936.030 3429.185 936.670 ;
        RECT 3428.585 792.330 3429.185 793.035 ;
      LAYER met4 ;
        RECT 3429.585 792.730 3434.235 936.270 ;
      LAYER met4 ;
        RECT 3434.635 936.030 3435.335 936.670 ;
        RECT 3434.635 792.330 3435.335 793.035 ;
        RECT 3388.535 790.990 3435.335 792.330 ;
      LAYER met4 ;
        RECT 3435.735 791.390 3436.065 967.910 ;
        RECT 3436.365 962.855 3439.345 1181.535 ;
      LAYER met4 ;
        RECT 3439.745 1157.670 3440.725 1181.935 ;
      LAYER met4 ;
        RECT 3439.645 1156.000 3440.825 1157.270 ;
      LAYER met4 ;
        RECT 3439.645 1015.000 3440.825 1156.000 ;
      LAYER met4 ;
        RECT 3439.645 1013.730 3440.825 1015.000 ;
      LAYER met4 ;
        RECT 3439.745 978.160 3440.725 1013.330 ;
      LAYER met4 ;
        RECT 3441.125 978.560 3444.105 1197.240 ;
      LAYER met4 ;
        RECT 3444.505 1189.310 3588.000 1197.640 ;
      LAYER met4 ;
        RECT 3444.405 1012.390 3444.735 1188.910 ;
      LAYER met4 ;
        RECT 3445.135 1157.670 3588.000 1189.310 ;
        RECT 3445.135 1157.030 3445.835 1157.670 ;
        RECT 3445.135 1015.000 3445.835 1156.000 ;
        RECT 3445.135 1013.330 3445.835 1014.035 ;
      LAYER met4 ;
        RECT 3446.235 1013.730 3450.685 1157.270 ;
      LAYER met4 ;
        RECT 3451.085 1157.030 3451.685 1157.670 ;
        RECT 3451.085 1015.000 3451.685 1156.000 ;
        RECT 3451.085 1013.330 3451.685 1014.035 ;
      LAYER met4 ;
        RECT 3452.085 1013.730 3456.535 1157.270 ;
      LAYER met4 ;
        RECT 3456.935 1157.030 3457.635 1157.670 ;
        RECT 3456.935 1015.000 3457.635 1156.000 ;
        RECT 3456.935 1013.330 3457.635 1014.035 ;
      LAYER met4 ;
        RECT 3458.035 1013.730 3483.000 1157.270 ;
      LAYER met4 ;
        RECT 3483.400 1157.030 3563.385 1157.670 ;
      LAYER met4 ;
        RECT 3563.785 1156.000 3588.000 1157.270 ;
      LAYER met4 ;
        RECT 3483.400 1015.000 3588.000 1156.000 ;
        RECT 3483.400 1013.330 3563.385 1014.035 ;
      LAYER met4 ;
        RECT 3563.785 1013.730 3588.000 1015.000 ;
      LAYER met4 ;
        RECT 3445.135 1011.990 3588.000 1013.330 ;
        RECT 3444.505 978.160 3588.000 1011.990 ;
        RECT 3439.745 976.640 3588.000 978.160 ;
        RECT 3439.745 962.455 3440.725 976.640 ;
        RECT 3436.465 960.935 3440.725 962.455 ;
        RECT 3388.535 747.310 3435.965 790.990 ;
        RECT 3388.535 715.670 3435.335 747.310 ;
        RECT 3388.535 715.030 3389.635 715.670 ;
        RECT 152.665 552.670 197.965 624.330 ;
        RECT 3388.535 570.330 3389.635 571.035 ;
      LAYER met4 ;
        RECT 3390.035 570.730 3395.485 715.270 ;
      LAYER met4 ;
        RECT 3395.885 715.030 3396.485 715.670 ;
        RECT 3401.935 715.430 3407.385 715.670 ;
        RECT 3395.885 570.330 3396.485 571.035 ;
      LAYER met4 ;
        RECT 3396.885 570.730 3401.535 715.270 ;
      LAYER met4 ;
        RECT 3401.935 715.030 3402.535 715.430 ;
        RECT 3406.785 715.030 3407.385 715.430 ;
      LAYER met4 ;
        RECT 3402.935 571.035 3406.385 715.030 ;
      LAYER met4 ;
        RECT 3401.935 570.635 3402.535 571.035 ;
        RECT 3406.785 570.635 3407.385 571.035 ;
      LAYER met4 ;
        RECT 3407.785 570.730 3412.435 715.270 ;
      LAYER met4 ;
        RECT 3412.835 715.030 3413.435 715.670 ;
        RECT 3401.935 570.330 3407.385 570.635 ;
        RECT 3412.835 570.330 3413.435 571.035 ;
      LAYER met4 ;
        RECT 3413.835 570.730 3418.485 715.270 ;
      LAYER met4 ;
        RECT 3418.885 715.030 3419.485 715.670 ;
        RECT 3418.885 570.330 3419.485 571.035 ;
      LAYER met4 ;
        RECT 3419.885 570.730 3423.335 715.270 ;
      LAYER met4 ;
        RECT 3423.735 715.030 3424.335 715.670 ;
        RECT 3423.735 570.330 3424.335 571.035 ;
      LAYER met4 ;
        RECT 3424.735 570.730 3428.185 715.270 ;
      LAYER met4 ;
        RECT 3428.585 715.030 3429.185 715.670 ;
        RECT 3428.585 570.330 3429.185 571.035 ;
      LAYER met4 ;
        RECT 3429.585 570.730 3434.235 715.270 ;
      LAYER met4 ;
        RECT 3434.635 715.030 3435.335 715.670 ;
        RECT 3434.635 570.330 3435.335 571.035 ;
        RECT 3388.535 568.990 3435.335 570.330 ;
      LAYER met4 ;
        RECT 3435.735 569.390 3436.065 746.910 ;
        RECT 3436.365 741.855 3439.345 960.535 ;
      LAYER met4 ;
        RECT 3439.745 936.670 3440.725 960.935 ;
      LAYER met4 ;
        RECT 3439.645 935.000 3440.825 936.270 ;
      LAYER met4 ;
        RECT 3439.645 794.000 3440.825 935.000 ;
      LAYER met4 ;
        RECT 3439.645 792.730 3440.825 794.000 ;
      LAYER met4 ;
        RECT 3439.745 757.160 3440.725 792.330 ;
      LAYER met4 ;
        RECT 3441.125 757.560 3444.105 976.240 ;
      LAYER met4 ;
        RECT 3444.505 968.310 3588.000 976.640 ;
      LAYER met4 ;
        RECT 3444.405 791.390 3444.735 967.910 ;
      LAYER met4 ;
        RECT 3445.135 936.670 3588.000 968.310 ;
        RECT 3445.135 936.030 3445.835 936.670 ;
        RECT 3445.135 794.000 3445.835 935.000 ;
        RECT 3445.135 792.330 3445.835 793.035 ;
      LAYER met4 ;
        RECT 3446.235 792.730 3450.685 936.270 ;
      LAYER met4 ;
        RECT 3451.085 936.030 3451.685 936.670 ;
        RECT 3451.085 794.000 3451.685 935.000 ;
        RECT 3451.085 792.330 3451.685 793.035 ;
      LAYER met4 ;
        RECT 3452.085 792.730 3456.535 936.270 ;
      LAYER met4 ;
        RECT 3456.935 936.030 3457.635 936.670 ;
        RECT 3456.935 794.000 3457.635 935.000 ;
        RECT 3456.935 792.330 3457.635 793.035 ;
      LAYER met4 ;
        RECT 3458.035 792.730 3483.000 936.270 ;
      LAYER met4 ;
        RECT 3483.400 936.030 3563.385 936.670 ;
      LAYER met4 ;
        RECT 3563.785 935.000 3588.000 936.270 ;
      LAYER met4 ;
        RECT 3483.400 794.000 3588.000 935.000 ;
        RECT 3483.400 792.330 3563.385 793.035 ;
      LAYER met4 ;
        RECT 3563.785 792.730 3588.000 794.000 ;
      LAYER met4 ;
        RECT 3445.135 790.990 3588.000 792.330 ;
        RECT 3444.505 757.160 3588.000 790.990 ;
        RECT 3439.745 755.640 3588.000 757.160 ;
        RECT 3439.745 741.455 3440.725 755.640 ;
        RECT 3436.465 739.935 3440.725 741.455 ;
        RECT 152.665 551.965 153.365 552.670 ;
        RECT 152.665 413.330 153.365 415.000 ;
      LAYER met4 ;
        RECT 153.765 413.730 158.415 552.270 ;
      LAYER met4 ;
        RECT 158.815 551.965 159.415 552.670 ;
        RECT 158.815 413.330 159.415 415.000 ;
      LAYER met4 ;
        RECT 159.815 413.730 163.265 552.270 ;
      LAYER met4 ;
        RECT 163.665 551.965 164.265 552.670 ;
        RECT 163.665 413.330 164.265 415.000 ;
      LAYER met4 ;
        RECT 164.665 413.730 168.115 552.270 ;
      LAYER met4 ;
        RECT 168.515 551.965 169.115 552.670 ;
        RECT 168.515 413.330 169.115 415.000 ;
      LAYER met4 ;
        RECT 169.515 413.730 174.165 552.270 ;
      LAYER met4 ;
        RECT 174.565 551.965 175.165 552.670 ;
        RECT 180.615 552.365 186.065 552.670 ;
        RECT 174.565 413.330 175.165 415.000 ;
      LAYER met4 ;
        RECT 175.565 413.730 180.215 552.270 ;
      LAYER met4 ;
        RECT 180.615 551.965 181.215 552.365 ;
        RECT 185.465 551.965 186.065 552.365 ;
        RECT 180.615 413.635 181.215 415.000 ;
      LAYER met4 ;
        RECT 181.615 414.035 185.065 551.965 ;
      LAYER met4 ;
        RECT 185.465 413.635 186.065 415.000 ;
      LAYER met4 ;
        RECT 186.465 413.730 191.115 552.270 ;
      LAYER met4 ;
        RECT 191.515 551.965 192.115 552.670 ;
        RECT 180.615 413.330 186.065 413.635 ;
        RECT 191.515 413.330 192.115 415.000 ;
      LAYER met4 ;
        RECT 192.515 413.730 197.965 552.270 ;
      LAYER met4 ;
        RECT 3388.535 525.310 3435.965 568.990 ;
        RECT 3388.535 493.670 3435.335 525.310 ;
        RECT 3388.535 493.030 3389.635 493.670 ;
        RECT 152.665 341.670 197.965 413.330 ;
        RECT 152.665 340.965 153.365 341.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 341.270 ;
      LAYER met4 ;
        RECT 158.815 340.965 159.415 341.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 341.270 ;
      LAYER met4 ;
        RECT 163.665 340.965 164.265 341.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 341.270 ;
      LAYER met4 ;
        RECT 168.515 340.965 169.115 341.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 341.270 ;
      LAYER met4 ;
        RECT 174.565 340.965 175.165 341.670 ;
        RECT 180.615 341.365 186.065 341.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 341.270 ;
      LAYER met4 ;
        RECT 180.615 340.965 181.215 341.365 ;
        RECT 185.465 340.965 186.065 341.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 340.965 ;
      LAYER met4 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
      LAYER met4 ;
        RECT 186.465 202.730 191.115 341.270 ;
      LAYER met4 ;
        RECT 191.515 340.965 192.115 341.670 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 341.270 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
        RECT 933.030 198.365 1011.035 199.465 ;
        RECT 1476.030 198.365 1554.035 199.465 ;
        RECT 1750.030 198.365 1828.035 199.465 ;
        RECT 2024.030 198.365 2102.035 199.465 ;
        RECT 2298.030 198.365 2376.035 199.465 ;
        RECT 2572.030 198.365 2650.035 199.465 ;
        RECT 3385.255 198.365 3389.635 200.000 ;
        RECT 152.665 192.115 197.250 198.365 ;
      LAYER met4 ;
        RECT 197.650 192.515 395.270 197.965 ;
      LAYER met4 ;
        RECT 395.670 192.115 467.330 197.965 ;
      LAYER met4 ;
        RECT 467.730 192.515 664.270 197.965 ;
      LAYER met4 ;
        RECT 664.670 192.115 736.330 197.965 ;
      LAYER met4 ;
        RECT 736.730 192.515 933.270 197.965 ;
      LAYER met4 ;
        RECT 933.670 192.115 1010.330 198.365 ;
      LAYER met4 ;
        RECT 1010.730 192.515 1207.270 197.965 ;
      LAYER met4 ;
        RECT 1207.670 192.115 1279.330 197.965 ;
      LAYER met4 ;
        RECT 1279.730 192.515 1476.270 197.965 ;
      LAYER met4 ;
        RECT 1476.670 192.115 1553.330 198.365 ;
      LAYER met4 ;
        RECT 1553.730 192.515 1750.270 197.965 ;
      LAYER met4 ;
        RECT 1750.670 192.115 1827.330 198.365 ;
      LAYER met4 ;
        RECT 1827.730 192.515 2024.270 197.965 ;
      LAYER met4 ;
        RECT 2024.670 192.115 2101.330 198.365 ;
      LAYER met4 ;
        RECT 2101.730 192.515 2298.270 197.965 ;
      LAYER met4 ;
        RECT 2298.670 192.115 2375.330 198.365 ;
      LAYER met4 ;
        RECT 2375.730 192.515 2572.270 197.965 ;
      LAYER met4 ;
        RECT 2572.670 192.115 2649.330 198.365 ;
      LAYER met4 ;
        RECT 2649.730 192.515 2846.270 197.965 ;
      LAYER met4 ;
        RECT 2846.670 192.115 2918.330 197.965 ;
      LAYER met4 ;
        RECT 2918.730 192.515 3115.270 197.965 ;
      LAYER met4 ;
        RECT 3115.670 192.115 3187.330 197.965 ;
      LAYER met4 ;
        RECT 3187.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 198.365 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 493.270 ;
      LAYER met4 ;
        RECT 3395.885 493.030 3396.485 493.670 ;
        RECT 3401.935 493.430 3407.385 493.670 ;
      LAYER met4 ;
        RECT 3396.885 351.000 3401.535 493.270 ;
      LAYER met4 ;
        RECT 3401.935 493.030 3402.535 493.430 ;
        RECT 3406.785 493.030 3407.385 493.430 ;
      LAYER met4 ;
        RECT 3402.935 346.000 3406.385 493.030 ;
      LAYER met4 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 346.000 ;
      LAYER met4 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 341.000 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 493.270 ;
      LAYER met4 ;
        RECT 3412.835 493.030 3413.435 493.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 493.270 ;
      LAYER met4 ;
        RECT 3418.885 493.030 3419.485 493.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 493.270 ;
      LAYER met4 ;
        RECT 3423.735 493.030 3424.335 493.670 ;
      LAYER met4 ;
        RECT 3424.735 346.000 3428.185 493.270 ;
      LAYER met4 ;
        RECT 3428.585 493.030 3429.185 493.670 ;
      LAYER met4 ;
        RECT 3429.585 351.000 3434.235 493.270 ;
      LAYER met4 ;
        RECT 3434.635 493.030 3435.335 493.670 ;
      LAYER met4 ;
        RECT 3435.735 346.000 3436.065 524.910 ;
        RECT 3436.365 519.855 3439.345 739.535 ;
      LAYER met4 ;
        RECT 3439.745 715.670 3440.725 739.935 ;
      LAYER met4 ;
        RECT 3439.645 714.000 3440.825 715.270 ;
      LAYER met4 ;
        RECT 3439.645 572.000 3440.825 714.000 ;
      LAYER met4 ;
        RECT 3439.645 570.730 3440.825 572.000 ;
      LAYER met4 ;
        RECT 3439.745 535.160 3440.725 570.330 ;
      LAYER met4 ;
        RECT 3441.125 535.560 3444.105 755.240 ;
      LAYER met4 ;
        RECT 3444.505 747.310 3588.000 755.640 ;
      LAYER met4 ;
        RECT 3444.405 569.390 3444.735 746.910 ;
      LAYER met4 ;
        RECT 3445.135 715.670 3588.000 747.310 ;
        RECT 3445.135 715.030 3445.835 715.670 ;
        RECT 3445.135 572.000 3445.835 714.000 ;
        RECT 3445.135 570.330 3445.835 571.035 ;
      LAYER met4 ;
        RECT 3446.235 570.730 3450.685 715.270 ;
      LAYER met4 ;
        RECT 3451.085 715.030 3451.685 715.670 ;
        RECT 3451.085 572.000 3451.685 714.000 ;
        RECT 3451.085 570.330 3451.685 571.035 ;
      LAYER met4 ;
        RECT 3452.085 570.730 3456.535 715.270 ;
      LAYER met4 ;
        RECT 3456.935 715.030 3457.635 715.670 ;
        RECT 3456.935 572.000 3457.635 714.000 ;
        RECT 3456.935 570.330 3457.635 571.035 ;
      LAYER met4 ;
        RECT 3458.035 570.730 3483.000 715.270 ;
      LAYER met4 ;
        RECT 3483.400 715.030 3563.385 715.670 ;
      LAYER met4 ;
        RECT 3563.785 714.000 3588.000 715.270 ;
      LAYER met4 ;
        RECT 3483.400 572.000 3588.000 714.000 ;
        RECT 3483.400 570.330 3563.385 571.035 ;
      LAYER met4 ;
        RECT 3563.785 570.730 3588.000 572.000 ;
      LAYER met4 ;
        RECT 3445.135 568.990 3588.000 570.330 ;
        RECT 3444.505 535.160 3588.000 568.990 ;
        RECT 3439.745 533.640 3588.000 535.160 ;
        RECT 3439.745 519.455 3440.725 533.640 ;
        RECT 3436.465 517.935 3440.725 519.455 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 341.000 ;
      LAYER met4 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 346.000 ;
      LAYER met4 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 394.965 191.515 468.035 192.115 ;
        RECT 663.965 191.515 737.035 192.115 ;
        RECT 933.030 191.515 1011.035 192.115 ;
        RECT 1206.000 191.515 1280.035 192.115 ;
        RECT 1476.030 191.515 1554.035 192.115 ;
        RECT 1750.030 191.515 1828.035 192.115 ;
        RECT 2024.030 191.515 2102.035 192.115 ;
        RECT 2298.030 191.515 2376.035 192.115 ;
        RECT 2572.030 191.515 2650.035 192.115 ;
        RECT 2845.965 191.515 2919.035 192.115 ;
        RECT 3114.965 191.515 3188.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 395.270 191.115 ;
      LAYER met4 ;
        RECT 395.670 186.065 467.330 191.515 ;
      LAYER met4 ;
        RECT 467.730 186.465 664.270 191.115 ;
      LAYER met4 ;
        RECT 664.670 186.065 736.330 191.515 ;
      LAYER met4 ;
        RECT 736.730 186.465 933.270 191.115 ;
      LAYER met4 ;
        RECT 933.670 186.065 1010.330 191.515 ;
      LAYER met4 ;
        RECT 1010.730 186.465 1207.270 191.115 ;
      LAYER met4 ;
        RECT 1207.670 186.065 1279.330 191.515 ;
      LAYER met4 ;
        RECT 1279.730 186.465 1476.270 191.115 ;
      LAYER met4 ;
        RECT 1476.670 186.065 1553.330 191.515 ;
      LAYER met4 ;
        RECT 1553.730 186.465 1750.270 191.115 ;
      LAYER met4 ;
        RECT 1750.670 186.065 1827.330 191.515 ;
      LAYER met4 ;
        RECT 1827.730 186.465 2024.270 191.115 ;
      LAYER met4 ;
        RECT 2024.670 186.065 2101.330 191.515 ;
      LAYER met4 ;
        RECT 2101.730 186.465 2298.270 191.115 ;
      LAYER met4 ;
        RECT 2298.670 186.065 2375.330 191.515 ;
      LAYER met4 ;
        RECT 2375.730 186.465 2572.270 191.115 ;
      LAYER met4 ;
        RECT 2572.670 186.065 2649.330 191.515 ;
      LAYER met4 ;
        RECT 2649.730 186.465 2846.270 191.115 ;
      LAYER met4 ;
        RECT 2846.670 186.065 2918.330 191.515 ;
      LAYER met4 ;
        RECT 2918.730 186.465 3115.270 191.115 ;
      LAYER met4 ;
        RECT 3115.670 186.065 3187.330 191.515 ;
      LAYER met4 ;
        RECT 3187.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 394.965 185.465 468.035 186.065 ;
        RECT 663.965 185.465 737.035 186.065 ;
        RECT 933.030 185.465 1011.035 186.065 ;
        RECT 1206.000 185.465 1280.035 186.065 ;
        RECT 1476.030 185.465 1554.035 186.065 ;
        RECT 1750.030 185.465 1828.035 186.065 ;
        RECT 2024.030 185.465 2102.035 186.065 ;
        RECT 2298.030 185.465 2376.035 186.065 ;
        RECT 2572.030 185.465 2650.035 186.065 ;
        RECT 2845.965 185.465 2919.035 186.065 ;
        RECT 3114.965 185.465 3188.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 394.965 185.065 ;
      LAYER met4 ;
        RECT 395.365 181.215 467.635 185.465 ;
        RECT 664.365 181.215 736.635 185.465 ;
      LAYER met4 ;
        RECT 737.035 181.615 933.030 185.065 ;
      LAYER met4 ;
        RECT 933.430 181.215 1010.635 185.465 ;
      LAYER met4 ;
        RECT 1011.035 181.615 1206.965 185.065 ;
      LAYER met4 ;
        RECT 1207.365 181.215 1279.635 185.465 ;
      LAYER met4 ;
        RECT 1280.035 181.615 1476.030 185.065 ;
      LAYER met4 ;
        RECT 1476.430 181.215 1553.635 185.465 ;
      LAYER met4 ;
        RECT 1554.035 181.615 1750.030 185.065 ;
      LAYER met4 ;
        RECT 1750.430 181.215 1827.635 185.465 ;
      LAYER met4 ;
        RECT 1828.035 181.615 2024.030 185.065 ;
      LAYER met4 ;
        RECT 2024.430 181.215 2101.635 185.465 ;
      LAYER met4 ;
        RECT 2102.035 181.615 2298.030 185.065 ;
      LAYER met4 ;
        RECT 2298.430 181.215 2375.635 185.465 ;
      LAYER met4 ;
        RECT 2376.035 181.615 2572.030 185.065 ;
      LAYER met4 ;
        RECT 2572.430 181.215 2649.635 185.465 ;
      LAYER met4 ;
        RECT 2650.035 181.615 2845.965 185.065 ;
      LAYER met4 ;
        RECT 2846.365 181.215 2918.635 185.465 ;
      LAYER met4 ;
        RECT 2919.035 181.615 3114.965 185.065 ;
      LAYER met4 ;
        RECT 3115.365 181.215 3187.635 185.465 ;
      LAYER met4 ;
        RECT 3188.035 181.615 3385.255 185.065 ;
      LAYER met4 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 394.965 180.615 468.035 181.215 ;
        RECT 663.965 180.615 737.035 181.215 ;
        RECT 933.030 180.615 1011.035 181.215 ;
        RECT 1206.000 180.615 1280.035 181.215 ;
        RECT 1476.030 180.615 1554.035 181.215 ;
        RECT 1750.030 180.615 1828.035 181.215 ;
        RECT 2024.030 180.615 2102.035 181.215 ;
        RECT 2298.030 180.615 2376.035 181.215 ;
        RECT 2572.030 180.615 2650.035 181.215 ;
        RECT 2845.965 180.615 2919.035 181.215 ;
        RECT 3114.965 180.615 3188.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 395.270 180.215 ;
      LAYER met4 ;
        RECT 395.670 175.165 467.330 180.615 ;
      LAYER met4 ;
        RECT 467.730 175.565 664.270 180.215 ;
      LAYER met4 ;
        RECT 664.670 175.165 736.330 180.615 ;
      LAYER met4 ;
        RECT 736.730 175.565 933.270 180.215 ;
      LAYER met4 ;
        RECT 933.670 175.165 1010.330 180.615 ;
      LAYER met4 ;
        RECT 1010.730 175.565 1207.270 180.215 ;
      LAYER met4 ;
        RECT 1207.670 175.165 1279.330 180.615 ;
      LAYER met4 ;
        RECT 1279.730 175.565 1476.270 180.215 ;
      LAYER met4 ;
        RECT 1476.670 175.165 1553.330 180.615 ;
      LAYER met4 ;
        RECT 1553.730 175.565 1750.270 180.215 ;
      LAYER met4 ;
        RECT 1750.670 175.165 1827.330 180.615 ;
      LAYER met4 ;
        RECT 1827.730 175.565 2024.270 180.215 ;
      LAYER met4 ;
        RECT 2024.670 175.165 2101.330 180.615 ;
      LAYER met4 ;
        RECT 2101.730 175.565 2298.270 180.215 ;
      LAYER met4 ;
        RECT 2298.670 175.165 2375.330 180.615 ;
      LAYER met4 ;
        RECT 2375.730 175.565 2572.270 180.215 ;
      LAYER met4 ;
        RECT 2572.670 175.165 2649.330 180.615 ;
      LAYER met4 ;
        RECT 2649.730 175.565 2846.270 180.215 ;
      LAYER met4 ;
        RECT 2846.670 175.165 2918.330 180.615 ;
      LAYER met4 ;
        RECT 2918.730 175.565 3115.270 180.215 ;
      LAYER met4 ;
        RECT 3115.670 175.165 3187.330 180.615 ;
      LAYER met4 ;
        RECT 3187.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 341.000 ;
      LAYER met4 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 517.535 ;
      LAYER met4 ;
        RECT 3439.745 493.670 3440.725 517.935 ;
      LAYER met4 ;
        RECT 3439.645 492.000 3440.825 493.270 ;
      LAYER met4 ;
        RECT 3439.645 346.000 3440.825 492.000 ;
        RECT 3439.645 200.000 3440.825 341.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 533.240 ;
      LAYER met4 ;
        RECT 3444.505 525.310 3588.000 533.640 ;
      LAYER met4 ;
        RECT 3444.405 346.000 3444.735 524.910 ;
      LAYER met4 ;
        RECT 3445.135 493.670 3588.000 525.310 ;
        RECT 3445.135 493.030 3445.835 493.670 ;
        RECT 3445.135 346.000 3445.835 492.000 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 341.000 ;
      LAYER met4 ;
        RECT 3445.135 197.975 3445.835 341.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 493.270 ;
      LAYER met4 ;
        RECT 3451.085 493.030 3451.685 493.670 ;
        RECT 3451.085 346.000 3451.685 492.000 ;
        RECT 3451.085 198.120 3451.685 341.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 493.270 ;
      LAYER met4 ;
        RECT 3456.935 493.030 3457.635 493.670 ;
        RECT 3456.935 346.000 3457.635 492.000 ;
        RECT 3456.935 198.120 3457.635 341.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 493.270 ;
      LAYER met4 ;
        RECT 3483.400 493.030 3563.385 493.670 ;
      LAYER met4 ;
        RECT 3563.785 492.000 3588.000 493.270 ;
      LAYER met4 ;
        RECT 3483.400 346.000 3588.000 492.000 ;
        RECT 3563.785 341.000 3588.000 346.000 ;
        RECT 3483.400 200.000 3588.000 341.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 394.965 174.565 468.035 175.165 ;
        RECT 663.965 174.565 737.035 175.165 ;
        RECT 933.030 174.565 1011.035 175.165 ;
        RECT 1206.000 174.565 1280.035 175.165 ;
        RECT 1476.030 174.565 1554.035 175.165 ;
        RECT 1750.030 174.565 1828.035 175.165 ;
        RECT 2024.030 174.565 2102.035 175.165 ;
        RECT 2298.030 174.565 2376.035 175.165 ;
        RECT 2572.030 174.565 2650.035 175.165 ;
        RECT 2845.965 174.565 2919.035 175.165 ;
        RECT 3114.965 174.565 3188.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 395.270 174.165 ;
      LAYER met4 ;
        RECT 395.670 169.115 467.330 174.565 ;
      LAYER met4 ;
        RECT 467.730 169.515 664.270 174.165 ;
      LAYER met4 ;
        RECT 664.670 169.115 736.330 174.565 ;
      LAYER met4 ;
        RECT 736.730 169.515 933.270 174.165 ;
      LAYER met4 ;
        RECT 933.670 169.115 1010.330 174.565 ;
      LAYER met4 ;
        RECT 1010.730 169.515 1207.270 174.165 ;
      LAYER met4 ;
        RECT 1207.670 169.115 1279.330 174.565 ;
      LAYER met4 ;
        RECT 1279.730 169.515 1476.270 174.165 ;
      LAYER met4 ;
        RECT 1476.670 169.115 1553.330 174.565 ;
      LAYER met4 ;
        RECT 1553.730 169.515 1750.270 174.165 ;
      LAYER met4 ;
        RECT 1750.670 169.115 1827.330 174.565 ;
      LAYER met4 ;
        RECT 1827.730 169.515 2024.270 174.165 ;
      LAYER met4 ;
        RECT 2024.670 169.115 2101.330 174.565 ;
      LAYER met4 ;
        RECT 2101.730 169.515 2298.270 174.165 ;
      LAYER met4 ;
        RECT 2298.670 169.115 2375.330 174.565 ;
      LAYER met4 ;
        RECT 2375.730 169.515 2572.270 174.165 ;
      LAYER met4 ;
        RECT 2572.670 169.115 2649.330 174.565 ;
      LAYER met4 ;
        RECT 2649.730 169.515 2846.270 174.165 ;
      LAYER met4 ;
        RECT 2846.670 169.115 2918.330 174.565 ;
      LAYER met4 ;
        RECT 2918.730 169.515 3115.270 174.165 ;
      LAYER met4 ;
        RECT 3115.670 169.115 3187.330 174.565 ;
      LAYER met4 ;
        RECT 3187.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 394.965 168.515 468.035 169.115 ;
        RECT 663.965 168.515 737.035 169.115 ;
        RECT 933.030 168.515 1011.035 169.115 ;
        RECT 1206.000 168.515 1280.035 169.115 ;
        RECT 1476.030 168.515 1554.035 169.115 ;
        RECT 1750.030 168.515 1828.035 169.115 ;
        RECT 2024.030 168.515 2102.035 169.115 ;
        RECT 2298.030 168.515 2376.035 169.115 ;
        RECT 2572.030 168.515 2650.035 169.115 ;
        RECT 2845.965 168.515 2919.035 169.115 ;
        RECT 3114.965 168.515 3188.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 395.270 168.115 ;
      LAYER met4 ;
        RECT 395.670 164.265 467.330 168.515 ;
      LAYER met4 ;
        RECT 467.730 164.665 664.270 168.115 ;
      LAYER met4 ;
        RECT 664.670 164.265 736.330 168.515 ;
      LAYER met4 ;
        RECT 736.730 164.665 933.270 168.115 ;
      LAYER met4 ;
        RECT 933.670 164.265 1010.330 168.515 ;
      LAYER met4 ;
        RECT 1010.730 164.665 1207.270 168.115 ;
      LAYER met4 ;
        RECT 1207.670 164.265 1279.330 168.515 ;
      LAYER met4 ;
        RECT 1279.730 164.665 1476.270 168.115 ;
      LAYER met4 ;
        RECT 1476.670 164.265 1553.330 168.515 ;
      LAYER met4 ;
        RECT 1553.730 164.665 1750.270 168.115 ;
      LAYER met4 ;
        RECT 1750.670 164.265 1827.330 168.515 ;
      LAYER met4 ;
        RECT 1827.730 164.665 2024.270 168.115 ;
      LAYER met4 ;
        RECT 2024.670 164.265 2101.330 168.515 ;
      LAYER met4 ;
        RECT 2101.730 164.665 2298.270 168.115 ;
      LAYER met4 ;
        RECT 2298.670 164.265 2375.330 168.515 ;
      LAYER met4 ;
        RECT 2375.730 164.665 2572.270 168.115 ;
      LAYER met4 ;
        RECT 2572.670 164.265 2649.330 168.515 ;
      LAYER met4 ;
        RECT 2649.730 164.665 2846.270 168.115 ;
      LAYER met4 ;
        RECT 2846.670 164.265 2918.330 168.515 ;
      LAYER met4 ;
        RECT 2918.730 164.665 3115.270 168.115 ;
      LAYER met4 ;
        RECT 3115.670 164.265 3187.330 168.515 ;
      LAYER met4 ;
        RECT 3187.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 394.965 163.665 468.035 164.265 ;
        RECT 663.965 163.665 737.035 164.265 ;
        RECT 933.030 163.665 1011.035 164.265 ;
        RECT 1206.000 163.665 1280.035 164.265 ;
        RECT 1476.030 163.665 1554.035 164.265 ;
        RECT 1750.030 163.665 1828.035 164.265 ;
        RECT 2024.030 163.665 2102.035 164.265 ;
        RECT 2298.030 163.665 2376.035 164.265 ;
        RECT 2572.030 163.665 2650.035 164.265 ;
        RECT 2845.965 163.665 2919.035 164.265 ;
        RECT 3114.965 163.665 3188.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
      LAYER met4 ;
        RECT 198.665 159.815 395.270 163.265 ;
      LAYER met4 ;
        RECT 395.670 159.415 467.330 163.665 ;
      LAYER met4 ;
        RECT 467.730 159.815 664.270 163.265 ;
      LAYER met4 ;
        RECT 664.670 159.415 736.330 163.665 ;
      LAYER met4 ;
        RECT 736.730 159.815 933.270 163.265 ;
      LAYER met4 ;
        RECT 933.670 159.415 1010.330 163.665 ;
      LAYER met4 ;
        RECT 1010.730 159.815 1207.270 163.265 ;
      LAYER met4 ;
        RECT 1207.670 159.415 1279.330 163.665 ;
      LAYER met4 ;
        RECT 1279.730 159.815 1476.270 163.265 ;
      LAYER met4 ;
        RECT 1476.670 159.415 1553.330 163.665 ;
      LAYER met4 ;
        RECT 1553.730 159.815 1750.270 163.265 ;
      LAYER met4 ;
        RECT 1750.670 159.415 1827.330 163.665 ;
      LAYER met4 ;
        RECT 1827.730 159.815 2024.270 163.265 ;
      LAYER met4 ;
        RECT 2024.670 159.415 2101.330 163.665 ;
      LAYER met4 ;
        RECT 2101.730 159.815 2298.270 163.265 ;
      LAYER met4 ;
        RECT 2298.670 159.415 2375.330 163.665 ;
      LAYER met4 ;
        RECT 2375.730 159.815 2572.270 163.265 ;
      LAYER met4 ;
        RECT 2572.670 159.415 2649.330 163.665 ;
      LAYER met4 ;
        RECT 2649.730 159.815 2846.270 163.265 ;
      LAYER met4 ;
        RECT 2846.670 159.415 2918.330 163.665 ;
      LAYER met4 ;
        RECT 2918.730 159.815 3115.270 163.265 ;
      LAYER met4 ;
        RECT 3115.670 159.415 3187.330 163.665 ;
      LAYER met4 ;
        RECT 3187.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 394.965 158.815 468.035 159.415 ;
        RECT 663.965 158.815 737.035 159.415 ;
        RECT 933.030 158.815 1011.035 159.415 ;
        RECT 1206.000 158.815 1280.035 159.415 ;
        RECT 1476.030 158.815 1554.035 159.415 ;
        RECT 1750.030 158.815 1828.035 159.415 ;
        RECT 2024.030 158.815 2102.035 159.415 ;
        RECT 2298.030 158.815 2376.035 159.415 ;
        RECT 2572.030 158.815 2650.035 159.415 ;
        RECT 2845.965 158.815 2919.035 159.415 ;
        RECT 3114.965 158.815 3188.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 395.270 158.415 ;
      LAYER met4 ;
        RECT 395.670 153.365 467.330 158.815 ;
        RECT 664.670 158.770 736.330 158.815 ;
        RECT 664.745 153.410 736.330 158.770 ;
      LAYER met4 ;
        RECT 736.730 153.765 933.270 158.415 ;
      LAYER met4 ;
        RECT 664.670 153.365 736.330 153.410 ;
        RECT 933.670 153.365 1010.330 158.815 ;
      LAYER met4 ;
        RECT 1010.730 153.765 1207.270 158.415 ;
      LAYER met4 ;
        RECT 1207.670 153.365 1279.330 158.815 ;
      LAYER met4 ;
        RECT 1279.730 153.765 1476.270 158.415 ;
      LAYER met4 ;
        RECT 1476.670 153.365 1553.330 158.815 ;
      LAYER met4 ;
        RECT 1553.730 153.765 1750.270 158.415 ;
      LAYER met4 ;
        RECT 1750.670 153.365 1827.330 158.815 ;
      LAYER met4 ;
        RECT 1827.730 153.765 2024.270 158.415 ;
      LAYER met4 ;
        RECT 2024.670 153.365 2101.330 158.815 ;
      LAYER met4 ;
        RECT 2101.730 153.765 2298.270 158.415 ;
      LAYER met4 ;
        RECT 2298.670 153.365 2375.330 158.815 ;
      LAYER met4 ;
        RECT 2375.730 153.765 2572.270 158.415 ;
      LAYER met4 ;
        RECT 2572.670 153.365 2649.330 158.815 ;
      LAYER met4 ;
        RECT 2649.730 153.765 2846.270 158.415 ;
      LAYER met4 ;
        RECT 2846.670 153.365 2918.330 158.815 ;
      LAYER met4 ;
        RECT 2918.730 153.765 3115.270 158.415 ;
      LAYER met4 ;
        RECT 3115.670 153.365 3187.330 158.815 ;
      LAYER met4 ;
        RECT 3187.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 394.965 152.665 468.035 153.365 ;
        RECT 663.965 152.665 737.035 153.365 ;
        RECT 933.030 152.665 1011.035 153.365 ;
        RECT 1206.000 152.665 1280.035 153.365 ;
        RECT 1476.030 152.665 1554.035 153.365 ;
        RECT 1750.030 152.665 1828.035 153.365 ;
        RECT 2024.030 152.665 2102.035 153.365 ;
        RECT 2298.030 152.665 2376.035 153.365 ;
        RECT 2572.030 152.665 2650.035 153.365 ;
        RECT 2845.965 152.665 2919.035 153.365 ;
        RECT 3114.965 152.665 3188.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 180.425 151.935 395.270 152.265 ;
      LAYER met4 ;
        RECT 395.670 152.035 467.330 152.665 ;
      LAYER met4 ;
        RECT 467.730 151.935 964.910 152.265 ;
      LAYER met4 ;
        RECT 965.310 152.035 1008.990 152.665 ;
      LAYER met4 ;
        RECT 1009.390 151.935 1507.910 152.265 ;
      LAYER met4 ;
        RECT 1508.310 152.035 1551.990 152.665 ;
      LAYER met4 ;
        RECT 1552.390 151.935 1781.910 152.265 ;
      LAYER met4 ;
        RECT 1782.310 152.035 1825.990 152.665 ;
      LAYER met4 ;
        RECT 1826.390 151.935 2055.910 152.265 ;
      LAYER met4 ;
        RECT 2056.310 152.035 2099.990 152.665 ;
      LAYER met4 ;
        RECT 2100.390 151.935 2329.910 152.265 ;
      LAYER met4 ;
        RECT 2330.310 152.035 2373.990 152.665 ;
      LAYER met4 ;
        RECT 2374.390 151.935 2603.910 152.265 ;
      LAYER met4 ;
        RECT 2604.310 152.035 2647.990 152.665 ;
      LAYER met4 ;
        RECT 2648.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 957.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 200.000 147.175 394.000 148.355 ;
      LAYER met4 ;
        RECT 394.000 147.175 395.270 148.355 ;
      LAYER met4 ;
        RECT 395.670 147.275 467.330 148.255 ;
      LAYER met4 ;
        RECT 467.730 147.175 469.000 148.355 ;
      LAYER met4 ;
        RECT 469.000 147.175 663.000 148.355 ;
      LAYER met4 ;
        RECT 663.000 147.175 664.270 148.355 ;
      LAYER met4 ;
        RECT 664.670 147.275 736.330 148.255 ;
      LAYER met4 ;
        RECT 736.730 147.175 738.000 148.355 ;
      LAYER met4 ;
        RECT 738.000 147.175 932.000 148.355 ;
      LAYER met4 ;
        RECT 932.000 147.175 933.270 148.355 ;
      LAYER met4 ;
        RECT 957.935 148.255 959.455 151.535 ;
      LAYER met4 ;
        RECT 959.855 148.655 1500.535 151.635 ;
      LAYER met4 ;
        RECT 933.670 147.275 1010.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 973.240 146.875 ;
        RECT 176.825 143.265 395.270 143.595 ;
      LAYER met4 ;
        RECT 973.640 143.495 975.160 147.275 ;
      LAYER met4 ;
        RECT 1010.730 147.175 1012.000 148.355 ;
      LAYER met4 ;
        RECT 1012.000 147.175 1206.000 148.355 ;
      LAYER met4 ;
        RECT 1206.000 147.175 1207.270 148.355 ;
      LAYER met4 ;
        RECT 1207.670 147.275 1279.330 148.255 ;
      LAYER met4 ;
        RECT 1279.730 147.175 1281.000 148.355 ;
      LAYER met4 ;
        RECT 1281.000 147.175 1475.000 148.355 ;
      LAYER met4 ;
        RECT 1475.000 147.175 1476.270 148.355 ;
      LAYER met4 ;
        RECT 1500.935 148.255 1502.455 151.535 ;
      LAYER met4 ;
        RECT 1502.855 148.655 1774.535 151.635 ;
      LAYER met4 ;
        RECT 1476.670 147.275 1553.330 148.255 ;
      LAYER met4 ;
        RECT 975.560 143.895 1516.240 146.875 ;
      LAYER met4 ;
        RECT 395.670 142.865 467.330 143.495 ;
        RECT 965.310 142.865 1008.990 143.495 ;
      LAYER met4 ;
        RECT 1009.390 143.265 1507.910 143.595 ;
      LAYER met4 ;
        RECT 1516.640 143.495 1518.160 147.275 ;
      LAYER met4 ;
        RECT 1553.730 147.175 1555.000 148.355 ;
      LAYER met4 ;
        RECT 1555.000 147.175 1749.000 148.355 ;
      LAYER met4 ;
        RECT 1749.000 147.175 1750.270 148.355 ;
      LAYER met4 ;
        RECT 1774.935 148.255 1776.455 151.535 ;
      LAYER met4 ;
        RECT 1776.855 148.655 2048.535 151.635 ;
      LAYER met4 ;
        RECT 1750.670 147.275 1827.330 148.255 ;
      LAYER met4 ;
        RECT 1518.560 143.895 1790.240 146.875 ;
      LAYER met4 ;
        RECT 1508.310 142.865 1551.990 143.495 ;
      LAYER met4 ;
        RECT 1552.390 143.265 1781.910 143.595 ;
      LAYER met4 ;
        RECT 1790.640 143.495 1792.160 147.275 ;
      LAYER met4 ;
        RECT 1827.730 147.175 1829.000 148.355 ;
      LAYER met4 ;
        RECT 1829.000 147.175 2023.000 148.355 ;
      LAYER met4 ;
        RECT 2023.000 147.175 2024.270 148.355 ;
      LAYER met4 ;
        RECT 2048.935 148.255 2050.455 151.535 ;
      LAYER met4 ;
        RECT 2050.855 148.655 2322.535 151.635 ;
      LAYER met4 ;
        RECT 2024.670 147.275 2101.330 148.255 ;
      LAYER met4 ;
        RECT 1792.560 143.895 2064.240 146.875 ;
      LAYER met4 ;
        RECT 1782.310 142.865 1825.990 143.495 ;
      LAYER met4 ;
        RECT 1826.390 143.265 2055.910 143.595 ;
      LAYER met4 ;
        RECT 2064.640 143.495 2066.160 147.275 ;
      LAYER met4 ;
        RECT 2101.730 147.175 2103.000 148.355 ;
      LAYER met4 ;
        RECT 2103.000 147.175 2297.000 148.355 ;
      LAYER met4 ;
        RECT 2297.000 147.175 2298.270 148.355 ;
      LAYER met4 ;
        RECT 2322.935 148.255 2324.455 151.535 ;
      LAYER met4 ;
        RECT 2324.855 148.655 2596.535 151.635 ;
      LAYER met4 ;
        RECT 2298.670 147.275 2375.330 148.255 ;
      LAYER met4 ;
        RECT 2066.560 143.895 2338.240 146.875 ;
      LAYER met4 ;
        RECT 2056.310 142.865 2099.990 143.495 ;
      LAYER met4 ;
        RECT 2100.390 143.265 2329.910 143.595 ;
      LAYER met4 ;
        RECT 2338.640 143.495 2340.160 147.275 ;
      LAYER met4 ;
        RECT 2375.730 147.175 2377.000 148.355 ;
      LAYER met4 ;
        RECT 2377.000 147.175 2571.000 148.355 ;
      LAYER met4 ;
        RECT 2571.000 147.175 2572.270 148.355 ;
      LAYER met4 ;
        RECT 2596.935 148.255 2598.455 151.535 ;
      LAYER met4 ;
        RECT 2598.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 2572.670 147.275 2649.330 148.255 ;
      LAYER met4 ;
        RECT 2340.560 143.895 2612.240 146.875 ;
      LAYER met4 ;
        RECT 2330.310 142.865 2373.990 143.495 ;
      LAYER met4 ;
        RECT 2374.390 143.265 2603.910 143.595 ;
      LAYER met4 ;
        RECT 2612.640 143.495 2614.160 147.275 ;
      LAYER met4 ;
        RECT 2649.730 147.175 2651.000 148.355 ;
      LAYER met4 ;
        RECT 2651.000 147.175 2845.000 148.355 ;
      LAYER met4 ;
        RECT 2845.000 147.175 2846.270 148.355 ;
      LAYER met4 ;
        RECT 2846.670 147.275 2918.330 148.255 ;
      LAYER met4 ;
        RECT 2918.730 147.175 2920.000 148.355 ;
      LAYER met4 ;
        RECT 2920.000 147.175 3114.000 148.355 ;
      LAYER met4 ;
        RECT 3114.000 147.175 3115.270 148.355 ;
      LAYER met4 ;
        RECT 3115.670 147.275 3187.330 148.255 ;
      LAYER met4 ;
        RECT 3187.730 147.175 3189.000 148.355 ;
      LAYER met4 ;
        RECT 3189.000 147.175 3384.000 148.355 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 2614.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 2604.310 142.865 2647.990 143.495 ;
      LAYER met4 ;
        RECT 2648.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 394.000 142.865 ;
        RECT 394.965 142.165 468.035 142.865 ;
        RECT 469.000 142.165 663.000 142.865 ;
        RECT 663.965 142.165 737.035 142.865 ;
        RECT 738.000 142.165 932.000 142.865 ;
        RECT 933.030 142.165 1011.035 142.865 ;
        RECT 1012.000 142.165 1280.035 142.865 ;
        RECT 1281.000 142.165 1475.000 142.865 ;
        RECT 1476.030 142.165 1554.035 142.865 ;
        RECT 1555.000 142.165 1749.000 142.865 ;
        RECT 1750.030 142.165 1828.035 142.865 ;
        RECT 1829.000 142.165 2023.000 142.865 ;
        RECT 2024.030 142.165 2102.035 142.865 ;
        RECT 2103.000 142.165 2297.000 142.865 ;
        RECT 2298.030 142.165 2376.035 142.865 ;
        RECT 2377.000 142.165 2571.000 142.865 ;
        RECT 2572.030 142.165 2650.035 142.865 ;
        RECT 2651.000 142.165 2845.000 142.865 ;
        RECT 2845.965 142.165 2919.035 142.865 ;
        RECT 2920.000 142.165 3114.000 142.865 ;
        RECT 3114.965 142.165 3188.035 142.865 ;
        RECT 3189.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 395.270 141.765 ;
      LAYER met4 ;
        RECT 395.670 136.915 467.330 142.165 ;
      LAYER met4 ;
        RECT 467.730 137.315 664.270 141.765 ;
      LAYER met4 ;
        RECT 664.670 136.915 736.330 142.165 ;
      LAYER met4 ;
        RECT 736.730 137.315 933.270 141.765 ;
      LAYER met4 ;
        RECT 933.670 136.915 1010.330 142.165 ;
      LAYER met4 ;
        RECT 1010.730 137.315 1207.270 141.765 ;
      LAYER met4 ;
        RECT 1207.670 136.915 1279.330 142.165 ;
      LAYER met4 ;
        RECT 1279.730 137.315 1476.270 141.765 ;
      LAYER met4 ;
        RECT 1476.670 136.915 1553.330 142.165 ;
      LAYER met4 ;
        RECT 1553.730 137.315 1750.270 141.765 ;
      LAYER met4 ;
        RECT 1750.670 136.915 1827.330 142.165 ;
      LAYER met4 ;
        RECT 1827.730 137.315 2024.270 141.765 ;
      LAYER met4 ;
        RECT 2024.670 136.915 2101.330 142.165 ;
      LAYER met4 ;
        RECT 2101.730 137.315 2298.270 141.765 ;
      LAYER met4 ;
        RECT 2298.670 136.915 2375.330 142.165 ;
      LAYER met4 ;
        RECT 2375.730 137.315 2572.270 141.765 ;
      LAYER met4 ;
        RECT 2572.670 136.915 2649.330 142.165 ;
      LAYER met4 ;
        RECT 2649.730 137.315 2846.270 141.765 ;
      LAYER met4 ;
        RECT 2846.670 136.915 2918.330 142.165 ;
      LAYER met4 ;
        RECT 2918.730 137.315 3115.270 141.765 ;
      LAYER met4 ;
        RECT 3115.670 136.915 3187.330 142.165 ;
      LAYER met4 ;
        RECT 3187.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 394.000 136.915 ;
        RECT 394.965 136.315 468.035 136.915 ;
        RECT 469.000 136.315 663.000 136.915 ;
        RECT 663.965 136.315 737.035 136.915 ;
        RECT 738.000 136.315 932.000 136.915 ;
        RECT 933.030 136.315 1011.035 136.915 ;
        RECT 1012.000 136.315 1280.035 136.915 ;
        RECT 1281.000 136.315 1475.000 136.915 ;
        RECT 1476.030 136.315 1554.035 136.915 ;
        RECT 1555.000 136.315 1749.000 136.915 ;
        RECT 1750.030 136.315 1828.035 136.915 ;
        RECT 1829.000 136.315 2023.000 136.915 ;
        RECT 2024.030 136.315 2102.035 136.915 ;
        RECT 2103.000 136.315 2297.000 136.915 ;
        RECT 2298.030 136.315 2376.035 136.915 ;
        RECT 2377.000 136.315 2571.000 136.915 ;
        RECT 2572.030 136.315 2650.035 136.915 ;
        RECT 2651.000 136.315 2845.000 136.915 ;
        RECT 2845.965 136.315 2919.035 136.915 ;
        RECT 2920.000 136.315 3114.000 136.915 ;
        RECT 3114.965 136.315 3188.035 136.915 ;
        RECT 3189.000 136.315 3384.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 395.270 135.915 ;
      LAYER met4 ;
        RECT 395.670 131.065 467.330 136.315 ;
      LAYER met4 ;
        RECT 467.730 131.465 664.270 135.915 ;
      LAYER met4 ;
        RECT 664.670 131.065 736.330 136.315 ;
      LAYER met4 ;
        RECT 736.730 131.465 933.270 135.915 ;
      LAYER met4 ;
        RECT 933.670 131.065 1010.330 136.315 ;
      LAYER met4 ;
        RECT 1010.730 131.465 1207.270 135.915 ;
      LAYER met4 ;
        RECT 1207.670 131.065 1279.330 136.315 ;
      LAYER met4 ;
        RECT 1279.730 131.465 1476.270 135.915 ;
      LAYER met4 ;
        RECT 1476.670 131.065 1553.330 136.315 ;
      LAYER met4 ;
        RECT 1553.730 131.465 1750.270 135.915 ;
      LAYER met4 ;
        RECT 1750.670 131.065 1827.330 136.315 ;
      LAYER met4 ;
        RECT 1827.730 131.465 2024.270 135.915 ;
      LAYER met4 ;
        RECT 2024.670 131.065 2101.330 136.315 ;
      LAYER met4 ;
        RECT 2101.730 131.465 2298.270 135.915 ;
      LAYER met4 ;
        RECT 2298.670 131.065 2375.330 136.315 ;
      LAYER met4 ;
        RECT 2375.730 131.465 2572.270 135.915 ;
      LAYER met4 ;
        RECT 2572.670 131.065 2649.330 136.315 ;
      LAYER met4 ;
        RECT 2649.730 131.465 2846.270 135.915 ;
      LAYER met4 ;
        RECT 2846.670 131.065 2918.330 136.315 ;
      LAYER met4 ;
        RECT 2918.730 131.465 3115.270 135.915 ;
      LAYER met4 ;
        RECT 3115.670 131.065 3187.330 136.315 ;
      LAYER met4 ;
        RECT 3187.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 394.000 131.065 ;
        RECT 394.965 130.365 468.035 131.065 ;
        RECT 469.000 130.365 663.000 131.065 ;
        RECT 663.965 130.365 737.035 131.065 ;
        RECT 738.000 130.365 932.000 131.065 ;
        RECT 933.030 130.365 1011.035 131.065 ;
        RECT 1012.000 130.365 1280.035 131.065 ;
        RECT 1281.000 130.365 1475.000 131.065 ;
        RECT 1476.030 130.365 1554.035 131.065 ;
        RECT 1555.000 130.365 1749.000 131.065 ;
        RECT 1750.030 130.365 1828.035 131.065 ;
        RECT 1829.000 130.365 2023.000 131.065 ;
        RECT 2024.030 130.365 2102.035 131.065 ;
        RECT 2103.000 130.365 2297.000 131.065 ;
        RECT 2298.030 130.365 2376.035 131.065 ;
        RECT 2377.000 130.365 2571.000 131.065 ;
        RECT 2572.030 130.365 2650.035 131.065 ;
        RECT 2651.000 130.365 2845.000 131.065 ;
        RECT 2845.965 130.365 2919.035 131.065 ;
        RECT 2920.000 130.365 3114.000 131.065 ;
        RECT 3114.965 130.365 3188.035 131.065 ;
        RECT 3189.000 130.365 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
      LAYER met4 ;
        RECT 197.355 105.000 395.270 129.965 ;
      LAYER met4 ;
        RECT 395.670 104.600 467.330 130.365 ;
      LAYER met4 ;
        RECT 467.730 105.000 664.270 129.965 ;
      LAYER met4 ;
        RECT 664.670 104.600 736.330 130.365 ;
      LAYER met4 ;
        RECT 736.730 105.000 933.270 129.965 ;
      LAYER met4 ;
        RECT 933.670 104.600 1010.330 130.365 ;
      LAYER met4 ;
        RECT 1010.730 105.000 1207.270 129.965 ;
      LAYER met4 ;
        RECT 1207.670 104.600 1279.330 130.365 ;
      LAYER met4 ;
        RECT 1279.730 105.000 1476.270 129.965 ;
      LAYER met4 ;
        RECT 1476.670 104.600 1553.330 130.365 ;
      LAYER met4 ;
        RECT 1553.730 105.000 1750.270 129.965 ;
      LAYER met4 ;
        RECT 1750.670 104.600 1827.330 130.365 ;
      LAYER met4 ;
        RECT 1827.730 105.000 2024.270 129.965 ;
      LAYER met4 ;
        RECT 2024.670 104.600 2101.330 130.365 ;
      LAYER met4 ;
        RECT 2101.730 105.000 2298.270 129.965 ;
      LAYER met4 ;
        RECT 2298.670 104.600 2375.330 130.365 ;
      LAYER met4 ;
        RECT 2375.730 105.000 2572.270 129.965 ;
      LAYER met4 ;
        RECT 2572.670 104.600 2649.330 130.365 ;
      LAYER met4 ;
        RECT 2649.730 105.000 2846.270 129.965 ;
      LAYER met4 ;
        RECT 2846.670 104.600 2918.330 130.365 ;
      LAYER met4 ;
        RECT 2918.730 105.000 3115.270 129.965 ;
      LAYER met4 ;
        RECT 3115.670 104.600 3187.330 130.365 ;
      LAYER met4 ;
        RECT 3187.730 105.000 3385.855 129.965 ;
      LAYER met4 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
        RECT 0.000 24.615 394.000 104.600 ;
        RECT 394.965 24.615 468.035 104.600 ;
        RECT 0.000 0.000 198.165 24.615 ;
      LAYER met4 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 394.000 24.615 ;
      LAYER met4 ;
        RECT 394.000 0.000 395.270 24.215 ;
      LAYER met4 ;
        RECT 395.670 0.000 467.330 24.615 ;
      LAYER met4 ;
        RECT 467.730 0.000 469.000 24.215 ;
      LAYER met4 ;
        RECT 469.000 0.000 663.000 104.600 ;
        RECT 663.965 24.615 737.035 104.600 ;
      LAYER met4 ;
        RECT 663.000 0.000 664.270 24.215 ;
      LAYER met4 ;
        RECT 664.670 0.000 736.330 24.615 ;
      LAYER met4 ;
        RECT 736.730 0.000 738.000 24.215 ;
      LAYER met4 ;
        RECT 738.000 0.000 932.000 104.600 ;
        RECT 933.030 24.615 1011.035 104.600 ;
        RECT 1012.000 24.615 1280.035 104.600 ;
      LAYER met4 ;
        RECT 932.000 0.000 933.270 24.215 ;
      LAYER met4 ;
        RECT 933.670 0.000 1010.330 24.615 ;
      LAYER met4 ;
        RECT 1010.730 0.000 1012.000 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.000 1206.000 24.615 ;
      LAYER met4 ;
        RECT 1206.000 0.000 1207.270 24.215 ;
      LAYER met4 ;
        RECT 1207.670 0.000 1279.330 24.615 ;
      LAYER met4 ;
        RECT 1279.730 0.000 1281.000 24.215 ;
      LAYER met4 ;
        RECT 1281.000 0.000 1475.000 104.600 ;
        RECT 1476.030 24.615 1554.035 104.600 ;
      LAYER met4 ;
        RECT 1475.000 0.000 1476.270 24.215 ;
      LAYER met4 ;
        RECT 1476.670 0.000 1553.330 24.615 ;
      LAYER met4 ;
        RECT 1553.730 0.000 1555.000 24.215 ;
      LAYER met4 ;
        RECT 1555.000 0.000 1749.000 104.600 ;
        RECT 1750.030 24.615 1828.035 104.600 ;
      LAYER met4 ;
        RECT 1749.000 0.000 1750.270 24.215 ;
      LAYER met4 ;
        RECT 1750.670 0.000 1827.330 24.615 ;
      LAYER met4 ;
        RECT 1827.730 0.000 1829.000 24.215 ;
      LAYER met4 ;
        RECT 1829.000 0.000 2023.000 104.600 ;
        RECT 2024.030 24.615 2102.035 104.600 ;
      LAYER met4 ;
        RECT 2023.000 0.000 2024.270 24.215 ;
      LAYER met4 ;
        RECT 2024.670 0.000 2101.330 24.615 ;
      LAYER met4 ;
        RECT 2101.730 0.000 2103.000 24.215 ;
      LAYER met4 ;
        RECT 2103.000 0.000 2297.000 104.600 ;
        RECT 2298.030 24.615 2376.035 104.600 ;
      LAYER met4 ;
        RECT 2297.000 0.000 2298.270 24.215 ;
      LAYER met4 ;
        RECT 2298.670 0.000 2375.330 24.615 ;
      LAYER met4 ;
        RECT 2375.730 0.000 2377.000 24.215 ;
      LAYER met4 ;
        RECT 2377.000 0.000 2571.000 104.600 ;
        RECT 2572.030 24.615 2650.035 104.600 ;
      LAYER met4 ;
        RECT 2571.000 0.000 2572.270 24.215 ;
      LAYER met4 ;
        RECT 2572.670 0.000 2649.330 24.615 ;
      LAYER met4 ;
        RECT 2649.730 0.000 2651.000 24.215 ;
      LAYER met4 ;
        RECT 2651.000 0.000 2845.000 104.600 ;
        RECT 2845.965 24.615 2919.035 104.600 ;
      LAYER met4 ;
        RECT 2845.000 0.000 2846.270 24.215 ;
      LAYER met4 ;
        RECT 2846.670 0.000 2918.330 24.615 ;
      LAYER met4 ;
        RECT 2918.730 0.000 2920.000 24.215 ;
      LAYER met4 ;
        RECT 2920.000 0.000 3114.000 104.600 ;
        RECT 3114.965 24.615 3188.035 104.600 ;
      LAYER met4 ;
        RECT 3114.000 0.000 3115.270 24.215 ;
      LAYER met4 ;
        RECT 3115.670 0.000 3187.330 24.615 ;
      LAYER met4 ;
        RECT 3187.730 0.000 3189.000 24.215 ;
      LAYER met4 ;
        RECT 3189.000 0.000 3384.000 104.600 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 376.270 5188.000 ;
      LAYER met5 ;
        RECT 377.870 5162.185 447.130 5188.000 ;
      LAYER met5 ;
        RECT 448.730 5163.785 616.270 5188.000 ;
      LAYER met5 ;
        RECT 617.870 5162.185 687.130 5188.000 ;
      LAYER met5 ;
        RECT 688.730 5163.785 856.270 5188.000 ;
      LAYER met5 ;
        RECT 857.870 5162.185 927.130 5188.000 ;
      LAYER met5 ;
        RECT 928.730 5163.785 1100.000 5188.000 ;
      LAYER met5 ;
        RECT 375.000 5155.545 450.000 5162.185 ;
        RECT 375.000 5091.520 380.450 5155.545 ;
        RECT 444.490 5091.520 450.000 5155.545 ;
        RECT 375.000 5084.585 450.000 5091.520 ;
        RECT 615.000 5155.545 690.000 5162.185 ;
        RECT 615.000 5091.520 620.450 5155.545 ;
        RECT 684.490 5091.520 690.000 5155.545 ;
        RECT 615.000 5084.585 690.000 5091.520 ;
        RECT 855.000 5155.545 930.000 5162.185 ;
        RECT 855.000 5091.520 860.450 5155.545 ;
        RECT 924.490 5091.520 930.000 5155.545 ;
        RECT 855.000 5084.585 930.000 5091.520 ;
        RECT 1100.000 5155.545 1269.000 5188.000 ;
      LAYER met5 ;
        RECT 1269.000 5163.785 1357.000 5188.000 ;
      LAYER met5 ;
        RECT 1100.000 5091.520 1152.450 5155.545 ;
        RECT 1216.490 5091.520 1269.000 5155.545 ;
        RECT 1100.000 5084.585 1269.000 5091.520 ;
        RECT 1357.000 5155.545 1526.000 5188.000 ;
      LAYER met5 ;
        RECT 1526.000 5163.785 1697.000 5188.000 ;
      LAYER met5 ;
        RECT 1357.000 5091.520 1409.450 5155.545 ;
        RECT 1473.490 5091.520 1526.000 5155.545 ;
        RECT 1357.000 5084.585 1526.000 5091.520 ;
        RECT 1697.000 5155.545 1772.000 5188.000 ;
      LAYER met5 ;
        RECT 1772.000 5163.785 2125.270 5188.000 ;
      LAYER met5 ;
        RECT 2126.870 5162.185 2196.130 5188.000 ;
      LAYER met5 ;
        RECT 2197.730 5163.785 2372.270 5188.000 ;
      LAYER met5 ;
        RECT 2373.870 5162.185 2443.130 5188.000 ;
      LAYER met5 ;
        RECT 2444.730 5163.785 2630.270 5188.000 ;
      LAYER met5 ;
        RECT 2631.870 5162.185 2701.130 5188.000 ;
      LAYER met5 ;
        RECT 2702.730 5163.785 2878.000 5188.000 ;
      LAYER met5 ;
        RECT 1697.000 5091.520 1702.450 5155.545 ;
        RECT 1766.490 5091.520 1772.000 5155.545 ;
        RECT 1697.000 5084.585 1772.000 5091.520 ;
        RECT 2124.000 5155.545 2199.000 5162.185 ;
        RECT 2124.000 5091.520 2129.450 5155.545 ;
        RECT 2193.490 5091.520 2199.000 5155.545 ;
        RECT 2124.000 5084.585 2199.000 5091.520 ;
        RECT 2371.000 5155.545 2446.000 5162.185 ;
        RECT 2371.000 5091.520 2376.450 5155.545 ;
        RECT 2440.490 5091.520 2446.000 5155.545 ;
        RECT 2371.000 5084.585 2446.000 5091.520 ;
        RECT 2629.000 5155.545 2704.000 5162.185 ;
        RECT 2629.000 5091.520 2634.450 5155.545 ;
        RECT 2698.490 5091.520 2704.000 5155.545 ;
        RECT 2629.000 5084.585 2704.000 5091.520 ;
        RECT 2878.000 5155.545 2953.000 5188.000 ;
      LAYER met5 ;
        RECT 2953.000 5163.785 3136.270 5188.000 ;
      LAYER met5 ;
        RECT 3137.870 5162.185 3207.130 5188.000 ;
      LAYER met5 ;
        RECT 3208.730 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 2878.000 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 2953.000 5155.545 ;
        RECT 2878.000 5084.585 2953.000 5091.520 ;
        RECT 3135.000 5155.545 3210.000 5162.185 ;
        RECT 3135.000 5091.520 3140.450 5155.545 ;
        RECT 3204.490 5091.520 3210.000 5155.545 ;
        RECT 3135.000 5084.585 3210.000 5091.520 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 376.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 376.270 5056.435 ;
        RECT 202.730 5046.335 376.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 376.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 376.270 5034.135 ;
        RECT 202.730 5024.840 376.270 5028.085 ;
      LAYER met5 ;
        RECT 377.870 5024.840 447.130 5084.585 ;
      LAYER met5 ;
        RECT 448.730 5058.035 616.270 5082.985 ;
        RECT 448.730 5052.185 616.270 5056.435 ;
        RECT 448.730 5046.335 616.270 5050.585 ;
        RECT 448.730 5035.735 616.270 5044.735 ;
        RECT 448.730 5029.685 616.270 5034.135 ;
        RECT 448.730 5024.840 616.270 5028.085 ;
      LAYER met5 ;
        RECT 617.870 5024.840 687.130 5084.585 ;
      LAYER met5 ;
        RECT 688.730 5058.035 856.270 5082.985 ;
        RECT 688.730 5052.185 856.270 5056.435 ;
        RECT 688.730 5046.335 856.270 5050.585 ;
        RECT 688.730 5035.735 856.270 5044.735 ;
        RECT 688.730 5029.685 856.270 5034.135 ;
        RECT 688.730 5024.840 856.270 5028.085 ;
      LAYER met5 ;
        RECT 857.870 5024.840 927.130 5084.585 ;
      LAYER met5 ;
        RECT 928.730 5058.035 1147.715 5082.985 ;
        RECT 928.730 5052.185 1147.715 5056.435 ;
        RECT 928.730 5046.335 1147.715 5050.585 ;
      LAYER met5 ;
        RECT 1149.315 5044.735 1224.285 5084.585 ;
      LAYER met5 ;
        RECT 1225.885 5058.035 1404.715 5082.985 ;
        RECT 1225.885 5052.185 1404.715 5056.435 ;
        RECT 1225.885 5046.335 1404.715 5050.585 ;
      LAYER met5 ;
        RECT 1406.315 5044.735 1481.285 5084.585 ;
      LAYER met5 ;
        RECT 1482.885 5058.035 1698.270 5082.985 ;
        RECT 1482.885 5052.185 1698.270 5056.435 ;
        RECT 1482.885 5046.335 1698.270 5050.585 ;
        RECT 928.730 5035.735 1147.240 5044.735 ;
      LAYER met5 ;
        RECT 1148.840 5035.735 1224.285 5044.735 ;
      LAYER met5 ;
        RECT 1225.885 5035.735 1404.240 5044.735 ;
      LAYER met5 ;
        RECT 1405.840 5035.735 1481.285 5044.735 ;
      LAYER met5 ;
        RECT 1482.885 5035.735 1698.270 5044.735 ;
        RECT 928.730 5029.685 1147.715 5034.135 ;
        RECT 928.730 5024.840 1147.715 5028.085 ;
        RECT 204.000 5024.835 375.000 5024.840 ;
      LAYER met5 ;
        RECT 375.000 5024.835 450.000 5024.840 ;
      LAYER met5 ;
        RECT 450.000 5024.835 615.000 5024.840 ;
      LAYER met5 ;
        RECT 615.000 5024.835 690.000 5024.840 ;
      LAYER met5 ;
        RECT 690.000 5024.835 855.000 5024.840 ;
      LAYER met5 ;
        RECT 855.000 5024.835 930.000 5024.840 ;
      LAYER met5 ;
        RECT 930.000 5024.835 1147.715 5024.840 ;
        RECT 202.730 5019.985 376.270 5023.235 ;
        RECT 202.730 5013.935 376.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4849.730 24.215 4988.000 ;
      LAYER met5 ;
        RECT 25.815 4848.130 103.415 4851.000 ;
      LAYER met5 ;
        RECT 105.015 4849.730 129.965 4990.645 ;
        RECT 131.565 4849.730 135.815 4989.480 ;
        RECT 137.415 4849.730 141.665 4989.625 ;
        RECT 143.265 4849.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 376.270 5012.335 ;
      LAYER met5 ;
        RECT 377.870 5006.285 447.130 5024.835 ;
      LAYER met5 ;
        RECT 448.730 5019.985 616.270 5023.235 ;
        RECT 448.730 5013.935 616.270 5018.385 ;
        RECT 448.730 5007.885 616.270 5012.335 ;
      LAYER met5 ;
        RECT 617.870 5006.285 687.130 5024.835 ;
      LAYER met5 ;
        RECT 688.730 5019.985 856.270 5023.235 ;
        RECT 688.730 5013.935 856.270 5018.385 ;
        RECT 688.730 5007.885 856.270 5012.335 ;
      LAYER met5 ;
        RECT 857.870 5006.285 927.130 5024.835 ;
      LAYER met5 ;
        RECT 928.730 5019.985 1147.715 5023.235 ;
        RECT 928.730 5013.935 1147.715 5018.385 ;
        RECT 928.730 5007.885 1147.715 5012.335 ;
      LAYER met5 ;
        RECT 1149.315 5007.885 1224.285 5035.735 ;
      LAYER met5 ;
        RECT 1225.885 5029.685 1404.715 5034.135 ;
        RECT 1225.885 5024.835 1404.715 5028.085 ;
        RECT 1225.885 5019.985 1404.715 5023.235 ;
        RECT 1225.885 5013.935 1404.715 5018.385 ;
        RECT 1225.885 5007.885 1404.715 5012.335 ;
      LAYER met5 ;
        RECT 1406.315 5007.885 1481.285 5035.735 ;
      LAYER met5 ;
        RECT 1482.885 5029.685 1698.270 5034.135 ;
        RECT 1482.885 5024.840 1698.270 5028.085 ;
      LAYER met5 ;
        RECT 1699.870 5024.840 1769.130 5084.585 ;
      LAYER met5 ;
        RECT 1770.730 5058.035 2125.270 5082.985 ;
        RECT 1770.730 5052.185 2125.270 5056.435 ;
        RECT 1770.730 5046.335 2125.270 5050.585 ;
        RECT 1770.730 5035.735 1943.000 5044.735 ;
        RECT 1948.000 5035.735 2125.270 5044.735 ;
        RECT 1770.730 5029.685 1948.000 5034.135 ;
        RECT 1953.000 5029.685 2125.270 5034.135 ;
        RECT 1770.730 5024.840 1943.000 5028.085 ;
        RECT 1482.885 5024.835 1697.000 5024.840 ;
      LAYER met5 ;
        RECT 1697.000 5024.835 1772.000 5024.840 ;
      LAYER met5 ;
        RECT 1772.000 5024.835 1943.000 5024.840 ;
        RECT 1948.000 5024.840 2125.270 5028.085 ;
      LAYER met5 ;
        RECT 2126.870 5024.840 2196.130 5084.585 ;
      LAYER met5 ;
        RECT 2197.730 5058.035 2372.270 5082.985 ;
        RECT 2197.730 5052.185 2372.270 5056.435 ;
        RECT 2197.730 5046.335 2372.270 5050.585 ;
        RECT 2197.730 5035.735 2372.270 5044.735 ;
        RECT 2197.730 5029.685 2372.270 5034.135 ;
        RECT 2197.730 5024.840 2372.270 5028.085 ;
      LAYER met5 ;
        RECT 2373.870 5024.840 2443.130 5084.585 ;
      LAYER met5 ;
        RECT 2444.730 5058.035 2630.270 5082.985 ;
        RECT 2444.730 5052.185 2630.270 5056.435 ;
        RECT 2444.730 5046.335 2630.270 5050.585 ;
        RECT 2444.730 5035.735 2630.270 5044.735 ;
        RECT 2444.730 5029.685 2630.270 5034.135 ;
        RECT 2444.730 5024.840 2630.270 5028.085 ;
      LAYER met5 ;
        RECT 2631.870 5024.840 2701.130 5084.585 ;
      LAYER met5 ;
        RECT 2702.730 5058.035 2879.270 5082.985 ;
        RECT 2702.730 5052.185 2879.270 5056.435 ;
        RECT 2702.730 5046.335 2879.270 5050.585 ;
        RECT 2702.730 5035.735 2879.270 5044.735 ;
        RECT 2702.730 5029.685 2879.270 5034.135 ;
        RECT 2702.730 5024.840 2879.270 5028.085 ;
      LAYER met5 ;
        RECT 2880.870 5024.840 2950.130 5084.585 ;
      LAYER met5 ;
        RECT 2951.730 5058.035 3136.270 5082.985 ;
        RECT 2951.730 5052.185 3136.270 5056.435 ;
        RECT 2951.730 5046.335 3136.270 5050.585 ;
        RECT 2951.730 5035.735 3136.270 5044.735 ;
        RECT 2951.730 5029.685 3136.270 5034.135 ;
        RECT 2951.730 5024.840 3136.270 5028.085 ;
      LAYER met5 ;
        RECT 3137.870 5024.840 3207.130 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 3208.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 3208.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 3208.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 3208.730 5024.840 3389.335 5028.085 ;
        RECT 1948.000 5024.835 2124.000 5024.840 ;
      LAYER met5 ;
        RECT 2124.000 5024.835 2199.000 5024.840 ;
      LAYER met5 ;
        RECT 2199.000 5024.835 2371.000 5024.840 ;
      LAYER met5 ;
        RECT 2371.000 5024.835 2446.000 5024.840 ;
      LAYER met5 ;
        RECT 2446.000 5024.835 2629.000 5024.840 ;
      LAYER met5 ;
        RECT 2629.000 5024.835 2704.000 5024.840 ;
      LAYER met5 ;
        RECT 2704.000 5024.835 2878.000 5024.840 ;
      LAYER met5 ;
        RECT 2878.000 5024.835 2953.000 5024.840 ;
      LAYER met5 ;
        RECT 2953.000 5024.835 3135.000 5024.840 ;
      LAYER met5 ;
        RECT 3135.000 5024.835 3210.000 5024.840 ;
      LAYER met5 ;
        RECT 3210.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 1482.885 5019.985 1698.270 5023.235 ;
        RECT 1482.885 5013.935 1698.270 5018.385 ;
        RECT 1482.885 5007.885 1698.270 5012.335 ;
      LAYER met5 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 375.965 5006.285 ;
      LAYER met5 ;
        RECT 377.565 5003.035 447.435 5006.285 ;
      LAYER met5 ;
        RECT 449.035 5003.035 615.965 5006.285 ;
      LAYER met5 ;
        RECT 617.565 5003.035 687.435 5006.285 ;
      LAYER met5 ;
        RECT 689.035 5003.035 855.965 5006.285 ;
      LAYER met5 ;
        RECT 857.565 5003.035 927.435 5006.285 ;
      LAYER met5 ;
        RECT 929.035 5003.035 1147.715 5006.285 ;
      LAYER met5 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 376.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4849.730 158.315 4989.475 ;
        RECT 159.915 4851.000 163.165 4989.335 ;
        RECT 159.915 4849.730 163.160 4851.000 ;
      LAYER met5 ;
        RECT 163.160 4848.130 163.165 4851.000 ;
      LAYER met5 ;
        RECT 164.765 4849.730 168.015 4989.385 ;
        RECT 169.615 4849.730 174.065 4989.600 ;
        RECT 175.665 4849.730 180.115 4989.525 ;
        RECT 181.715 4850.035 184.965 4989.470 ;
        RECT 186.565 4849.730 191.015 4991.785 ;
        RECT 192.615 4849.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4988.535 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 376.270 4995.385 ;
      LAYER met5 ;
        RECT 377.870 4990.135 447.130 5003.035 ;
      LAYER met5 ;
        RECT 448.730 4996.985 616.270 5001.435 ;
        RECT 448.730 4990.135 616.270 4995.385 ;
      LAYER met5 ;
        RECT 617.870 4990.135 687.130 5003.035 ;
      LAYER met5 ;
        RECT 688.730 4996.985 856.270 5001.435 ;
        RECT 688.730 4990.135 856.270 4995.385 ;
      LAYER met5 ;
        RECT 857.870 4990.135 927.130 5003.035 ;
        RECT 1149.315 5001.435 1219.605 5007.885 ;
      LAYER met5 ;
        RECT 1221.205 5003.035 1404.715 5006.285 ;
      LAYER met5 ;
        RECT 1406.315 5001.435 1476.605 5007.885 ;
        RECT 1699.870 5006.285 1769.130 5024.835 ;
      LAYER met5 ;
        RECT 1770.730 5019.985 2125.270 5023.235 ;
        RECT 1770.730 5013.935 2125.270 5018.385 ;
        RECT 1770.730 5007.885 2125.270 5012.335 ;
      LAYER met5 ;
        RECT 2126.870 5006.285 2196.130 5024.835 ;
      LAYER met5 ;
        RECT 2197.730 5019.985 2372.270 5023.235 ;
        RECT 2197.730 5013.935 2372.270 5018.385 ;
        RECT 2197.730 5007.885 2372.270 5012.335 ;
      LAYER met5 ;
        RECT 2373.870 5006.285 2443.130 5024.835 ;
      LAYER met5 ;
        RECT 2444.730 5019.985 2630.270 5023.235 ;
        RECT 2444.730 5013.935 2630.270 5018.385 ;
        RECT 2444.730 5007.885 2630.270 5012.335 ;
      LAYER met5 ;
        RECT 2631.870 5006.285 2701.130 5024.835 ;
      LAYER met5 ;
        RECT 2702.730 5019.985 2879.270 5023.235 ;
        RECT 2702.730 5013.935 2879.270 5018.385 ;
        RECT 2702.730 5007.885 2879.270 5012.335 ;
      LAYER met5 ;
        RECT 2880.870 5006.285 2950.130 5024.835 ;
      LAYER met5 ;
        RECT 2951.730 5019.985 3136.270 5023.235 ;
        RECT 2951.730 5013.935 3136.270 5018.385 ;
        RECT 2951.730 5007.885 3136.270 5012.335 ;
      LAYER met5 ;
        RECT 3137.870 5006.285 3207.130 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 3208.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
      LAYER met5 ;
        RECT 1478.205 5003.035 1697.965 5006.285 ;
      LAYER met5 ;
        RECT 1699.565 5003.035 1769.435 5006.285 ;
      LAYER met5 ;
        RECT 1771.035 5003.035 1943.000 5006.285 ;
        RECT 1948.000 5003.035 2124.965 5006.285 ;
      LAYER met5 ;
        RECT 2126.565 5003.035 2196.435 5006.285 ;
      LAYER met5 ;
        RECT 2198.035 5003.035 2371.965 5006.285 ;
      LAYER met5 ;
        RECT 2373.565 5003.035 2443.435 5006.285 ;
      LAYER met5 ;
        RECT 2445.035 5003.035 2629.965 5006.285 ;
      LAYER met5 ;
        RECT 2631.565 5003.035 2701.435 5006.285 ;
      LAYER met5 ;
        RECT 2703.035 5003.035 2878.965 5006.285 ;
      LAYER met5 ;
        RECT 2880.565 5003.035 2950.435 5006.285 ;
      LAYER met5 ;
        RECT 2952.035 5003.035 3135.965 5006.285 ;
      LAYER met5 ;
        RECT 3137.565 5003.035 3207.435 5006.285 ;
      LAYER met5 ;
        RECT 3209.035 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
      LAYER met5 ;
        RECT 928.730 4996.985 1147.715 5001.435 ;
        RECT 928.730 4990.135 1147.715 4995.385 ;
      LAYER met5 ;
        RECT 1149.315 4990.135 1224.285 5001.435 ;
      LAYER met5 ;
        RECT 1225.885 4996.985 1404.715 5001.435 ;
        RECT 1225.885 4990.135 1404.715 4995.385 ;
      LAYER met5 ;
        RECT 1406.315 4990.135 1481.285 5001.435 ;
      LAYER met5 ;
        RECT 1482.885 4996.985 1698.270 5001.435 ;
        RECT 1482.885 4990.135 1698.270 4995.385 ;
      LAYER met5 ;
        RECT 1699.870 4990.135 1769.130 5003.035 ;
      LAYER met5 ;
        RECT 1770.730 4996.985 1948.000 5001.435 ;
        RECT 1953.000 4996.985 2125.270 5001.435 ;
        RECT 1770.730 4990.135 2125.270 4995.385 ;
      LAYER met5 ;
        RECT 2126.870 4990.135 2196.130 5003.035 ;
      LAYER met5 ;
        RECT 2197.730 4996.985 2372.270 5001.435 ;
        RECT 2197.730 4990.135 2372.270 4995.385 ;
      LAYER met5 ;
        RECT 2373.870 4990.135 2443.130 5003.035 ;
      LAYER met5 ;
        RECT 2444.730 4996.985 2630.270 5001.435 ;
        RECT 2444.730 4990.135 2630.270 4995.385 ;
      LAYER met5 ;
        RECT 2631.870 4990.135 2701.130 5003.035 ;
      LAYER met5 ;
        RECT 2702.730 4996.985 2879.270 5001.435 ;
        RECT 2702.730 4990.135 2879.270 4995.385 ;
      LAYER met5 ;
        RECT 2880.870 4990.135 2950.130 5003.035 ;
      LAYER met5 ;
        RECT 2951.730 4996.985 3136.270 5001.435 ;
        RECT 2951.730 4990.135 3136.270 4995.385 ;
      LAYER met5 ;
        RECT 3137.870 4990.135 3207.130 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4848.130 184.965 4848.435 ;
        RECT 0.000 4845.490 197.865 4848.130 ;
        RECT 0.000 4781.450 32.455 4845.490 ;
        RECT 96.480 4781.450 197.865 4845.490 ;
      LAYER met5 ;
        RECT 3390.135 4794.285 3395.385 4985.270 ;
        RECT 3396.985 4794.285 3401.435 4985.270 ;
        RECT 3403.035 4794.285 3406.285 4985.255 ;
        RECT 3407.885 4794.285 3412.335 4985.270 ;
        RECT 3413.935 4794.285 3418.385 4985.270 ;
        RECT 3419.985 4794.285 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4794.285 3428.085 4984.000 ;
        RECT 3429.685 4794.285 3434.135 4985.270 ;
        RECT 3435.735 4794.760 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4794.285 3450.585 4985.270 ;
        RECT 3452.185 4794.285 3456.435 4985.270 ;
        RECT 3458.035 4794.285 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
      LAYER met5 ;
        RECT 3563.785 4842.000 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 3435.735 4792.685 3444.735 4793.160 ;
        RECT 3484.585 4792.685 3588.000 4842.000 ;
        RECT 0.000 4778.870 197.865 4781.450 ;
        RECT 3390.135 4789.550 3588.000 4792.685 ;
      LAYER met5 ;
        RECT 0.000 4640.000 24.215 4777.270 ;
      LAYER met5 ;
        RECT 25.815 4776.000 103.415 4778.870 ;
        RECT 0.000 4637.130 103.415 4640.000 ;
      LAYER met5 ;
        RECT 105.015 4638.730 129.965 4777.270 ;
        RECT 131.565 4638.730 135.815 4777.270 ;
        RECT 137.415 4638.730 141.665 4777.270 ;
        RECT 143.265 4638.730 152.265 4777.270 ;
        RECT 153.865 4638.730 158.315 4777.270 ;
        RECT 159.915 4776.000 163.160 4777.270 ;
      LAYER met5 ;
        RECT 163.160 4776.000 163.165 4778.870 ;
        RECT 181.715 4778.565 184.965 4778.870 ;
      LAYER met5 ;
        RECT 159.915 4640.000 163.165 4776.000 ;
        RECT 159.915 4638.730 163.160 4640.000 ;
        RECT 164.765 4638.730 168.015 4777.270 ;
        RECT 169.615 4638.730 174.065 4777.270 ;
        RECT 175.665 4638.730 180.115 4777.270 ;
        RECT 181.715 4639.035 184.965 4776.965 ;
        RECT 186.565 4638.730 191.015 4777.270 ;
        RECT 192.615 4638.730 197.865 4777.270 ;
      LAYER met5 ;
        RECT 3390.135 4725.510 3491.520 4789.550 ;
        RECT 3555.545 4725.510 3588.000 4789.550 ;
        RECT 3390.135 4722.395 3588.000 4725.510 ;
        RECT 3390.135 4717.715 3401.435 4722.395 ;
        RECT 181.715 4637.130 184.965 4637.435 ;
        RECT 0.000 4631.270 197.865 4637.130 ;
        RECT 0.000 4573.670 29.235 4631.270 ;
        RECT 99.700 4573.670 197.865 4631.270 ;
        RECT 0.000 4567.870 197.865 4573.670 ;
        RECT 0.000 4565.000 103.415 4567.870 ;
        RECT 181.715 4567.565 184.965 4567.870 ;
      LAYER met5 ;
        RECT 0.000 4429.000 24.215 4565.000 ;
      LAYER met5 ;
        RECT 0.000 4426.130 103.415 4429.000 ;
      LAYER met5 ;
        RECT 105.015 4427.730 129.965 4566.270 ;
        RECT 131.565 4427.730 135.815 4566.270 ;
        RECT 137.415 4427.730 141.665 4566.270 ;
        RECT 143.265 4427.730 152.265 4566.270 ;
        RECT 153.865 4427.730 158.315 4566.270 ;
        RECT 159.915 4565.000 163.160 4566.270 ;
        RECT 159.915 4429.000 163.165 4565.000 ;
        RECT 159.915 4427.730 163.160 4429.000 ;
      LAYER met5 ;
        RECT 163.160 4426.130 163.165 4429.000 ;
      LAYER met5 ;
        RECT 164.765 4427.730 168.015 4566.270 ;
        RECT 169.615 4427.730 174.065 4566.270 ;
        RECT 175.665 4427.730 180.115 4566.270 ;
        RECT 181.715 4428.035 184.965 4565.965 ;
        RECT 186.565 4427.730 191.015 4566.270 ;
        RECT 192.615 4427.730 197.865 4566.270 ;
        RECT 3390.135 4530.730 3395.385 4716.115 ;
        RECT 3396.985 4530.730 3401.435 4716.115 ;
        RECT 3403.035 4531.035 3406.285 4720.795 ;
      LAYER met5 ;
        RECT 3407.885 4717.715 3588.000 4722.395 ;
      LAYER met5 ;
        RECT 3407.885 4530.730 3412.335 4716.115 ;
        RECT 3413.935 4530.730 3418.385 4716.115 ;
        RECT 3419.985 4530.730 3423.235 4716.115 ;
        RECT 3424.835 4532.000 3428.085 4716.115 ;
        RECT 3424.840 4530.730 3428.085 4532.000 ;
        RECT 3429.685 4530.730 3434.135 4716.115 ;
        RECT 3435.735 4530.730 3444.735 4716.115 ;
        RECT 3446.335 4530.730 3450.585 4716.115 ;
        RECT 3452.185 4530.730 3456.435 4716.115 ;
        RECT 3458.035 4530.730 3482.985 4716.115 ;
      LAYER met5 ;
        RECT 3484.585 4673.000 3588.000 4717.715 ;
      LAYER met5 ;
        RECT 3563.785 4532.000 3588.000 4673.000 ;
      LAYER met5 ;
        RECT 3403.035 4529.130 3406.285 4529.435 ;
        RECT 3484.585 4529.130 3588.000 4532.000 ;
        RECT 3390.135 4523.330 3588.000 4529.130 ;
        RECT 3390.135 4465.730 3488.300 4523.330 ;
        RECT 3558.765 4465.730 3588.000 4523.330 ;
        RECT 3390.135 4459.870 3588.000 4465.730 ;
        RECT 3403.035 4459.565 3406.285 4459.870 ;
        RECT 181.715 4426.130 184.965 4426.435 ;
        RECT 0.000 4423.490 197.865 4426.130 ;
        RECT 0.000 4359.450 32.455 4423.490 ;
        RECT 96.480 4359.450 197.865 4423.490 ;
        RECT 0.000 4356.870 197.865 4359.450 ;
        RECT 0.000 4354.000 103.415 4356.870 ;
      LAYER met5 ;
        RECT 0.000 4217.000 24.215 4354.000 ;
      LAYER met5 ;
        RECT 0.000 4214.130 103.415 4217.000 ;
      LAYER met5 ;
        RECT 105.015 4215.730 129.965 4355.270 ;
        RECT 131.565 4215.730 135.815 4355.270 ;
        RECT 137.415 4215.730 141.665 4355.270 ;
        RECT 143.265 4215.730 152.265 4355.270 ;
        RECT 153.865 4215.730 158.315 4355.270 ;
        RECT 159.915 4354.000 163.160 4355.270 ;
      LAYER met5 ;
        RECT 163.160 4354.000 163.165 4356.870 ;
        RECT 181.715 4356.565 184.965 4356.870 ;
      LAYER met5 ;
        RECT 159.915 4217.000 163.165 4354.000 ;
        RECT 159.915 4215.730 163.160 4217.000 ;
      LAYER met5 ;
        RECT 163.160 4214.130 163.165 4217.000 ;
      LAYER met5 ;
        RECT 164.765 4215.730 168.015 4355.270 ;
        RECT 169.615 4215.730 174.065 4355.270 ;
        RECT 175.665 4215.730 180.115 4355.270 ;
        RECT 181.715 4216.035 184.965 4354.965 ;
        RECT 186.565 4215.730 191.015 4355.270 ;
        RECT 192.615 4215.730 197.865 4355.270 ;
        RECT 3390.135 4313.730 3395.385 4458.270 ;
        RECT 3396.985 4313.730 3401.435 4458.270 ;
        RECT 3403.035 4314.035 3406.285 4457.965 ;
        RECT 3407.885 4313.730 3412.335 4458.270 ;
        RECT 3413.935 4313.730 3418.385 4458.270 ;
        RECT 3419.985 4313.730 3423.235 4458.270 ;
        RECT 3424.840 4457.000 3428.085 4458.270 ;
        RECT 3424.835 4315.000 3428.085 4457.000 ;
        RECT 3424.840 4313.730 3428.085 4315.000 ;
        RECT 3429.685 4313.730 3434.135 4458.270 ;
        RECT 3435.735 4313.730 3444.735 4458.270 ;
        RECT 3446.335 4313.730 3450.585 4458.270 ;
        RECT 3452.185 4313.730 3456.435 4458.270 ;
        RECT 3458.035 4313.730 3482.985 4458.270 ;
      LAYER met5 ;
        RECT 3484.585 4457.000 3588.000 4459.870 ;
      LAYER met5 ;
        RECT 3563.785 4315.000 3588.000 4457.000 ;
      LAYER met5 ;
        RECT 3403.035 4312.130 3406.285 4312.435 ;
        RECT 3484.585 4312.130 3588.000 4315.000 ;
        RECT 3390.135 4305.500 3588.000 4312.130 ;
        RECT 3390.135 4239.600 3490.960 4305.500 ;
        RECT 3556.610 4239.600 3588.000 4305.500 ;
        RECT 3390.135 4237.870 3588.000 4239.600 ;
        RECT 3403.035 4237.630 3406.285 4237.870 ;
        RECT 181.715 4214.130 184.965 4214.435 ;
        RECT 0.000 4211.490 197.865 4214.130 ;
        RECT 0.000 4147.450 32.455 4211.490 ;
        RECT 96.480 4147.450 197.865 4211.490 ;
        RECT 0.000 4144.870 197.865 4147.450 ;
        RECT 0.000 4142.000 103.415 4144.870 ;
      LAYER met5 ;
        RECT 0.000 4006.000 24.215 4142.000 ;
      LAYER met5 ;
        RECT 0.000 4003.130 103.415 4006.000 ;
      LAYER met5 ;
        RECT 105.015 4004.730 129.965 4143.270 ;
        RECT 131.565 4004.730 135.815 4143.270 ;
        RECT 137.415 4004.730 141.665 4143.270 ;
        RECT 143.265 4004.730 152.265 4143.270 ;
        RECT 153.865 4004.730 158.315 4143.270 ;
        RECT 159.915 4142.000 163.160 4143.270 ;
      LAYER met5 ;
        RECT 163.160 4142.000 163.165 4144.870 ;
        RECT 181.715 4144.565 184.965 4144.870 ;
      LAYER met5 ;
        RECT 159.915 4006.000 163.165 4142.000 ;
        RECT 159.915 4004.730 163.160 4006.000 ;
        RECT 164.765 4004.730 168.015 4143.270 ;
        RECT 169.615 4004.730 174.065 4143.270 ;
        RECT 175.665 4004.730 180.115 4143.270 ;
        RECT 181.715 4004.970 184.965 4142.965 ;
        RECT 186.565 4004.730 191.015 4143.270 ;
        RECT 192.615 4004.730 197.865 4143.270 ;
        RECT 3390.135 4092.730 3395.385 4236.270 ;
        RECT 3396.985 4092.730 3401.435 4236.270 ;
        RECT 3403.035 4093.035 3406.285 4236.030 ;
        RECT 3407.885 4092.730 3412.335 4236.270 ;
        RECT 3413.935 4092.730 3418.385 4236.270 ;
        RECT 3419.985 4092.730 3423.235 4236.270 ;
        RECT 3424.840 4235.000 3428.085 4236.270 ;
        RECT 3424.835 4094.000 3428.085 4235.000 ;
      LAYER met5 ;
        RECT 3403.035 4091.130 3406.285 4091.435 ;
        RECT 3424.835 4091.130 3424.840 4094.000 ;
      LAYER met5 ;
        RECT 3424.840 4092.730 3428.085 4094.000 ;
        RECT 3429.685 4092.730 3434.135 4236.270 ;
        RECT 3435.735 4092.730 3444.735 4236.270 ;
        RECT 3446.335 4092.730 3450.585 4236.270 ;
        RECT 3452.185 4092.730 3456.435 4236.270 ;
        RECT 3458.035 4092.730 3482.985 4236.270 ;
      LAYER met5 ;
        RECT 3484.585 4235.000 3588.000 4237.870 ;
      LAYER met5 ;
        RECT 3563.785 4094.000 3588.000 4235.000 ;
      LAYER met5 ;
        RECT 3484.585 4091.130 3588.000 4094.000 ;
        RECT 3390.135 4088.550 3588.000 4091.130 ;
        RECT 3390.135 4024.510 3491.520 4088.550 ;
        RECT 3555.545 4024.510 3588.000 4088.550 ;
        RECT 3390.135 4021.870 3588.000 4024.510 ;
        RECT 3403.035 4021.565 3406.285 4021.870 ;
        RECT 181.715 4003.130 184.965 4003.370 ;
        RECT 0.000 4001.400 197.865 4003.130 ;
        RECT 0.000 3935.500 31.390 4001.400 ;
        RECT 97.040 3935.500 197.865 4001.400 ;
        RECT 0.000 3928.870 197.865 3935.500 ;
        RECT 0.000 3926.000 103.415 3928.870 ;
        RECT 181.715 3928.565 184.965 3928.870 ;
      LAYER met5 ;
        RECT 0.000 3790.000 24.215 3926.000 ;
      LAYER met5 ;
        RECT 0.000 3787.130 103.415 3790.000 ;
      LAYER met5 ;
        RECT 105.015 3788.730 129.965 3927.270 ;
        RECT 131.565 3788.730 135.815 3927.270 ;
        RECT 137.415 3788.730 141.665 3927.270 ;
        RECT 143.265 3788.730 152.265 3927.270 ;
        RECT 153.865 3788.730 158.315 3927.270 ;
        RECT 159.915 3926.000 163.160 3927.270 ;
        RECT 159.915 3790.000 163.165 3926.000 ;
        RECT 159.915 3788.730 163.160 3790.000 ;
        RECT 164.765 3788.730 168.015 3927.270 ;
        RECT 169.615 3788.730 174.065 3927.270 ;
        RECT 175.665 3788.730 180.115 3927.270 ;
        RECT 181.715 3788.970 184.965 3926.965 ;
        RECT 186.565 3788.730 191.015 3927.270 ;
        RECT 192.615 3788.730 197.865 3927.270 ;
        RECT 3390.135 3876.730 3395.385 4020.270 ;
        RECT 3396.985 3876.730 3401.435 4020.270 ;
        RECT 3403.035 3877.035 3406.285 4019.965 ;
        RECT 3407.885 3876.730 3412.335 4020.270 ;
        RECT 3413.935 3876.730 3418.385 4020.270 ;
        RECT 3419.985 3876.730 3423.235 4020.270 ;
      LAYER met5 ;
        RECT 3424.835 4019.000 3424.840 4021.870 ;
      LAYER met5 ;
        RECT 3424.840 4019.000 3428.085 4020.270 ;
        RECT 3424.835 3878.000 3428.085 4019.000 ;
        RECT 3424.840 3876.730 3428.085 3878.000 ;
        RECT 3429.685 3876.730 3434.135 4020.270 ;
        RECT 3435.735 3876.730 3444.735 4020.270 ;
        RECT 3446.335 3876.730 3450.585 4020.270 ;
        RECT 3452.185 3876.730 3456.435 4020.270 ;
        RECT 3458.035 3876.730 3482.985 4020.270 ;
      LAYER met5 ;
        RECT 3484.585 4019.000 3588.000 4021.870 ;
      LAYER met5 ;
        RECT 3563.785 3878.000 3588.000 4019.000 ;
      LAYER met5 ;
        RECT 3403.035 3875.130 3406.285 3875.435 ;
        RECT 3484.585 3875.130 3588.000 3878.000 ;
        RECT 3390.135 3868.500 3588.000 3875.130 ;
        RECT 3390.135 3802.600 3490.960 3868.500 ;
        RECT 3556.610 3802.600 3588.000 3868.500 ;
        RECT 3390.135 3800.870 3588.000 3802.600 ;
        RECT 3403.035 3800.630 3406.285 3800.870 ;
        RECT 181.715 3787.130 184.965 3787.370 ;
        RECT 0.000 3785.400 197.865 3787.130 ;
        RECT 0.000 3719.500 31.390 3785.400 ;
        RECT 97.040 3719.500 197.865 3785.400 ;
        RECT 0.000 3712.870 197.865 3719.500 ;
        RECT 0.000 3710.000 103.415 3712.870 ;
        RECT 181.715 3712.565 184.965 3712.870 ;
      LAYER met5 ;
        RECT 0.000 3574.000 24.215 3710.000 ;
      LAYER met5 ;
        RECT 0.000 3571.130 103.415 3574.000 ;
      LAYER met5 ;
        RECT 105.015 3572.730 129.965 3711.270 ;
        RECT 131.565 3572.730 135.815 3711.270 ;
        RECT 137.415 3572.730 141.665 3711.270 ;
        RECT 143.265 3572.730 152.265 3711.270 ;
        RECT 153.865 3572.730 158.315 3711.270 ;
        RECT 159.915 3710.000 163.160 3711.270 ;
        RECT 159.915 3574.000 163.165 3710.000 ;
        RECT 159.915 3572.730 163.160 3574.000 ;
        RECT 164.765 3572.730 168.015 3711.270 ;
        RECT 169.615 3572.730 174.065 3711.270 ;
        RECT 175.665 3572.730 180.115 3711.270 ;
        RECT 181.715 3572.970 184.965 3710.965 ;
        RECT 186.565 3572.730 191.015 3711.270 ;
        RECT 192.615 3572.730 197.865 3711.270 ;
        RECT 3390.135 3654.730 3395.385 3799.270 ;
        RECT 3396.985 3654.730 3401.435 3799.270 ;
        RECT 3403.035 3655.035 3406.285 3799.030 ;
        RECT 3407.885 3654.730 3412.335 3799.270 ;
        RECT 3413.935 3654.730 3418.385 3799.270 ;
        RECT 3419.985 3654.730 3423.235 3799.270 ;
        RECT 3424.840 3798.000 3428.085 3799.270 ;
        RECT 3424.835 3656.000 3428.085 3798.000 ;
        RECT 3424.840 3654.730 3428.085 3656.000 ;
        RECT 3429.685 3654.730 3434.135 3799.270 ;
        RECT 3435.735 3654.730 3444.735 3799.270 ;
        RECT 3446.335 3654.730 3450.585 3799.270 ;
        RECT 3452.185 3654.730 3456.435 3799.270 ;
        RECT 3458.035 3654.730 3482.985 3799.270 ;
      LAYER met5 ;
        RECT 3484.585 3798.000 3588.000 3800.870 ;
      LAYER met5 ;
        RECT 3563.785 3656.000 3588.000 3798.000 ;
      LAYER met5 ;
        RECT 3403.035 3653.130 3406.285 3653.435 ;
        RECT 3484.585 3653.130 3588.000 3656.000 ;
        RECT 3390.135 3646.500 3588.000 3653.130 ;
        RECT 3390.135 3580.600 3490.960 3646.500 ;
        RECT 3556.610 3580.600 3588.000 3646.500 ;
        RECT 3390.135 3578.870 3588.000 3580.600 ;
        RECT 3403.035 3578.630 3406.285 3578.870 ;
        RECT 181.715 3571.130 184.965 3571.370 ;
        RECT 0.000 3569.400 197.865 3571.130 ;
        RECT 0.000 3503.500 31.390 3569.400 ;
        RECT 97.040 3503.500 197.865 3569.400 ;
        RECT 0.000 3496.870 197.865 3503.500 ;
        RECT 0.000 3494.000 103.415 3496.870 ;
        RECT 181.715 3496.565 184.965 3496.870 ;
      LAYER met5 ;
        RECT 0.000 3357.000 24.215 3494.000 ;
      LAYER met5 ;
        RECT 0.000 3354.130 103.415 3357.000 ;
      LAYER met5 ;
        RECT 105.015 3355.730 129.965 3495.270 ;
        RECT 131.565 3355.730 135.815 3495.270 ;
        RECT 137.415 3355.730 141.665 3495.270 ;
        RECT 143.265 3355.730 152.265 3495.270 ;
        RECT 153.865 3355.730 158.315 3495.270 ;
        RECT 159.915 3494.000 163.160 3495.270 ;
        RECT 159.915 3357.000 163.165 3494.000 ;
        RECT 159.915 3355.730 163.160 3357.000 ;
        RECT 164.765 3355.730 168.015 3495.270 ;
        RECT 169.615 3355.730 174.065 3495.270 ;
        RECT 175.665 3355.730 180.115 3495.270 ;
        RECT 181.715 3355.970 184.965 3494.965 ;
        RECT 186.565 3355.730 191.015 3495.270 ;
        RECT 192.615 3355.730 197.865 3495.270 ;
        RECT 3390.135 3433.730 3395.385 3577.270 ;
        RECT 3396.985 3433.730 3401.435 3577.270 ;
        RECT 3403.035 3434.035 3406.285 3577.030 ;
        RECT 3407.885 3433.730 3412.335 3577.270 ;
        RECT 3413.935 3433.730 3418.385 3577.270 ;
        RECT 3419.985 3433.730 3423.235 3577.270 ;
        RECT 3424.840 3576.000 3428.085 3577.270 ;
        RECT 3424.835 3435.000 3428.085 3576.000 ;
        RECT 3424.840 3433.730 3428.085 3435.000 ;
        RECT 3429.685 3433.730 3434.135 3577.270 ;
        RECT 3435.735 3433.730 3444.735 3577.270 ;
        RECT 3446.335 3433.730 3450.585 3577.270 ;
        RECT 3452.185 3433.730 3456.435 3577.270 ;
        RECT 3458.035 3433.730 3482.985 3577.270 ;
      LAYER met5 ;
        RECT 3484.585 3576.000 3588.000 3578.870 ;
      LAYER met5 ;
        RECT 3563.785 3435.000 3588.000 3576.000 ;
      LAYER met5 ;
        RECT 3403.035 3432.130 3406.285 3432.435 ;
        RECT 3484.585 3432.130 3588.000 3435.000 ;
        RECT 3390.135 3425.500 3588.000 3432.130 ;
        RECT 3390.135 3359.600 3490.960 3425.500 ;
        RECT 3556.610 3359.600 3588.000 3425.500 ;
        RECT 3390.135 3357.870 3588.000 3359.600 ;
        RECT 3403.035 3357.630 3406.285 3357.870 ;
        RECT 181.715 3354.130 184.965 3354.370 ;
        RECT 0.000 3352.400 197.865 3354.130 ;
        RECT 0.000 3286.500 31.390 3352.400 ;
        RECT 97.040 3286.500 197.865 3352.400 ;
        RECT 0.000 3279.870 197.865 3286.500 ;
        RECT 0.000 3277.000 103.415 3279.870 ;
        RECT 181.715 3279.565 184.965 3279.870 ;
      LAYER met5 ;
        RECT 0.000 3141.000 24.215 3277.000 ;
      LAYER met5 ;
        RECT 0.000 3138.130 103.415 3141.000 ;
      LAYER met5 ;
        RECT 105.015 3139.730 129.965 3278.270 ;
        RECT 131.565 3139.730 135.815 3278.270 ;
        RECT 137.415 3139.730 141.665 3278.270 ;
        RECT 143.265 3139.730 152.265 3278.270 ;
        RECT 153.865 3139.730 158.315 3278.270 ;
        RECT 159.915 3277.000 163.160 3278.270 ;
        RECT 159.915 3141.000 163.165 3277.000 ;
        RECT 159.915 3139.730 163.160 3141.000 ;
        RECT 164.765 3139.730 168.015 3278.270 ;
        RECT 169.615 3139.730 174.065 3278.270 ;
        RECT 175.665 3139.730 180.115 3278.270 ;
        RECT 181.715 3139.970 184.965 3277.965 ;
        RECT 186.565 3139.730 191.015 3278.270 ;
        RECT 192.615 3139.730 197.865 3278.270 ;
        RECT 3390.135 3212.730 3395.385 3356.270 ;
        RECT 3396.985 3212.730 3401.435 3356.270 ;
        RECT 3403.035 3213.035 3406.285 3356.030 ;
        RECT 3407.885 3212.730 3412.335 3356.270 ;
        RECT 3413.935 3212.730 3418.385 3356.270 ;
        RECT 3419.985 3212.730 3423.235 3356.270 ;
        RECT 3424.840 3355.000 3428.085 3356.270 ;
        RECT 3424.835 3214.000 3428.085 3355.000 ;
        RECT 3424.840 3212.730 3428.085 3214.000 ;
        RECT 3429.685 3212.730 3434.135 3356.270 ;
        RECT 3435.735 3212.730 3444.735 3356.270 ;
        RECT 3446.335 3212.730 3450.585 3356.270 ;
        RECT 3452.185 3212.730 3456.435 3356.270 ;
        RECT 3458.035 3212.730 3482.985 3356.270 ;
      LAYER met5 ;
        RECT 3484.585 3355.000 3588.000 3357.870 ;
      LAYER met5 ;
        RECT 3563.785 3214.000 3588.000 3355.000 ;
      LAYER met5 ;
        RECT 3403.035 3211.130 3406.285 3211.435 ;
        RECT 3484.585 3211.130 3588.000 3214.000 ;
        RECT 3390.135 3204.500 3588.000 3211.130 ;
        RECT 3390.135 3138.600 3490.960 3204.500 ;
        RECT 3556.610 3138.600 3588.000 3204.500 ;
        RECT 181.715 3138.130 184.965 3138.370 ;
        RECT 0.000 3136.400 197.865 3138.130 ;
        RECT 3390.135 3136.870 3588.000 3138.600 ;
        RECT 3403.035 3136.630 3406.285 3136.870 ;
        RECT 0.000 3070.500 31.390 3136.400 ;
        RECT 97.040 3070.500 197.865 3136.400 ;
        RECT 0.000 3063.870 197.865 3070.500 ;
        RECT 0.000 3061.000 103.415 3063.870 ;
        RECT 181.715 3063.565 184.965 3063.870 ;
      LAYER met5 ;
        RECT 0.000 2925.000 24.215 3061.000 ;
      LAYER met5 ;
        RECT 0.000 2922.130 103.415 2925.000 ;
      LAYER met5 ;
        RECT 105.015 2923.730 129.965 3062.270 ;
        RECT 131.565 2923.730 135.815 3062.270 ;
        RECT 137.415 2923.730 141.665 3062.270 ;
        RECT 143.265 2923.730 152.265 3062.270 ;
        RECT 153.865 2923.730 158.315 3062.270 ;
        RECT 159.915 3061.000 163.160 3062.270 ;
        RECT 159.915 2925.000 163.165 3061.000 ;
        RECT 159.915 2923.730 163.160 2925.000 ;
        RECT 164.765 2923.730 168.015 3062.270 ;
        RECT 169.615 2923.730 174.065 3062.270 ;
        RECT 175.665 2923.730 180.115 3062.270 ;
        RECT 181.715 2923.970 184.965 3061.965 ;
        RECT 186.565 2923.730 191.015 3062.270 ;
        RECT 192.615 2923.730 197.865 3062.270 ;
        RECT 3390.135 2990.730 3395.385 3135.270 ;
        RECT 3396.985 2990.730 3401.435 3135.270 ;
        RECT 3403.035 2991.035 3406.285 3135.030 ;
        RECT 3407.885 2990.730 3412.335 3135.270 ;
        RECT 3413.935 2990.730 3418.385 3135.270 ;
        RECT 3419.985 2990.730 3423.235 3135.270 ;
        RECT 3424.840 3134.000 3428.085 3135.270 ;
        RECT 3424.835 2992.000 3428.085 3134.000 ;
        RECT 3424.840 2990.730 3428.085 2992.000 ;
        RECT 3429.685 2990.730 3434.135 3135.270 ;
        RECT 3435.735 2990.730 3444.735 3135.270 ;
        RECT 3446.335 2990.730 3450.585 3135.270 ;
        RECT 3452.185 2990.730 3456.435 3135.270 ;
        RECT 3458.035 2990.730 3482.985 3135.270 ;
      LAYER met5 ;
        RECT 3484.585 3134.000 3588.000 3136.870 ;
      LAYER met5 ;
        RECT 3563.785 2992.000 3588.000 3134.000 ;
      LAYER met5 ;
        RECT 3403.035 2989.130 3406.285 2989.435 ;
        RECT 3484.585 2989.130 3588.000 2992.000 ;
        RECT 3390.135 2982.500 3588.000 2989.130 ;
        RECT 181.715 2922.130 184.965 2922.370 ;
        RECT 0.000 2920.400 197.865 2922.130 ;
        RECT 0.000 2854.500 31.390 2920.400 ;
        RECT 97.040 2854.500 197.865 2920.400 ;
        RECT 3390.135 2916.600 3490.960 2982.500 ;
        RECT 3556.610 2916.600 3588.000 2982.500 ;
        RECT 3390.135 2914.870 3588.000 2916.600 ;
        RECT 3403.035 2914.630 3406.285 2914.870 ;
        RECT 0.000 2847.870 197.865 2854.500 ;
        RECT 0.000 2845.000 103.415 2847.870 ;
        RECT 181.715 2847.565 184.965 2847.870 ;
      LAYER met5 ;
        RECT 0.000 2709.000 24.215 2845.000 ;
      LAYER met5 ;
        RECT 0.000 2706.130 103.415 2709.000 ;
      LAYER met5 ;
        RECT 105.015 2707.730 129.965 2846.270 ;
        RECT 131.565 2707.730 135.815 2846.270 ;
        RECT 137.415 2707.730 141.665 2846.270 ;
        RECT 143.265 2707.730 152.265 2846.270 ;
        RECT 153.865 2707.730 158.315 2846.270 ;
        RECT 159.915 2845.000 163.160 2846.270 ;
        RECT 159.915 2709.000 163.165 2845.000 ;
        RECT 159.915 2707.730 163.160 2709.000 ;
        RECT 164.765 2707.730 168.015 2846.270 ;
        RECT 169.615 2707.730 174.065 2846.270 ;
        RECT 175.665 2707.730 180.115 2846.270 ;
        RECT 181.715 2707.970 184.965 2845.965 ;
        RECT 186.565 2707.730 191.015 2846.270 ;
        RECT 192.615 2707.730 197.865 2846.270 ;
        RECT 3390.135 2769.730 3395.385 2913.270 ;
        RECT 3396.985 2769.730 3401.435 2913.270 ;
        RECT 3403.035 2770.035 3406.285 2913.030 ;
        RECT 3407.885 2769.730 3412.335 2913.270 ;
        RECT 3413.935 2769.730 3418.385 2913.270 ;
        RECT 3419.985 2769.730 3423.235 2913.270 ;
        RECT 3424.840 2912.000 3428.085 2913.270 ;
        RECT 3424.835 2771.000 3428.085 2912.000 ;
        RECT 3424.840 2769.730 3428.085 2771.000 ;
        RECT 3429.685 2769.730 3434.135 2913.270 ;
        RECT 3435.735 2769.730 3444.735 2913.270 ;
        RECT 3446.335 2769.730 3450.585 2913.270 ;
        RECT 3452.185 2769.730 3456.435 2913.270 ;
        RECT 3458.035 2769.730 3482.985 2913.270 ;
      LAYER met5 ;
        RECT 3484.585 2912.000 3588.000 2914.870 ;
      LAYER met5 ;
        RECT 3563.785 2771.000 3588.000 2912.000 ;
      LAYER met5 ;
        RECT 3403.035 2768.130 3406.285 2768.435 ;
        RECT 3484.585 2768.130 3588.000 2771.000 ;
        RECT 3390.135 2761.500 3588.000 2768.130 ;
        RECT 181.715 2706.130 184.965 2706.370 ;
        RECT 0.000 2704.400 197.865 2706.130 ;
        RECT 0.000 2638.500 31.390 2704.400 ;
        RECT 97.040 2638.500 197.865 2704.400 ;
        RECT 3390.135 2695.600 3490.960 2761.500 ;
        RECT 3556.610 2695.600 3588.000 2761.500 ;
        RECT 3390.135 2693.870 3588.000 2695.600 ;
        RECT 3403.035 2693.630 3406.285 2693.870 ;
        RECT 0.000 2631.870 197.865 2638.500 ;
        RECT 0.000 2629.000 103.415 2631.870 ;
        RECT 181.715 2631.565 184.965 2631.870 ;
      LAYER met5 ;
        RECT 0.000 2492.000 24.215 2629.000 ;
      LAYER met5 ;
        RECT 0.000 2489.130 103.415 2492.000 ;
      LAYER met5 ;
        RECT 105.015 2490.730 129.965 2630.270 ;
        RECT 131.565 2490.730 135.815 2630.270 ;
        RECT 137.415 2490.730 141.665 2630.270 ;
        RECT 143.265 2490.730 152.265 2630.270 ;
        RECT 153.865 2490.730 158.315 2630.270 ;
        RECT 159.915 2629.000 163.160 2630.270 ;
        RECT 159.915 2492.000 163.165 2629.000 ;
        RECT 159.915 2490.730 163.160 2492.000 ;
      LAYER met5 ;
        RECT 163.160 2489.130 163.165 2492.000 ;
      LAYER met5 ;
        RECT 164.765 2490.730 168.015 2630.270 ;
        RECT 169.615 2490.730 174.065 2630.270 ;
        RECT 175.665 2490.730 180.115 2630.270 ;
        RECT 181.715 2491.035 184.965 2629.965 ;
        RECT 186.565 2490.730 191.015 2630.270 ;
        RECT 192.615 2490.730 197.865 2630.270 ;
        RECT 3390.135 2548.730 3395.385 2692.270 ;
        RECT 3396.985 2548.730 3401.435 2692.270 ;
        RECT 3403.035 2549.035 3406.285 2692.030 ;
        RECT 3407.885 2548.730 3412.335 2692.270 ;
        RECT 3413.935 2548.730 3418.385 2692.270 ;
        RECT 3419.985 2548.730 3423.235 2692.270 ;
        RECT 3424.840 2691.000 3428.085 2692.270 ;
        RECT 3424.835 2550.000 3428.085 2691.000 ;
      LAYER met5 ;
        RECT 3403.035 2547.130 3406.285 2547.435 ;
        RECT 3424.835 2547.130 3424.840 2550.000 ;
      LAYER met5 ;
        RECT 3424.840 2548.730 3428.085 2550.000 ;
        RECT 3429.685 2548.730 3434.135 2692.270 ;
        RECT 3435.735 2548.730 3444.735 2692.270 ;
        RECT 3446.335 2548.730 3450.585 2692.270 ;
        RECT 3452.185 2548.730 3456.435 2692.270 ;
        RECT 3458.035 2548.730 3482.985 2692.270 ;
      LAYER met5 ;
        RECT 3484.585 2691.000 3588.000 2693.870 ;
      LAYER met5 ;
        RECT 3563.785 2550.000 3588.000 2691.000 ;
      LAYER met5 ;
        RECT 3484.585 2547.130 3588.000 2550.000 ;
        RECT 3390.135 2544.550 3588.000 2547.130 ;
        RECT 181.715 2489.130 184.965 2489.435 ;
        RECT 0.000 2486.490 197.865 2489.130 ;
        RECT 0.000 2422.450 32.455 2486.490 ;
        RECT 96.480 2422.450 197.865 2486.490 ;
        RECT 3390.135 2480.510 3491.520 2544.550 ;
        RECT 3555.545 2480.510 3588.000 2544.550 ;
        RECT 3390.135 2477.870 3588.000 2480.510 ;
        RECT 3403.035 2477.565 3406.285 2477.870 ;
        RECT 0.000 2419.870 197.865 2422.450 ;
        RECT 0.000 2417.000 103.415 2419.870 ;
      LAYER met5 ;
        RECT 0.000 2281.000 24.215 2417.000 ;
      LAYER met5 ;
        RECT 0.000 2278.130 103.415 2281.000 ;
      LAYER met5 ;
        RECT 105.015 2279.730 129.965 2418.270 ;
        RECT 131.565 2279.730 135.815 2418.270 ;
        RECT 137.415 2279.730 141.665 2418.270 ;
        RECT 143.265 2279.730 152.265 2418.270 ;
        RECT 153.865 2279.730 158.315 2418.270 ;
        RECT 159.915 2417.000 163.160 2418.270 ;
      LAYER met5 ;
        RECT 163.160 2417.000 163.165 2419.870 ;
        RECT 181.715 2419.565 184.965 2419.870 ;
      LAYER met5 ;
        RECT 159.915 2281.000 163.165 2417.000 ;
        RECT 159.915 2279.730 163.160 2281.000 ;
        RECT 164.765 2279.730 168.015 2418.270 ;
        RECT 169.615 2279.730 174.065 2418.270 ;
        RECT 175.665 2279.730 180.115 2418.270 ;
        RECT 181.715 2280.035 184.965 2417.965 ;
        RECT 186.565 2279.730 191.015 2418.270 ;
        RECT 192.615 2279.730 197.865 2418.270 ;
        RECT 3390.135 2331.730 3395.385 2476.270 ;
        RECT 3396.985 2331.730 3401.435 2476.270 ;
        RECT 3403.035 2332.035 3406.285 2475.965 ;
        RECT 3407.885 2331.730 3412.335 2476.270 ;
        RECT 3413.935 2331.730 3418.385 2476.270 ;
        RECT 3419.985 2331.730 3423.235 2476.270 ;
      LAYER met5 ;
        RECT 3424.835 2475.000 3424.840 2477.870 ;
      LAYER met5 ;
        RECT 3424.840 2475.000 3428.085 2476.270 ;
        RECT 3424.835 2333.000 3428.085 2475.000 ;
        RECT 3424.840 2331.730 3428.085 2333.000 ;
        RECT 3429.685 2331.730 3434.135 2476.270 ;
        RECT 3435.735 2331.730 3444.735 2476.270 ;
        RECT 3446.335 2331.730 3450.585 2476.270 ;
        RECT 3452.185 2331.730 3456.435 2476.270 ;
        RECT 3458.035 2331.730 3482.985 2476.270 ;
      LAYER met5 ;
        RECT 3484.585 2475.000 3588.000 2477.870 ;
      LAYER met5 ;
        RECT 3563.785 2333.000 3588.000 2475.000 ;
      LAYER met5 ;
        RECT 3403.035 2330.130 3406.285 2330.435 ;
        RECT 3484.585 2330.130 3588.000 2333.000 ;
        RECT 3390.135 2324.330 3588.000 2330.130 ;
        RECT 181.715 2278.130 184.965 2278.435 ;
        RECT 0.000 2272.270 197.865 2278.130 ;
        RECT 0.000 2214.670 29.235 2272.270 ;
        RECT 99.700 2214.670 197.865 2272.270 ;
        RECT 3390.135 2266.730 3488.300 2324.330 ;
        RECT 3558.765 2266.730 3588.000 2324.330 ;
        RECT 3390.135 2260.870 3588.000 2266.730 ;
        RECT 3403.035 2260.565 3406.285 2260.870 ;
        RECT 0.000 2208.870 197.865 2214.670 ;
        RECT 0.000 2206.000 103.415 2208.870 ;
        RECT 181.715 2208.565 184.965 2208.870 ;
      LAYER met5 ;
        RECT 0.000 2070.000 24.215 2206.000 ;
      LAYER met5 ;
        RECT 0.000 2067.130 103.415 2070.000 ;
      LAYER met5 ;
        RECT 105.015 2068.730 129.965 2207.270 ;
        RECT 131.565 2068.730 135.815 2207.270 ;
        RECT 137.415 2068.730 141.665 2207.270 ;
        RECT 143.265 2068.730 152.265 2207.270 ;
        RECT 153.865 2068.730 158.315 2207.270 ;
        RECT 159.915 2206.000 163.160 2207.270 ;
        RECT 159.915 2070.000 163.165 2206.000 ;
        RECT 159.915 2068.730 163.160 2070.000 ;
        RECT 164.765 2068.730 168.015 2207.270 ;
        RECT 169.615 2068.730 174.065 2207.270 ;
        RECT 175.665 2068.730 180.115 2207.270 ;
        RECT 181.715 2068.970 184.965 2206.965 ;
        RECT 186.565 2068.730 191.015 2207.270 ;
        RECT 192.615 2068.730 197.865 2207.270 ;
        RECT 3390.135 2115.730 3395.385 2259.270 ;
        RECT 3396.985 2115.730 3401.435 2259.270 ;
        RECT 3403.035 2116.035 3406.285 2258.965 ;
        RECT 3407.885 2115.730 3412.335 2259.270 ;
        RECT 3413.935 2115.730 3418.385 2259.270 ;
        RECT 3419.985 2115.730 3423.235 2259.270 ;
        RECT 3424.840 2258.000 3428.085 2259.270 ;
        RECT 3424.835 2117.000 3428.085 2258.000 ;
      LAYER met5 ;
        RECT 3403.035 2114.130 3406.285 2114.435 ;
        RECT 3424.835 2114.130 3424.840 2117.000 ;
      LAYER met5 ;
        RECT 3424.840 2115.730 3428.085 2117.000 ;
        RECT 3429.685 2115.730 3434.135 2259.270 ;
        RECT 3435.735 2115.730 3444.735 2259.270 ;
        RECT 3446.335 2115.730 3450.585 2259.270 ;
        RECT 3452.185 2115.730 3456.435 2259.270 ;
        RECT 3458.035 2115.730 3482.985 2259.270 ;
      LAYER met5 ;
        RECT 3484.585 2258.000 3588.000 2260.870 ;
      LAYER met5 ;
        RECT 3563.785 2117.000 3588.000 2258.000 ;
      LAYER met5 ;
        RECT 3484.585 2114.130 3588.000 2117.000 ;
        RECT 3390.135 2111.550 3588.000 2114.130 ;
        RECT 181.715 2067.130 184.965 2067.370 ;
        RECT 0.000 2065.400 197.865 2067.130 ;
        RECT 0.000 1999.500 31.390 2065.400 ;
        RECT 97.040 1999.500 197.865 2065.400 ;
        RECT 3390.135 2047.510 3491.520 2111.550 ;
        RECT 3555.545 2047.510 3588.000 2111.550 ;
        RECT 3390.135 2044.870 3588.000 2047.510 ;
        RECT 3403.035 2044.565 3406.285 2044.870 ;
        RECT 0.000 1992.870 197.865 1999.500 ;
        RECT 0.000 1990.000 103.415 1992.870 ;
        RECT 181.715 1992.565 184.965 1992.870 ;
      LAYER met5 ;
        RECT 0.000 1854.000 24.215 1990.000 ;
      LAYER met5 ;
        RECT 0.000 1851.130 103.415 1854.000 ;
      LAYER met5 ;
        RECT 105.015 1852.730 129.965 1991.270 ;
        RECT 131.565 1852.730 135.815 1991.270 ;
        RECT 137.415 1852.730 141.665 1991.270 ;
        RECT 143.265 1852.730 152.265 1991.270 ;
        RECT 153.865 1852.730 158.315 1991.270 ;
        RECT 159.915 1990.000 163.160 1991.270 ;
        RECT 159.915 1854.000 163.165 1990.000 ;
        RECT 159.915 1852.730 163.160 1854.000 ;
        RECT 164.765 1852.730 168.015 1991.270 ;
        RECT 169.615 1852.730 174.065 1991.270 ;
        RECT 175.665 1852.730 180.115 1991.270 ;
        RECT 181.715 1852.970 184.965 1990.965 ;
        RECT 186.565 1852.730 191.015 1991.270 ;
        RECT 192.615 1852.730 197.865 1991.270 ;
        RECT 3390.135 1898.730 3395.385 2043.270 ;
        RECT 3396.985 1898.730 3401.435 2043.270 ;
        RECT 3403.035 1899.035 3406.285 2042.965 ;
        RECT 3407.885 1898.730 3412.335 2043.270 ;
        RECT 3413.935 1898.730 3418.385 2043.270 ;
        RECT 3419.985 1898.730 3423.235 2043.270 ;
      LAYER met5 ;
        RECT 3424.835 2042.000 3424.840 2044.870 ;
      LAYER met5 ;
        RECT 3424.840 2042.000 3428.085 2043.270 ;
        RECT 3424.835 1900.000 3428.085 2042.000 ;
        RECT 3424.840 1898.730 3428.085 1900.000 ;
        RECT 3429.685 1898.730 3434.135 2043.270 ;
        RECT 3435.735 1898.730 3444.735 2043.270 ;
        RECT 3446.335 1898.730 3450.585 2043.270 ;
        RECT 3452.185 1898.730 3456.435 2043.270 ;
        RECT 3458.035 1898.730 3482.985 2043.270 ;
      LAYER met5 ;
        RECT 3484.585 2042.000 3588.000 2044.870 ;
      LAYER met5 ;
        RECT 3563.785 1900.000 3588.000 2042.000 ;
      LAYER met5 ;
        RECT 3403.035 1897.130 3406.285 1897.435 ;
        RECT 3484.585 1897.130 3588.000 1900.000 ;
        RECT 3390.135 1890.500 3588.000 1897.130 ;
        RECT 181.715 1851.130 184.965 1851.370 ;
        RECT 0.000 1849.400 197.865 1851.130 ;
        RECT 0.000 1783.500 31.390 1849.400 ;
        RECT 97.040 1783.500 197.865 1849.400 ;
        RECT 3390.135 1824.600 3490.960 1890.500 ;
        RECT 3556.610 1824.600 3588.000 1890.500 ;
        RECT 3390.135 1822.870 3588.000 1824.600 ;
        RECT 3403.035 1822.630 3406.285 1822.870 ;
        RECT 0.000 1776.870 197.865 1783.500 ;
        RECT 0.000 1774.000 103.415 1776.870 ;
        RECT 181.715 1776.565 184.965 1776.870 ;
      LAYER met5 ;
        RECT 0.000 1637.000 24.215 1774.000 ;
      LAYER met5 ;
        RECT 0.000 1634.130 103.415 1637.000 ;
      LAYER met5 ;
        RECT 105.015 1635.730 129.965 1775.270 ;
        RECT 131.565 1635.730 135.815 1775.270 ;
        RECT 137.415 1635.730 141.665 1775.270 ;
        RECT 143.265 1635.730 152.265 1775.270 ;
        RECT 153.865 1635.730 158.315 1775.270 ;
        RECT 159.915 1774.000 163.160 1775.270 ;
        RECT 159.915 1637.000 163.165 1774.000 ;
        RECT 159.915 1635.730 163.160 1637.000 ;
        RECT 164.765 1635.730 168.015 1775.270 ;
        RECT 169.615 1635.730 174.065 1775.270 ;
        RECT 175.665 1635.730 180.115 1775.270 ;
        RECT 181.715 1635.970 184.965 1774.965 ;
        RECT 186.565 1635.730 191.015 1775.270 ;
        RECT 192.615 1635.730 197.865 1775.270 ;
        RECT 3390.135 1677.730 3395.385 1821.270 ;
        RECT 3396.985 1677.730 3401.435 1821.270 ;
        RECT 3403.035 1678.035 3406.285 1821.030 ;
        RECT 3407.885 1677.730 3412.335 1821.270 ;
        RECT 3413.935 1677.730 3418.385 1821.270 ;
        RECT 3419.985 1677.730 3423.235 1821.270 ;
        RECT 3424.840 1820.000 3428.085 1821.270 ;
        RECT 3424.835 1679.000 3428.085 1820.000 ;
        RECT 3424.840 1677.730 3428.085 1679.000 ;
        RECT 3429.685 1677.730 3434.135 1821.270 ;
        RECT 3435.735 1677.730 3444.735 1821.270 ;
        RECT 3446.335 1677.730 3450.585 1821.270 ;
        RECT 3452.185 1677.730 3456.435 1821.270 ;
        RECT 3458.035 1677.730 3482.985 1821.270 ;
      LAYER met5 ;
        RECT 3484.585 1820.000 3588.000 1822.870 ;
      LAYER met5 ;
        RECT 3563.785 1679.000 3588.000 1820.000 ;
      LAYER met5 ;
        RECT 3403.035 1676.130 3406.285 1676.435 ;
        RECT 3484.585 1676.130 3588.000 1679.000 ;
        RECT 3390.135 1669.500 3588.000 1676.130 ;
        RECT 181.715 1634.130 184.965 1634.370 ;
        RECT 0.000 1632.400 197.865 1634.130 ;
        RECT 0.000 1566.500 31.390 1632.400 ;
        RECT 97.040 1566.500 197.865 1632.400 ;
        RECT 3390.135 1603.600 3490.960 1669.500 ;
        RECT 3556.610 1603.600 3588.000 1669.500 ;
        RECT 3390.135 1601.870 3588.000 1603.600 ;
        RECT 3403.035 1601.630 3406.285 1601.870 ;
        RECT 0.000 1559.870 197.865 1566.500 ;
        RECT 0.000 1557.000 103.415 1559.870 ;
        RECT 181.715 1559.565 184.965 1559.870 ;
      LAYER met5 ;
        RECT 0.000 1421.000 24.215 1557.000 ;
      LAYER met5 ;
        RECT 0.000 1418.130 103.415 1421.000 ;
      LAYER met5 ;
        RECT 105.015 1419.730 129.965 1558.270 ;
        RECT 131.565 1419.730 135.815 1558.270 ;
        RECT 137.415 1419.730 141.665 1558.270 ;
        RECT 143.265 1419.730 152.265 1558.270 ;
        RECT 153.865 1419.730 158.315 1558.270 ;
        RECT 159.915 1557.000 163.160 1558.270 ;
        RECT 159.915 1421.000 163.165 1557.000 ;
        RECT 159.915 1419.730 163.160 1421.000 ;
        RECT 164.765 1419.730 168.015 1558.270 ;
        RECT 169.615 1419.730 174.065 1558.270 ;
        RECT 175.665 1419.730 180.115 1558.270 ;
        RECT 181.715 1419.970 184.965 1557.965 ;
        RECT 186.565 1419.730 191.015 1558.270 ;
        RECT 192.615 1419.730 197.865 1558.270 ;
        RECT 3390.135 1456.730 3395.385 1600.270 ;
        RECT 3396.985 1456.730 3401.435 1600.270 ;
        RECT 3403.035 1457.035 3406.285 1600.030 ;
        RECT 3407.885 1456.730 3412.335 1600.270 ;
        RECT 3413.935 1456.730 3418.385 1600.270 ;
        RECT 3419.985 1456.730 3423.235 1600.270 ;
        RECT 3424.840 1599.000 3428.085 1600.270 ;
        RECT 3424.835 1458.000 3428.085 1599.000 ;
        RECT 3424.840 1456.730 3428.085 1458.000 ;
        RECT 3429.685 1456.730 3434.135 1600.270 ;
        RECT 3435.735 1456.730 3444.735 1600.270 ;
        RECT 3446.335 1456.730 3450.585 1600.270 ;
        RECT 3452.185 1456.730 3456.435 1600.270 ;
        RECT 3458.035 1456.730 3482.985 1600.270 ;
      LAYER met5 ;
        RECT 3484.585 1599.000 3588.000 1601.870 ;
      LAYER met5 ;
        RECT 3563.785 1458.000 3588.000 1599.000 ;
      LAYER met5 ;
        RECT 3403.035 1455.130 3406.285 1455.435 ;
        RECT 3484.585 1455.130 3588.000 1458.000 ;
        RECT 3390.135 1448.500 3588.000 1455.130 ;
        RECT 181.715 1418.130 184.965 1418.370 ;
        RECT 0.000 1416.400 197.865 1418.130 ;
        RECT 0.000 1350.500 31.390 1416.400 ;
        RECT 97.040 1350.500 197.865 1416.400 ;
        RECT 3390.135 1382.600 3490.960 1448.500 ;
        RECT 3556.610 1382.600 3588.000 1448.500 ;
        RECT 3390.135 1380.870 3588.000 1382.600 ;
        RECT 3403.035 1380.630 3406.285 1380.870 ;
        RECT 0.000 1343.870 197.865 1350.500 ;
        RECT 0.000 1341.000 103.415 1343.870 ;
        RECT 181.715 1343.565 184.965 1343.870 ;
      LAYER met5 ;
        RECT 0.000 1205.000 24.215 1341.000 ;
      LAYER met5 ;
        RECT 0.000 1202.130 103.415 1205.000 ;
      LAYER met5 ;
        RECT 105.015 1203.730 129.965 1342.270 ;
        RECT 131.565 1203.730 135.815 1342.270 ;
        RECT 137.415 1203.730 141.665 1342.270 ;
        RECT 143.265 1203.730 152.265 1342.270 ;
        RECT 153.865 1203.730 158.315 1342.270 ;
        RECT 159.915 1341.000 163.160 1342.270 ;
        RECT 159.915 1205.000 163.165 1341.000 ;
        RECT 159.915 1203.730 163.160 1205.000 ;
        RECT 164.765 1203.730 168.015 1342.270 ;
        RECT 169.615 1203.730 174.065 1342.270 ;
        RECT 175.665 1203.730 180.115 1342.270 ;
        RECT 181.715 1203.970 184.965 1341.965 ;
        RECT 186.565 1203.730 191.015 1342.270 ;
        RECT 192.615 1203.730 197.865 1342.270 ;
        RECT 3390.135 1234.730 3395.385 1379.270 ;
        RECT 3396.985 1234.730 3401.435 1379.270 ;
        RECT 3403.035 1235.035 3406.285 1379.030 ;
        RECT 3407.885 1234.730 3412.335 1379.270 ;
        RECT 3413.935 1234.730 3418.385 1379.270 ;
        RECT 3419.985 1234.730 3423.235 1379.270 ;
        RECT 3424.840 1378.000 3428.085 1379.270 ;
        RECT 3424.835 1236.000 3428.085 1378.000 ;
        RECT 3424.840 1234.730 3428.085 1236.000 ;
        RECT 3429.685 1234.730 3434.135 1379.270 ;
        RECT 3435.735 1234.730 3444.735 1379.270 ;
        RECT 3446.335 1234.730 3450.585 1379.270 ;
        RECT 3452.185 1234.730 3456.435 1379.270 ;
        RECT 3458.035 1234.730 3482.985 1379.270 ;
      LAYER met5 ;
        RECT 3484.585 1378.000 3588.000 1380.870 ;
      LAYER met5 ;
        RECT 3563.785 1236.000 3588.000 1378.000 ;
      LAYER met5 ;
        RECT 3403.035 1233.130 3406.285 1233.435 ;
        RECT 3484.585 1233.130 3588.000 1236.000 ;
        RECT 3390.135 1226.500 3588.000 1233.130 ;
        RECT 181.715 1202.130 184.965 1202.370 ;
        RECT 0.000 1200.400 197.865 1202.130 ;
        RECT 0.000 1134.500 31.390 1200.400 ;
        RECT 97.040 1134.500 197.865 1200.400 ;
        RECT 3390.135 1160.600 3490.960 1226.500 ;
        RECT 3556.610 1160.600 3588.000 1226.500 ;
        RECT 3390.135 1158.870 3588.000 1160.600 ;
        RECT 3403.035 1158.630 3406.285 1158.870 ;
        RECT 0.000 1127.870 197.865 1134.500 ;
        RECT 0.000 1125.000 103.415 1127.870 ;
        RECT 181.715 1127.565 184.965 1127.870 ;
      LAYER met5 ;
        RECT 0.000 989.000 24.215 1125.000 ;
      LAYER met5 ;
        RECT 0.000 986.130 103.415 989.000 ;
      LAYER met5 ;
        RECT 105.015 987.730 129.965 1126.270 ;
        RECT 131.565 987.730 135.815 1126.270 ;
        RECT 137.415 987.730 141.665 1126.270 ;
        RECT 143.265 987.730 152.265 1126.270 ;
        RECT 153.865 987.730 158.315 1126.270 ;
        RECT 159.915 1125.000 163.160 1126.270 ;
        RECT 159.915 989.000 163.165 1125.000 ;
        RECT 159.915 987.730 163.160 989.000 ;
        RECT 164.765 987.730 168.015 1126.270 ;
        RECT 169.615 987.730 174.065 1126.270 ;
        RECT 175.665 987.730 180.115 1126.270 ;
        RECT 181.715 987.970 184.965 1125.965 ;
        RECT 186.565 987.730 191.015 1126.270 ;
        RECT 192.615 987.730 197.865 1126.270 ;
        RECT 3390.135 1013.730 3395.385 1157.270 ;
        RECT 3396.985 1013.730 3401.435 1157.270 ;
        RECT 3403.035 1014.035 3406.285 1157.030 ;
        RECT 3407.885 1013.730 3412.335 1157.270 ;
        RECT 3413.935 1013.730 3418.385 1157.270 ;
        RECT 3419.985 1013.730 3423.235 1157.270 ;
        RECT 3424.840 1156.000 3428.085 1157.270 ;
        RECT 3424.835 1015.000 3428.085 1156.000 ;
        RECT 3424.840 1013.730 3428.085 1015.000 ;
        RECT 3429.685 1013.730 3434.135 1157.270 ;
        RECT 3435.735 1013.730 3444.735 1157.270 ;
        RECT 3446.335 1013.730 3450.585 1157.270 ;
        RECT 3452.185 1013.730 3456.435 1157.270 ;
        RECT 3458.035 1013.730 3482.985 1157.270 ;
      LAYER met5 ;
        RECT 3484.585 1156.000 3588.000 1158.870 ;
      LAYER met5 ;
        RECT 3563.785 1015.000 3588.000 1156.000 ;
      LAYER met5 ;
        RECT 3403.035 1012.130 3406.285 1012.435 ;
        RECT 3484.585 1012.130 3588.000 1015.000 ;
        RECT 3390.135 1005.500 3588.000 1012.130 ;
        RECT 181.715 986.130 184.965 986.370 ;
        RECT 0.000 984.400 197.865 986.130 ;
        RECT 0.000 918.500 31.390 984.400 ;
        RECT 97.040 918.500 197.865 984.400 ;
        RECT 3390.135 939.600 3490.960 1005.500 ;
        RECT 3556.610 939.600 3588.000 1005.500 ;
        RECT 3390.135 937.870 3588.000 939.600 ;
        RECT 3403.035 937.630 3406.285 937.870 ;
        RECT 0.000 911.870 197.865 918.500 ;
        RECT 0.000 909.000 103.415 911.870 ;
        RECT 181.715 911.565 184.965 911.870 ;
      LAYER met5 ;
        RECT 0.000 626.000 24.215 909.000 ;
      LAYER met5 ;
        RECT 0.000 623.130 103.415 626.000 ;
      LAYER met5 ;
        RECT 105.015 624.730 129.965 910.270 ;
        RECT 131.565 624.730 135.815 910.270 ;
        RECT 137.415 624.730 141.665 910.270 ;
        RECT 143.265 767.000 152.265 910.270 ;
        RECT 153.865 772.000 158.315 910.270 ;
        RECT 159.915 909.000 163.160 910.270 ;
        RECT 159.915 767.000 163.165 909.000 ;
        RECT 143.265 624.730 152.265 762.000 ;
        RECT 153.865 624.730 158.315 767.000 ;
        RECT 159.915 626.000 163.165 762.000 ;
        RECT 159.915 624.730 163.160 626.000 ;
      LAYER met5 ;
        RECT 163.160 623.130 163.165 626.000 ;
      LAYER met5 ;
        RECT 164.765 624.730 168.015 910.270 ;
        RECT 169.615 624.730 174.065 910.270 ;
        RECT 175.665 624.730 180.115 910.270 ;
        RECT 181.715 767.000 184.965 909.965 ;
        RECT 186.565 772.000 191.015 910.270 ;
        RECT 181.715 625.035 184.965 762.000 ;
        RECT 186.565 624.730 191.015 767.000 ;
        RECT 192.615 624.730 197.865 910.270 ;
        RECT 3390.135 792.730 3395.385 936.270 ;
        RECT 3396.985 792.730 3401.435 936.270 ;
        RECT 3403.035 793.035 3406.285 936.030 ;
        RECT 3407.885 792.730 3412.335 936.270 ;
        RECT 3413.935 792.730 3418.385 936.270 ;
        RECT 3419.985 792.730 3423.235 936.270 ;
        RECT 3424.840 935.000 3428.085 936.270 ;
        RECT 3424.835 794.000 3428.085 935.000 ;
        RECT 3424.840 792.730 3428.085 794.000 ;
        RECT 3429.685 792.730 3434.135 936.270 ;
        RECT 3435.735 792.730 3444.735 936.270 ;
        RECT 3446.335 792.730 3450.585 936.270 ;
        RECT 3452.185 792.730 3456.435 936.270 ;
        RECT 3458.035 792.730 3482.985 936.270 ;
      LAYER met5 ;
        RECT 3484.585 935.000 3588.000 937.870 ;
      LAYER met5 ;
        RECT 3563.785 794.000 3588.000 935.000 ;
      LAYER met5 ;
        RECT 3403.035 791.130 3406.285 791.435 ;
        RECT 3484.585 791.130 3588.000 794.000 ;
        RECT 3390.135 784.500 3588.000 791.130 ;
        RECT 3390.135 718.600 3490.960 784.500 ;
        RECT 3556.610 718.600 3588.000 784.500 ;
        RECT 3390.135 716.870 3588.000 718.600 ;
        RECT 3403.035 716.630 3406.285 716.870 ;
        RECT 181.715 623.130 184.965 623.435 ;
        RECT 0.000 620.490 197.865 623.130 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 556.450 197.865 620.490 ;
      LAYER met5 ;
        RECT 3390.135 570.730 3395.385 715.270 ;
        RECT 3396.985 570.730 3401.435 715.270 ;
        RECT 3403.035 571.035 3406.285 715.030 ;
        RECT 3407.885 570.730 3412.335 715.270 ;
        RECT 3413.935 570.730 3418.385 715.270 ;
        RECT 3419.985 570.730 3423.235 715.270 ;
        RECT 3424.840 714.000 3428.085 715.270 ;
        RECT 3424.835 572.000 3428.085 714.000 ;
        RECT 3424.840 570.730 3428.085 572.000 ;
        RECT 3429.685 570.730 3434.135 715.270 ;
        RECT 3435.735 570.730 3444.735 715.270 ;
        RECT 3446.335 570.730 3450.585 715.270 ;
        RECT 3452.185 570.730 3456.435 715.270 ;
        RECT 3458.035 570.730 3482.985 715.270 ;
      LAYER met5 ;
        RECT 3484.585 714.000 3588.000 716.870 ;
      LAYER met5 ;
        RECT 3563.785 572.000 3588.000 714.000 ;
      LAYER met5 ;
        RECT 3403.035 569.130 3406.285 569.435 ;
        RECT 3484.585 569.130 3588.000 572.000 ;
        RECT 0.000 553.870 197.865 556.450 ;
        RECT 3390.135 562.500 3588.000 569.130 ;
        RECT 0.000 551.000 103.415 553.870 ;
      LAYER met5 ;
        RECT 0.000 415.000 24.215 551.000 ;
      LAYER met5 ;
        RECT 0.000 412.130 103.415 415.000 ;
      LAYER met5 ;
        RECT 105.015 413.730 129.965 552.270 ;
        RECT 131.565 413.730 135.815 552.270 ;
        RECT 137.415 413.730 141.665 552.270 ;
        RECT 143.265 413.730 152.265 552.270 ;
        RECT 153.865 413.730 158.315 552.270 ;
        RECT 159.915 551.000 163.160 552.270 ;
      LAYER met5 ;
        RECT 163.160 551.000 163.165 553.870 ;
        RECT 181.715 553.565 184.965 553.870 ;
      LAYER met5 ;
        RECT 159.915 415.000 163.165 551.000 ;
        RECT 159.915 413.730 163.160 415.000 ;
      LAYER met5 ;
        RECT 163.160 412.130 163.165 415.000 ;
      LAYER met5 ;
        RECT 164.765 413.730 168.015 552.270 ;
        RECT 169.615 413.730 174.065 552.270 ;
        RECT 175.665 413.730 180.115 552.270 ;
        RECT 181.715 414.035 184.965 551.965 ;
        RECT 186.565 413.730 191.015 552.270 ;
        RECT 192.615 413.730 197.865 552.270 ;
      LAYER met5 ;
        RECT 3390.135 496.600 3490.960 562.500 ;
        RECT 3556.610 496.600 3588.000 562.500 ;
        RECT 3390.135 494.870 3588.000 496.600 ;
        RECT 3403.035 494.630 3406.285 494.870 ;
        RECT 181.715 412.130 184.965 412.435 ;
        RECT 0.000 406.270 197.865 412.130 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 197.865 406.270 ;
        RECT 0.000 342.870 197.865 348.670 ;
        RECT 0.000 340.000 103.415 342.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 340.000 ;
      LAYER met5 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 341.270 ;
        RECT 131.565 202.730 135.815 341.270 ;
        RECT 137.415 202.730 141.665 341.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 341.270 ;
        RECT 153.865 202.730 158.315 341.270 ;
        RECT 159.915 340.000 163.160 341.270 ;
      LAYER met5 ;
        RECT 163.160 340.000 163.165 342.870 ;
        RECT 181.715 342.565 184.965 342.870 ;
      LAYER met5 ;
        RECT 159.915 204.000 163.165 340.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 341.270 ;
        RECT 169.615 202.730 174.065 341.270 ;
        RECT 175.665 202.730 180.115 341.270 ;
        RECT 181.715 202.745 184.965 340.965 ;
        RECT 186.565 202.730 191.015 341.270 ;
        RECT 192.615 202.730 197.865 341.270 ;
      LAYER met5 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
      LAYER met5 ;
        RECT 197.650 192.615 395.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 237.000 191.015 357.000 192.615 ;
        RECT 196.215 186.565 395.270 191.015 ;
      LAYER met5 ;
        RECT 396.870 184.965 466.130 197.865 ;
      LAYER met5 ;
        RECT 467.730 192.615 664.270 197.865 ;
        RECT 506.000 191.015 626.000 192.615 ;
        RECT 467.730 186.565 664.270 191.015 ;
      LAYER met5 ;
        RECT 665.870 184.965 735.130 197.865 ;
      LAYER met5 ;
        RECT 736.730 192.615 933.270 197.865 ;
        RECT 775.000 191.015 895.000 192.615 ;
        RECT 736.730 186.565 933.270 191.015 ;
      LAYER met5 ;
        RECT 934.870 184.965 1009.130 197.865 ;
      LAYER met5 ;
        RECT 1010.730 192.615 1207.270 197.865 ;
        RECT 1049.000 191.015 1169.000 192.615 ;
        RECT 1010.730 186.565 1207.270 191.015 ;
      LAYER met5 ;
        RECT 1208.870 184.965 1278.130 197.865 ;
      LAYER met5 ;
        RECT 1279.730 192.615 1476.270 197.865 ;
        RECT 1318.000 191.015 1438.000 192.615 ;
        RECT 1279.730 186.565 1476.270 191.015 ;
      LAYER met5 ;
        RECT 1477.870 184.965 1552.130 197.865 ;
      LAYER met5 ;
        RECT 1553.730 192.615 1750.270 197.865 ;
        RECT 1592.000 191.015 1712.000 192.615 ;
        RECT 1553.730 186.565 1750.270 191.015 ;
      LAYER met5 ;
        RECT 1751.870 184.965 1826.130 197.865 ;
      LAYER met5 ;
        RECT 1827.730 192.615 2024.270 197.865 ;
        RECT 1866.000 191.015 1986.000 192.615 ;
        RECT 1827.730 186.565 2024.270 191.015 ;
      LAYER met5 ;
        RECT 2025.870 184.965 2100.130 197.865 ;
      LAYER met5 ;
        RECT 2101.730 192.615 2298.270 197.865 ;
        RECT 2140.000 191.015 2260.000 192.615 ;
        RECT 2101.730 186.565 2298.270 191.015 ;
      LAYER met5 ;
        RECT 2299.870 184.965 2374.130 197.865 ;
      LAYER met5 ;
        RECT 2375.730 192.615 2572.270 197.865 ;
        RECT 2414.000 191.015 2534.000 192.615 ;
        RECT 2375.730 186.565 2572.270 191.015 ;
      LAYER met5 ;
        RECT 2573.870 184.965 2648.130 197.865 ;
      LAYER met5 ;
        RECT 2649.730 192.615 2846.270 197.865 ;
        RECT 2688.000 191.015 2808.000 192.615 ;
        RECT 2649.730 186.565 2846.270 191.015 ;
      LAYER met5 ;
        RECT 2847.870 184.965 2917.130 197.865 ;
      LAYER met5 ;
        RECT 2918.730 192.615 3115.270 197.865 ;
        RECT 2957.000 191.015 3077.000 192.615 ;
        RECT 2918.730 186.565 3115.270 191.015 ;
      LAYER met5 ;
        RECT 3116.870 184.965 3186.130 197.865 ;
      LAYER met5 ;
        RECT 3187.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 199.465 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 493.270 ;
        RECT 3396.985 351.000 3401.435 493.270 ;
        RECT 3403.035 346.000 3406.285 493.030 ;
        RECT 3396.985 196.215 3401.435 346.000 ;
        RECT 3403.035 198.530 3406.285 341.000 ;
        RECT 3407.885 198.475 3412.335 493.270 ;
        RECT 3413.935 198.400 3418.385 493.270 ;
        RECT 3419.985 198.615 3423.235 493.270 ;
        RECT 3424.840 492.000 3428.085 493.270 ;
        RECT 3424.835 346.000 3428.085 492.000 ;
        RECT 3429.685 351.000 3434.135 493.270 ;
        RECT 3435.735 346.000 3444.735 493.270 ;
        RECT 3424.835 198.665 3428.085 341.000 ;
        RECT 3429.685 198.525 3434.135 346.000 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 3226.000 191.015 3346.000 192.615 ;
        RECT 3187.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 394.965 184.965 ;
      LAYER met5 ;
        RECT 396.565 181.715 466.435 184.965 ;
      LAYER met5 ;
        RECT 468.035 181.715 663.965 184.965 ;
      LAYER met5 ;
        RECT 665.565 181.715 735.435 184.965 ;
      LAYER met5 ;
        RECT 737.035 181.715 933.030 184.965 ;
      LAYER met5 ;
        RECT 934.630 181.715 1009.435 184.965 ;
      LAYER met5 ;
        RECT 1011.035 181.715 1206.965 184.965 ;
      LAYER met5 ;
        RECT 1208.565 181.715 1278.435 184.965 ;
      LAYER met5 ;
        RECT 1280.035 181.715 1476.030 184.965 ;
      LAYER met5 ;
        RECT 1477.630 181.715 1552.435 184.965 ;
      LAYER met5 ;
        RECT 1554.035 181.715 1750.030 184.965 ;
      LAYER met5 ;
        RECT 1751.630 181.715 1826.435 184.965 ;
      LAYER met5 ;
        RECT 1828.035 181.715 2024.030 184.965 ;
      LAYER met5 ;
        RECT 2025.630 181.715 2100.435 184.965 ;
      LAYER met5 ;
        RECT 2102.035 181.715 2298.030 184.965 ;
      LAYER met5 ;
        RECT 2299.630 181.715 2374.435 184.965 ;
      LAYER met5 ;
        RECT 2376.035 181.715 2572.030 184.965 ;
      LAYER met5 ;
        RECT 2573.630 181.715 2648.435 184.965 ;
      LAYER met5 ;
        RECT 2650.035 181.715 2845.965 184.965 ;
      LAYER met5 ;
        RECT 2847.565 181.715 2917.435 184.965 ;
      LAYER met5 ;
        RECT 2919.035 181.715 3114.965 184.965 ;
      LAYER met5 ;
        RECT 3116.565 181.715 3186.435 184.965 ;
      LAYER met5 ;
        RECT 3188.035 181.715 3385.255 184.965 ;
      LAYER met5 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 395.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 395.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 395.270 168.015 ;
      LAYER met5 ;
        RECT 396.870 163.165 466.130 181.715 ;
      LAYER met5 ;
        RECT 467.730 175.665 664.270 180.115 ;
        RECT 467.730 169.615 664.270 174.065 ;
        RECT 467.730 164.765 664.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
      LAYER met5 ;
        RECT 198.665 163.160 394.000 163.165 ;
      LAYER met5 ;
        RECT 394.000 163.160 469.000 163.165 ;
      LAYER met5 ;
        RECT 469.000 163.160 663.000 163.165 ;
        RECT 198.665 159.915 395.270 163.160 ;
      LAYER met5 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 395.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
      LAYER met5 ;
        RECT 176.845 143.265 395.270 152.265 ;
      LAYER met5 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 395.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 395.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 395.270 129.965 ;
      LAYER met5 ;
        RECT 396.870 103.415 466.130 163.160 ;
      LAYER met5 ;
        RECT 467.730 159.915 664.270 163.160 ;
        RECT 467.730 153.865 664.270 158.315 ;
        RECT 467.730 143.265 664.270 152.265 ;
        RECT 467.730 137.415 664.270 141.665 ;
        RECT 467.730 131.565 664.270 135.815 ;
        RECT 467.730 105.015 664.270 129.965 ;
      LAYER met5 ;
        RECT 665.870 103.415 735.130 181.715 ;
      LAYER met5 ;
        RECT 736.730 175.665 933.270 180.115 ;
        RECT 736.730 169.615 933.270 174.065 ;
        RECT 736.730 164.765 933.270 168.015 ;
        RECT 738.000 163.160 932.000 163.165 ;
        RECT 736.730 159.915 933.270 163.160 ;
        RECT 736.730 153.865 933.270 158.315 ;
        RECT 736.730 143.265 933.270 152.265 ;
        RECT 736.730 137.415 933.270 141.665 ;
        RECT 736.730 131.565 933.270 135.815 ;
        RECT 736.730 105.015 933.270 129.965 ;
      LAYER met5 ;
        RECT 934.870 103.415 1009.130 181.715 ;
      LAYER met5 ;
        RECT 1010.730 175.665 1207.270 180.115 ;
        RECT 1010.730 169.615 1207.270 174.065 ;
        RECT 1010.730 164.765 1207.270 168.015 ;
      LAYER met5 ;
        RECT 1208.870 163.165 1278.130 181.715 ;
      LAYER met5 ;
        RECT 1279.730 175.665 1476.270 180.115 ;
        RECT 1279.730 169.615 1476.270 174.065 ;
        RECT 1279.730 164.765 1476.270 168.015 ;
        RECT 1012.000 163.160 1206.000 163.165 ;
      LAYER met5 ;
        RECT 1206.000 163.160 1281.000 163.165 ;
      LAYER met5 ;
        RECT 1281.000 163.160 1475.000 163.165 ;
        RECT 1010.730 159.915 1207.270 163.160 ;
        RECT 1010.730 153.865 1207.270 158.315 ;
        RECT 1010.730 143.265 1207.270 152.265 ;
        RECT 1010.730 137.415 1207.270 141.665 ;
        RECT 1010.730 131.565 1207.270 135.815 ;
        RECT 1010.730 105.015 1207.270 129.965 ;
      LAYER met5 ;
        RECT 1208.870 103.415 1278.130 163.160 ;
      LAYER met5 ;
        RECT 1279.730 159.915 1476.270 163.160 ;
        RECT 1279.730 153.865 1476.270 158.315 ;
        RECT 1279.730 143.265 1476.270 152.265 ;
        RECT 1279.730 137.415 1476.270 141.665 ;
        RECT 1279.730 131.565 1476.270 135.815 ;
        RECT 1279.730 105.015 1476.270 129.965 ;
      LAYER met5 ;
        RECT 1477.870 103.415 1552.130 181.715 ;
      LAYER met5 ;
        RECT 1553.730 175.665 1750.270 180.115 ;
        RECT 1553.730 169.615 1750.270 174.065 ;
        RECT 1553.730 164.765 1750.270 168.015 ;
        RECT 1555.000 163.160 1749.000 163.165 ;
        RECT 1553.730 159.915 1750.270 163.160 ;
        RECT 1553.730 153.865 1750.270 158.315 ;
        RECT 1553.730 143.265 1750.270 152.265 ;
        RECT 1553.730 137.415 1750.270 141.665 ;
        RECT 1553.730 131.565 1750.270 135.815 ;
        RECT 1553.730 105.015 1750.270 129.965 ;
      LAYER met5 ;
        RECT 1751.870 103.415 1826.130 181.715 ;
      LAYER met5 ;
        RECT 1827.730 175.665 2024.270 180.115 ;
        RECT 1827.730 169.615 2024.270 174.065 ;
        RECT 1827.730 164.765 2024.270 168.015 ;
        RECT 1829.000 163.160 2023.000 163.165 ;
        RECT 1827.730 159.915 2024.270 163.160 ;
        RECT 1827.730 153.865 2024.270 158.315 ;
        RECT 1827.730 143.265 2024.270 152.265 ;
        RECT 1827.730 137.415 2024.270 141.665 ;
        RECT 1827.730 131.565 2024.270 135.815 ;
        RECT 1827.730 105.015 2024.270 129.965 ;
      LAYER met5 ;
        RECT 2025.870 103.415 2100.130 181.715 ;
      LAYER met5 ;
        RECT 2101.730 175.665 2298.270 180.115 ;
        RECT 2101.730 169.615 2298.270 174.065 ;
        RECT 2101.730 164.765 2298.270 168.015 ;
        RECT 2103.000 163.160 2297.000 163.165 ;
        RECT 2101.730 159.915 2298.270 163.160 ;
        RECT 2101.730 153.865 2298.270 158.315 ;
        RECT 2101.730 143.265 2298.270 152.265 ;
        RECT 2101.730 137.415 2298.270 141.665 ;
        RECT 2101.730 131.565 2298.270 135.815 ;
        RECT 2101.730 105.015 2298.270 129.965 ;
      LAYER met5 ;
        RECT 2299.870 103.415 2374.130 181.715 ;
      LAYER met5 ;
        RECT 2375.730 175.665 2572.270 180.115 ;
        RECT 2375.730 169.615 2572.270 174.065 ;
        RECT 2375.730 164.765 2572.270 168.015 ;
        RECT 2377.000 163.160 2571.000 163.165 ;
        RECT 2375.730 159.915 2572.270 163.160 ;
        RECT 2375.730 153.865 2572.270 158.315 ;
        RECT 2375.730 143.265 2572.270 152.265 ;
        RECT 2375.730 137.415 2572.270 141.665 ;
        RECT 2375.730 131.565 2572.270 135.815 ;
        RECT 2375.730 105.015 2572.270 129.965 ;
      LAYER met5 ;
        RECT 2573.870 103.415 2648.130 181.715 ;
      LAYER met5 ;
        RECT 2649.730 175.665 2846.270 180.115 ;
        RECT 2649.730 169.615 2846.270 174.065 ;
        RECT 2649.730 164.765 2846.270 168.015 ;
      LAYER met5 ;
        RECT 2847.870 163.165 2917.130 181.715 ;
      LAYER met5 ;
        RECT 2918.730 175.665 3115.270 180.115 ;
        RECT 2918.730 169.615 3115.270 174.065 ;
        RECT 2918.730 164.765 3115.270 168.015 ;
      LAYER met5 ;
        RECT 3116.870 163.165 3186.130 181.715 ;
      LAYER met5 ;
        RECT 3187.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 341.000 ;
        RECT 3446.335 198.375 3450.585 493.270 ;
        RECT 3452.185 198.520 3456.435 493.270 ;
        RECT 3458.035 197.355 3482.985 493.270 ;
      LAYER met5 ;
        RECT 3484.585 492.000 3588.000 494.870 ;
      LAYER met5 ;
        RECT 3563.785 200.000 3588.000 492.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 3187.730 169.615 3385.270 174.065 ;
        RECT 3187.730 164.765 3385.270 168.015 ;
        RECT 2651.000 163.160 2845.000 163.165 ;
      LAYER met5 ;
        RECT 2845.000 163.160 2920.000 163.165 ;
      LAYER met5 ;
        RECT 2920.000 163.160 3114.000 163.165 ;
      LAYER met5 ;
        RECT 3114.000 163.160 3189.000 163.165 ;
      LAYER met5 ;
        RECT 3189.000 163.160 3384.000 163.165 ;
        RECT 2649.730 159.915 2846.270 163.160 ;
        RECT 2649.730 153.865 2846.270 158.315 ;
        RECT 2649.730 143.265 2846.270 152.265 ;
        RECT 2649.730 137.415 2846.270 141.665 ;
        RECT 2649.730 131.565 2846.270 135.815 ;
        RECT 2649.730 105.015 2846.270 129.965 ;
      LAYER met5 ;
        RECT 2847.870 103.415 2917.130 163.160 ;
      LAYER met5 ;
        RECT 2918.730 159.915 3115.270 163.160 ;
        RECT 2918.730 153.865 3115.270 158.315 ;
        RECT 2918.730 143.265 3115.270 152.265 ;
        RECT 2918.730 137.415 3115.270 141.665 ;
        RECT 2918.730 131.565 3115.270 135.815 ;
        RECT 2918.730 105.015 3115.270 129.965 ;
      LAYER met5 ;
        RECT 3116.870 103.415 3186.130 163.160 ;
      LAYER met5 ;
        RECT 3187.730 159.915 3385.270 163.160 ;
        RECT 3187.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 3187.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 3187.730 137.415 3385.270 141.665 ;
        RECT 3187.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 3187.730 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 394.000 96.480 469.000 103.415 ;
        RECT 394.000 32.455 399.510 96.480 ;
        RECT 463.550 32.455 469.000 96.480 ;
      LAYER met5 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met5 ;
        RECT 394.000 0.000 469.000 32.455 ;
        RECT 663.000 93.145 738.000 103.415 ;
        RECT 663.000 34.115 681.965 93.145 ;
        RECT 722.350 34.115 738.000 93.145 ;
        RECT 663.000 25.815 738.000 34.115 ;
        RECT 932.000 97.040 1012.000 103.415 ;
        RECT 932.000 31.390 936.600 97.040 ;
        RECT 1002.500 31.390 1012.000 97.040 ;
      LAYER met5 ;
        RECT 469.000 0.000 664.270 24.215 ;
      LAYER met5 ;
        RECT 665.870 0.000 735.130 25.815 ;
      LAYER met5 ;
        RECT 736.730 0.000 932.000 24.215 ;
      LAYER met5 ;
        RECT 932.000 0.000 1012.000 31.390 ;
        RECT 1206.000 99.700 1281.000 103.415 ;
        RECT 1206.000 29.235 1214.730 99.700 ;
        RECT 1272.330 29.235 1281.000 99.700 ;
      LAYER met5 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met5 ;
        RECT 1206.000 0.000 1281.000 29.235 ;
        RECT 1475.000 97.040 1555.000 103.415 ;
        RECT 1475.000 31.390 1479.600 97.040 ;
        RECT 1545.500 31.390 1555.000 97.040 ;
      LAYER met5 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met5 ;
        RECT 1475.000 0.000 1555.000 31.390 ;
        RECT 1749.000 97.040 1829.000 103.415 ;
        RECT 1749.000 31.390 1753.600 97.040 ;
        RECT 1819.500 31.390 1829.000 97.040 ;
      LAYER met5 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met5 ;
        RECT 1749.000 0.000 1829.000 31.390 ;
        RECT 2023.000 97.040 2103.000 103.415 ;
        RECT 2023.000 31.390 2027.600 97.040 ;
        RECT 2093.500 31.390 2103.000 97.040 ;
      LAYER met5 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met5 ;
        RECT 2023.000 0.000 2103.000 31.390 ;
        RECT 2297.000 97.040 2377.000 103.415 ;
        RECT 2297.000 31.390 2301.600 97.040 ;
        RECT 2367.500 31.390 2377.000 97.040 ;
      LAYER met5 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met5 ;
        RECT 2297.000 0.000 2377.000 31.390 ;
        RECT 2571.000 97.040 2651.000 103.415 ;
        RECT 2571.000 31.390 2575.600 97.040 ;
        RECT 2641.500 31.390 2651.000 97.040 ;
      LAYER met5 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met5 ;
        RECT 2571.000 0.000 2651.000 31.390 ;
        RECT 2845.000 96.480 2920.000 103.415 ;
        RECT 2845.000 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 2920.000 96.480 ;
      LAYER met5 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met5 ;
        RECT 2845.000 0.000 2920.000 32.455 ;
        RECT 3114.000 96.480 3189.000 103.415 ;
        RECT 3114.000 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3189.000 96.480 ;
      LAYER met5 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met5 ;
        RECT 3114.000 0.000 3189.000 32.455 ;
      LAYER met5 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io_alt
END LIBRARY

