magic
tech sky130A
magscale 1 2
timestamp 1622552488
<< obsli1 >>
rect 1104 85 198812 29155
<< obsm1 >>
rect 106 8 199810 29164
<< metal2 >>
rect 294 28400 350 29600
rect 846 28400 902 29600
rect 1398 28400 1454 29600
rect 2042 28400 2098 29600
rect 2594 28400 2650 29600
rect 3146 28400 3202 29600
rect 3790 28400 3846 29600
rect 4342 28400 4398 29600
rect 4986 28400 5042 29600
rect 5538 28400 5594 29600
rect 6090 28400 6146 29600
rect 6734 28400 6790 29600
rect 7286 28400 7342 29600
rect 7930 28400 7986 29600
rect 8482 28400 8538 29600
rect 9034 28400 9090 29600
rect 9678 28400 9734 29600
rect 10230 28400 10286 29600
rect 10874 28400 10930 29600
rect 11426 28400 11482 29600
rect 11978 28400 12034 29600
rect 12622 28400 12678 29600
rect 13174 28400 13230 29600
rect 13818 28400 13874 29600
rect 14370 28400 14426 29600
rect 14922 28400 14978 29600
rect 15566 28400 15622 29600
rect 16118 28400 16174 29600
rect 16762 28400 16818 29600
rect 17314 28400 17370 29600
rect 17866 28400 17922 29600
rect 18510 28400 18566 29600
rect 19062 28400 19118 29600
rect 19706 28400 19762 29600
rect 20258 28400 20314 29600
rect 20810 28400 20866 29600
rect 21454 28400 21510 29600
rect 22006 28400 22062 29600
rect 22558 28400 22614 29600
rect 23202 28400 23258 29600
rect 23754 28400 23810 29600
rect 24398 28400 24454 29600
rect 24950 28400 25006 29600
rect 25502 28400 25558 29600
rect 26146 28400 26202 29600
rect 26698 28400 26754 29600
rect 27342 28400 27398 29600
rect 27894 28400 27950 29600
rect 28446 28400 28502 29600
rect 29090 28400 29146 29600
rect 29642 28400 29698 29600
rect 30286 28400 30342 29600
rect 30838 28400 30894 29600
rect 31390 28400 31446 29600
rect 32034 28400 32090 29600
rect 32586 28400 32642 29600
rect 33230 28400 33286 29600
rect 33782 28400 33838 29600
rect 34334 28400 34390 29600
rect 34978 28400 35034 29600
rect 35530 28400 35586 29600
rect 36174 28400 36230 29600
rect 36726 28400 36782 29600
rect 37278 28400 37334 29600
rect 37922 28400 37978 29600
rect 38474 28400 38530 29600
rect 39118 28400 39174 29600
rect 39670 28400 39726 29600
rect 40222 28400 40278 29600
rect 40866 28400 40922 29600
rect 41418 28400 41474 29600
rect 41970 28400 42026 29600
rect 42614 28400 42670 29600
rect 43166 28400 43222 29600
rect 43810 28400 43866 29600
rect 44362 28400 44418 29600
rect 44914 28400 44970 29600
rect 45558 28400 45614 29600
rect 46110 28400 46166 29600
rect 46754 28400 46810 29600
rect 47306 28400 47362 29600
rect 47858 28400 47914 29600
rect 48502 28400 48558 29600
rect 49054 28400 49110 29600
rect 49698 28400 49754 29600
rect 50250 28400 50306 29600
rect 50802 28400 50858 29600
rect 51446 28400 51502 29600
rect 51998 28400 52054 29600
rect 52642 28400 52698 29600
rect 53194 28400 53250 29600
rect 53746 28400 53802 29600
rect 54390 28400 54446 29600
rect 54942 28400 54998 29600
rect 55586 28400 55642 29600
rect 56138 28400 56194 29600
rect 56690 28400 56746 29600
rect 57334 28400 57390 29600
rect 57886 28400 57942 29600
rect 58530 28400 58586 29600
rect 59082 28400 59138 29600
rect 59634 28400 59690 29600
rect 60278 28400 60334 29600
rect 60830 28400 60886 29600
rect 61382 28400 61438 29600
rect 62026 28400 62082 29600
rect 62578 28400 62634 29600
rect 63222 28400 63278 29600
rect 63774 28400 63830 29600
rect 64326 28400 64382 29600
rect 64970 28400 65026 29600
rect 65522 28400 65578 29600
rect 66166 28400 66222 29600
rect 66718 28400 66774 29600
rect 67270 28400 67326 29600
rect 67914 28400 67970 29600
rect 68466 28400 68522 29600
rect 69110 28400 69166 29600
rect 69662 28400 69718 29600
rect 70214 28400 70270 29600
rect 70858 28400 70914 29600
rect 71410 28400 71466 29600
rect 72054 28400 72110 29600
rect 72606 28400 72662 29600
rect 73158 28400 73214 29600
rect 73802 28400 73858 29600
rect 74354 28400 74410 29600
rect 74998 28400 75054 29600
rect 75550 28400 75606 29600
rect 76102 28400 76158 29600
rect 76746 28400 76802 29600
rect 77298 28400 77354 29600
rect 77942 28400 77998 29600
rect 78494 28400 78550 29600
rect 79046 28400 79102 29600
rect 79690 28400 79746 29600
rect 80242 28400 80298 29600
rect 80794 28400 80850 29600
rect 81438 28400 81494 29600
rect 81990 28400 82046 29600
rect 82634 28400 82690 29600
rect 83186 28400 83242 29600
rect 83738 28400 83794 29600
rect 84382 28400 84438 29600
rect 84934 28400 84990 29600
rect 85578 28400 85634 29600
rect 86130 28400 86186 29600
rect 86682 28400 86738 29600
rect 87326 28400 87382 29600
rect 87878 28400 87934 29600
rect 88522 28400 88578 29600
rect 89074 28400 89130 29600
rect 89626 28400 89682 29600
rect 90270 28400 90326 29600
rect 90822 28400 90878 29600
rect 91466 28400 91522 29600
rect 92018 28400 92074 29600
rect 92570 28400 92626 29600
rect 93214 28400 93270 29600
rect 93766 28400 93822 29600
rect 94410 28400 94466 29600
rect 94962 28400 95018 29600
rect 95514 28400 95570 29600
rect 96158 28400 96214 29600
rect 96710 28400 96766 29600
rect 97354 28400 97410 29600
rect 97906 28400 97962 29600
rect 98458 28400 98514 29600
rect 99102 28400 99158 29600
rect 99654 28400 99710 29600
rect 100298 28400 100354 29600
rect 100850 28400 100906 29600
rect 101402 28400 101458 29600
rect 102046 28400 102102 29600
rect 102598 28400 102654 29600
rect 103150 28400 103206 29600
rect 103794 28400 103850 29600
rect 104346 28400 104402 29600
rect 104990 28400 105046 29600
rect 105542 28400 105598 29600
rect 106094 28400 106150 29600
rect 106738 28400 106794 29600
rect 107290 28400 107346 29600
rect 107934 28400 107990 29600
rect 108486 28400 108542 29600
rect 109038 28400 109094 29600
rect 109682 28400 109738 29600
rect 110234 28400 110290 29600
rect 110878 28400 110934 29600
rect 111430 28400 111486 29600
rect 111982 28400 112038 29600
rect 112626 28400 112682 29600
rect 113178 28400 113234 29600
rect 113822 28400 113878 29600
rect 114374 28400 114430 29600
rect 114926 28400 114982 29600
rect 115570 28400 115626 29600
rect 116122 28400 116178 29600
rect 116766 28400 116822 29600
rect 117318 28400 117374 29600
rect 117870 28400 117926 29600
rect 118514 28400 118570 29600
rect 119066 28400 119122 29600
rect 119710 28400 119766 29600
rect 120262 28400 120318 29600
rect 120814 28400 120870 29600
rect 121458 28400 121514 29600
rect 122010 28400 122066 29600
rect 122562 28400 122618 29600
rect 123206 28400 123262 29600
rect 123758 28400 123814 29600
rect 124402 28400 124458 29600
rect 124954 28400 125010 29600
rect 125506 28400 125562 29600
rect 126150 28400 126206 29600
rect 126702 28400 126758 29600
rect 127346 28400 127402 29600
rect 127898 28400 127954 29600
rect 128450 28400 128506 29600
rect 129094 28400 129150 29600
rect 129646 28400 129702 29600
rect 130290 28400 130346 29600
rect 130842 28400 130898 29600
rect 131394 28400 131450 29600
rect 132038 28400 132094 29600
rect 132590 28400 132646 29600
rect 133234 28400 133290 29600
rect 133786 28400 133842 29600
rect 134338 28400 134394 29600
rect 134982 28400 135038 29600
rect 135534 28400 135590 29600
rect 136178 28400 136234 29600
rect 136730 28400 136786 29600
rect 137282 28400 137338 29600
rect 137926 28400 137982 29600
rect 138478 28400 138534 29600
rect 139122 28400 139178 29600
rect 139674 28400 139730 29600
rect 140226 28400 140282 29600
rect 140870 28400 140926 29600
rect 141422 28400 141478 29600
rect 141974 28400 142030 29600
rect 142618 28400 142674 29600
rect 143170 28400 143226 29600
rect 143814 28400 143870 29600
rect 144366 28400 144422 29600
rect 144918 28400 144974 29600
rect 145562 28400 145618 29600
rect 146114 28400 146170 29600
rect 146758 28400 146814 29600
rect 147310 28400 147366 29600
rect 147862 28400 147918 29600
rect 148506 28400 148562 29600
rect 149058 28400 149114 29600
rect 149702 28400 149758 29600
rect 150254 28400 150310 29600
rect 150806 28400 150862 29600
rect 151450 28400 151506 29600
rect 152002 28400 152058 29600
rect 152646 28400 152702 29600
rect 153198 28400 153254 29600
rect 153750 28400 153806 29600
rect 154394 28400 154450 29600
rect 154946 28400 155002 29600
rect 155590 28400 155646 29600
rect 156142 28400 156198 29600
rect 156694 28400 156750 29600
rect 157338 28400 157394 29600
rect 157890 28400 157946 29600
rect 158534 28400 158590 29600
rect 159086 28400 159142 29600
rect 159638 28400 159694 29600
rect 160282 28400 160338 29600
rect 160834 28400 160890 29600
rect 161386 28400 161442 29600
rect 162030 28400 162086 29600
rect 162582 28400 162638 29600
rect 163226 28400 163282 29600
rect 163778 28400 163834 29600
rect 164330 28400 164386 29600
rect 164974 28400 165030 29600
rect 165526 28400 165582 29600
rect 166170 28400 166226 29600
rect 166722 28400 166778 29600
rect 167274 28400 167330 29600
rect 167918 28400 167974 29600
rect 168470 28400 168526 29600
rect 169114 28400 169170 29600
rect 169666 28400 169722 29600
rect 170218 28400 170274 29600
rect 170862 28400 170918 29600
rect 171414 28400 171470 29600
rect 172058 28400 172114 29600
rect 172610 28400 172666 29600
rect 173162 28400 173218 29600
rect 173806 28400 173862 29600
rect 174358 28400 174414 29600
rect 175002 28400 175058 29600
rect 175554 28400 175610 29600
rect 176106 28400 176162 29600
rect 176750 28400 176806 29600
rect 177302 28400 177358 29600
rect 177946 28400 178002 29600
rect 178498 28400 178554 29600
rect 179050 28400 179106 29600
rect 179694 28400 179750 29600
rect 180246 28400 180302 29600
rect 180798 28400 180854 29600
rect 181442 28400 181498 29600
rect 181994 28400 182050 29600
rect 182638 28400 182694 29600
rect 183190 28400 183246 29600
rect 183742 28400 183798 29600
rect 184386 28400 184442 29600
rect 184938 28400 184994 29600
rect 185582 28400 185638 29600
rect 186134 28400 186190 29600
rect 186686 28400 186742 29600
rect 187330 28400 187386 29600
rect 187882 28400 187938 29600
rect 188526 28400 188582 29600
rect 189078 28400 189134 29600
rect 189630 28400 189686 29600
rect 190274 28400 190330 29600
rect 190826 28400 190882 29600
rect 191470 28400 191526 29600
rect 192022 28400 192078 29600
rect 192574 28400 192630 29600
rect 193218 28400 193274 29600
rect 193770 28400 193826 29600
rect 194414 28400 194470 29600
rect 194966 28400 195022 29600
rect 195518 28400 195574 29600
rect 196162 28400 196218 29600
rect 196714 28400 196770 29600
rect 197358 28400 197414 29600
rect 197910 28400 197966 29600
rect 198462 28400 198518 29600
rect 199106 28400 199162 29600
rect 199658 28400 199714 29600
rect 110 -400 166 800
rect 386 -400 442 800
rect 662 -400 718 800
rect 938 -400 994 800
rect 1214 -400 1270 800
rect 1490 -400 1546 800
rect 1766 -400 1822 800
rect 2042 -400 2098 800
rect 2318 -400 2374 800
rect 2594 -400 2650 800
rect 2870 -400 2926 800
rect 3146 -400 3202 800
rect 3422 -400 3478 800
rect 3698 -400 3754 800
rect 3974 -400 4030 800
rect 4250 -400 4306 800
rect 4526 -400 4582 800
rect 4802 -400 4858 800
rect 5078 -400 5134 800
rect 5354 -400 5410 800
rect 5630 -400 5686 800
rect 5906 -400 5962 800
rect 6182 -400 6238 800
rect 6458 -400 6514 800
rect 6734 -400 6790 800
rect 7102 -400 7158 800
rect 7378 -400 7434 800
rect 7654 -400 7710 800
rect 7930 -400 7986 800
rect 8206 -400 8262 800
rect 8482 -400 8538 800
rect 8758 -400 8814 800
rect 9034 -400 9090 800
rect 9310 -400 9366 800
rect 9586 -400 9642 800
rect 9862 -400 9918 800
rect 10138 -400 10194 800
rect 10414 -400 10470 800
rect 10690 -400 10746 800
rect 10966 -400 11022 800
rect 11242 -400 11298 800
rect 11518 -400 11574 800
rect 11794 -400 11850 800
rect 12070 -400 12126 800
rect 12346 -400 12402 800
rect 12622 -400 12678 800
rect 12898 -400 12954 800
rect 13174 -400 13230 800
rect 13450 -400 13506 800
rect 13726 -400 13782 800
rect 14094 -400 14150 800
rect 14370 -400 14426 800
rect 14646 -400 14702 800
rect 14922 -400 14978 800
rect 15198 -400 15254 800
rect 15474 -400 15530 800
rect 15750 -400 15806 800
rect 16026 -400 16082 800
rect 16302 -400 16358 800
rect 16578 -400 16634 800
rect 16854 -400 16910 800
rect 17130 -400 17186 800
rect 17406 -400 17462 800
rect 17682 -400 17738 800
rect 17958 -400 18014 800
rect 18234 -400 18290 800
rect 18510 -400 18566 800
rect 18786 -400 18842 800
rect 19062 -400 19118 800
rect 19338 -400 19394 800
rect 19614 -400 19670 800
rect 19890 -400 19946 800
rect 20166 -400 20222 800
rect 20442 -400 20498 800
rect 20810 -400 20866 800
rect 21086 -400 21142 800
rect 21362 -400 21418 800
rect 21638 -400 21694 800
rect 21914 -400 21970 800
rect 22190 -400 22246 800
rect 22466 -400 22522 800
rect 22742 -400 22798 800
rect 23018 -400 23074 800
rect 23294 -400 23350 800
rect 23570 -400 23626 800
rect 23846 -400 23902 800
rect 24122 -400 24178 800
rect 24398 -400 24454 800
rect 24674 -400 24730 800
rect 24950 -400 25006 800
rect 25226 -400 25282 800
rect 25502 -400 25558 800
rect 25778 -400 25834 800
rect 26054 -400 26110 800
rect 26330 -400 26386 800
rect 26606 -400 26662 800
rect 26882 -400 26938 800
rect 27158 -400 27214 800
rect 27434 -400 27490 800
rect 27802 -400 27858 800
rect 28078 -400 28134 800
rect 28354 -400 28410 800
rect 28630 -400 28686 800
rect 28906 -400 28962 800
rect 29182 -400 29238 800
rect 29458 -400 29514 800
rect 29734 -400 29790 800
rect 30010 -400 30066 800
rect 30286 -400 30342 800
rect 30562 -400 30618 800
rect 30838 -400 30894 800
rect 31114 -400 31170 800
rect 31390 -400 31446 800
rect 31666 -400 31722 800
rect 31942 -400 31998 800
rect 32218 -400 32274 800
rect 32494 -400 32550 800
rect 32770 -400 32826 800
rect 33046 -400 33102 800
rect 33322 -400 33378 800
rect 33598 -400 33654 800
rect 33874 -400 33930 800
rect 34150 -400 34206 800
rect 34426 -400 34482 800
rect 34794 -400 34850 800
rect 35070 -400 35126 800
rect 35346 -400 35402 800
rect 35622 -400 35678 800
rect 35898 -400 35954 800
rect 36174 -400 36230 800
rect 36450 -400 36506 800
rect 36726 -400 36782 800
rect 37002 -400 37058 800
rect 37278 -400 37334 800
rect 37554 -400 37610 800
rect 37830 -400 37886 800
rect 38106 -400 38162 800
rect 38382 -400 38438 800
rect 38658 -400 38714 800
rect 38934 -400 38990 800
rect 39210 -400 39266 800
rect 39486 -400 39542 800
rect 39762 -400 39818 800
rect 40038 -400 40094 800
rect 40314 -400 40370 800
rect 40590 -400 40646 800
rect 40866 -400 40922 800
rect 41142 -400 41198 800
rect 41510 -400 41566 800
rect 41786 -400 41842 800
rect 42062 -400 42118 800
rect 42338 -400 42394 800
rect 42614 -400 42670 800
rect 42890 -400 42946 800
rect 43166 -400 43222 800
rect 43442 -400 43498 800
rect 43718 -400 43774 800
rect 43994 -400 44050 800
rect 44270 -400 44326 800
rect 44546 -400 44602 800
rect 44822 -400 44878 800
rect 45098 -400 45154 800
rect 45374 -400 45430 800
rect 45650 -400 45706 800
rect 45926 -400 45982 800
rect 46202 -400 46258 800
rect 46478 -400 46534 800
rect 46754 -400 46810 800
rect 47030 -400 47086 800
rect 47306 -400 47362 800
rect 47582 -400 47638 800
rect 47858 -400 47914 800
rect 48134 -400 48190 800
rect 48502 -400 48558 800
rect 48778 -400 48834 800
rect 49054 -400 49110 800
rect 49330 -400 49386 800
rect 49606 -400 49662 800
rect 49882 -400 49938 800
rect 50158 -400 50214 800
rect 50434 -400 50490 800
rect 50710 -400 50766 800
rect 50986 -400 51042 800
rect 51262 -400 51318 800
rect 51538 -400 51594 800
rect 51814 -400 51870 800
rect 52090 -400 52146 800
rect 52366 -400 52422 800
rect 52642 -400 52698 800
rect 52918 -400 52974 800
rect 53194 -400 53250 800
rect 53470 -400 53526 800
rect 53746 -400 53802 800
rect 54022 -400 54078 800
rect 54298 -400 54354 800
rect 54574 -400 54630 800
rect 54850 -400 54906 800
rect 55126 -400 55182 800
rect 55494 -400 55550 800
rect 55770 -400 55826 800
rect 56046 -400 56102 800
rect 56322 -400 56378 800
rect 56598 -400 56654 800
rect 56874 -400 56930 800
rect 57150 -400 57206 800
rect 57426 -400 57482 800
rect 57702 -400 57758 800
rect 57978 -400 58034 800
rect 58254 -400 58310 800
rect 58530 -400 58586 800
rect 58806 -400 58862 800
rect 59082 -400 59138 800
rect 59358 -400 59414 800
rect 59634 -400 59690 800
rect 59910 -400 59966 800
rect 60186 -400 60242 800
rect 60462 -400 60518 800
rect 60738 -400 60794 800
rect 61014 -400 61070 800
rect 61290 -400 61346 800
rect 61566 -400 61622 800
rect 61842 -400 61898 800
rect 62210 -400 62266 800
rect 62486 -400 62542 800
rect 62762 -400 62818 800
rect 63038 -400 63094 800
rect 63314 -400 63370 800
rect 63590 -400 63646 800
rect 63866 -400 63922 800
rect 64142 -400 64198 800
rect 64418 -400 64474 800
rect 64694 -400 64750 800
rect 64970 -400 65026 800
rect 65246 -400 65302 800
rect 65522 -400 65578 800
rect 65798 -400 65854 800
rect 66074 -400 66130 800
rect 66350 -400 66406 800
rect 66626 -400 66682 800
rect 66902 -400 66958 800
rect 67178 -400 67234 800
rect 67454 -400 67510 800
rect 67730 -400 67786 800
rect 68006 -400 68062 800
rect 68282 -400 68338 800
rect 68558 -400 68614 800
rect 68834 -400 68890 800
rect 69202 -400 69258 800
rect 69478 -400 69534 800
rect 69754 -400 69810 800
rect 70030 -400 70086 800
rect 70306 -400 70362 800
rect 70582 -400 70638 800
rect 70858 -400 70914 800
rect 71134 -400 71190 800
rect 71410 -400 71466 800
rect 71686 -400 71742 800
rect 71962 -400 72018 800
rect 72238 -400 72294 800
rect 72514 -400 72570 800
rect 72790 -400 72846 800
rect 73066 -400 73122 800
rect 73342 -400 73398 800
rect 73618 -400 73674 800
rect 73894 -400 73950 800
rect 74170 -400 74226 800
rect 74446 -400 74502 800
rect 74722 -400 74778 800
rect 74998 -400 75054 800
rect 75274 -400 75330 800
rect 75550 -400 75606 800
rect 75826 -400 75882 800
rect 76194 -400 76250 800
rect 76470 -400 76526 800
rect 76746 -400 76802 800
rect 77022 -400 77078 800
rect 77298 -400 77354 800
rect 77574 -400 77630 800
rect 77850 -400 77906 800
rect 78126 -400 78182 800
rect 78402 -400 78458 800
rect 78678 -400 78734 800
rect 78954 -400 79010 800
rect 79230 -400 79286 800
rect 79506 -400 79562 800
rect 79782 -400 79838 800
rect 80058 -400 80114 800
rect 80334 -400 80390 800
rect 80610 -400 80666 800
rect 80886 -400 80942 800
rect 81162 -400 81218 800
rect 81438 -400 81494 800
rect 81714 -400 81770 800
rect 81990 -400 82046 800
rect 82266 -400 82322 800
rect 82542 -400 82598 800
rect 82910 -400 82966 800
rect 83186 -400 83242 800
rect 83462 -400 83518 800
rect 83738 -400 83794 800
rect 84014 -400 84070 800
rect 84290 -400 84346 800
rect 84566 -400 84622 800
rect 84842 -400 84898 800
rect 85118 -400 85174 800
rect 85394 -400 85450 800
rect 85670 -400 85726 800
rect 85946 -400 86002 800
rect 86222 -400 86278 800
rect 86498 -400 86554 800
rect 86774 -400 86830 800
rect 87050 -400 87106 800
rect 87326 -400 87382 800
rect 87602 -400 87658 800
rect 87878 -400 87934 800
rect 88154 -400 88210 800
rect 88430 -400 88486 800
rect 88706 -400 88762 800
rect 88982 -400 89038 800
rect 89258 -400 89314 800
rect 89534 -400 89590 800
rect 89902 -400 89958 800
rect 90178 -400 90234 800
rect 90454 -400 90510 800
rect 90730 -400 90786 800
rect 91006 -400 91062 800
rect 91282 -400 91338 800
rect 91558 -400 91614 800
rect 91834 -400 91890 800
rect 92110 -400 92166 800
rect 92386 -400 92442 800
rect 92662 -400 92718 800
rect 92938 -400 92994 800
rect 93214 -400 93270 800
rect 93490 -400 93546 800
rect 93766 -400 93822 800
rect 94042 -400 94098 800
rect 94318 -400 94374 800
rect 94594 -400 94650 800
rect 94870 -400 94926 800
rect 95146 -400 95202 800
rect 95422 -400 95478 800
rect 95698 -400 95754 800
rect 95974 -400 96030 800
rect 96250 -400 96306 800
rect 96526 -400 96582 800
rect 96894 -400 96950 800
rect 97170 -400 97226 800
rect 97446 -400 97502 800
rect 97722 -400 97778 800
rect 97998 -400 98054 800
rect 98274 -400 98330 800
rect 98550 -400 98606 800
rect 98826 -400 98882 800
rect 99102 -400 99158 800
rect 99378 -400 99434 800
rect 99654 -400 99710 800
rect 99930 -400 99986 800
rect 100206 -400 100262 800
rect 100482 -400 100538 800
rect 100758 -400 100814 800
rect 101034 -400 101090 800
rect 101310 -400 101366 800
rect 101586 -400 101642 800
rect 101862 -400 101918 800
rect 102138 -400 102194 800
rect 102414 -400 102470 800
rect 102690 -400 102746 800
rect 102966 -400 103022 800
rect 103242 -400 103298 800
rect 103610 -400 103666 800
rect 103886 -400 103942 800
rect 104162 -400 104218 800
rect 104438 -400 104494 800
rect 104714 -400 104770 800
rect 104990 -400 105046 800
rect 105266 -400 105322 800
rect 105542 -400 105598 800
rect 105818 -400 105874 800
rect 106094 -400 106150 800
rect 106370 -400 106426 800
rect 106646 -400 106702 800
rect 106922 -400 106978 800
rect 107198 -400 107254 800
rect 107474 -400 107530 800
rect 107750 -400 107806 800
rect 108026 -400 108082 800
rect 108302 -400 108358 800
rect 108578 -400 108634 800
rect 108854 -400 108910 800
rect 109130 -400 109186 800
rect 109406 -400 109462 800
rect 109682 -400 109738 800
rect 109958 -400 110014 800
rect 110234 -400 110290 800
rect 110602 -400 110658 800
rect 110878 -400 110934 800
rect 111154 -400 111210 800
rect 111430 -400 111486 800
rect 111706 -400 111762 800
rect 111982 -400 112038 800
rect 112258 -400 112314 800
rect 112534 -400 112590 800
rect 112810 -400 112866 800
rect 113086 -400 113142 800
rect 113362 -400 113418 800
rect 113638 -400 113694 800
rect 113914 -400 113970 800
rect 114190 -400 114246 800
rect 114466 -400 114522 800
rect 114742 -400 114798 800
rect 115018 -400 115074 800
rect 115294 -400 115350 800
rect 115570 -400 115626 800
rect 115846 -400 115902 800
rect 116122 -400 116178 800
rect 116398 -400 116454 800
rect 116674 -400 116730 800
rect 116950 -400 117006 800
rect 117226 -400 117282 800
rect 117594 -400 117650 800
rect 117870 -400 117926 800
rect 118146 -400 118202 800
rect 118422 -400 118478 800
rect 118698 -400 118754 800
rect 118974 -400 119030 800
rect 119250 -400 119306 800
rect 119526 -400 119582 800
rect 119802 -400 119858 800
rect 120078 -400 120134 800
rect 120354 -400 120410 800
rect 120630 -400 120686 800
rect 120906 -400 120962 800
rect 121182 -400 121238 800
rect 121458 -400 121514 800
rect 121734 -400 121790 800
rect 122010 -400 122066 800
rect 122286 -400 122342 800
rect 122562 -400 122618 800
rect 122838 -400 122894 800
rect 123114 -400 123170 800
rect 123390 -400 123446 800
rect 123666 -400 123722 800
rect 123942 -400 123998 800
rect 124310 -400 124366 800
rect 124586 -400 124642 800
rect 124862 -400 124918 800
rect 125138 -400 125194 800
rect 125414 -400 125470 800
rect 125690 -400 125746 800
rect 125966 -400 126022 800
rect 126242 -400 126298 800
rect 126518 -400 126574 800
rect 126794 -400 126850 800
rect 127070 -400 127126 800
rect 127346 -400 127402 800
rect 127622 -400 127678 800
rect 127898 -400 127954 800
rect 128174 -400 128230 800
rect 128450 -400 128506 800
rect 128726 -400 128782 800
rect 129002 -400 129058 800
rect 129278 -400 129334 800
rect 129554 -400 129610 800
rect 129830 -400 129886 800
rect 130106 -400 130162 800
rect 130382 -400 130438 800
rect 130658 -400 130714 800
rect 130934 -400 130990 800
rect 131302 -400 131358 800
rect 131578 -400 131634 800
rect 131854 -400 131910 800
rect 132130 -400 132186 800
rect 132406 -400 132462 800
rect 132682 -400 132738 800
rect 132958 -400 133014 800
rect 133234 -400 133290 800
rect 133510 -400 133566 800
rect 133786 -400 133842 800
rect 134062 -400 134118 800
rect 134338 -400 134394 800
rect 134614 -400 134670 800
rect 134890 -400 134946 800
rect 135166 -400 135222 800
rect 135442 -400 135498 800
rect 135718 -400 135774 800
rect 135994 -400 136050 800
rect 136270 -400 136326 800
rect 136546 -400 136602 800
rect 136822 -400 136878 800
rect 137098 -400 137154 800
rect 137374 -400 137430 800
rect 137650 -400 137706 800
rect 137926 -400 137982 800
rect 138294 -400 138350 800
rect 138570 -400 138626 800
rect 138846 -400 138902 800
rect 139122 -400 139178 800
rect 139398 -400 139454 800
rect 139674 -400 139730 800
rect 139950 -400 140006 800
rect 140226 -400 140282 800
rect 140502 -400 140558 800
rect 140778 -400 140834 800
rect 141054 -400 141110 800
rect 141330 -400 141386 800
rect 141606 -400 141662 800
rect 141882 -400 141938 800
rect 142158 -400 142214 800
rect 142434 -400 142490 800
rect 142710 -400 142766 800
rect 142986 -400 143042 800
rect 143262 -400 143318 800
rect 143538 -400 143594 800
rect 143814 -400 143870 800
rect 144090 -400 144146 800
rect 144366 -400 144422 800
rect 144642 -400 144698 800
rect 145010 -400 145066 800
rect 145286 -400 145342 800
rect 145562 -400 145618 800
rect 145838 -400 145894 800
rect 146114 -400 146170 800
rect 146390 -400 146446 800
rect 146666 -400 146722 800
rect 146942 -400 146998 800
rect 147218 -400 147274 800
rect 147494 -400 147550 800
rect 147770 -400 147826 800
rect 148046 -400 148102 800
rect 148322 -400 148378 800
rect 148598 -400 148654 800
rect 148874 -400 148930 800
rect 149150 -400 149206 800
rect 149426 -400 149482 800
rect 149702 -400 149758 800
rect 149978 -400 150034 800
rect 150254 -400 150310 800
rect 150530 -400 150586 800
rect 150806 -400 150862 800
rect 151082 -400 151138 800
rect 151358 -400 151414 800
rect 151634 -400 151690 800
rect 152002 -400 152058 800
rect 152278 -400 152334 800
rect 152554 -400 152610 800
rect 152830 -400 152886 800
rect 153106 -400 153162 800
rect 153382 -400 153438 800
rect 153658 -400 153714 800
rect 153934 -400 153990 800
rect 154210 -400 154266 800
rect 154486 -400 154542 800
rect 154762 -400 154818 800
rect 155038 -400 155094 800
rect 155314 -400 155370 800
rect 155590 -400 155646 800
rect 155866 -400 155922 800
rect 156142 -400 156198 800
rect 156418 -400 156474 800
rect 156694 -400 156750 800
rect 156970 -400 157026 800
rect 157246 -400 157302 800
rect 157522 -400 157578 800
rect 157798 -400 157854 800
rect 158074 -400 158130 800
rect 158350 -400 158406 800
rect 158626 -400 158682 800
rect 158994 -400 159050 800
rect 159270 -400 159326 800
rect 159546 -400 159602 800
rect 159822 -400 159878 800
rect 160098 -400 160154 800
rect 160374 -400 160430 800
rect 160650 -400 160706 800
rect 160926 -400 160982 800
rect 161202 -400 161258 800
rect 161478 -400 161534 800
rect 161754 -400 161810 800
rect 162030 -400 162086 800
rect 162306 -400 162362 800
rect 162582 -400 162638 800
rect 162858 -400 162914 800
rect 163134 -400 163190 800
rect 163410 -400 163466 800
rect 163686 -400 163742 800
rect 163962 -400 164018 800
rect 164238 -400 164294 800
rect 164514 -400 164570 800
rect 164790 -400 164846 800
rect 165066 -400 165122 800
rect 165342 -400 165398 800
rect 165710 -400 165766 800
rect 165986 -400 166042 800
rect 166262 -400 166318 800
rect 166538 -400 166594 800
rect 166814 -400 166870 800
rect 167090 -400 167146 800
rect 167366 -400 167422 800
rect 167642 -400 167698 800
rect 167918 -400 167974 800
rect 168194 -400 168250 800
rect 168470 -400 168526 800
rect 168746 -400 168802 800
rect 169022 -400 169078 800
rect 169298 -400 169354 800
rect 169574 -400 169630 800
rect 169850 -400 169906 800
rect 170126 -400 170182 800
rect 170402 -400 170458 800
rect 170678 -400 170734 800
rect 170954 -400 171010 800
rect 171230 -400 171286 800
rect 171506 -400 171562 800
rect 171782 -400 171838 800
rect 172058 -400 172114 800
rect 172334 -400 172390 800
rect 172702 -400 172758 800
rect 172978 -400 173034 800
rect 173254 -400 173310 800
rect 173530 -400 173586 800
rect 173806 -400 173862 800
rect 174082 -400 174138 800
rect 174358 -400 174414 800
rect 174634 -400 174690 800
rect 174910 -400 174966 800
rect 175186 -400 175242 800
rect 175462 -400 175518 800
rect 175738 -400 175794 800
rect 176014 -400 176070 800
rect 176290 -400 176346 800
rect 176566 -400 176622 800
rect 176842 -400 176898 800
rect 177118 -400 177174 800
rect 177394 -400 177450 800
rect 177670 -400 177726 800
rect 177946 -400 178002 800
rect 178222 -400 178278 800
rect 178498 -400 178554 800
rect 178774 -400 178830 800
rect 179050 -400 179106 800
rect 179326 -400 179382 800
rect 179694 -400 179750 800
rect 179970 -400 180026 800
rect 180246 -400 180302 800
rect 180522 -400 180578 800
rect 180798 -400 180854 800
rect 181074 -400 181130 800
rect 181350 -400 181406 800
rect 181626 -400 181682 800
rect 181902 -400 181958 800
rect 182178 -400 182234 800
rect 182454 -400 182510 800
rect 182730 -400 182786 800
rect 183006 -400 183062 800
rect 183282 -400 183338 800
rect 183558 -400 183614 800
rect 183834 -400 183890 800
rect 184110 -400 184166 800
rect 184386 -400 184442 800
rect 184662 -400 184718 800
rect 184938 -400 184994 800
rect 185214 -400 185270 800
rect 185490 -400 185546 800
rect 185766 -400 185822 800
rect 186042 -400 186098 800
rect 186410 -400 186466 800
rect 186686 -400 186742 800
rect 186962 -400 187018 800
rect 187238 -400 187294 800
rect 187514 -400 187570 800
rect 187790 -400 187846 800
rect 188066 -400 188122 800
rect 188342 -400 188398 800
rect 188618 -400 188674 800
rect 188894 -400 188950 800
rect 189170 -400 189226 800
rect 189446 -400 189502 800
rect 189722 -400 189778 800
rect 189998 -400 190054 800
rect 190274 -400 190330 800
rect 190550 -400 190606 800
rect 190826 -400 190882 800
rect 191102 -400 191158 800
rect 191378 -400 191434 800
rect 191654 -400 191710 800
rect 191930 -400 191986 800
rect 192206 -400 192262 800
rect 192482 -400 192538 800
rect 192758 -400 192814 800
rect 193034 -400 193090 800
rect 193402 -400 193458 800
rect 193678 -400 193734 800
rect 193954 -400 194010 800
rect 194230 -400 194286 800
rect 194506 -400 194562 800
rect 194782 -400 194838 800
rect 195058 -400 195114 800
rect 195334 -400 195390 800
rect 195610 -400 195666 800
rect 195886 -400 195942 800
rect 196162 -400 196218 800
rect 196438 -400 196494 800
rect 196714 -400 196770 800
rect 196990 -400 197046 800
rect 197266 -400 197322 800
rect 197542 -400 197598 800
rect 197818 -400 197874 800
rect 198094 -400 198150 800
rect 198370 -400 198426 800
rect 198646 -400 198702 800
rect 198922 -400 198978 800
rect 199198 -400 199254 800
rect 199474 -400 199530 800
rect 199750 -400 199806 800
<< obsm2 >>
rect 112 28344 238 29170
rect 406 28344 790 29170
rect 958 28344 1342 29170
rect 1510 28344 1986 29170
rect 2154 28344 2538 29170
rect 2706 28344 3090 29170
rect 3258 28344 3734 29170
rect 3902 28344 4286 29170
rect 4454 28344 4930 29170
rect 5098 28344 5482 29170
rect 5650 28344 6034 29170
rect 6202 28344 6678 29170
rect 6846 28344 7230 29170
rect 7398 28344 7874 29170
rect 8042 28344 8426 29170
rect 8594 28344 8978 29170
rect 9146 28344 9622 29170
rect 9790 28344 10174 29170
rect 10342 28344 10818 29170
rect 10986 28344 11370 29170
rect 11538 28344 11922 29170
rect 12090 28344 12566 29170
rect 12734 28344 13118 29170
rect 13286 28344 13762 29170
rect 13930 28344 14314 29170
rect 14482 28344 14866 29170
rect 15034 28344 15510 29170
rect 15678 28344 16062 29170
rect 16230 28344 16706 29170
rect 16874 28344 17258 29170
rect 17426 28344 17810 29170
rect 17978 28344 18454 29170
rect 18622 28344 19006 29170
rect 19174 28344 19650 29170
rect 19818 28344 20202 29170
rect 20370 28344 20754 29170
rect 20922 28344 21398 29170
rect 21566 28344 21950 29170
rect 22118 28344 22502 29170
rect 22670 28344 23146 29170
rect 23314 28344 23698 29170
rect 23866 28344 24342 29170
rect 24510 28344 24894 29170
rect 25062 28344 25446 29170
rect 25614 28344 26090 29170
rect 26258 28344 26642 29170
rect 26810 28344 27286 29170
rect 27454 28344 27838 29170
rect 28006 28344 28390 29170
rect 28558 28344 29034 29170
rect 29202 28344 29586 29170
rect 29754 28344 30230 29170
rect 30398 28344 30782 29170
rect 30950 28344 31334 29170
rect 31502 28344 31978 29170
rect 32146 28344 32530 29170
rect 32698 28344 33174 29170
rect 33342 28344 33726 29170
rect 33894 28344 34278 29170
rect 34446 28344 34922 29170
rect 35090 28344 35474 29170
rect 35642 28344 36118 29170
rect 36286 28344 36670 29170
rect 36838 28344 37222 29170
rect 37390 28344 37866 29170
rect 38034 28344 38418 29170
rect 38586 28344 39062 29170
rect 39230 28344 39614 29170
rect 39782 28344 40166 29170
rect 40334 28344 40810 29170
rect 40978 28344 41362 29170
rect 41530 28344 41914 29170
rect 42082 28344 42558 29170
rect 42726 28344 43110 29170
rect 43278 28344 43754 29170
rect 43922 28344 44306 29170
rect 44474 28344 44858 29170
rect 45026 28344 45502 29170
rect 45670 28344 46054 29170
rect 46222 28344 46698 29170
rect 46866 28344 47250 29170
rect 47418 28344 47802 29170
rect 47970 28344 48446 29170
rect 48614 28344 48998 29170
rect 49166 28344 49642 29170
rect 49810 28344 50194 29170
rect 50362 28344 50746 29170
rect 50914 28344 51390 29170
rect 51558 28344 51942 29170
rect 52110 28344 52586 29170
rect 52754 28344 53138 29170
rect 53306 28344 53690 29170
rect 53858 28344 54334 29170
rect 54502 28344 54886 29170
rect 55054 28344 55530 29170
rect 55698 28344 56082 29170
rect 56250 28344 56634 29170
rect 56802 28344 57278 29170
rect 57446 28344 57830 29170
rect 57998 28344 58474 29170
rect 58642 28344 59026 29170
rect 59194 28344 59578 29170
rect 59746 28344 60222 29170
rect 60390 28344 60774 29170
rect 60942 28344 61326 29170
rect 61494 28344 61970 29170
rect 62138 28344 62522 29170
rect 62690 28344 63166 29170
rect 63334 28344 63718 29170
rect 63886 28344 64270 29170
rect 64438 28344 64914 29170
rect 65082 28344 65466 29170
rect 65634 28344 66110 29170
rect 66278 28344 66662 29170
rect 66830 28344 67214 29170
rect 67382 28344 67858 29170
rect 68026 28344 68410 29170
rect 68578 28344 69054 29170
rect 69222 28344 69606 29170
rect 69774 28344 70158 29170
rect 70326 28344 70802 29170
rect 70970 28344 71354 29170
rect 71522 28344 71998 29170
rect 72166 28344 72550 29170
rect 72718 28344 73102 29170
rect 73270 28344 73746 29170
rect 73914 28344 74298 29170
rect 74466 28344 74942 29170
rect 75110 28344 75494 29170
rect 75662 28344 76046 29170
rect 76214 28344 76690 29170
rect 76858 28344 77242 29170
rect 77410 28344 77886 29170
rect 78054 28344 78438 29170
rect 78606 28344 78990 29170
rect 79158 28344 79634 29170
rect 79802 28344 80186 29170
rect 80354 28344 80738 29170
rect 80906 28344 81382 29170
rect 81550 28344 81934 29170
rect 82102 28344 82578 29170
rect 82746 28344 83130 29170
rect 83298 28344 83682 29170
rect 83850 28344 84326 29170
rect 84494 28344 84878 29170
rect 85046 28344 85522 29170
rect 85690 28344 86074 29170
rect 86242 28344 86626 29170
rect 86794 28344 87270 29170
rect 87438 28344 87822 29170
rect 87990 28344 88466 29170
rect 88634 28344 89018 29170
rect 89186 28344 89570 29170
rect 89738 28344 90214 29170
rect 90382 28344 90766 29170
rect 90934 28344 91410 29170
rect 91578 28344 91962 29170
rect 92130 28344 92514 29170
rect 92682 28344 93158 29170
rect 93326 28344 93710 29170
rect 93878 28344 94354 29170
rect 94522 28344 94906 29170
rect 95074 28344 95458 29170
rect 95626 28344 96102 29170
rect 96270 28344 96654 29170
rect 96822 28344 97298 29170
rect 97466 28344 97850 29170
rect 98018 28344 98402 29170
rect 98570 28344 99046 29170
rect 99214 28344 99598 29170
rect 99766 28344 100242 29170
rect 100410 28344 100794 29170
rect 100962 28344 101346 29170
rect 101514 28344 101990 29170
rect 102158 28344 102542 29170
rect 102710 28344 103094 29170
rect 103262 28344 103738 29170
rect 103906 28344 104290 29170
rect 104458 28344 104934 29170
rect 105102 28344 105486 29170
rect 105654 28344 106038 29170
rect 106206 28344 106682 29170
rect 106850 28344 107234 29170
rect 107402 28344 107878 29170
rect 108046 28344 108430 29170
rect 108598 28344 108982 29170
rect 109150 28344 109626 29170
rect 109794 28344 110178 29170
rect 110346 28344 110822 29170
rect 110990 28344 111374 29170
rect 111542 28344 111926 29170
rect 112094 28344 112570 29170
rect 112738 28344 113122 29170
rect 113290 28344 113766 29170
rect 113934 28344 114318 29170
rect 114486 28344 114870 29170
rect 115038 28344 115514 29170
rect 115682 28344 116066 29170
rect 116234 28344 116710 29170
rect 116878 28344 117262 29170
rect 117430 28344 117814 29170
rect 117982 28344 118458 29170
rect 118626 28344 119010 29170
rect 119178 28344 119654 29170
rect 119822 28344 120206 29170
rect 120374 28344 120758 29170
rect 120926 28344 121402 29170
rect 121570 28344 121954 29170
rect 122122 28344 122506 29170
rect 122674 28344 123150 29170
rect 123318 28344 123702 29170
rect 123870 28344 124346 29170
rect 124514 28344 124898 29170
rect 125066 28344 125450 29170
rect 125618 28344 126094 29170
rect 126262 28344 126646 29170
rect 126814 28344 127290 29170
rect 127458 28344 127842 29170
rect 128010 28344 128394 29170
rect 128562 28344 129038 29170
rect 129206 28344 129590 29170
rect 129758 28344 130234 29170
rect 130402 28344 130786 29170
rect 130954 28344 131338 29170
rect 131506 28344 131982 29170
rect 132150 28344 132534 29170
rect 132702 28344 133178 29170
rect 133346 28344 133730 29170
rect 133898 28344 134282 29170
rect 134450 28344 134926 29170
rect 135094 28344 135478 29170
rect 135646 28344 136122 29170
rect 136290 28344 136674 29170
rect 136842 28344 137226 29170
rect 137394 28344 137870 29170
rect 138038 28344 138422 29170
rect 138590 28344 139066 29170
rect 139234 28344 139618 29170
rect 139786 28344 140170 29170
rect 140338 28344 140814 29170
rect 140982 28344 141366 29170
rect 141534 28344 141918 29170
rect 142086 28344 142562 29170
rect 142730 28344 143114 29170
rect 143282 28344 143758 29170
rect 143926 28344 144310 29170
rect 144478 28344 144862 29170
rect 145030 28344 145506 29170
rect 145674 28344 146058 29170
rect 146226 28344 146702 29170
rect 146870 28344 147254 29170
rect 147422 28344 147806 29170
rect 147974 28344 148450 29170
rect 148618 28344 149002 29170
rect 149170 28344 149646 29170
rect 149814 28344 150198 29170
rect 150366 28344 150750 29170
rect 150918 28344 151394 29170
rect 151562 28344 151946 29170
rect 152114 28344 152590 29170
rect 152758 28344 153142 29170
rect 153310 28344 153694 29170
rect 153862 28344 154338 29170
rect 154506 28344 154890 29170
rect 155058 28344 155534 29170
rect 155702 28344 156086 29170
rect 156254 28344 156638 29170
rect 156806 28344 157282 29170
rect 157450 28344 157834 29170
rect 158002 28344 158478 29170
rect 158646 28344 159030 29170
rect 159198 28344 159582 29170
rect 159750 28344 160226 29170
rect 160394 28344 160778 29170
rect 160946 28344 161330 29170
rect 161498 28344 161974 29170
rect 162142 28344 162526 29170
rect 162694 28344 163170 29170
rect 163338 28344 163722 29170
rect 163890 28344 164274 29170
rect 164442 28344 164918 29170
rect 165086 28344 165470 29170
rect 165638 28344 166114 29170
rect 166282 28344 166666 29170
rect 166834 28344 167218 29170
rect 167386 28344 167862 29170
rect 168030 28344 168414 29170
rect 168582 28344 169058 29170
rect 169226 28344 169610 29170
rect 169778 28344 170162 29170
rect 170330 28344 170806 29170
rect 170974 28344 171358 29170
rect 171526 28344 172002 29170
rect 172170 28344 172554 29170
rect 172722 28344 173106 29170
rect 173274 28344 173750 29170
rect 173918 28344 174302 29170
rect 174470 28344 174946 29170
rect 175114 28344 175498 29170
rect 175666 28344 176050 29170
rect 176218 28344 176694 29170
rect 176862 28344 177246 29170
rect 177414 28344 177890 29170
rect 178058 28344 178442 29170
rect 178610 28344 178994 29170
rect 179162 28344 179638 29170
rect 179806 28344 180190 29170
rect 180358 28344 180742 29170
rect 180910 28344 181386 29170
rect 181554 28344 181938 29170
rect 182106 28344 182582 29170
rect 182750 28344 183134 29170
rect 183302 28344 183686 29170
rect 183854 28344 184330 29170
rect 184498 28344 184882 29170
rect 185050 28344 185526 29170
rect 185694 28344 186078 29170
rect 186246 28344 186630 29170
rect 186798 28344 187274 29170
rect 187442 28344 187826 29170
rect 187994 28344 188470 29170
rect 188638 28344 189022 29170
rect 189190 28344 189574 29170
rect 189742 28344 190218 29170
rect 190386 28344 190770 29170
rect 190938 28344 191414 29170
rect 191582 28344 191966 29170
rect 192134 28344 192518 29170
rect 192686 28344 193162 29170
rect 193330 28344 193714 29170
rect 193882 28344 194358 29170
rect 194526 28344 194910 29170
rect 195078 28344 195462 29170
rect 195630 28344 196106 29170
rect 196274 28344 196658 29170
rect 196826 28344 197302 29170
rect 197470 28344 197854 29170
rect 198022 28344 198406 29170
rect 198574 28344 199050 29170
rect 199218 28344 199602 29170
rect 199770 28344 199804 29170
rect 112 856 199804 28344
rect 222 2 330 856
rect 498 2 606 856
rect 774 2 882 856
rect 1050 2 1158 856
rect 1326 2 1434 856
rect 1602 2 1710 856
rect 1878 2 1986 856
rect 2154 2 2262 856
rect 2430 2 2538 856
rect 2706 2 2814 856
rect 2982 2 3090 856
rect 3258 2 3366 856
rect 3534 2 3642 856
rect 3810 2 3918 856
rect 4086 2 4194 856
rect 4362 2 4470 856
rect 4638 2 4746 856
rect 4914 2 5022 856
rect 5190 2 5298 856
rect 5466 2 5574 856
rect 5742 2 5850 856
rect 6018 2 6126 856
rect 6294 2 6402 856
rect 6570 2 6678 856
rect 6846 2 7046 856
rect 7214 2 7322 856
rect 7490 2 7598 856
rect 7766 2 7874 856
rect 8042 2 8150 856
rect 8318 2 8426 856
rect 8594 2 8702 856
rect 8870 2 8978 856
rect 9146 2 9254 856
rect 9422 2 9530 856
rect 9698 2 9806 856
rect 9974 2 10082 856
rect 10250 2 10358 856
rect 10526 2 10634 856
rect 10802 2 10910 856
rect 11078 2 11186 856
rect 11354 2 11462 856
rect 11630 2 11738 856
rect 11906 2 12014 856
rect 12182 2 12290 856
rect 12458 2 12566 856
rect 12734 2 12842 856
rect 13010 2 13118 856
rect 13286 2 13394 856
rect 13562 2 13670 856
rect 13838 2 14038 856
rect 14206 2 14314 856
rect 14482 2 14590 856
rect 14758 2 14866 856
rect 15034 2 15142 856
rect 15310 2 15418 856
rect 15586 2 15694 856
rect 15862 2 15970 856
rect 16138 2 16246 856
rect 16414 2 16522 856
rect 16690 2 16798 856
rect 16966 2 17074 856
rect 17242 2 17350 856
rect 17518 2 17626 856
rect 17794 2 17902 856
rect 18070 2 18178 856
rect 18346 2 18454 856
rect 18622 2 18730 856
rect 18898 2 19006 856
rect 19174 2 19282 856
rect 19450 2 19558 856
rect 19726 2 19834 856
rect 20002 2 20110 856
rect 20278 2 20386 856
rect 20554 2 20754 856
rect 20922 2 21030 856
rect 21198 2 21306 856
rect 21474 2 21582 856
rect 21750 2 21858 856
rect 22026 2 22134 856
rect 22302 2 22410 856
rect 22578 2 22686 856
rect 22854 2 22962 856
rect 23130 2 23238 856
rect 23406 2 23514 856
rect 23682 2 23790 856
rect 23958 2 24066 856
rect 24234 2 24342 856
rect 24510 2 24618 856
rect 24786 2 24894 856
rect 25062 2 25170 856
rect 25338 2 25446 856
rect 25614 2 25722 856
rect 25890 2 25998 856
rect 26166 2 26274 856
rect 26442 2 26550 856
rect 26718 2 26826 856
rect 26994 2 27102 856
rect 27270 2 27378 856
rect 27546 2 27746 856
rect 27914 2 28022 856
rect 28190 2 28298 856
rect 28466 2 28574 856
rect 28742 2 28850 856
rect 29018 2 29126 856
rect 29294 2 29402 856
rect 29570 2 29678 856
rect 29846 2 29954 856
rect 30122 2 30230 856
rect 30398 2 30506 856
rect 30674 2 30782 856
rect 30950 2 31058 856
rect 31226 2 31334 856
rect 31502 2 31610 856
rect 31778 2 31886 856
rect 32054 2 32162 856
rect 32330 2 32438 856
rect 32606 2 32714 856
rect 32882 2 32990 856
rect 33158 2 33266 856
rect 33434 2 33542 856
rect 33710 2 33818 856
rect 33986 2 34094 856
rect 34262 2 34370 856
rect 34538 2 34738 856
rect 34906 2 35014 856
rect 35182 2 35290 856
rect 35458 2 35566 856
rect 35734 2 35842 856
rect 36010 2 36118 856
rect 36286 2 36394 856
rect 36562 2 36670 856
rect 36838 2 36946 856
rect 37114 2 37222 856
rect 37390 2 37498 856
rect 37666 2 37774 856
rect 37942 2 38050 856
rect 38218 2 38326 856
rect 38494 2 38602 856
rect 38770 2 38878 856
rect 39046 2 39154 856
rect 39322 2 39430 856
rect 39598 2 39706 856
rect 39874 2 39982 856
rect 40150 2 40258 856
rect 40426 2 40534 856
rect 40702 2 40810 856
rect 40978 2 41086 856
rect 41254 2 41454 856
rect 41622 2 41730 856
rect 41898 2 42006 856
rect 42174 2 42282 856
rect 42450 2 42558 856
rect 42726 2 42834 856
rect 43002 2 43110 856
rect 43278 2 43386 856
rect 43554 2 43662 856
rect 43830 2 43938 856
rect 44106 2 44214 856
rect 44382 2 44490 856
rect 44658 2 44766 856
rect 44934 2 45042 856
rect 45210 2 45318 856
rect 45486 2 45594 856
rect 45762 2 45870 856
rect 46038 2 46146 856
rect 46314 2 46422 856
rect 46590 2 46698 856
rect 46866 2 46974 856
rect 47142 2 47250 856
rect 47418 2 47526 856
rect 47694 2 47802 856
rect 47970 2 48078 856
rect 48246 2 48446 856
rect 48614 2 48722 856
rect 48890 2 48998 856
rect 49166 2 49274 856
rect 49442 2 49550 856
rect 49718 2 49826 856
rect 49994 2 50102 856
rect 50270 2 50378 856
rect 50546 2 50654 856
rect 50822 2 50930 856
rect 51098 2 51206 856
rect 51374 2 51482 856
rect 51650 2 51758 856
rect 51926 2 52034 856
rect 52202 2 52310 856
rect 52478 2 52586 856
rect 52754 2 52862 856
rect 53030 2 53138 856
rect 53306 2 53414 856
rect 53582 2 53690 856
rect 53858 2 53966 856
rect 54134 2 54242 856
rect 54410 2 54518 856
rect 54686 2 54794 856
rect 54962 2 55070 856
rect 55238 2 55438 856
rect 55606 2 55714 856
rect 55882 2 55990 856
rect 56158 2 56266 856
rect 56434 2 56542 856
rect 56710 2 56818 856
rect 56986 2 57094 856
rect 57262 2 57370 856
rect 57538 2 57646 856
rect 57814 2 57922 856
rect 58090 2 58198 856
rect 58366 2 58474 856
rect 58642 2 58750 856
rect 58918 2 59026 856
rect 59194 2 59302 856
rect 59470 2 59578 856
rect 59746 2 59854 856
rect 60022 2 60130 856
rect 60298 2 60406 856
rect 60574 2 60682 856
rect 60850 2 60958 856
rect 61126 2 61234 856
rect 61402 2 61510 856
rect 61678 2 61786 856
rect 61954 2 62154 856
rect 62322 2 62430 856
rect 62598 2 62706 856
rect 62874 2 62982 856
rect 63150 2 63258 856
rect 63426 2 63534 856
rect 63702 2 63810 856
rect 63978 2 64086 856
rect 64254 2 64362 856
rect 64530 2 64638 856
rect 64806 2 64914 856
rect 65082 2 65190 856
rect 65358 2 65466 856
rect 65634 2 65742 856
rect 65910 2 66018 856
rect 66186 2 66294 856
rect 66462 2 66570 856
rect 66738 2 66846 856
rect 67014 2 67122 856
rect 67290 2 67398 856
rect 67566 2 67674 856
rect 67842 2 67950 856
rect 68118 2 68226 856
rect 68394 2 68502 856
rect 68670 2 68778 856
rect 68946 2 69146 856
rect 69314 2 69422 856
rect 69590 2 69698 856
rect 69866 2 69974 856
rect 70142 2 70250 856
rect 70418 2 70526 856
rect 70694 2 70802 856
rect 70970 2 71078 856
rect 71246 2 71354 856
rect 71522 2 71630 856
rect 71798 2 71906 856
rect 72074 2 72182 856
rect 72350 2 72458 856
rect 72626 2 72734 856
rect 72902 2 73010 856
rect 73178 2 73286 856
rect 73454 2 73562 856
rect 73730 2 73838 856
rect 74006 2 74114 856
rect 74282 2 74390 856
rect 74558 2 74666 856
rect 74834 2 74942 856
rect 75110 2 75218 856
rect 75386 2 75494 856
rect 75662 2 75770 856
rect 75938 2 76138 856
rect 76306 2 76414 856
rect 76582 2 76690 856
rect 76858 2 76966 856
rect 77134 2 77242 856
rect 77410 2 77518 856
rect 77686 2 77794 856
rect 77962 2 78070 856
rect 78238 2 78346 856
rect 78514 2 78622 856
rect 78790 2 78898 856
rect 79066 2 79174 856
rect 79342 2 79450 856
rect 79618 2 79726 856
rect 79894 2 80002 856
rect 80170 2 80278 856
rect 80446 2 80554 856
rect 80722 2 80830 856
rect 80998 2 81106 856
rect 81274 2 81382 856
rect 81550 2 81658 856
rect 81826 2 81934 856
rect 82102 2 82210 856
rect 82378 2 82486 856
rect 82654 2 82854 856
rect 83022 2 83130 856
rect 83298 2 83406 856
rect 83574 2 83682 856
rect 83850 2 83958 856
rect 84126 2 84234 856
rect 84402 2 84510 856
rect 84678 2 84786 856
rect 84954 2 85062 856
rect 85230 2 85338 856
rect 85506 2 85614 856
rect 85782 2 85890 856
rect 86058 2 86166 856
rect 86334 2 86442 856
rect 86610 2 86718 856
rect 86886 2 86994 856
rect 87162 2 87270 856
rect 87438 2 87546 856
rect 87714 2 87822 856
rect 87990 2 88098 856
rect 88266 2 88374 856
rect 88542 2 88650 856
rect 88818 2 88926 856
rect 89094 2 89202 856
rect 89370 2 89478 856
rect 89646 2 89846 856
rect 90014 2 90122 856
rect 90290 2 90398 856
rect 90566 2 90674 856
rect 90842 2 90950 856
rect 91118 2 91226 856
rect 91394 2 91502 856
rect 91670 2 91778 856
rect 91946 2 92054 856
rect 92222 2 92330 856
rect 92498 2 92606 856
rect 92774 2 92882 856
rect 93050 2 93158 856
rect 93326 2 93434 856
rect 93602 2 93710 856
rect 93878 2 93986 856
rect 94154 2 94262 856
rect 94430 2 94538 856
rect 94706 2 94814 856
rect 94982 2 95090 856
rect 95258 2 95366 856
rect 95534 2 95642 856
rect 95810 2 95918 856
rect 96086 2 96194 856
rect 96362 2 96470 856
rect 96638 2 96838 856
rect 97006 2 97114 856
rect 97282 2 97390 856
rect 97558 2 97666 856
rect 97834 2 97942 856
rect 98110 2 98218 856
rect 98386 2 98494 856
rect 98662 2 98770 856
rect 98938 2 99046 856
rect 99214 2 99322 856
rect 99490 2 99598 856
rect 99766 2 99874 856
rect 100042 2 100150 856
rect 100318 2 100426 856
rect 100594 2 100702 856
rect 100870 2 100978 856
rect 101146 2 101254 856
rect 101422 2 101530 856
rect 101698 2 101806 856
rect 101974 2 102082 856
rect 102250 2 102358 856
rect 102526 2 102634 856
rect 102802 2 102910 856
rect 103078 2 103186 856
rect 103354 2 103554 856
rect 103722 2 103830 856
rect 103998 2 104106 856
rect 104274 2 104382 856
rect 104550 2 104658 856
rect 104826 2 104934 856
rect 105102 2 105210 856
rect 105378 2 105486 856
rect 105654 2 105762 856
rect 105930 2 106038 856
rect 106206 2 106314 856
rect 106482 2 106590 856
rect 106758 2 106866 856
rect 107034 2 107142 856
rect 107310 2 107418 856
rect 107586 2 107694 856
rect 107862 2 107970 856
rect 108138 2 108246 856
rect 108414 2 108522 856
rect 108690 2 108798 856
rect 108966 2 109074 856
rect 109242 2 109350 856
rect 109518 2 109626 856
rect 109794 2 109902 856
rect 110070 2 110178 856
rect 110346 2 110546 856
rect 110714 2 110822 856
rect 110990 2 111098 856
rect 111266 2 111374 856
rect 111542 2 111650 856
rect 111818 2 111926 856
rect 112094 2 112202 856
rect 112370 2 112478 856
rect 112646 2 112754 856
rect 112922 2 113030 856
rect 113198 2 113306 856
rect 113474 2 113582 856
rect 113750 2 113858 856
rect 114026 2 114134 856
rect 114302 2 114410 856
rect 114578 2 114686 856
rect 114854 2 114962 856
rect 115130 2 115238 856
rect 115406 2 115514 856
rect 115682 2 115790 856
rect 115958 2 116066 856
rect 116234 2 116342 856
rect 116510 2 116618 856
rect 116786 2 116894 856
rect 117062 2 117170 856
rect 117338 2 117538 856
rect 117706 2 117814 856
rect 117982 2 118090 856
rect 118258 2 118366 856
rect 118534 2 118642 856
rect 118810 2 118918 856
rect 119086 2 119194 856
rect 119362 2 119470 856
rect 119638 2 119746 856
rect 119914 2 120022 856
rect 120190 2 120298 856
rect 120466 2 120574 856
rect 120742 2 120850 856
rect 121018 2 121126 856
rect 121294 2 121402 856
rect 121570 2 121678 856
rect 121846 2 121954 856
rect 122122 2 122230 856
rect 122398 2 122506 856
rect 122674 2 122782 856
rect 122950 2 123058 856
rect 123226 2 123334 856
rect 123502 2 123610 856
rect 123778 2 123886 856
rect 124054 2 124254 856
rect 124422 2 124530 856
rect 124698 2 124806 856
rect 124974 2 125082 856
rect 125250 2 125358 856
rect 125526 2 125634 856
rect 125802 2 125910 856
rect 126078 2 126186 856
rect 126354 2 126462 856
rect 126630 2 126738 856
rect 126906 2 127014 856
rect 127182 2 127290 856
rect 127458 2 127566 856
rect 127734 2 127842 856
rect 128010 2 128118 856
rect 128286 2 128394 856
rect 128562 2 128670 856
rect 128838 2 128946 856
rect 129114 2 129222 856
rect 129390 2 129498 856
rect 129666 2 129774 856
rect 129942 2 130050 856
rect 130218 2 130326 856
rect 130494 2 130602 856
rect 130770 2 130878 856
rect 131046 2 131246 856
rect 131414 2 131522 856
rect 131690 2 131798 856
rect 131966 2 132074 856
rect 132242 2 132350 856
rect 132518 2 132626 856
rect 132794 2 132902 856
rect 133070 2 133178 856
rect 133346 2 133454 856
rect 133622 2 133730 856
rect 133898 2 134006 856
rect 134174 2 134282 856
rect 134450 2 134558 856
rect 134726 2 134834 856
rect 135002 2 135110 856
rect 135278 2 135386 856
rect 135554 2 135662 856
rect 135830 2 135938 856
rect 136106 2 136214 856
rect 136382 2 136490 856
rect 136658 2 136766 856
rect 136934 2 137042 856
rect 137210 2 137318 856
rect 137486 2 137594 856
rect 137762 2 137870 856
rect 138038 2 138238 856
rect 138406 2 138514 856
rect 138682 2 138790 856
rect 138958 2 139066 856
rect 139234 2 139342 856
rect 139510 2 139618 856
rect 139786 2 139894 856
rect 140062 2 140170 856
rect 140338 2 140446 856
rect 140614 2 140722 856
rect 140890 2 140998 856
rect 141166 2 141274 856
rect 141442 2 141550 856
rect 141718 2 141826 856
rect 141994 2 142102 856
rect 142270 2 142378 856
rect 142546 2 142654 856
rect 142822 2 142930 856
rect 143098 2 143206 856
rect 143374 2 143482 856
rect 143650 2 143758 856
rect 143926 2 144034 856
rect 144202 2 144310 856
rect 144478 2 144586 856
rect 144754 2 144954 856
rect 145122 2 145230 856
rect 145398 2 145506 856
rect 145674 2 145782 856
rect 145950 2 146058 856
rect 146226 2 146334 856
rect 146502 2 146610 856
rect 146778 2 146886 856
rect 147054 2 147162 856
rect 147330 2 147438 856
rect 147606 2 147714 856
rect 147882 2 147990 856
rect 148158 2 148266 856
rect 148434 2 148542 856
rect 148710 2 148818 856
rect 148986 2 149094 856
rect 149262 2 149370 856
rect 149538 2 149646 856
rect 149814 2 149922 856
rect 150090 2 150198 856
rect 150366 2 150474 856
rect 150642 2 150750 856
rect 150918 2 151026 856
rect 151194 2 151302 856
rect 151470 2 151578 856
rect 151746 2 151946 856
rect 152114 2 152222 856
rect 152390 2 152498 856
rect 152666 2 152774 856
rect 152942 2 153050 856
rect 153218 2 153326 856
rect 153494 2 153602 856
rect 153770 2 153878 856
rect 154046 2 154154 856
rect 154322 2 154430 856
rect 154598 2 154706 856
rect 154874 2 154982 856
rect 155150 2 155258 856
rect 155426 2 155534 856
rect 155702 2 155810 856
rect 155978 2 156086 856
rect 156254 2 156362 856
rect 156530 2 156638 856
rect 156806 2 156914 856
rect 157082 2 157190 856
rect 157358 2 157466 856
rect 157634 2 157742 856
rect 157910 2 158018 856
rect 158186 2 158294 856
rect 158462 2 158570 856
rect 158738 2 158938 856
rect 159106 2 159214 856
rect 159382 2 159490 856
rect 159658 2 159766 856
rect 159934 2 160042 856
rect 160210 2 160318 856
rect 160486 2 160594 856
rect 160762 2 160870 856
rect 161038 2 161146 856
rect 161314 2 161422 856
rect 161590 2 161698 856
rect 161866 2 161974 856
rect 162142 2 162250 856
rect 162418 2 162526 856
rect 162694 2 162802 856
rect 162970 2 163078 856
rect 163246 2 163354 856
rect 163522 2 163630 856
rect 163798 2 163906 856
rect 164074 2 164182 856
rect 164350 2 164458 856
rect 164626 2 164734 856
rect 164902 2 165010 856
rect 165178 2 165286 856
rect 165454 2 165654 856
rect 165822 2 165930 856
rect 166098 2 166206 856
rect 166374 2 166482 856
rect 166650 2 166758 856
rect 166926 2 167034 856
rect 167202 2 167310 856
rect 167478 2 167586 856
rect 167754 2 167862 856
rect 168030 2 168138 856
rect 168306 2 168414 856
rect 168582 2 168690 856
rect 168858 2 168966 856
rect 169134 2 169242 856
rect 169410 2 169518 856
rect 169686 2 169794 856
rect 169962 2 170070 856
rect 170238 2 170346 856
rect 170514 2 170622 856
rect 170790 2 170898 856
rect 171066 2 171174 856
rect 171342 2 171450 856
rect 171618 2 171726 856
rect 171894 2 172002 856
rect 172170 2 172278 856
rect 172446 2 172646 856
rect 172814 2 172922 856
rect 173090 2 173198 856
rect 173366 2 173474 856
rect 173642 2 173750 856
rect 173918 2 174026 856
rect 174194 2 174302 856
rect 174470 2 174578 856
rect 174746 2 174854 856
rect 175022 2 175130 856
rect 175298 2 175406 856
rect 175574 2 175682 856
rect 175850 2 175958 856
rect 176126 2 176234 856
rect 176402 2 176510 856
rect 176678 2 176786 856
rect 176954 2 177062 856
rect 177230 2 177338 856
rect 177506 2 177614 856
rect 177782 2 177890 856
rect 178058 2 178166 856
rect 178334 2 178442 856
rect 178610 2 178718 856
rect 178886 2 178994 856
rect 179162 2 179270 856
rect 179438 2 179638 856
rect 179806 2 179914 856
rect 180082 2 180190 856
rect 180358 2 180466 856
rect 180634 2 180742 856
rect 180910 2 181018 856
rect 181186 2 181294 856
rect 181462 2 181570 856
rect 181738 2 181846 856
rect 182014 2 182122 856
rect 182290 2 182398 856
rect 182566 2 182674 856
rect 182842 2 182950 856
rect 183118 2 183226 856
rect 183394 2 183502 856
rect 183670 2 183778 856
rect 183946 2 184054 856
rect 184222 2 184330 856
rect 184498 2 184606 856
rect 184774 2 184882 856
rect 185050 2 185158 856
rect 185326 2 185434 856
rect 185602 2 185710 856
rect 185878 2 185986 856
rect 186154 2 186354 856
rect 186522 2 186630 856
rect 186798 2 186906 856
rect 187074 2 187182 856
rect 187350 2 187458 856
rect 187626 2 187734 856
rect 187902 2 188010 856
rect 188178 2 188286 856
rect 188454 2 188562 856
rect 188730 2 188838 856
rect 189006 2 189114 856
rect 189282 2 189390 856
rect 189558 2 189666 856
rect 189834 2 189942 856
rect 190110 2 190218 856
rect 190386 2 190494 856
rect 190662 2 190770 856
rect 190938 2 191046 856
rect 191214 2 191322 856
rect 191490 2 191598 856
rect 191766 2 191874 856
rect 192042 2 192150 856
rect 192318 2 192426 856
rect 192594 2 192702 856
rect 192870 2 192978 856
rect 193146 2 193346 856
rect 193514 2 193622 856
rect 193790 2 193898 856
rect 194066 2 194174 856
rect 194342 2 194450 856
rect 194618 2 194726 856
rect 194894 2 195002 856
rect 195170 2 195278 856
rect 195446 2 195554 856
rect 195722 2 195830 856
rect 195998 2 196106 856
rect 196274 2 196382 856
rect 196550 2 196658 856
rect 196826 2 196934 856
rect 197102 2 197210 856
rect 197378 2 197486 856
rect 197654 2 197762 856
rect 197930 2 198038 856
rect 198206 2 198314 856
rect 198482 2 198590 856
rect 198758 2 198866 856
rect 199034 2 199142 856
rect 199310 2 199418 856
rect 199586 2 199694 856
<< metal3 >>
rect -2762 31430 202678 31610
rect -2498 31166 202414 31346
rect -2234 30902 202150 31082
rect -1970 30638 201886 30818
rect -1706 30374 201622 30554
rect -1442 30110 201358 30290
rect -1178 29846 201094 30026
rect -914 29582 200830 29762
rect -650 29318 200566 29498
rect -386 29054 200302 29234
rect -400 24216 800 24336
rect -400 14424 800 14544
rect -400 4768 800 4888
rect -386 -402 200302 -222
rect -650 -666 200566 -486
rect -914 -930 200830 -750
rect -1178 -1194 201094 -1014
rect -1442 -1458 201358 -1278
rect -1706 -1722 201622 -1542
rect -1970 -1986 201886 -1806
rect -2234 -2250 202150 -2070
rect -2498 -2514 202414 -2334
rect -2762 -2778 202678 -2598
<< obsm3 >>
rect 800 24416 197728 28933
rect 880 24136 197728 24416
rect 800 14624 197728 24136
rect 880 14344 197728 14624
rect 800 4968 197728 14344
rect 880 4688 197728 4968
rect 800 35 197728 4688
<< metal4 >>
rect -2762 -2778 -2582 31610
rect -2498 -2514 -2318 31346
rect -2234 -2250 -2054 31082
rect -1970 -1986 -1790 30818
rect -1706 -1722 -1526 30554
rect -1442 -1458 -1262 30290
rect -1178 -1194 -998 30026
rect -914 -930 -734 29762
rect -650 -666 -470 29498
rect -386 -402 -206 29234
rect 4014 -666 4194 29498
rect 4834 -1194 5014 30026
rect 5654 -1722 5834 30554
rect 6474 -2250 6654 31082
rect 7294 -2778 7474 31610
rect 18514 -666 18694 29498
rect 19334 -1194 19514 30026
rect 20154 -1722 20334 30554
rect 20974 -2250 21154 31082
rect 21794 -2778 21974 31610
rect 33014 -666 33194 29498
rect 33834 -1194 34014 30026
rect 34654 -1722 34834 30554
rect 35474 -2250 35654 31082
rect 36294 -2778 36474 31610
rect 47514 -666 47694 29498
rect 48334 -1194 48514 30026
rect 49154 -1722 49334 30554
rect 49974 -2250 50154 31082
rect 50794 -2778 50974 31610
rect 62014 -666 62194 29498
rect 62834 -1194 63014 30026
rect 63654 -1722 63834 30554
rect 64474 -2250 64654 31082
rect 65294 -2778 65474 31610
rect 76514 -666 76694 29498
rect 77334 -1194 77514 30026
rect 78154 -1722 78334 30554
rect 78974 -2250 79154 31082
rect 79794 -2778 79974 31610
rect 91014 -666 91194 29498
rect 91834 -1194 92014 30026
rect 92654 -1722 92834 30554
rect 93474 -2250 93654 31082
rect 94294 -2778 94474 31610
rect 105514 -666 105694 29498
rect 106334 -1194 106514 30026
rect 107154 -1722 107334 30554
rect 107974 -2250 108154 31082
rect 108794 -2778 108974 31610
rect 120014 -666 120194 29498
rect 120834 -1194 121014 30026
rect 121654 -1722 121834 30554
rect 122474 -2250 122654 31082
rect 123294 -2778 123474 31610
rect 134514 -666 134694 29498
rect 135334 -1194 135514 30026
rect 136154 -1722 136334 30554
rect 136974 -2250 137154 31082
rect 137794 -2778 137974 31610
rect 149014 -666 149194 29498
rect 149834 -1194 150014 30026
rect 150654 -1722 150834 30554
rect 151474 -2250 151654 31082
rect 152294 -2778 152474 31610
rect 163514 -666 163694 29498
rect 164334 -1194 164514 30026
rect 165154 -1722 165334 30554
rect 165974 -2250 166154 31082
rect 166794 -2778 166974 31610
rect 178014 -666 178194 29498
rect 178834 -1194 179014 30026
rect 179654 -1722 179834 30554
rect 180474 -2250 180654 31082
rect 181294 -2778 181474 31610
rect 192514 -666 192694 29498
rect 193334 -1194 193514 30026
rect 194154 -1722 194334 30554
rect 194974 -2250 195154 31082
rect 195794 -2778 195974 31610
rect 200122 -402 200302 29234
rect 200386 -666 200566 29498
rect 200650 -930 200830 29762
rect 200914 -1194 201094 30026
rect 201178 -1458 201358 30290
rect 201442 -1722 201622 30554
rect 201706 -1986 201886 30818
rect 201970 -2250 202150 31082
rect 202234 -2514 202414 31346
rect 202498 -2778 202678 31610
<< obsm4 >>
rect 5211 851 5574 28933
rect 5914 851 6394 28933
rect 6734 851 7214 28933
rect 7554 851 18434 28933
rect 18774 851 19254 28933
rect 19594 851 20074 28933
rect 20414 851 20894 28933
rect 21234 851 21714 28933
rect 22054 851 32934 28933
rect 33274 851 33754 28933
rect 34094 851 34574 28933
rect 34914 851 35394 28933
rect 35734 851 36214 28933
rect 36554 851 47434 28933
rect 47774 851 48254 28933
rect 48594 851 49074 28933
rect 49414 851 49894 28933
rect 50234 851 50714 28933
rect 51054 851 61934 28933
rect 62274 851 62754 28933
rect 63094 851 63574 28933
rect 63914 851 64394 28933
rect 64734 851 65214 28933
rect 65554 851 76434 28933
rect 76774 851 77254 28933
rect 77594 851 78074 28933
rect 78414 851 78894 28933
rect 79234 851 79714 28933
rect 80054 851 90934 28933
rect 91274 851 91754 28933
rect 92094 851 92574 28933
rect 92914 851 93394 28933
rect 93734 851 94214 28933
rect 94554 851 105434 28933
rect 105774 851 106254 28933
rect 106594 851 107074 28933
rect 107414 851 107894 28933
rect 108234 851 108714 28933
rect 109054 851 119934 28933
rect 120274 851 120754 28933
rect 121094 851 121574 28933
rect 121914 851 122394 28933
rect 122734 851 123214 28933
rect 123554 851 134434 28933
rect 134774 851 135254 28933
rect 135594 851 136074 28933
rect 136414 851 136894 28933
rect 137234 851 137714 28933
rect 138054 851 148934 28933
rect 149274 851 149754 28933
rect 150094 851 150574 28933
rect 150914 851 151394 28933
rect 151734 851 152214 28933
rect 152554 851 163434 28933
rect 163774 851 164254 28933
rect 164594 851 165074 28933
rect 165414 851 165894 28933
rect 166234 851 166714 28933
rect 167054 851 177934 28933
rect 178274 851 178754 28933
rect 179094 851 179574 28933
rect 179914 851 180394 28933
rect 180734 851 181214 28933
rect 181554 851 192434 28933
rect 192774 851 193254 28933
rect 193594 851 194074 28933
rect 194414 851 194894 28933
rect 195234 851 195533 28933
<< labels >>
rlabel metal3 s -400 4768 800 4888 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s -400 14424 800 14544 6 caravel_clk2
port 2 nsew signal input
rlabel metal3 s -400 24216 800 24336 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 7930 28400 7986 29600 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 66718 28400 66774 29600 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 67270 28400 67326 29600 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 67914 28400 67970 29600 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 68466 28400 68522 29600 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 69110 28400 69166 29600 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 69662 28400 69718 29600 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 70214 28400 70270 29600 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 70858 28400 70914 29600 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 71410 28400 71466 29600 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 72054 28400 72110 29600 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 13818 28400 13874 29600 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 72606 28400 72662 29600 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 73158 28400 73214 29600 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 73802 28400 73858 29600 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 74354 28400 74410 29600 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 74998 28400 75054 29600 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 75550 28400 75606 29600 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 76102 28400 76158 29600 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 76746 28400 76802 29600 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 77298 28400 77354 29600 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 77942 28400 77998 29600 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 14370 28400 14426 29600 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 78494 28400 78550 29600 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 79046 28400 79102 29600 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 79690 28400 79746 29600 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 80242 28400 80298 29600 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 80794 28400 80850 29600 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 81438 28400 81494 29600 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 81990 28400 82046 29600 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 82634 28400 82690 29600 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 14922 28400 14978 29600 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 15566 28400 15622 29600 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 16118 28400 16174 29600 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 16762 28400 16818 29600 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 17314 28400 17370 29600 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 17866 28400 17922 29600 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 18510 28400 18566 29600 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 19062 28400 19118 29600 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 8482 28400 8538 29600 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 19706 28400 19762 29600 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 20258 28400 20314 29600 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 20810 28400 20866 29600 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 21454 28400 21510 29600 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 22006 28400 22062 29600 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 22558 28400 22614 29600 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 23202 28400 23258 29600 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 23754 28400 23810 29600 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 24398 28400 24454 29600 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 24950 28400 25006 29600 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 9034 28400 9090 29600 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 25502 28400 25558 29600 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 26146 28400 26202 29600 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 26698 28400 26754 29600 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 27342 28400 27398 29600 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 27894 28400 27950 29600 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 28446 28400 28502 29600 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 29090 28400 29146 29600 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 29642 28400 29698 29600 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 30286 28400 30342 29600 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 30838 28400 30894 29600 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 9678 28400 9734 29600 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 31390 28400 31446 29600 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 32034 28400 32090 29600 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 32586 28400 32642 29600 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 33230 28400 33286 29600 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 33782 28400 33838 29600 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 34334 28400 34390 29600 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 34978 28400 35034 29600 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 35530 28400 35586 29600 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 36174 28400 36230 29600 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 36726 28400 36782 29600 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 10230 28400 10286 29600 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 37278 28400 37334 29600 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 37922 28400 37978 29600 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 38474 28400 38530 29600 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 39118 28400 39174 29600 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 39670 28400 39726 29600 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 40222 28400 40278 29600 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 40866 28400 40922 29600 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 41418 28400 41474 29600 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 41970 28400 42026 29600 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 42614 28400 42670 29600 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 10874 28400 10930 29600 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 43166 28400 43222 29600 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 43810 28400 43866 29600 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 44362 28400 44418 29600 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 44914 28400 44970 29600 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 45558 28400 45614 29600 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 46110 28400 46166 29600 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 46754 28400 46810 29600 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 47306 28400 47362 29600 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 47858 28400 47914 29600 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 48502 28400 48558 29600 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 11426 28400 11482 29600 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 49054 28400 49110 29600 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 49698 28400 49754 29600 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 50250 28400 50306 29600 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 50802 28400 50858 29600 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 51446 28400 51502 29600 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 51998 28400 52054 29600 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 52642 28400 52698 29600 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 53194 28400 53250 29600 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 53746 28400 53802 29600 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 54390 28400 54446 29600 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 11978 28400 12034 29600 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 54942 28400 54998 29600 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 55586 28400 55642 29600 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 56138 28400 56194 29600 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 56690 28400 56746 29600 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 57334 28400 57390 29600 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 57886 28400 57942 29600 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 58530 28400 58586 29600 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 59082 28400 59138 29600 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 59634 28400 59690 29600 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 60278 28400 60334 29600 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 12622 28400 12678 29600 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 60830 28400 60886 29600 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 61382 28400 61438 29600 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 62026 28400 62082 29600 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 62578 28400 62634 29600 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 63222 28400 63278 29600 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 63774 28400 63830 29600 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 64326 28400 64382 29600 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 64970 28400 65026 29600 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 65522 28400 65578 29600 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 66166 28400 66222 29600 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 13174 28400 13230 29600 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 35898 -400 35954 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 63866 -400 63922 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 64142 -400 64198 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 64418 -400 64474 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 64694 -400 64750 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 64970 -400 65026 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 65246 -400 65302 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 65522 -400 65578 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 65798 -400 65854 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 66074 -400 66130 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 66350 -400 66406 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 38658 -400 38714 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 66626 -400 66682 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 66902 -400 66958 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 67178 -400 67234 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 67454 -400 67510 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 67730 -400 67786 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 68006 -400 68062 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 68282 -400 68338 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 68558 -400 68614 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 68834 -400 68890 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 69202 -400 69258 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 38934 -400 38990 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 69478 -400 69534 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 69754 -400 69810 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 70030 -400 70086 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 70306 -400 70362 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 70582 -400 70638 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 70858 -400 70914 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 71134 -400 71190 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 71410 -400 71466 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 39210 -400 39266 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 39486 -400 39542 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 39762 -400 39818 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 40038 -400 40094 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 40314 -400 40370 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 40590 -400 40646 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 40866 -400 40922 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 41142 -400 41198 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 36174 -400 36230 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 41510 -400 41566 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 41786 -400 41842 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 42062 -400 42118 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 42338 -400 42394 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 42614 -400 42670 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 42890 -400 42946 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 43166 -400 43222 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 43442 -400 43498 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 43718 -400 43774 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 43994 -400 44050 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 36450 -400 36506 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 44270 -400 44326 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 44546 -400 44602 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 44822 -400 44878 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 45098 -400 45154 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 45374 -400 45430 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 45650 -400 45706 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 45926 -400 45982 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 46202 -400 46258 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 46478 -400 46534 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 46754 -400 46810 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 36726 -400 36782 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 47030 -400 47086 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 47306 -400 47362 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 47582 -400 47638 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 47858 -400 47914 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 48134 -400 48190 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 48502 -400 48558 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 48778 -400 48834 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 49054 -400 49110 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 49330 -400 49386 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 49606 -400 49662 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 37002 -400 37058 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 49882 -400 49938 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 50158 -400 50214 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 50434 -400 50490 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 50710 -400 50766 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 50986 -400 51042 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 51262 -400 51318 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 51538 -400 51594 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 51814 -400 51870 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 52090 -400 52146 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 52366 -400 52422 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 37278 -400 37334 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 52642 -400 52698 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 52918 -400 52974 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 53194 -400 53250 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 53470 -400 53526 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 53746 -400 53802 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 54022 -400 54078 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 54298 -400 54354 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 54574 -400 54630 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 54850 -400 54906 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 55126 -400 55182 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 37554 -400 37610 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 55494 -400 55550 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 55770 -400 55826 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 56046 -400 56102 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 56322 -400 56378 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 56598 -400 56654 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 56874 -400 56930 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 57150 -400 57206 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 57426 -400 57482 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 57702 -400 57758 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 57978 -400 58034 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 37830 -400 37886 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 58254 -400 58310 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 58530 -400 58586 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 58806 -400 58862 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 59082 -400 59138 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 59358 -400 59414 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 59634 -400 59690 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 59910 -400 59966 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 60186 -400 60242 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 60462 -400 60518 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 60738 -400 60794 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 38106 -400 38162 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 61014 -400 61070 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 61290 -400 61346 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 61566 -400 61622 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 61842 -400 61898 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 62210 -400 62266 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 62486 -400 62542 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 62762 -400 62818 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 63038 -400 63094 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 63314 -400 63370 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 63590 -400 63646 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 38382 -400 38438 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 83186 28400 83242 29600 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 141974 28400 142030 29600 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 142618 28400 142674 29600 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 143170 28400 143226 29600 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 143814 28400 143870 29600 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 144366 28400 144422 29600 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 144918 28400 144974 29600 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 145562 28400 145618 29600 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 146114 28400 146170 29600 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 146758 28400 146814 29600 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 147310 28400 147366 29600 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 89074 28400 89130 29600 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 147862 28400 147918 29600 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 148506 28400 148562 29600 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 149058 28400 149114 29600 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 149702 28400 149758 29600 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 150254 28400 150310 29600 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 150806 28400 150862 29600 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 151450 28400 151506 29600 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 152002 28400 152058 29600 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 152646 28400 152702 29600 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 153198 28400 153254 29600 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 89626 28400 89682 29600 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 153750 28400 153806 29600 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 154394 28400 154450 29600 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 154946 28400 155002 29600 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 155590 28400 155646 29600 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 156142 28400 156198 29600 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 156694 28400 156750 29600 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 157338 28400 157394 29600 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 157890 28400 157946 29600 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 90270 28400 90326 29600 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 90822 28400 90878 29600 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 91466 28400 91522 29600 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 92018 28400 92074 29600 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 92570 28400 92626 29600 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 93214 28400 93270 29600 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 93766 28400 93822 29600 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 94410 28400 94466 29600 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 83738 28400 83794 29600 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 94962 28400 95018 29600 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 95514 28400 95570 29600 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 96158 28400 96214 29600 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 96710 28400 96766 29600 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 97354 28400 97410 29600 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 97906 28400 97962 29600 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 98458 28400 98514 29600 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 99102 28400 99158 29600 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 99654 28400 99710 29600 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 100298 28400 100354 29600 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 84382 28400 84438 29600 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 100850 28400 100906 29600 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 101402 28400 101458 29600 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 102046 28400 102102 29600 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 102598 28400 102654 29600 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 103150 28400 103206 29600 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 103794 28400 103850 29600 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 104346 28400 104402 29600 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 104990 28400 105046 29600 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 105542 28400 105598 29600 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 106094 28400 106150 29600 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 84934 28400 84990 29600 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 106738 28400 106794 29600 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 107290 28400 107346 29600 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 107934 28400 107990 29600 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 108486 28400 108542 29600 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 109038 28400 109094 29600 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 109682 28400 109738 29600 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 110234 28400 110290 29600 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 110878 28400 110934 29600 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 111430 28400 111486 29600 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 111982 28400 112038 29600 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 85578 28400 85634 29600 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 112626 28400 112682 29600 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 113178 28400 113234 29600 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 113822 28400 113878 29600 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 114374 28400 114430 29600 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 114926 28400 114982 29600 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 115570 28400 115626 29600 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 116122 28400 116178 29600 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 116766 28400 116822 29600 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 117318 28400 117374 29600 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 117870 28400 117926 29600 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 86130 28400 86186 29600 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 118514 28400 118570 29600 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 119066 28400 119122 29600 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 119710 28400 119766 29600 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 120262 28400 120318 29600 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 120814 28400 120870 29600 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 121458 28400 121514 29600 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 122010 28400 122066 29600 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 122562 28400 122618 29600 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 123206 28400 123262 29600 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 123758 28400 123814 29600 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 86682 28400 86738 29600 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 124402 28400 124458 29600 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 124954 28400 125010 29600 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 125506 28400 125562 29600 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 126150 28400 126206 29600 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 126702 28400 126758 29600 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 127346 28400 127402 29600 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 127898 28400 127954 29600 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 128450 28400 128506 29600 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 129094 28400 129150 29600 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 129646 28400 129702 29600 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 87326 28400 87382 29600 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 130290 28400 130346 29600 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 130842 28400 130898 29600 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 131394 28400 131450 29600 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 132038 28400 132094 29600 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 132590 28400 132646 29600 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 133234 28400 133290 29600 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 133786 28400 133842 29600 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 134338 28400 134394 29600 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 134982 28400 135038 29600 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 135534 28400 135590 29600 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 87878 28400 87934 29600 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 136178 28400 136234 29600 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 136730 28400 136786 29600 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 137282 28400 137338 29600 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 137926 28400 137982 29600 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 138478 28400 138534 29600 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 139122 28400 139178 29600 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 139674 28400 139730 29600 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 140226 28400 140282 29600 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 140870 28400 140926 29600 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 141422 28400 141478 29600 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 88522 28400 88578 29600 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 110 -400 166 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 28078 -400 28134 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 28354 -400 28410 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 28630 -400 28686 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 28906 -400 28962 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 29182 -400 29238 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 29458 -400 29514 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 29734 -400 29790 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 30010 -400 30066 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 30286 -400 30342 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 30562 -400 30618 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 2870 -400 2926 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 30838 -400 30894 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 31114 -400 31170 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 31390 -400 31446 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 31666 -400 31722 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 31942 -400 31998 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 32218 -400 32274 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 32494 -400 32550 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 32770 -400 32826 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 33046 -400 33102 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 33322 -400 33378 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 3146 -400 3202 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 33598 -400 33654 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 33874 -400 33930 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 34150 -400 34206 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 34426 -400 34482 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 34794 -400 34850 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 35070 -400 35126 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 35346 -400 35402 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 35622 -400 35678 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 3422 -400 3478 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 3698 -400 3754 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 3974 -400 4030 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 4250 -400 4306 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 4526 -400 4582 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 4802 -400 4858 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 5078 -400 5134 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 5354 -400 5410 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 386 -400 442 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 5630 -400 5686 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 5906 -400 5962 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 6182 -400 6238 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 6458 -400 6514 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 6734 -400 6790 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 7102 -400 7158 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 7378 -400 7434 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 7654 -400 7710 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 7930 -400 7986 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 8206 -400 8262 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 662 -400 718 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 8482 -400 8538 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 8758 -400 8814 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 9034 -400 9090 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 9310 -400 9366 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 9586 -400 9642 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 9862 -400 9918 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 10138 -400 10194 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 10414 -400 10470 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 10690 -400 10746 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 10966 -400 11022 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 938 -400 994 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 11242 -400 11298 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 11518 -400 11574 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 11794 -400 11850 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 12070 -400 12126 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 12346 -400 12402 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 12622 -400 12678 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 12898 -400 12954 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 13174 -400 13230 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 13450 -400 13506 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 13726 -400 13782 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 1214 -400 1270 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 14094 -400 14150 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 14370 -400 14426 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 14646 -400 14702 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 14922 -400 14978 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 15198 -400 15254 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 15474 -400 15530 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 15750 -400 15806 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 16026 -400 16082 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 16302 -400 16358 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 16578 -400 16634 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 1490 -400 1546 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 16854 -400 16910 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 17130 -400 17186 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 17406 -400 17462 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 17682 -400 17738 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 17958 -400 18014 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 18234 -400 18290 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 18510 -400 18566 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 18786 -400 18842 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 19062 -400 19118 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 19338 -400 19394 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 1766 -400 1822 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 19614 -400 19670 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 19890 -400 19946 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 20166 -400 20222 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 20442 -400 20498 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 20810 -400 20866 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 21086 -400 21142 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 21362 -400 21418 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 21638 -400 21694 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 21914 -400 21970 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 22190 -400 22246 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 2042 -400 2098 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 22466 -400 22522 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 22742 -400 22798 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 23018 -400 23074 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 23294 -400 23350 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 23570 -400 23626 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 23846 -400 23902 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 24122 -400 24178 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 24398 -400 24454 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 24674 -400 24730 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 24950 -400 25006 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 2318 -400 2374 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 25226 -400 25282 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 25502 -400 25558 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 25778 -400 25834 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 26054 -400 26110 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 26330 -400 26386 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 26606 -400 26662 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 26882 -400 26938 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 27158 -400 27214 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 27434 -400 27490 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 27802 -400 27858 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 2594 -400 2650 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 107474 -400 107530 800 6 la_iena_mprj[0]
port 516 nsew signal input
rlabel metal2 s 135442 -400 135498 800 6 la_iena_mprj[100]
port 517 nsew signal input
rlabel metal2 s 135718 -400 135774 800 6 la_iena_mprj[101]
port 518 nsew signal input
rlabel metal2 s 135994 -400 136050 800 6 la_iena_mprj[102]
port 519 nsew signal input
rlabel metal2 s 136270 -400 136326 800 6 la_iena_mprj[103]
port 520 nsew signal input
rlabel metal2 s 136546 -400 136602 800 6 la_iena_mprj[104]
port 521 nsew signal input
rlabel metal2 s 136822 -400 136878 800 6 la_iena_mprj[105]
port 522 nsew signal input
rlabel metal2 s 137098 -400 137154 800 6 la_iena_mprj[106]
port 523 nsew signal input
rlabel metal2 s 137374 -400 137430 800 6 la_iena_mprj[107]
port 524 nsew signal input
rlabel metal2 s 137650 -400 137706 800 6 la_iena_mprj[108]
port 525 nsew signal input
rlabel metal2 s 137926 -400 137982 800 6 la_iena_mprj[109]
port 526 nsew signal input
rlabel metal2 s 110234 -400 110290 800 6 la_iena_mprj[10]
port 527 nsew signal input
rlabel metal2 s 138294 -400 138350 800 6 la_iena_mprj[110]
port 528 nsew signal input
rlabel metal2 s 138570 -400 138626 800 6 la_iena_mprj[111]
port 529 nsew signal input
rlabel metal2 s 138846 -400 138902 800 6 la_iena_mprj[112]
port 530 nsew signal input
rlabel metal2 s 139122 -400 139178 800 6 la_iena_mprj[113]
port 531 nsew signal input
rlabel metal2 s 139398 -400 139454 800 6 la_iena_mprj[114]
port 532 nsew signal input
rlabel metal2 s 139674 -400 139730 800 6 la_iena_mprj[115]
port 533 nsew signal input
rlabel metal2 s 139950 -400 140006 800 6 la_iena_mprj[116]
port 534 nsew signal input
rlabel metal2 s 140226 -400 140282 800 6 la_iena_mprj[117]
port 535 nsew signal input
rlabel metal2 s 140502 -400 140558 800 6 la_iena_mprj[118]
port 536 nsew signal input
rlabel metal2 s 140778 -400 140834 800 6 la_iena_mprj[119]
port 537 nsew signal input
rlabel metal2 s 110602 -400 110658 800 6 la_iena_mprj[11]
port 538 nsew signal input
rlabel metal2 s 141054 -400 141110 800 6 la_iena_mprj[120]
port 539 nsew signal input
rlabel metal2 s 141330 -400 141386 800 6 la_iena_mprj[121]
port 540 nsew signal input
rlabel metal2 s 141606 -400 141662 800 6 la_iena_mprj[122]
port 541 nsew signal input
rlabel metal2 s 141882 -400 141938 800 6 la_iena_mprj[123]
port 542 nsew signal input
rlabel metal2 s 142158 -400 142214 800 6 la_iena_mprj[124]
port 543 nsew signal input
rlabel metal2 s 142434 -400 142490 800 6 la_iena_mprj[125]
port 544 nsew signal input
rlabel metal2 s 142710 -400 142766 800 6 la_iena_mprj[126]
port 545 nsew signal input
rlabel metal2 s 142986 -400 143042 800 6 la_iena_mprj[127]
port 546 nsew signal input
rlabel metal2 s 110878 -400 110934 800 6 la_iena_mprj[12]
port 547 nsew signal input
rlabel metal2 s 111154 -400 111210 800 6 la_iena_mprj[13]
port 548 nsew signal input
rlabel metal2 s 111430 -400 111486 800 6 la_iena_mprj[14]
port 549 nsew signal input
rlabel metal2 s 111706 -400 111762 800 6 la_iena_mprj[15]
port 550 nsew signal input
rlabel metal2 s 111982 -400 112038 800 6 la_iena_mprj[16]
port 551 nsew signal input
rlabel metal2 s 112258 -400 112314 800 6 la_iena_mprj[17]
port 552 nsew signal input
rlabel metal2 s 112534 -400 112590 800 6 la_iena_mprj[18]
port 553 nsew signal input
rlabel metal2 s 112810 -400 112866 800 6 la_iena_mprj[19]
port 554 nsew signal input
rlabel metal2 s 107750 -400 107806 800 6 la_iena_mprj[1]
port 555 nsew signal input
rlabel metal2 s 113086 -400 113142 800 6 la_iena_mprj[20]
port 556 nsew signal input
rlabel metal2 s 113362 -400 113418 800 6 la_iena_mprj[21]
port 557 nsew signal input
rlabel metal2 s 113638 -400 113694 800 6 la_iena_mprj[22]
port 558 nsew signal input
rlabel metal2 s 113914 -400 113970 800 6 la_iena_mprj[23]
port 559 nsew signal input
rlabel metal2 s 114190 -400 114246 800 6 la_iena_mprj[24]
port 560 nsew signal input
rlabel metal2 s 114466 -400 114522 800 6 la_iena_mprj[25]
port 561 nsew signal input
rlabel metal2 s 114742 -400 114798 800 6 la_iena_mprj[26]
port 562 nsew signal input
rlabel metal2 s 115018 -400 115074 800 6 la_iena_mprj[27]
port 563 nsew signal input
rlabel metal2 s 115294 -400 115350 800 6 la_iena_mprj[28]
port 564 nsew signal input
rlabel metal2 s 115570 -400 115626 800 6 la_iena_mprj[29]
port 565 nsew signal input
rlabel metal2 s 108026 -400 108082 800 6 la_iena_mprj[2]
port 566 nsew signal input
rlabel metal2 s 115846 -400 115902 800 6 la_iena_mprj[30]
port 567 nsew signal input
rlabel metal2 s 116122 -400 116178 800 6 la_iena_mprj[31]
port 568 nsew signal input
rlabel metal2 s 116398 -400 116454 800 6 la_iena_mprj[32]
port 569 nsew signal input
rlabel metal2 s 116674 -400 116730 800 6 la_iena_mprj[33]
port 570 nsew signal input
rlabel metal2 s 116950 -400 117006 800 6 la_iena_mprj[34]
port 571 nsew signal input
rlabel metal2 s 117226 -400 117282 800 6 la_iena_mprj[35]
port 572 nsew signal input
rlabel metal2 s 117594 -400 117650 800 6 la_iena_mprj[36]
port 573 nsew signal input
rlabel metal2 s 117870 -400 117926 800 6 la_iena_mprj[37]
port 574 nsew signal input
rlabel metal2 s 118146 -400 118202 800 6 la_iena_mprj[38]
port 575 nsew signal input
rlabel metal2 s 118422 -400 118478 800 6 la_iena_mprj[39]
port 576 nsew signal input
rlabel metal2 s 108302 -400 108358 800 6 la_iena_mprj[3]
port 577 nsew signal input
rlabel metal2 s 118698 -400 118754 800 6 la_iena_mprj[40]
port 578 nsew signal input
rlabel metal2 s 118974 -400 119030 800 6 la_iena_mprj[41]
port 579 nsew signal input
rlabel metal2 s 119250 -400 119306 800 6 la_iena_mprj[42]
port 580 nsew signal input
rlabel metal2 s 119526 -400 119582 800 6 la_iena_mprj[43]
port 581 nsew signal input
rlabel metal2 s 119802 -400 119858 800 6 la_iena_mprj[44]
port 582 nsew signal input
rlabel metal2 s 120078 -400 120134 800 6 la_iena_mprj[45]
port 583 nsew signal input
rlabel metal2 s 120354 -400 120410 800 6 la_iena_mprj[46]
port 584 nsew signal input
rlabel metal2 s 120630 -400 120686 800 6 la_iena_mprj[47]
port 585 nsew signal input
rlabel metal2 s 120906 -400 120962 800 6 la_iena_mprj[48]
port 586 nsew signal input
rlabel metal2 s 121182 -400 121238 800 6 la_iena_mprj[49]
port 587 nsew signal input
rlabel metal2 s 108578 -400 108634 800 6 la_iena_mprj[4]
port 588 nsew signal input
rlabel metal2 s 121458 -400 121514 800 6 la_iena_mprj[50]
port 589 nsew signal input
rlabel metal2 s 121734 -400 121790 800 6 la_iena_mprj[51]
port 590 nsew signal input
rlabel metal2 s 122010 -400 122066 800 6 la_iena_mprj[52]
port 591 nsew signal input
rlabel metal2 s 122286 -400 122342 800 6 la_iena_mprj[53]
port 592 nsew signal input
rlabel metal2 s 122562 -400 122618 800 6 la_iena_mprj[54]
port 593 nsew signal input
rlabel metal2 s 122838 -400 122894 800 6 la_iena_mprj[55]
port 594 nsew signal input
rlabel metal2 s 123114 -400 123170 800 6 la_iena_mprj[56]
port 595 nsew signal input
rlabel metal2 s 123390 -400 123446 800 6 la_iena_mprj[57]
port 596 nsew signal input
rlabel metal2 s 123666 -400 123722 800 6 la_iena_mprj[58]
port 597 nsew signal input
rlabel metal2 s 123942 -400 123998 800 6 la_iena_mprj[59]
port 598 nsew signal input
rlabel metal2 s 108854 -400 108910 800 6 la_iena_mprj[5]
port 599 nsew signal input
rlabel metal2 s 124310 -400 124366 800 6 la_iena_mprj[60]
port 600 nsew signal input
rlabel metal2 s 124586 -400 124642 800 6 la_iena_mprj[61]
port 601 nsew signal input
rlabel metal2 s 124862 -400 124918 800 6 la_iena_mprj[62]
port 602 nsew signal input
rlabel metal2 s 125138 -400 125194 800 6 la_iena_mprj[63]
port 603 nsew signal input
rlabel metal2 s 125414 -400 125470 800 6 la_iena_mprj[64]
port 604 nsew signal input
rlabel metal2 s 125690 -400 125746 800 6 la_iena_mprj[65]
port 605 nsew signal input
rlabel metal2 s 125966 -400 126022 800 6 la_iena_mprj[66]
port 606 nsew signal input
rlabel metal2 s 126242 -400 126298 800 6 la_iena_mprj[67]
port 607 nsew signal input
rlabel metal2 s 126518 -400 126574 800 6 la_iena_mprj[68]
port 608 nsew signal input
rlabel metal2 s 126794 -400 126850 800 6 la_iena_mprj[69]
port 609 nsew signal input
rlabel metal2 s 109130 -400 109186 800 6 la_iena_mprj[6]
port 610 nsew signal input
rlabel metal2 s 127070 -400 127126 800 6 la_iena_mprj[70]
port 611 nsew signal input
rlabel metal2 s 127346 -400 127402 800 6 la_iena_mprj[71]
port 612 nsew signal input
rlabel metal2 s 127622 -400 127678 800 6 la_iena_mprj[72]
port 613 nsew signal input
rlabel metal2 s 127898 -400 127954 800 6 la_iena_mprj[73]
port 614 nsew signal input
rlabel metal2 s 128174 -400 128230 800 6 la_iena_mprj[74]
port 615 nsew signal input
rlabel metal2 s 128450 -400 128506 800 6 la_iena_mprj[75]
port 616 nsew signal input
rlabel metal2 s 128726 -400 128782 800 6 la_iena_mprj[76]
port 617 nsew signal input
rlabel metal2 s 129002 -400 129058 800 6 la_iena_mprj[77]
port 618 nsew signal input
rlabel metal2 s 129278 -400 129334 800 6 la_iena_mprj[78]
port 619 nsew signal input
rlabel metal2 s 129554 -400 129610 800 6 la_iena_mprj[79]
port 620 nsew signal input
rlabel metal2 s 109406 -400 109462 800 6 la_iena_mprj[7]
port 621 nsew signal input
rlabel metal2 s 129830 -400 129886 800 6 la_iena_mprj[80]
port 622 nsew signal input
rlabel metal2 s 130106 -400 130162 800 6 la_iena_mprj[81]
port 623 nsew signal input
rlabel metal2 s 130382 -400 130438 800 6 la_iena_mprj[82]
port 624 nsew signal input
rlabel metal2 s 130658 -400 130714 800 6 la_iena_mprj[83]
port 625 nsew signal input
rlabel metal2 s 130934 -400 130990 800 6 la_iena_mprj[84]
port 626 nsew signal input
rlabel metal2 s 131302 -400 131358 800 6 la_iena_mprj[85]
port 627 nsew signal input
rlabel metal2 s 131578 -400 131634 800 6 la_iena_mprj[86]
port 628 nsew signal input
rlabel metal2 s 131854 -400 131910 800 6 la_iena_mprj[87]
port 629 nsew signal input
rlabel metal2 s 132130 -400 132186 800 6 la_iena_mprj[88]
port 630 nsew signal input
rlabel metal2 s 132406 -400 132462 800 6 la_iena_mprj[89]
port 631 nsew signal input
rlabel metal2 s 109682 -400 109738 800 6 la_iena_mprj[8]
port 632 nsew signal input
rlabel metal2 s 132682 -400 132738 800 6 la_iena_mprj[90]
port 633 nsew signal input
rlabel metal2 s 132958 -400 133014 800 6 la_iena_mprj[91]
port 634 nsew signal input
rlabel metal2 s 133234 -400 133290 800 6 la_iena_mprj[92]
port 635 nsew signal input
rlabel metal2 s 133510 -400 133566 800 6 la_iena_mprj[93]
port 636 nsew signal input
rlabel metal2 s 133786 -400 133842 800 6 la_iena_mprj[94]
port 637 nsew signal input
rlabel metal2 s 134062 -400 134118 800 6 la_iena_mprj[95]
port 638 nsew signal input
rlabel metal2 s 134338 -400 134394 800 6 la_iena_mprj[96]
port 639 nsew signal input
rlabel metal2 s 134614 -400 134670 800 6 la_iena_mprj[97]
port 640 nsew signal input
rlabel metal2 s 134890 -400 134946 800 6 la_iena_mprj[98]
port 641 nsew signal input
rlabel metal2 s 135166 -400 135222 800 6 la_iena_mprj[99]
port 642 nsew signal input
rlabel metal2 s 109958 -400 110014 800 6 la_iena_mprj[9]
port 643 nsew signal input
rlabel metal2 s 143262 -400 143318 800 6 la_oenb_core[0]
port 644 nsew signal output
rlabel metal2 s 171230 -400 171286 800 6 la_oenb_core[100]
port 645 nsew signal output
rlabel metal2 s 171506 -400 171562 800 6 la_oenb_core[101]
port 646 nsew signal output
rlabel metal2 s 171782 -400 171838 800 6 la_oenb_core[102]
port 647 nsew signal output
rlabel metal2 s 172058 -400 172114 800 6 la_oenb_core[103]
port 648 nsew signal output
rlabel metal2 s 172334 -400 172390 800 6 la_oenb_core[104]
port 649 nsew signal output
rlabel metal2 s 172702 -400 172758 800 6 la_oenb_core[105]
port 650 nsew signal output
rlabel metal2 s 172978 -400 173034 800 6 la_oenb_core[106]
port 651 nsew signal output
rlabel metal2 s 173254 -400 173310 800 6 la_oenb_core[107]
port 652 nsew signal output
rlabel metal2 s 173530 -400 173586 800 6 la_oenb_core[108]
port 653 nsew signal output
rlabel metal2 s 173806 -400 173862 800 6 la_oenb_core[109]
port 654 nsew signal output
rlabel metal2 s 146114 -400 146170 800 6 la_oenb_core[10]
port 655 nsew signal output
rlabel metal2 s 174082 -400 174138 800 6 la_oenb_core[110]
port 656 nsew signal output
rlabel metal2 s 174358 -400 174414 800 6 la_oenb_core[111]
port 657 nsew signal output
rlabel metal2 s 174634 -400 174690 800 6 la_oenb_core[112]
port 658 nsew signal output
rlabel metal2 s 174910 -400 174966 800 6 la_oenb_core[113]
port 659 nsew signal output
rlabel metal2 s 175186 -400 175242 800 6 la_oenb_core[114]
port 660 nsew signal output
rlabel metal2 s 175462 -400 175518 800 6 la_oenb_core[115]
port 661 nsew signal output
rlabel metal2 s 175738 -400 175794 800 6 la_oenb_core[116]
port 662 nsew signal output
rlabel metal2 s 176014 -400 176070 800 6 la_oenb_core[117]
port 663 nsew signal output
rlabel metal2 s 176290 -400 176346 800 6 la_oenb_core[118]
port 664 nsew signal output
rlabel metal2 s 176566 -400 176622 800 6 la_oenb_core[119]
port 665 nsew signal output
rlabel metal2 s 146390 -400 146446 800 6 la_oenb_core[11]
port 666 nsew signal output
rlabel metal2 s 176842 -400 176898 800 6 la_oenb_core[120]
port 667 nsew signal output
rlabel metal2 s 177118 -400 177174 800 6 la_oenb_core[121]
port 668 nsew signal output
rlabel metal2 s 177394 -400 177450 800 6 la_oenb_core[122]
port 669 nsew signal output
rlabel metal2 s 177670 -400 177726 800 6 la_oenb_core[123]
port 670 nsew signal output
rlabel metal2 s 177946 -400 178002 800 6 la_oenb_core[124]
port 671 nsew signal output
rlabel metal2 s 178222 -400 178278 800 6 la_oenb_core[125]
port 672 nsew signal output
rlabel metal2 s 178498 -400 178554 800 6 la_oenb_core[126]
port 673 nsew signal output
rlabel metal2 s 178774 -400 178830 800 6 la_oenb_core[127]
port 674 nsew signal output
rlabel metal2 s 146666 -400 146722 800 6 la_oenb_core[12]
port 675 nsew signal output
rlabel metal2 s 146942 -400 146998 800 6 la_oenb_core[13]
port 676 nsew signal output
rlabel metal2 s 147218 -400 147274 800 6 la_oenb_core[14]
port 677 nsew signal output
rlabel metal2 s 147494 -400 147550 800 6 la_oenb_core[15]
port 678 nsew signal output
rlabel metal2 s 147770 -400 147826 800 6 la_oenb_core[16]
port 679 nsew signal output
rlabel metal2 s 148046 -400 148102 800 6 la_oenb_core[17]
port 680 nsew signal output
rlabel metal2 s 148322 -400 148378 800 6 la_oenb_core[18]
port 681 nsew signal output
rlabel metal2 s 148598 -400 148654 800 6 la_oenb_core[19]
port 682 nsew signal output
rlabel metal2 s 143538 -400 143594 800 6 la_oenb_core[1]
port 683 nsew signal output
rlabel metal2 s 148874 -400 148930 800 6 la_oenb_core[20]
port 684 nsew signal output
rlabel metal2 s 149150 -400 149206 800 6 la_oenb_core[21]
port 685 nsew signal output
rlabel metal2 s 149426 -400 149482 800 6 la_oenb_core[22]
port 686 nsew signal output
rlabel metal2 s 149702 -400 149758 800 6 la_oenb_core[23]
port 687 nsew signal output
rlabel metal2 s 149978 -400 150034 800 6 la_oenb_core[24]
port 688 nsew signal output
rlabel metal2 s 150254 -400 150310 800 6 la_oenb_core[25]
port 689 nsew signal output
rlabel metal2 s 150530 -400 150586 800 6 la_oenb_core[26]
port 690 nsew signal output
rlabel metal2 s 150806 -400 150862 800 6 la_oenb_core[27]
port 691 nsew signal output
rlabel metal2 s 151082 -400 151138 800 6 la_oenb_core[28]
port 692 nsew signal output
rlabel metal2 s 151358 -400 151414 800 6 la_oenb_core[29]
port 693 nsew signal output
rlabel metal2 s 143814 -400 143870 800 6 la_oenb_core[2]
port 694 nsew signal output
rlabel metal2 s 151634 -400 151690 800 6 la_oenb_core[30]
port 695 nsew signal output
rlabel metal2 s 152002 -400 152058 800 6 la_oenb_core[31]
port 696 nsew signal output
rlabel metal2 s 152278 -400 152334 800 6 la_oenb_core[32]
port 697 nsew signal output
rlabel metal2 s 152554 -400 152610 800 6 la_oenb_core[33]
port 698 nsew signal output
rlabel metal2 s 152830 -400 152886 800 6 la_oenb_core[34]
port 699 nsew signal output
rlabel metal2 s 153106 -400 153162 800 6 la_oenb_core[35]
port 700 nsew signal output
rlabel metal2 s 153382 -400 153438 800 6 la_oenb_core[36]
port 701 nsew signal output
rlabel metal2 s 153658 -400 153714 800 6 la_oenb_core[37]
port 702 nsew signal output
rlabel metal2 s 153934 -400 153990 800 6 la_oenb_core[38]
port 703 nsew signal output
rlabel metal2 s 154210 -400 154266 800 6 la_oenb_core[39]
port 704 nsew signal output
rlabel metal2 s 144090 -400 144146 800 6 la_oenb_core[3]
port 705 nsew signal output
rlabel metal2 s 154486 -400 154542 800 6 la_oenb_core[40]
port 706 nsew signal output
rlabel metal2 s 154762 -400 154818 800 6 la_oenb_core[41]
port 707 nsew signal output
rlabel metal2 s 155038 -400 155094 800 6 la_oenb_core[42]
port 708 nsew signal output
rlabel metal2 s 155314 -400 155370 800 6 la_oenb_core[43]
port 709 nsew signal output
rlabel metal2 s 155590 -400 155646 800 6 la_oenb_core[44]
port 710 nsew signal output
rlabel metal2 s 155866 -400 155922 800 6 la_oenb_core[45]
port 711 nsew signal output
rlabel metal2 s 156142 -400 156198 800 6 la_oenb_core[46]
port 712 nsew signal output
rlabel metal2 s 156418 -400 156474 800 6 la_oenb_core[47]
port 713 nsew signal output
rlabel metal2 s 156694 -400 156750 800 6 la_oenb_core[48]
port 714 nsew signal output
rlabel metal2 s 156970 -400 157026 800 6 la_oenb_core[49]
port 715 nsew signal output
rlabel metal2 s 144366 -400 144422 800 6 la_oenb_core[4]
port 716 nsew signal output
rlabel metal2 s 157246 -400 157302 800 6 la_oenb_core[50]
port 717 nsew signal output
rlabel metal2 s 157522 -400 157578 800 6 la_oenb_core[51]
port 718 nsew signal output
rlabel metal2 s 157798 -400 157854 800 6 la_oenb_core[52]
port 719 nsew signal output
rlabel metal2 s 158074 -400 158130 800 6 la_oenb_core[53]
port 720 nsew signal output
rlabel metal2 s 158350 -400 158406 800 6 la_oenb_core[54]
port 721 nsew signal output
rlabel metal2 s 158626 -400 158682 800 6 la_oenb_core[55]
port 722 nsew signal output
rlabel metal2 s 158994 -400 159050 800 6 la_oenb_core[56]
port 723 nsew signal output
rlabel metal2 s 159270 -400 159326 800 6 la_oenb_core[57]
port 724 nsew signal output
rlabel metal2 s 159546 -400 159602 800 6 la_oenb_core[58]
port 725 nsew signal output
rlabel metal2 s 159822 -400 159878 800 6 la_oenb_core[59]
port 726 nsew signal output
rlabel metal2 s 144642 -400 144698 800 6 la_oenb_core[5]
port 727 nsew signal output
rlabel metal2 s 160098 -400 160154 800 6 la_oenb_core[60]
port 728 nsew signal output
rlabel metal2 s 160374 -400 160430 800 6 la_oenb_core[61]
port 729 nsew signal output
rlabel metal2 s 160650 -400 160706 800 6 la_oenb_core[62]
port 730 nsew signal output
rlabel metal2 s 160926 -400 160982 800 6 la_oenb_core[63]
port 731 nsew signal output
rlabel metal2 s 161202 -400 161258 800 6 la_oenb_core[64]
port 732 nsew signal output
rlabel metal2 s 161478 -400 161534 800 6 la_oenb_core[65]
port 733 nsew signal output
rlabel metal2 s 161754 -400 161810 800 6 la_oenb_core[66]
port 734 nsew signal output
rlabel metal2 s 162030 -400 162086 800 6 la_oenb_core[67]
port 735 nsew signal output
rlabel metal2 s 162306 -400 162362 800 6 la_oenb_core[68]
port 736 nsew signal output
rlabel metal2 s 162582 -400 162638 800 6 la_oenb_core[69]
port 737 nsew signal output
rlabel metal2 s 145010 -400 145066 800 6 la_oenb_core[6]
port 738 nsew signal output
rlabel metal2 s 162858 -400 162914 800 6 la_oenb_core[70]
port 739 nsew signal output
rlabel metal2 s 163134 -400 163190 800 6 la_oenb_core[71]
port 740 nsew signal output
rlabel metal2 s 163410 -400 163466 800 6 la_oenb_core[72]
port 741 nsew signal output
rlabel metal2 s 163686 -400 163742 800 6 la_oenb_core[73]
port 742 nsew signal output
rlabel metal2 s 163962 -400 164018 800 6 la_oenb_core[74]
port 743 nsew signal output
rlabel metal2 s 164238 -400 164294 800 6 la_oenb_core[75]
port 744 nsew signal output
rlabel metal2 s 164514 -400 164570 800 6 la_oenb_core[76]
port 745 nsew signal output
rlabel metal2 s 164790 -400 164846 800 6 la_oenb_core[77]
port 746 nsew signal output
rlabel metal2 s 165066 -400 165122 800 6 la_oenb_core[78]
port 747 nsew signal output
rlabel metal2 s 165342 -400 165398 800 6 la_oenb_core[79]
port 748 nsew signal output
rlabel metal2 s 145286 -400 145342 800 6 la_oenb_core[7]
port 749 nsew signal output
rlabel metal2 s 165710 -400 165766 800 6 la_oenb_core[80]
port 750 nsew signal output
rlabel metal2 s 165986 -400 166042 800 6 la_oenb_core[81]
port 751 nsew signal output
rlabel metal2 s 166262 -400 166318 800 6 la_oenb_core[82]
port 752 nsew signal output
rlabel metal2 s 166538 -400 166594 800 6 la_oenb_core[83]
port 753 nsew signal output
rlabel metal2 s 166814 -400 166870 800 6 la_oenb_core[84]
port 754 nsew signal output
rlabel metal2 s 167090 -400 167146 800 6 la_oenb_core[85]
port 755 nsew signal output
rlabel metal2 s 167366 -400 167422 800 6 la_oenb_core[86]
port 756 nsew signal output
rlabel metal2 s 167642 -400 167698 800 6 la_oenb_core[87]
port 757 nsew signal output
rlabel metal2 s 167918 -400 167974 800 6 la_oenb_core[88]
port 758 nsew signal output
rlabel metal2 s 168194 -400 168250 800 6 la_oenb_core[89]
port 759 nsew signal output
rlabel metal2 s 145562 -400 145618 800 6 la_oenb_core[8]
port 760 nsew signal output
rlabel metal2 s 168470 -400 168526 800 6 la_oenb_core[90]
port 761 nsew signal output
rlabel metal2 s 168746 -400 168802 800 6 la_oenb_core[91]
port 762 nsew signal output
rlabel metal2 s 169022 -400 169078 800 6 la_oenb_core[92]
port 763 nsew signal output
rlabel metal2 s 169298 -400 169354 800 6 la_oenb_core[93]
port 764 nsew signal output
rlabel metal2 s 169574 -400 169630 800 6 la_oenb_core[94]
port 765 nsew signal output
rlabel metal2 s 169850 -400 169906 800 6 la_oenb_core[95]
port 766 nsew signal output
rlabel metal2 s 170126 -400 170182 800 6 la_oenb_core[96]
port 767 nsew signal output
rlabel metal2 s 170402 -400 170458 800 6 la_oenb_core[97]
port 768 nsew signal output
rlabel metal2 s 170678 -400 170734 800 6 la_oenb_core[98]
port 769 nsew signal output
rlabel metal2 s 170954 -400 171010 800 6 la_oenb_core[99]
port 770 nsew signal output
rlabel metal2 s 145838 -400 145894 800 6 la_oenb_core[9]
port 771 nsew signal output
rlabel metal2 s 71686 -400 71742 800 6 la_oenb_mprj[0]
port 772 nsew signal input
rlabel metal2 s 99654 -400 99710 800 6 la_oenb_mprj[100]
port 773 nsew signal input
rlabel metal2 s 99930 -400 99986 800 6 la_oenb_mprj[101]
port 774 nsew signal input
rlabel metal2 s 100206 -400 100262 800 6 la_oenb_mprj[102]
port 775 nsew signal input
rlabel metal2 s 100482 -400 100538 800 6 la_oenb_mprj[103]
port 776 nsew signal input
rlabel metal2 s 100758 -400 100814 800 6 la_oenb_mprj[104]
port 777 nsew signal input
rlabel metal2 s 101034 -400 101090 800 6 la_oenb_mprj[105]
port 778 nsew signal input
rlabel metal2 s 101310 -400 101366 800 6 la_oenb_mprj[106]
port 779 nsew signal input
rlabel metal2 s 101586 -400 101642 800 6 la_oenb_mprj[107]
port 780 nsew signal input
rlabel metal2 s 101862 -400 101918 800 6 la_oenb_mprj[108]
port 781 nsew signal input
rlabel metal2 s 102138 -400 102194 800 6 la_oenb_mprj[109]
port 782 nsew signal input
rlabel metal2 s 74446 -400 74502 800 6 la_oenb_mprj[10]
port 783 nsew signal input
rlabel metal2 s 102414 -400 102470 800 6 la_oenb_mprj[110]
port 784 nsew signal input
rlabel metal2 s 102690 -400 102746 800 6 la_oenb_mprj[111]
port 785 nsew signal input
rlabel metal2 s 102966 -400 103022 800 6 la_oenb_mprj[112]
port 786 nsew signal input
rlabel metal2 s 103242 -400 103298 800 6 la_oenb_mprj[113]
port 787 nsew signal input
rlabel metal2 s 103610 -400 103666 800 6 la_oenb_mprj[114]
port 788 nsew signal input
rlabel metal2 s 103886 -400 103942 800 6 la_oenb_mprj[115]
port 789 nsew signal input
rlabel metal2 s 104162 -400 104218 800 6 la_oenb_mprj[116]
port 790 nsew signal input
rlabel metal2 s 104438 -400 104494 800 6 la_oenb_mprj[117]
port 791 nsew signal input
rlabel metal2 s 104714 -400 104770 800 6 la_oenb_mprj[118]
port 792 nsew signal input
rlabel metal2 s 104990 -400 105046 800 6 la_oenb_mprj[119]
port 793 nsew signal input
rlabel metal2 s 74722 -400 74778 800 6 la_oenb_mprj[11]
port 794 nsew signal input
rlabel metal2 s 105266 -400 105322 800 6 la_oenb_mprj[120]
port 795 nsew signal input
rlabel metal2 s 105542 -400 105598 800 6 la_oenb_mprj[121]
port 796 nsew signal input
rlabel metal2 s 105818 -400 105874 800 6 la_oenb_mprj[122]
port 797 nsew signal input
rlabel metal2 s 106094 -400 106150 800 6 la_oenb_mprj[123]
port 798 nsew signal input
rlabel metal2 s 106370 -400 106426 800 6 la_oenb_mprj[124]
port 799 nsew signal input
rlabel metal2 s 106646 -400 106702 800 6 la_oenb_mprj[125]
port 800 nsew signal input
rlabel metal2 s 106922 -400 106978 800 6 la_oenb_mprj[126]
port 801 nsew signal input
rlabel metal2 s 107198 -400 107254 800 6 la_oenb_mprj[127]
port 802 nsew signal input
rlabel metal2 s 74998 -400 75054 800 6 la_oenb_mprj[12]
port 803 nsew signal input
rlabel metal2 s 75274 -400 75330 800 6 la_oenb_mprj[13]
port 804 nsew signal input
rlabel metal2 s 75550 -400 75606 800 6 la_oenb_mprj[14]
port 805 nsew signal input
rlabel metal2 s 75826 -400 75882 800 6 la_oenb_mprj[15]
port 806 nsew signal input
rlabel metal2 s 76194 -400 76250 800 6 la_oenb_mprj[16]
port 807 nsew signal input
rlabel metal2 s 76470 -400 76526 800 6 la_oenb_mprj[17]
port 808 nsew signal input
rlabel metal2 s 76746 -400 76802 800 6 la_oenb_mprj[18]
port 809 nsew signal input
rlabel metal2 s 77022 -400 77078 800 6 la_oenb_mprj[19]
port 810 nsew signal input
rlabel metal2 s 71962 -400 72018 800 6 la_oenb_mprj[1]
port 811 nsew signal input
rlabel metal2 s 77298 -400 77354 800 6 la_oenb_mprj[20]
port 812 nsew signal input
rlabel metal2 s 77574 -400 77630 800 6 la_oenb_mprj[21]
port 813 nsew signal input
rlabel metal2 s 77850 -400 77906 800 6 la_oenb_mprj[22]
port 814 nsew signal input
rlabel metal2 s 78126 -400 78182 800 6 la_oenb_mprj[23]
port 815 nsew signal input
rlabel metal2 s 78402 -400 78458 800 6 la_oenb_mprj[24]
port 816 nsew signal input
rlabel metal2 s 78678 -400 78734 800 6 la_oenb_mprj[25]
port 817 nsew signal input
rlabel metal2 s 78954 -400 79010 800 6 la_oenb_mprj[26]
port 818 nsew signal input
rlabel metal2 s 79230 -400 79286 800 6 la_oenb_mprj[27]
port 819 nsew signal input
rlabel metal2 s 79506 -400 79562 800 6 la_oenb_mprj[28]
port 820 nsew signal input
rlabel metal2 s 79782 -400 79838 800 6 la_oenb_mprj[29]
port 821 nsew signal input
rlabel metal2 s 72238 -400 72294 800 6 la_oenb_mprj[2]
port 822 nsew signal input
rlabel metal2 s 80058 -400 80114 800 6 la_oenb_mprj[30]
port 823 nsew signal input
rlabel metal2 s 80334 -400 80390 800 6 la_oenb_mprj[31]
port 824 nsew signal input
rlabel metal2 s 80610 -400 80666 800 6 la_oenb_mprj[32]
port 825 nsew signal input
rlabel metal2 s 80886 -400 80942 800 6 la_oenb_mprj[33]
port 826 nsew signal input
rlabel metal2 s 81162 -400 81218 800 6 la_oenb_mprj[34]
port 827 nsew signal input
rlabel metal2 s 81438 -400 81494 800 6 la_oenb_mprj[35]
port 828 nsew signal input
rlabel metal2 s 81714 -400 81770 800 6 la_oenb_mprj[36]
port 829 nsew signal input
rlabel metal2 s 81990 -400 82046 800 6 la_oenb_mprj[37]
port 830 nsew signal input
rlabel metal2 s 82266 -400 82322 800 6 la_oenb_mprj[38]
port 831 nsew signal input
rlabel metal2 s 82542 -400 82598 800 6 la_oenb_mprj[39]
port 832 nsew signal input
rlabel metal2 s 72514 -400 72570 800 6 la_oenb_mprj[3]
port 833 nsew signal input
rlabel metal2 s 82910 -400 82966 800 6 la_oenb_mprj[40]
port 834 nsew signal input
rlabel metal2 s 83186 -400 83242 800 6 la_oenb_mprj[41]
port 835 nsew signal input
rlabel metal2 s 83462 -400 83518 800 6 la_oenb_mprj[42]
port 836 nsew signal input
rlabel metal2 s 83738 -400 83794 800 6 la_oenb_mprj[43]
port 837 nsew signal input
rlabel metal2 s 84014 -400 84070 800 6 la_oenb_mprj[44]
port 838 nsew signal input
rlabel metal2 s 84290 -400 84346 800 6 la_oenb_mprj[45]
port 839 nsew signal input
rlabel metal2 s 84566 -400 84622 800 6 la_oenb_mprj[46]
port 840 nsew signal input
rlabel metal2 s 84842 -400 84898 800 6 la_oenb_mprj[47]
port 841 nsew signal input
rlabel metal2 s 85118 -400 85174 800 6 la_oenb_mprj[48]
port 842 nsew signal input
rlabel metal2 s 85394 -400 85450 800 6 la_oenb_mprj[49]
port 843 nsew signal input
rlabel metal2 s 72790 -400 72846 800 6 la_oenb_mprj[4]
port 844 nsew signal input
rlabel metal2 s 85670 -400 85726 800 6 la_oenb_mprj[50]
port 845 nsew signal input
rlabel metal2 s 85946 -400 86002 800 6 la_oenb_mprj[51]
port 846 nsew signal input
rlabel metal2 s 86222 -400 86278 800 6 la_oenb_mprj[52]
port 847 nsew signal input
rlabel metal2 s 86498 -400 86554 800 6 la_oenb_mprj[53]
port 848 nsew signal input
rlabel metal2 s 86774 -400 86830 800 6 la_oenb_mprj[54]
port 849 nsew signal input
rlabel metal2 s 87050 -400 87106 800 6 la_oenb_mprj[55]
port 850 nsew signal input
rlabel metal2 s 87326 -400 87382 800 6 la_oenb_mprj[56]
port 851 nsew signal input
rlabel metal2 s 87602 -400 87658 800 6 la_oenb_mprj[57]
port 852 nsew signal input
rlabel metal2 s 87878 -400 87934 800 6 la_oenb_mprj[58]
port 853 nsew signal input
rlabel metal2 s 88154 -400 88210 800 6 la_oenb_mprj[59]
port 854 nsew signal input
rlabel metal2 s 73066 -400 73122 800 6 la_oenb_mprj[5]
port 855 nsew signal input
rlabel metal2 s 88430 -400 88486 800 6 la_oenb_mprj[60]
port 856 nsew signal input
rlabel metal2 s 88706 -400 88762 800 6 la_oenb_mprj[61]
port 857 nsew signal input
rlabel metal2 s 88982 -400 89038 800 6 la_oenb_mprj[62]
port 858 nsew signal input
rlabel metal2 s 89258 -400 89314 800 6 la_oenb_mprj[63]
port 859 nsew signal input
rlabel metal2 s 89534 -400 89590 800 6 la_oenb_mprj[64]
port 860 nsew signal input
rlabel metal2 s 89902 -400 89958 800 6 la_oenb_mprj[65]
port 861 nsew signal input
rlabel metal2 s 90178 -400 90234 800 6 la_oenb_mprj[66]
port 862 nsew signal input
rlabel metal2 s 90454 -400 90510 800 6 la_oenb_mprj[67]
port 863 nsew signal input
rlabel metal2 s 90730 -400 90786 800 6 la_oenb_mprj[68]
port 864 nsew signal input
rlabel metal2 s 91006 -400 91062 800 6 la_oenb_mprj[69]
port 865 nsew signal input
rlabel metal2 s 73342 -400 73398 800 6 la_oenb_mprj[6]
port 866 nsew signal input
rlabel metal2 s 91282 -400 91338 800 6 la_oenb_mprj[70]
port 867 nsew signal input
rlabel metal2 s 91558 -400 91614 800 6 la_oenb_mprj[71]
port 868 nsew signal input
rlabel metal2 s 91834 -400 91890 800 6 la_oenb_mprj[72]
port 869 nsew signal input
rlabel metal2 s 92110 -400 92166 800 6 la_oenb_mprj[73]
port 870 nsew signal input
rlabel metal2 s 92386 -400 92442 800 6 la_oenb_mprj[74]
port 871 nsew signal input
rlabel metal2 s 92662 -400 92718 800 6 la_oenb_mprj[75]
port 872 nsew signal input
rlabel metal2 s 92938 -400 92994 800 6 la_oenb_mprj[76]
port 873 nsew signal input
rlabel metal2 s 93214 -400 93270 800 6 la_oenb_mprj[77]
port 874 nsew signal input
rlabel metal2 s 93490 -400 93546 800 6 la_oenb_mprj[78]
port 875 nsew signal input
rlabel metal2 s 93766 -400 93822 800 6 la_oenb_mprj[79]
port 876 nsew signal input
rlabel metal2 s 73618 -400 73674 800 6 la_oenb_mprj[7]
port 877 nsew signal input
rlabel metal2 s 94042 -400 94098 800 6 la_oenb_mprj[80]
port 878 nsew signal input
rlabel metal2 s 94318 -400 94374 800 6 la_oenb_mprj[81]
port 879 nsew signal input
rlabel metal2 s 94594 -400 94650 800 6 la_oenb_mprj[82]
port 880 nsew signal input
rlabel metal2 s 94870 -400 94926 800 6 la_oenb_mprj[83]
port 881 nsew signal input
rlabel metal2 s 95146 -400 95202 800 6 la_oenb_mprj[84]
port 882 nsew signal input
rlabel metal2 s 95422 -400 95478 800 6 la_oenb_mprj[85]
port 883 nsew signal input
rlabel metal2 s 95698 -400 95754 800 6 la_oenb_mprj[86]
port 884 nsew signal input
rlabel metal2 s 95974 -400 96030 800 6 la_oenb_mprj[87]
port 885 nsew signal input
rlabel metal2 s 96250 -400 96306 800 6 la_oenb_mprj[88]
port 886 nsew signal input
rlabel metal2 s 96526 -400 96582 800 6 la_oenb_mprj[89]
port 887 nsew signal input
rlabel metal2 s 73894 -400 73950 800 6 la_oenb_mprj[8]
port 888 nsew signal input
rlabel metal2 s 96894 -400 96950 800 6 la_oenb_mprj[90]
port 889 nsew signal input
rlabel metal2 s 97170 -400 97226 800 6 la_oenb_mprj[91]
port 890 nsew signal input
rlabel metal2 s 97446 -400 97502 800 6 la_oenb_mprj[92]
port 891 nsew signal input
rlabel metal2 s 97722 -400 97778 800 6 la_oenb_mprj[93]
port 892 nsew signal input
rlabel metal2 s 97998 -400 98054 800 6 la_oenb_mprj[94]
port 893 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 la_oenb_mprj[95]
port 894 nsew signal input
rlabel metal2 s 98550 -400 98606 800 6 la_oenb_mprj[96]
port 895 nsew signal input
rlabel metal2 s 98826 -400 98882 800 6 la_oenb_mprj[97]
port 896 nsew signal input
rlabel metal2 s 99102 -400 99158 800 6 la_oenb_mprj[98]
port 897 nsew signal input
rlabel metal2 s 99378 -400 99434 800 6 la_oenb_mprj[99]
port 898 nsew signal input
rlabel metal2 s 74170 -400 74226 800 6 la_oenb_mprj[9]
port 899 nsew signal input
rlabel metal2 s 179970 -400 180026 800 6 mprj_adr_o_core[0]
port 900 nsew signal input
rlabel metal2 s 186686 -400 186742 800 6 mprj_adr_o_core[10]
port 901 nsew signal input
rlabel metal2 s 187238 -400 187294 800 6 mprj_adr_o_core[11]
port 902 nsew signal input
rlabel metal2 s 187790 -400 187846 800 6 mprj_adr_o_core[12]
port 903 nsew signal input
rlabel metal2 s 188342 -400 188398 800 6 mprj_adr_o_core[13]
port 904 nsew signal input
rlabel metal2 s 188894 -400 188950 800 6 mprj_adr_o_core[14]
port 905 nsew signal input
rlabel metal2 s 189446 -400 189502 800 6 mprj_adr_o_core[15]
port 906 nsew signal input
rlabel metal2 s 189998 -400 190054 800 6 mprj_adr_o_core[16]
port 907 nsew signal input
rlabel metal2 s 190550 -400 190606 800 6 mprj_adr_o_core[17]
port 908 nsew signal input
rlabel metal2 s 191102 -400 191158 800 6 mprj_adr_o_core[18]
port 909 nsew signal input
rlabel metal2 s 191654 -400 191710 800 6 mprj_adr_o_core[19]
port 910 nsew signal input
rlabel metal2 s 180798 -400 180854 800 6 mprj_adr_o_core[1]
port 911 nsew signal input
rlabel metal2 s 192206 -400 192262 800 6 mprj_adr_o_core[20]
port 912 nsew signal input
rlabel metal2 s 192758 -400 192814 800 6 mprj_adr_o_core[21]
port 913 nsew signal input
rlabel metal2 s 193402 -400 193458 800 6 mprj_adr_o_core[22]
port 914 nsew signal input
rlabel metal2 s 193954 -400 194010 800 6 mprj_adr_o_core[23]
port 915 nsew signal input
rlabel metal2 s 194506 -400 194562 800 6 mprj_adr_o_core[24]
port 916 nsew signal input
rlabel metal2 s 195058 -400 195114 800 6 mprj_adr_o_core[25]
port 917 nsew signal input
rlabel metal2 s 195610 -400 195666 800 6 mprj_adr_o_core[26]
port 918 nsew signal input
rlabel metal2 s 196162 -400 196218 800 6 mprj_adr_o_core[27]
port 919 nsew signal input
rlabel metal2 s 196714 -400 196770 800 6 mprj_adr_o_core[28]
port 920 nsew signal input
rlabel metal2 s 197266 -400 197322 800 6 mprj_adr_o_core[29]
port 921 nsew signal input
rlabel metal2 s 181626 -400 181682 800 6 mprj_adr_o_core[2]
port 922 nsew signal input
rlabel metal2 s 197818 -400 197874 800 6 mprj_adr_o_core[30]
port 923 nsew signal input
rlabel metal2 s 198370 -400 198426 800 6 mprj_adr_o_core[31]
port 924 nsew signal input
rlabel metal2 s 182454 -400 182510 800 6 mprj_adr_o_core[3]
port 925 nsew signal input
rlabel metal2 s 183282 -400 183338 800 6 mprj_adr_o_core[4]
port 926 nsew signal input
rlabel metal2 s 183834 -400 183890 800 6 mprj_adr_o_core[5]
port 927 nsew signal input
rlabel metal2 s 184386 -400 184442 800 6 mprj_adr_o_core[6]
port 928 nsew signal input
rlabel metal2 s 184938 -400 184994 800 6 mprj_adr_o_core[7]
port 929 nsew signal input
rlabel metal2 s 185490 -400 185546 800 6 mprj_adr_o_core[8]
port 930 nsew signal input
rlabel metal2 s 186042 -400 186098 800 6 mprj_adr_o_core[9]
port 931 nsew signal input
rlabel metal2 s 160282 28400 160338 29600 6 mprj_adr_o_user[0]
port 932 nsew signal output
rlabel metal2 s 174358 28400 174414 29600 6 mprj_adr_o_user[10]
port 933 nsew signal output
rlabel metal2 s 175554 28400 175610 29600 6 mprj_adr_o_user[11]
port 934 nsew signal output
rlabel metal2 s 176750 28400 176806 29600 6 mprj_adr_o_user[12]
port 935 nsew signal output
rlabel metal2 s 177946 28400 178002 29600 6 mprj_adr_o_user[13]
port 936 nsew signal output
rlabel metal2 s 179050 28400 179106 29600 6 mprj_adr_o_user[14]
port 937 nsew signal output
rlabel metal2 s 180246 28400 180302 29600 6 mprj_adr_o_user[15]
port 938 nsew signal output
rlabel metal2 s 181442 28400 181498 29600 6 mprj_adr_o_user[16]
port 939 nsew signal output
rlabel metal2 s 182638 28400 182694 29600 6 mprj_adr_o_user[17]
port 940 nsew signal output
rlabel metal2 s 183742 28400 183798 29600 6 mprj_adr_o_user[18]
port 941 nsew signal output
rlabel metal2 s 184938 28400 184994 29600 6 mprj_adr_o_user[19]
port 942 nsew signal output
rlabel metal2 s 162030 28400 162086 29600 6 mprj_adr_o_user[1]
port 943 nsew signal output
rlabel metal2 s 186134 28400 186190 29600 6 mprj_adr_o_user[20]
port 944 nsew signal output
rlabel metal2 s 187330 28400 187386 29600 6 mprj_adr_o_user[21]
port 945 nsew signal output
rlabel metal2 s 188526 28400 188582 29600 6 mprj_adr_o_user[22]
port 946 nsew signal output
rlabel metal2 s 189630 28400 189686 29600 6 mprj_adr_o_user[23]
port 947 nsew signal output
rlabel metal2 s 190826 28400 190882 29600 6 mprj_adr_o_user[24]
port 948 nsew signal output
rlabel metal2 s 192022 28400 192078 29600 6 mprj_adr_o_user[25]
port 949 nsew signal output
rlabel metal2 s 193218 28400 193274 29600 6 mprj_adr_o_user[26]
port 950 nsew signal output
rlabel metal2 s 194414 28400 194470 29600 6 mprj_adr_o_user[27]
port 951 nsew signal output
rlabel metal2 s 195518 28400 195574 29600 6 mprj_adr_o_user[28]
port 952 nsew signal output
rlabel metal2 s 196714 28400 196770 29600 6 mprj_adr_o_user[29]
port 953 nsew signal output
rlabel metal2 s 163778 28400 163834 29600 6 mprj_adr_o_user[2]
port 954 nsew signal output
rlabel metal2 s 197910 28400 197966 29600 6 mprj_adr_o_user[30]
port 955 nsew signal output
rlabel metal2 s 199106 28400 199162 29600 6 mprj_adr_o_user[31]
port 956 nsew signal output
rlabel metal2 s 165526 28400 165582 29600 6 mprj_adr_o_user[3]
port 957 nsew signal output
rlabel metal2 s 167274 28400 167330 29600 6 mprj_adr_o_user[4]
port 958 nsew signal output
rlabel metal2 s 168470 28400 168526 29600 6 mprj_adr_o_user[5]
port 959 nsew signal output
rlabel metal2 s 169666 28400 169722 29600 6 mprj_adr_o_user[6]
port 960 nsew signal output
rlabel metal2 s 170862 28400 170918 29600 6 mprj_adr_o_user[7]
port 961 nsew signal output
rlabel metal2 s 172058 28400 172114 29600 6 mprj_adr_o_user[8]
port 962 nsew signal output
rlabel metal2 s 173162 28400 173218 29600 6 mprj_adr_o_user[9]
port 963 nsew signal output
rlabel metal2 s 179050 -400 179106 800 6 mprj_cyc_o_core
port 964 nsew signal input
rlabel metal2 s 158534 28400 158590 29600 6 mprj_cyc_o_user
port 965 nsew signal output
rlabel metal2 s 180246 -400 180302 800 6 mprj_dat_o_core[0]
port 966 nsew signal input
rlabel metal2 s 186962 -400 187018 800 6 mprj_dat_o_core[10]
port 967 nsew signal input
rlabel metal2 s 187514 -400 187570 800 6 mprj_dat_o_core[11]
port 968 nsew signal input
rlabel metal2 s 188066 -400 188122 800 6 mprj_dat_o_core[12]
port 969 nsew signal input
rlabel metal2 s 188618 -400 188674 800 6 mprj_dat_o_core[13]
port 970 nsew signal input
rlabel metal2 s 189170 -400 189226 800 6 mprj_dat_o_core[14]
port 971 nsew signal input
rlabel metal2 s 189722 -400 189778 800 6 mprj_dat_o_core[15]
port 972 nsew signal input
rlabel metal2 s 190274 -400 190330 800 6 mprj_dat_o_core[16]
port 973 nsew signal input
rlabel metal2 s 190826 -400 190882 800 6 mprj_dat_o_core[17]
port 974 nsew signal input
rlabel metal2 s 191378 -400 191434 800 6 mprj_dat_o_core[18]
port 975 nsew signal input
rlabel metal2 s 191930 -400 191986 800 6 mprj_dat_o_core[19]
port 976 nsew signal input
rlabel metal2 s 181074 -400 181130 800 6 mprj_dat_o_core[1]
port 977 nsew signal input
rlabel metal2 s 192482 -400 192538 800 6 mprj_dat_o_core[20]
port 978 nsew signal input
rlabel metal2 s 193034 -400 193090 800 6 mprj_dat_o_core[21]
port 979 nsew signal input
rlabel metal2 s 193678 -400 193734 800 6 mprj_dat_o_core[22]
port 980 nsew signal input
rlabel metal2 s 194230 -400 194286 800 6 mprj_dat_o_core[23]
port 981 nsew signal input
rlabel metal2 s 194782 -400 194838 800 6 mprj_dat_o_core[24]
port 982 nsew signal input
rlabel metal2 s 195334 -400 195390 800 6 mprj_dat_o_core[25]
port 983 nsew signal input
rlabel metal2 s 195886 -400 195942 800 6 mprj_dat_o_core[26]
port 984 nsew signal input
rlabel metal2 s 196438 -400 196494 800 6 mprj_dat_o_core[27]
port 985 nsew signal input
rlabel metal2 s 196990 -400 197046 800 6 mprj_dat_o_core[28]
port 986 nsew signal input
rlabel metal2 s 197542 -400 197598 800 6 mprj_dat_o_core[29]
port 987 nsew signal input
rlabel metal2 s 181902 -400 181958 800 6 mprj_dat_o_core[2]
port 988 nsew signal input
rlabel metal2 s 198094 -400 198150 800 6 mprj_dat_o_core[30]
port 989 nsew signal input
rlabel metal2 s 198646 -400 198702 800 6 mprj_dat_o_core[31]
port 990 nsew signal input
rlabel metal2 s 182730 -400 182786 800 6 mprj_dat_o_core[3]
port 991 nsew signal input
rlabel metal2 s 183558 -400 183614 800 6 mprj_dat_o_core[4]
port 992 nsew signal input
rlabel metal2 s 184110 -400 184166 800 6 mprj_dat_o_core[5]
port 993 nsew signal input
rlabel metal2 s 184662 -400 184718 800 6 mprj_dat_o_core[6]
port 994 nsew signal input
rlabel metal2 s 185214 -400 185270 800 6 mprj_dat_o_core[7]
port 995 nsew signal input
rlabel metal2 s 185766 -400 185822 800 6 mprj_dat_o_core[8]
port 996 nsew signal input
rlabel metal2 s 186410 -400 186466 800 6 mprj_dat_o_core[9]
port 997 nsew signal input
rlabel metal2 s 160834 28400 160890 29600 6 mprj_dat_o_user[0]
port 998 nsew signal output
rlabel metal2 s 175002 28400 175058 29600 6 mprj_dat_o_user[10]
port 999 nsew signal output
rlabel metal2 s 176106 28400 176162 29600 6 mprj_dat_o_user[11]
port 1000 nsew signal output
rlabel metal2 s 177302 28400 177358 29600 6 mprj_dat_o_user[12]
port 1001 nsew signal output
rlabel metal2 s 178498 28400 178554 29600 6 mprj_dat_o_user[13]
port 1002 nsew signal output
rlabel metal2 s 179694 28400 179750 29600 6 mprj_dat_o_user[14]
port 1003 nsew signal output
rlabel metal2 s 180798 28400 180854 29600 6 mprj_dat_o_user[15]
port 1004 nsew signal output
rlabel metal2 s 181994 28400 182050 29600 6 mprj_dat_o_user[16]
port 1005 nsew signal output
rlabel metal2 s 183190 28400 183246 29600 6 mprj_dat_o_user[17]
port 1006 nsew signal output
rlabel metal2 s 184386 28400 184442 29600 6 mprj_dat_o_user[18]
port 1007 nsew signal output
rlabel metal2 s 185582 28400 185638 29600 6 mprj_dat_o_user[19]
port 1008 nsew signal output
rlabel metal2 s 162582 28400 162638 29600 6 mprj_dat_o_user[1]
port 1009 nsew signal output
rlabel metal2 s 186686 28400 186742 29600 6 mprj_dat_o_user[20]
port 1010 nsew signal output
rlabel metal2 s 187882 28400 187938 29600 6 mprj_dat_o_user[21]
port 1011 nsew signal output
rlabel metal2 s 189078 28400 189134 29600 6 mprj_dat_o_user[22]
port 1012 nsew signal output
rlabel metal2 s 190274 28400 190330 29600 6 mprj_dat_o_user[23]
port 1013 nsew signal output
rlabel metal2 s 191470 28400 191526 29600 6 mprj_dat_o_user[24]
port 1014 nsew signal output
rlabel metal2 s 192574 28400 192630 29600 6 mprj_dat_o_user[25]
port 1015 nsew signal output
rlabel metal2 s 193770 28400 193826 29600 6 mprj_dat_o_user[26]
port 1016 nsew signal output
rlabel metal2 s 194966 28400 195022 29600 6 mprj_dat_o_user[27]
port 1017 nsew signal output
rlabel metal2 s 196162 28400 196218 29600 6 mprj_dat_o_user[28]
port 1018 nsew signal output
rlabel metal2 s 197358 28400 197414 29600 6 mprj_dat_o_user[29]
port 1019 nsew signal output
rlabel metal2 s 164330 28400 164386 29600 6 mprj_dat_o_user[2]
port 1020 nsew signal output
rlabel metal2 s 198462 28400 198518 29600 6 mprj_dat_o_user[30]
port 1021 nsew signal output
rlabel metal2 s 199658 28400 199714 29600 6 mprj_dat_o_user[31]
port 1022 nsew signal output
rlabel metal2 s 166170 28400 166226 29600 6 mprj_dat_o_user[3]
port 1023 nsew signal output
rlabel metal2 s 167918 28400 167974 29600 6 mprj_dat_o_user[4]
port 1024 nsew signal output
rlabel metal2 s 169114 28400 169170 29600 6 mprj_dat_o_user[5]
port 1025 nsew signal output
rlabel metal2 s 170218 28400 170274 29600 6 mprj_dat_o_user[6]
port 1026 nsew signal output
rlabel metal2 s 171414 28400 171470 29600 6 mprj_dat_o_user[7]
port 1027 nsew signal output
rlabel metal2 s 172610 28400 172666 29600 6 mprj_dat_o_user[8]
port 1028 nsew signal output
rlabel metal2 s 173806 28400 173862 29600 6 mprj_dat_o_user[9]
port 1029 nsew signal output
rlabel metal2 s 180522 -400 180578 800 6 mprj_sel_o_core[0]
port 1030 nsew signal input
rlabel metal2 s 181350 -400 181406 800 6 mprj_sel_o_core[1]
port 1031 nsew signal input
rlabel metal2 s 182178 -400 182234 800 6 mprj_sel_o_core[2]
port 1032 nsew signal input
rlabel metal2 s 183006 -400 183062 800 6 mprj_sel_o_core[3]
port 1033 nsew signal input
rlabel metal2 s 161386 28400 161442 29600 6 mprj_sel_o_user[0]
port 1034 nsew signal output
rlabel metal2 s 163226 28400 163282 29600 6 mprj_sel_o_user[1]
port 1035 nsew signal output
rlabel metal2 s 164974 28400 165030 29600 6 mprj_sel_o_user[2]
port 1036 nsew signal output
rlabel metal2 s 166722 28400 166778 29600 6 mprj_sel_o_user[3]
port 1037 nsew signal output
rlabel metal2 s 179326 -400 179382 800 6 mprj_stb_o_core
port 1038 nsew signal input
rlabel metal2 s 159086 28400 159142 29600 6 mprj_stb_o_user
port 1039 nsew signal output
rlabel metal2 s 179694 -400 179750 800 6 mprj_we_o_core
port 1040 nsew signal input
rlabel metal2 s 159638 28400 159694 29600 6 mprj_we_o_user
port 1041 nsew signal output
rlabel metal2 s 198922 -400 198978 800 6 user1_vcc_powergood
port 1042 nsew signal output
rlabel metal2 s 199198 -400 199254 800 6 user1_vdd_powergood
port 1043 nsew signal output
rlabel metal2 s 199474 -400 199530 800 6 user2_vcc_powergood
port 1044 nsew signal output
rlabel metal2 s 199750 -400 199806 800 6 user2_vdd_powergood
port 1045 nsew signal output
rlabel metal2 s 294 28400 350 29600 6 user_clock
port 1046 nsew signal output
rlabel metal2 s 846 28400 902 29600 6 user_clock2
port 1047 nsew signal output
rlabel metal2 s 2594 28400 2650 29600 6 user_irq[0]
port 1048 nsew signal output
rlabel metal2 s 4342 28400 4398 29600 6 user_irq[1]
port 1049 nsew signal output
rlabel metal2 s 6090 28400 6146 29600 6 user_irq[2]
port 1050 nsew signal output
rlabel metal2 s 3146 28400 3202 29600 6 user_irq_core[0]
port 1051 nsew signal input
rlabel metal2 s 4986 28400 5042 29600 6 user_irq_core[1]
port 1052 nsew signal input
rlabel metal2 s 6734 28400 6790 29600 6 user_irq_core[2]
port 1053 nsew signal input
rlabel metal2 s 3790 28400 3846 29600 6 user_irq_ena[0]
port 1054 nsew signal input
rlabel metal2 s 5538 28400 5594 29600 6 user_irq_ena[1]
port 1055 nsew signal input
rlabel metal2 s 7286 28400 7342 29600 6 user_irq_ena[2]
port 1056 nsew signal input
rlabel metal2 s 1398 28400 1454 29600 6 user_reset
port 1057 nsew signal output
rlabel metal2 s 2042 28400 2098 29600 6 user_resetn
port 1058 nsew signal output
rlabel metal3 s -386 29054 200302 29234 6 vccd
port 1059 nsew power bidirectional
rlabel metal3 s -386 -402 200302 -222 8 vccd
port 1060 nsew power bidirectional
rlabel metal4 s 178014 -666 178194 29498 6 vccd
port 1061 nsew power bidirectional
rlabel metal4 s 149014 -666 149194 29498 6 vccd
port 1062 nsew power bidirectional
rlabel metal4 s 120014 -666 120194 29498 6 vccd
port 1063 nsew power bidirectional
rlabel metal4 s 91014 -666 91194 29498 6 vccd
port 1064 nsew power bidirectional
rlabel metal4 s 62014 -666 62194 29498 6 vccd
port 1065 nsew power bidirectional
rlabel metal4 s 33014 -666 33194 29498 6 vccd
port 1066 nsew power bidirectional
rlabel metal4 s 4014 -666 4194 29498 6 vccd
port 1067 nsew power bidirectional
rlabel metal4 s 200122 -402 200302 29234 6 vccd
port 1068 nsew power bidirectional
rlabel metal4 s -386 -402 -206 29234 4 vccd
port 1069 nsew power bidirectional
rlabel metal3 s -650 29318 200566 29498 6 vssd
port 1070 nsew ground bidirectional
rlabel metal3 s -650 -666 200566 -486 8 vssd
port 1071 nsew ground bidirectional
rlabel metal4 s 200386 -666 200566 29498 6 vssd
port 1072 nsew ground bidirectional
rlabel metal4 s 192514 -666 192694 29498 6 vssd
port 1073 nsew ground bidirectional
rlabel metal4 s 163514 -666 163694 29498 6 vssd
port 1074 nsew ground bidirectional
rlabel metal4 s 134514 -666 134694 29498 6 vssd
port 1075 nsew ground bidirectional
rlabel metal4 s 105514 -666 105694 29498 6 vssd
port 1076 nsew ground bidirectional
rlabel metal4 s 76514 -666 76694 29498 6 vssd
port 1077 nsew ground bidirectional
rlabel metal4 s 47514 -666 47694 29498 6 vssd
port 1078 nsew ground bidirectional
rlabel metal4 s 18514 -666 18694 29498 6 vssd
port 1079 nsew ground bidirectional
rlabel metal4 s -650 -666 -470 29498 4 vssd
port 1080 nsew ground bidirectional
rlabel metal3 s -914 29582 200830 29762 6 vccd1
port 1081 nsew power bidirectional
rlabel metal3 s -914 -930 200830 -750 8 vccd1
port 1082 nsew power bidirectional
rlabel metal4 s 178834 -1194 179014 30026 6 vccd1
port 1083 nsew power bidirectional
rlabel metal4 s 149834 -1194 150014 30026 6 vccd1
port 1084 nsew power bidirectional
rlabel metal4 s 120834 -1194 121014 30026 6 vccd1
port 1085 nsew power bidirectional
rlabel metal4 s 91834 -1194 92014 30026 6 vccd1
port 1086 nsew power bidirectional
rlabel metal4 s 62834 -1194 63014 30026 6 vccd1
port 1087 nsew power bidirectional
rlabel metal4 s 33834 -1194 34014 30026 6 vccd1
port 1088 nsew power bidirectional
rlabel metal4 s 4834 -1194 5014 30026 6 vccd1
port 1089 nsew power bidirectional
rlabel metal4 s 200650 -930 200830 29762 6 vccd1
port 1090 nsew power bidirectional
rlabel metal4 s -914 -930 -734 29762 4 vccd1
port 1091 nsew power bidirectional
rlabel metal3 s -1178 29846 201094 30026 6 vssd1
port 1092 nsew ground bidirectional
rlabel metal3 s -1178 -1194 201094 -1014 8 vssd1
port 1093 nsew ground bidirectional
rlabel metal4 s 200914 -1194 201094 30026 6 vssd1
port 1094 nsew ground bidirectional
rlabel metal4 s 193334 -1194 193514 30026 6 vssd1
port 1095 nsew ground bidirectional
rlabel metal4 s 164334 -1194 164514 30026 6 vssd1
port 1096 nsew ground bidirectional
rlabel metal4 s 135334 -1194 135514 30026 6 vssd1
port 1097 nsew ground bidirectional
rlabel metal4 s 106334 -1194 106514 30026 6 vssd1
port 1098 nsew ground bidirectional
rlabel metal4 s 77334 -1194 77514 30026 6 vssd1
port 1099 nsew ground bidirectional
rlabel metal4 s 48334 -1194 48514 30026 6 vssd1
port 1100 nsew ground bidirectional
rlabel metal4 s 19334 -1194 19514 30026 6 vssd1
port 1101 nsew ground bidirectional
rlabel metal4 s -1178 -1194 -998 30026 4 vssd1
port 1102 nsew ground bidirectional
rlabel metal3 s -1442 30110 201358 30290 6 vccd2
port 1103 nsew power bidirectional
rlabel metal3 s -1442 -1458 201358 -1278 8 vccd2
port 1104 nsew power bidirectional
rlabel metal4 s 179654 -1722 179834 30554 6 vccd2
port 1105 nsew power bidirectional
rlabel metal4 s 150654 -1722 150834 30554 6 vccd2
port 1106 nsew power bidirectional
rlabel metal4 s 121654 -1722 121834 30554 6 vccd2
port 1107 nsew power bidirectional
rlabel metal4 s 92654 -1722 92834 30554 6 vccd2
port 1108 nsew power bidirectional
rlabel metal4 s 63654 -1722 63834 30554 6 vccd2
port 1109 nsew power bidirectional
rlabel metal4 s 34654 -1722 34834 30554 6 vccd2
port 1110 nsew power bidirectional
rlabel metal4 s 5654 -1722 5834 30554 6 vccd2
port 1111 nsew power bidirectional
rlabel metal4 s 201178 -1458 201358 30290 6 vccd2
port 1112 nsew power bidirectional
rlabel metal4 s -1442 -1458 -1262 30290 4 vccd2
port 1113 nsew power bidirectional
rlabel metal3 s -1706 30374 201622 30554 6 vssd2
port 1114 nsew ground bidirectional
rlabel metal3 s -1706 -1722 201622 -1542 8 vssd2
port 1115 nsew ground bidirectional
rlabel metal4 s 201442 -1722 201622 30554 6 vssd2
port 1116 nsew ground bidirectional
rlabel metal4 s 194154 -1722 194334 30554 6 vssd2
port 1117 nsew ground bidirectional
rlabel metal4 s 165154 -1722 165334 30554 6 vssd2
port 1118 nsew ground bidirectional
rlabel metal4 s 136154 -1722 136334 30554 6 vssd2
port 1119 nsew ground bidirectional
rlabel metal4 s 107154 -1722 107334 30554 6 vssd2
port 1120 nsew ground bidirectional
rlabel metal4 s 78154 -1722 78334 30554 6 vssd2
port 1121 nsew ground bidirectional
rlabel metal4 s 49154 -1722 49334 30554 6 vssd2
port 1122 nsew ground bidirectional
rlabel metal4 s 20154 -1722 20334 30554 6 vssd2
port 1123 nsew ground bidirectional
rlabel metal4 s -1706 -1722 -1526 30554 4 vssd2
port 1124 nsew ground bidirectional
rlabel metal3 s -1970 30638 201886 30818 6 vdda1
port 1125 nsew power bidirectional
rlabel metal3 s -1970 -1986 201886 -1806 8 vdda1
port 1126 nsew power bidirectional
rlabel metal4 s 180474 -2250 180654 31082 6 vdda1
port 1127 nsew power bidirectional
rlabel metal4 s 151474 -2250 151654 31082 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 122474 -2250 122654 31082 6 vdda1
port 1129 nsew power bidirectional
rlabel metal4 s 93474 -2250 93654 31082 6 vdda1
port 1130 nsew power bidirectional
rlabel metal4 s 64474 -2250 64654 31082 6 vdda1
port 1131 nsew power bidirectional
rlabel metal4 s 35474 -2250 35654 31082 6 vdda1
port 1132 nsew power bidirectional
rlabel metal4 s 6474 -2250 6654 31082 6 vdda1
port 1133 nsew power bidirectional
rlabel metal4 s 201706 -1986 201886 30818 6 vdda1
port 1134 nsew power bidirectional
rlabel metal4 s -1970 -1986 -1790 30818 4 vdda1
port 1135 nsew power bidirectional
rlabel metal3 s -2234 30902 202150 31082 6 vssa1
port 1136 nsew ground bidirectional
rlabel metal3 s -2234 -2250 202150 -2070 8 vssa1
port 1137 nsew ground bidirectional
rlabel metal4 s 201970 -2250 202150 31082 6 vssa1
port 1138 nsew ground bidirectional
rlabel metal4 s 194974 -2250 195154 31082 6 vssa1
port 1139 nsew ground bidirectional
rlabel metal4 s 165974 -2250 166154 31082 6 vssa1
port 1140 nsew ground bidirectional
rlabel metal4 s 136974 -2250 137154 31082 6 vssa1
port 1141 nsew ground bidirectional
rlabel metal4 s 107974 -2250 108154 31082 6 vssa1
port 1142 nsew ground bidirectional
rlabel metal4 s 78974 -2250 79154 31082 6 vssa1
port 1143 nsew ground bidirectional
rlabel metal4 s 49974 -2250 50154 31082 6 vssa1
port 1144 nsew ground bidirectional
rlabel metal4 s 20974 -2250 21154 31082 6 vssa1
port 1145 nsew ground bidirectional
rlabel metal4 s -2234 -2250 -2054 31082 4 vssa1
port 1146 nsew ground bidirectional
rlabel metal3 s -2498 31166 202414 31346 6 vdda2
port 1147 nsew power bidirectional
rlabel metal3 s -2498 -2514 202414 -2334 8 vdda2
port 1148 nsew power bidirectional
rlabel metal4 s 181294 -2778 181474 31610 6 vdda2
port 1149 nsew power bidirectional
rlabel metal4 s 152294 -2778 152474 31610 6 vdda2
port 1150 nsew power bidirectional
rlabel metal4 s 123294 -2778 123474 31610 6 vdda2
port 1151 nsew power bidirectional
rlabel metal4 s 94294 -2778 94474 31610 6 vdda2
port 1152 nsew power bidirectional
rlabel metal4 s 65294 -2778 65474 31610 6 vdda2
port 1153 nsew power bidirectional
rlabel metal4 s 36294 -2778 36474 31610 6 vdda2
port 1154 nsew power bidirectional
rlabel metal4 s 7294 -2778 7474 31610 6 vdda2
port 1155 nsew power bidirectional
rlabel metal4 s 202234 -2514 202414 31346 6 vdda2
port 1156 nsew power bidirectional
rlabel metal4 s -2498 -2514 -2318 31346 4 vdda2
port 1157 nsew power bidirectional
rlabel metal3 s -2762 31430 202678 31610 6 vssa2
port 1158 nsew ground bidirectional
rlabel metal3 s -2762 -2778 202678 -2598 8 vssa2
port 1159 nsew ground bidirectional
rlabel metal4 s 202498 -2778 202678 31610 6 vssa2
port 1160 nsew ground bidirectional
rlabel metal4 s 195794 -2778 195974 31610 6 vssa2
port 1161 nsew ground bidirectional
rlabel metal4 s 166794 -2778 166974 31610 6 vssa2
port 1162 nsew ground bidirectional
rlabel metal4 s 137794 -2778 137974 31610 6 vssa2
port 1163 nsew ground bidirectional
rlabel metal4 s 108794 -2778 108974 31610 6 vssa2
port 1164 nsew ground bidirectional
rlabel metal4 s 79794 -2778 79974 31610 6 vssa2
port 1165 nsew ground bidirectional
rlabel metal4 s 50794 -2778 50974 31610 6 vssa2
port 1166 nsew ground bidirectional
rlabel metal4 s 21794 -2778 21974 31610 6 vssa2
port 1167 nsew ground bidirectional
rlabel metal4 s -2762 -2778 -2582 31610 4 vssa2
port 1168 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 29200
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_protect/runs/mgmt_protect/results/magic/mgmt_protect.gds
string GDS_END 7442798
string GDS_START 634152
<< end >>

