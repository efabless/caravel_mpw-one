sram_1rw1r_32_256_8_sky130.extracted.spice