magic
tech micross
magscale 1 2
timestamp 1611856895
<< checkpaint >>
rect 0 0 717600 1037600
<< pi1 >>
tri 80700 1027696 81760 1028756 se
rect 81760 1027696 87640 1028756
tri 87640 1027696 88700 1028756 sw
rect 80700 1021816 88700 1027696
tri 80700 1020756 81760 1021816 ne
rect 81760 1020756 87640 1021816
tri 87640 1020756 88700 1021816 nw
tri 132100 1027696 133160 1028756 se
rect 133160 1027696 139040 1028756
tri 139040 1027696 140100 1028756 sw
rect 132100 1021816 140100 1027696
tri 132100 1020756 133160 1021816 ne
rect 133160 1020756 139040 1021816
tri 139040 1020756 140100 1021816 nw
tri 183500 1027696 184560 1028756 se
rect 184560 1027696 190440 1028756
tri 190440 1027696 191500 1028756 sw
rect 183500 1021816 191500 1027696
tri 183500 1020756 184560 1021816 ne
rect 184560 1020756 190440 1021816
tri 190440 1020756 191500 1021816 nw
tri 234900 1027696 235960 1028756 se
rect 235960 1027696 241840 1028756
tri 241840 1027696 242900 1028756 sw
rect 234900 1021816 242900 1027696
tri 234900 1020756 235960 1021816 ne
rect 235960 1020756 241840 1021816
tri 241840 1020756 242900 1021816 nw
tri 286500 1027696 287560 1028756 se
rect 287560 1027696 293440 1028756
tri 293440 1027696 294500 1028756 sw
rect 286500 1021816 294500 1027696
tri 286500 1020756 287560 1021816 ne
rect 287560 1020756 293440 1021816
tri 293440 1020756 294500 1021816 nw
tri 336900 1027696 337960 1028756 se
rect 337960 1027696 343840 1028756
tri 343840 1027696 344900 1028756 sw
rect 336900 1021816 344900 1027696
tri 336900 1020756 337960 1021816 ne
rect 337960 1020756 343840 1021816
tri 343840 1020756 344900 1021816 nw
tri 388300 1027696 389360 1028756 se
rect 389360 1027696 395240 1028756
tri 395240 1027696 396300 1028756 sw
rect 388300 1021816 396300 1027696
tri 388300 1020756 389360 1021816 ne
rect 389360 1020756 395240 1021816
tri 395240 1020756 396300 1021816 nw
tri 477300 1027696 478360 1028756 se
rect 478360 1027696 484240 1028756
tri 484240 1027696 485300 1028756 sw
rect 477300 1021816 485300 1027696
tri 477300 1020756 478360 1021816 ne
rect 478360 1020756 484240 1021816
tri 484240 1020756 485300 1021816 nw
tri 528700 1027696 529760 1028756 se
rect 529760 1027696 535640 1028756
tri 535640 1027696 536700 1028756 sw
rect 528700 1021816 536700 1027696
tri 528700 1020756 529760 1021816 ne
rect 529760 1020756 535640 1021816
tri 535640 1020756 536700 1021816 nw
tri 579100 1027696 580160 1028756 se
rect 580160 1027696 586040 1028756
tri 586040 1027696 587100 1028756 sw
rect 579100 1021816 587100 1027696
tri 579100 1020756 580160 1021816 ne
rect 580160 1020756 586040 1021816
tri 586040 1020756 587100 1021816 nw
tri 630500 1027696 631560 1028756 se
rect 631560 1027696 637440 1028756
tri 637440 1027696 638500 1028756 sw
rect 630500 1021816 638500 1027696
tri 630500 1020756 631560 1021816 ne
rect 631560 1020756 637440 1021816
tri 637440 1020756 638500 1021816 nw
tri 8920 965640 9980 966700 se
rect 9980 965640 15860 966700
tri 15860 965640 16920 966700 sw
rect 8920 959760 16920 965640
tri 8920 958700 9980 959760 ne
rect 9980 958700 15860 959760
tri 15860 958700 16920 959760 nw
tri 700756 962040 701816 963100 se
rect 701816 962040 707696 963100
tri 707696 962040 708756 963100 sw
rect 700756 956160 708756 962040
tri 700756 955100 701816 956160 ne
rect 701816 955100 707696 956160
tri 707696 955100 708756 956160 nw
tri 8920 922440 9980 923500 se
rect 9980 922440 15860 923500
tri 15860 922440 16920 923500 sw
rect 8920 916560 16920 922440
tri 8920 915500 9980 916560 ne
rect 9980 915500 15860 916560
tri 15860 915500 16920 916560 nw
tri 700756 918040 701816 919100 se
rect 701816 918040 707696 919100
tri 707696 918040 708756 919100 sw
rect 700756 912160 708756 918040
tri 700756 911100 701816 912160 ne
rect 701816 911100 707696 912160
tri 707696 911100 708756 912160 nw
tri 8920 880240 9980 881300 se
rect 9980 880240 15860 881300
tri 15860 880240 16920 881300 sw
rect 8920 874360 16920 880240
tri 8920 873300 9980 874360 ne
rect 9980 873300 15860 874360
tri 15860 873300 16920 874360 nw
tri 700756 872840 701816 873900 se
rect 701816 872840 707696 873900
tri 707696 872840 708756 873900 sw
rect 700756 866960 708756 872840
tri 700756 865900 701816 866960 ne
rect 701816 865900 707696 866960
tri 707696 865900 708756 866960 nw
tri 8920 838040 9980 839100 se
rect 9980 838040 15860 839100
tri 15860 838040 16920 839100 sw
rect 8920 832160 16920 838040
tri 8920 831100 9980 832160 ne
rect 9980 831100 15860 832160
tri 15860 831100 16920 832160 nw
tri 700756 828840 701816 829900 se
rect 701816 828840 707696 829900
tri 707696 828840 708756 829900 sw
rect 700756 822960 708756 828840
tri 700756 821900 701816 822960 ne
rect 701816 821900 707696 822960
tri 707696 821900 708756 822960 nw
tri 8920 795840 9980 796900 se
rect 9980 795840 15860 796900
tri 15860 795840 16920 796900 sw
rect 8920 789960 16920 795840
tri 8920 788900 9980 789960 ne
rect 9980 788900 15860 789960
tri 15860 788900 16920 789960 nw
tri 700756 783640 701816 784700 se
rect 701816 783640 707696 784700
tri 707696 783640 708756 784700 sw
rect 700756 777760 708756 783640
tri 700756 776700 701816 777760 ne
rect 701816 776700 707696 777760
tri 707696 776700 708756 777760 nw
tri 8920 752640 9980 753700 se
rect 9980 752640 15860 753700
tri 15860 752640 16920 753700 sw
rect 8920 746760 16920 752640
tri 8920 745700 9980 746760 ne
rect 9980 745700 15860 746760
tri 15860 745700 16920 746760 nw
tri 700756 738640 701816 739700 se
rect 701816 738640 707696 739700
tri 707696 738640 708756 739700 sw
rect 700756 732760 708756 738640
tri 700756 731700 701816 732760 ne
rect 701816 731700 707696 732760
tri 707696 731700 708756 732760 nw
tri 8920 709440 9980 710500 se
rect 9980 709440 15860 710500
tri 15860 709440 16920 710500 sw
rect 8920 703560 16920 709440
tri 8920 702500 9980 703560 ne
rect 9980 702500 15860 703560
tri 15860 702500 16920 703560 nw
tri 700756 693640 701816 694700 se
rect 701816 693640 707696 694700
tri 707696 693640 708756 694700 sw
rect 700756 687760 708756 693640
tri 700756 686700 701816 687760 ne
rect 701816 686700 707696 687760
tri 707696 686700 708756 687760 nw
tri 8920 666240 9980 667300 se
rect 9980 666240 15860 667300
tri 15860 666240 16920 667300 sw
rect 8920 660360 16920 666240
tri 8920 659300 9980 660360 ne
rect 9980 659300 15860 660360
tri 15860 659300 16920 660360 nw
tri 700756 648440 701816 649500 se
rect 701816 648440 707696 649500
tri 707696 648440 708756 649500 sw
rect 700756 642560 708756 648440
tri 700756 641500 701816 642560 ne
rect 701816 641500 707696 642560
tri 707696 641500 708756 642560 nw
tri 8920 623040 9980 624100 se
rect 9980 623040 15860 624100
tri 15860 623040 16920 624100 sw
rect 8920 617160 16920 623040
tri 8920 616100 9980 617160 ne
rect 9980 616100 15860 617160
tri 15860 616100 16920 617160 nw
tri 700756 603440 701816 604500 se
rect 701816 603440 707696 604500
tri 707696 603440 708756 604500 sw
rect 700756 597560 708756 603440
tri 700756 596500 701816 597560 ne
rect 701816 596500 707696 597560
tri 707696 596500 708756 597560 nw
tri 8920 579840 9980 580900 se
rect 9980 579840 15860 580900
tri 15860 579840 16920 580900 sw
rect 8920 573960 16920 579840
tri 8920 572900 9980 573960 ne
rect 9980 572900 15860 573960
tri 15860 572900 16920 573960 nw
tri 700756 558240 701816 559300 se
rect 701816 558240 707696 559300
tri 707696 558240 708756 559300 sw
rect 700756 552360 708756 558240
tri 700756 551300 701816 552360 ne
rect 701816 551300 707696 552360
tri 707696 551300 708756 552360 nw
tri 8920 536640 9980 537700 se
rect 9980 536640 15860 537700
tri 15860 536640 16920 537700 sw
rect 8920 530760 16920 536640
tri 8920 529700 9980 530760 ne
rect 9980 529700 15860 530760
tri 15860 529700 16920 530760 nw
tri 700756 514240 701816 515300 se
rect 701816 514240 707696 515300
tri 707696 514240 708756 515300 sw
rect 700756 508360 708756 514240
tri 700756 507300 701816 508360 ne
rect 701816 507300 707696 508360
tri 707696 507300 708756 508360 nw
tri 8920 493440 9980 494500 se
rect 9980 493440 15860 494500
tri 15860 493440 16920 494500 sw
rect 8920 487560 16920 493440
tri 8920 486500 9980 487560 ne
rect 9980 486500 15860 487560
tri 15860 486500 16920 487560 nw
tri 700756 470240 701816 471300 se
rect 701816 470240 707696 471300
tri 707696 470240 708756 471300 sw
rect 700756 464360 708756 470240
tri 700756 463300 701816 464360 ne
rect 701816 463300 707696 464360
tri 707696 463300 708756 464360 nw
tri 8920 451240 9980 452300 se
rect 9980 451240 15860 452300
tri 15860 451240 16920 452300 sw
rect 8920 445360 16920 451240
tri 8920 444300 9980 445360 ne
rect 9980 444300 15860 445360
tri 15860 444300 16920 445360 nw
tri 700756 426040 701816 427100 se
rect 701816 426040 707696 427100
tri 707696 426040 708756 427100 sw
rect 700756 420160 708756 426040
tri 700756 419100 701816 420160 ne
rect 701816 419100 707696 420160
tri 707696 419100 708756 420160 nw
tri 8920 409040 9980 410100 se
rect 9980 409040 15860 410100
tri 15860 409040 16920 410100 sw
rect 8920 403160 16920 409040
tri 8920 402100 9980 403160 ne
rect 9980 402100 15860 403160
tri 15860 402100 16920 403160 nw
tri 700756 381040 701816 382100 se
rect 701816 381040 707696 382100
tri 707696 381040 708756 382100 sw
rect 700756 375160 708756 381040
tri 700756 374100 701816 375160 ne
rect 701816 374100 707696 375160
tri 707696 374100 708756 375160 nw
tri 8920 365840 9980 366900 se
rect 9980 365840 15860 366900
tri 15860 365840 16920 366900 sw
rect 8920 359960 16920 365840
tri 8920 358900 9980 359960 ne
rect 9980 358900 15860 359960
tri 15860 358900 16920 359960 nw
tri 700756 335840 701816 336900 se
rect 701816 335840 707696 336900
tri 707696 335840 708756 336900 sw
rect 700756 329960 708756 335840
tri 700756 328900 701816 329960 ne
rect 701816 328900 707696 329960
tri 707696 328900 708756 329960 nw
tri 8920 322640 9980 323700 se
rect 9980 322640 15860 323700
tri 15860 322640 16920 323700 sw
rect 8920 316760 16920 322640
tri 8920 315700 9980 316760 ne
rect 9980 315700 15860 316760
tri 15860 315700 16920 316760 nw
tri 700756 290840 701816 291900 se
rect 701816 290840 707696 291900
tri 707696 290840 708756 291900 sw
rect 700756 284960 708756 290840
tri 700756 283900 701816 284960 ne
rect 701816 283900 707696 284960
tri 707696 283900 708756 284960 nw
tri 8920 279440 9980 280500 se
rect 9980 279440 15860 280500
tri 15860 279440 16920 280500 sw
rect 8920 273560 16920 279440
tri 8920 272500 9980 273560 ne
rect 9980 272500 15860 273560
tri 15860 272500 16920 273560 nw
tri 700756 245840 701816 246900 se
rect 701816 245840 707696 246900
tri 707696 245840 708756 246900 sw
rect 700756 239960 708756 245840
tri 700756 238900 701816 239960 ne
rect 701816 238900 707696 239960
tri 707696 238900 708756 239960 nw
tri 8920 236240 9980 237300 se
rect 9980 236240 15860 237300
tri 15860 236240 16920 237300 sw
rect 8920 230360 16920 236240
tri 8920 229300 9980 230360 ne
rect 9980 229300 15860 230360
tri 15860 229300 16920 230360 nw
tri 700756 200640 701816 201700 se
rect 701816 200640 707696 201700
tri 707696 200640 708756 201700 sw
rect 700756 194760 708756 200640
tri 8920 193040 9980 194100 se
rect 9980 193040 15860 194100
tri 15860 193040 16920 194100 sw
tri 700756 193700 701816 194760 ne
rect 701816 193700 707696 194760
tri 707696 193700 708756 194760 nw
rect 8920 187160 16920 193040
tri 8920 186100 9980 187160 ne
rect 9980 186100 15860 187160
tri 15860 186100 16920 187160 nw
tri 700756 155640 701816 156700 se
rect 701816 155640 707696 156700
tri 707696 155640 708756 156700 sw
rect 700756 149760 708756 155640
tri 700756 148700 701816 149760 ne
rect 701816 148700 707696 149760
tri 707696 148700 708756 149760 nw
tri 8920 120640 9980 121700 se
rect 9980 120640 15860 121700
tri 15860 120640 16920 121700 sw
rect 8920 114760 16920 120640
tri 8920 113700 9980 114760 ne
rect 9980 113700 15860 114760
tri 15860 113700 16920 114760 nw
tri 700756 110440 701816 111500 se
rect 701816 110440 707696 111500
tri 707696 110440 708756 111500 sw
rect 700756 104560 708756 110440
tri 700756 103500 701816 104560 ne
rect 701816 103500 707696 104560
tri 707696 103500 708756 104560 nw
tri 8920 78440 9980 79500 se
rect 9980 78440 15860 79500
tri 15860 78440 16920 79500 sw
rect 8920 72560 16920 78440
tri 8920 71500 9980 72560 ne
rect 9980 71500 15860 72560
tri 15860 71500 16920 72560 nw
tri 82300 15860 83360 16920 se
rect 83360 15860 89240 16920
tri 89240 15860 90300 16920 sw
rect 82300 9980 90300 15860
tri 82300 8920 83360 9980 ne
rect 83360 8920 89240 9980
tri 89240 8920 90300 9980 nw
tri 136100 15860 137160 16920 se
rect 137160 15860 143040 16920
tri 143040 15860 144100 16920 sw
rect 136100 9980 144100 15860
tri 136100 8920 137160 9980 ne
rect 137160 8920 143040 9980
tri 143040 8920 144100 9980 nw
tri 189900 15860 190960 16920 se
rect 190960 15860 196840 16920
tri 196840 15860 197900 16920 sw
rect 189900 9980 197900 15860
tri 189900 8920 190960 9980 ne
rect 190960 8920 196840 9980
tri 196840 8920 197900 9980 nw
tri 244700 15860 245760 16920 se
rect 245760 15860 251640 16920
tri 251640 15860 252700 16920 sw
rect 244700 9980 252700 15860
tri 244700 8920 245760 9980 ne
rect 245760 8920 251640 9980
tri 251640 8920 252700 9980 nw
tri 298500 15860 299560 16920 se
rect 299560 15860 305440 16920
tri 305440 15860 306500 16920 sw
rect 298500 9980 306500 15860
tri 298500 8920 299560 9980 ne
rect 299560 8920 305440 9980
tri 305440 8920 306500 9980 nw
tri 353300 15860 354360 16920 se
rect 354360 15860 360240 16920
tri 360240 15860 361300 16920 sw
rect 353300 9980 361300 15860
tri 353300 8920 354360 9980 ne
rect 354360 8920 360240 9980
tri 360240 8920 361300 9980 nw
tri 408100 15860 409160 16920 se
rect 409160 15860 415040 16920
tri 415040 15860 416100 16920 sw
rect 408100 9980 416100 15860
tri 408100 8920 409160 9980 ne
rect 409160 8920 415040 9980
tri 415040 8920 416100 9980 nw
tri 462900 15860 463960 16920 se
rect 463960 15860 469840 16920
tri 469840 15860 470900 16920 sw
rect 462900 9980 470900 15860
tri 462900 8920 463960 9980 ne
rect 463960 8920 469840 9980
tri 469840 8920 470900 9980 nw
tri 517700 15860 518760 16920 se
rect 518760 15860 524640 16920
tri 524640 15860 525700 16920 sw
rect 517700 9980 525700 15860
tri 517700 8920 518760 9980 ne
rect 518760 8920 524640 9980
tri 524640 8920 525700 9980 nw
tri 572500 15860 573560 16920 se
rect 573560 15860 579440 16920
tri 579440 15860 580500 16920 sw
rect 572500 9980 580500 15860
tri 572500 8920 573560 9980 ne
rect 573560 8920 579440 9980
tri 579440 8920 580500 9980 nw
tri 626300 15860 627360 16920 se
rect 627360 15860 633240 16920
tri 633240 15860 634300 16920 sw
rect 626300 9980 634300 15860
tri 626300 8920 627360 9980 ne
rect 627360 8920 633240 9980
tri 633240 8920 634300 9980 nw
<< rdl >>
tri 79757 1030399 80114 1030756 se
rect 80114 1030399 89286 1030756
tri 89286 1030399 89643 1030756 sw
tri 131166 1030408 131514 1030756 se
rect 131514 1030408 140686 1030756
tri 140686 1030408 141034 1030756 sw
tri 182571 1030413 182914 1030756 se
rect 182914 1030413 192086 1030756
tri 192086 1030413 192429 1030756 sw
tri 79057 1029699 79757 1030399 se
rect 79757 1029699 89643 1030399
tri 78700 1029342 79057 1029699 se
rect 79057 1029342 89643 1029699
tri 89643 1029342 90700 1030399 sw
tri 130448 1029690 131166 1030408 se
rect 131166 1029690 141034 1030408
rect 78700 1028756 90700 1029342
rect 78700 1020756 80700 1028756
tri 80700 1027696 81760 1028756 nw
tri 87640 1027696 88700 1028756 ne
rect 88700 1024362 90700 1028756
tri 130100 1029342 130448 1029690 se
rect 130448 1029342 141034 1029690
tri 141034 1029342 142100 1030408 sw
tri 181843 1029685 182571 1030413 se
rect 182571 1029685 192429 1030413
rect 130100 1028756 142100 1029342
tri 90700 1024362 91249 1024839 sw
tri 80700 1020756 81760 1021816 sw
tri 87640 1020756 88700 1021816 se
rect 88700 1020756 91249 1024362
rect 78700 1020170 91249 1020756
tri 78700 1019813 79057 1020170 ne
rect 79057 1019822 91249 1020170
tri 91249 1019822 96470 1024362 sw
rect 130100 1020756 132100 1028756
tri 132100 1027696 133160 1028756 nw
tri 139040 1027696 140100 1028756 ne
rect 140100 1024530 142100 1028756
tri 181500 1029342 181843 1029685 se
rect 181843 1029591 192429 1029685
tri 192429 1029591 193251 1030413 sw
tri 233969 1030411 234314 1030756 se
rect 234314 1030411 243486 1030756
tri 243486 1030411 243831 1030756 sw
tri 233245 1029687 233969 1030411 se
rect 233969 1029964 243831 1030411
tri 243831 1029964 244278 1030411 sw
tri 285558 1030400 285914 1030756 se
rect 285914 1030400 295086 1030756
tri 295086 1030400 295442 1030756 sw
rect 233969 1029687 244278 1029964
rect 181843 1029342 193251 1029591
tri 193251 1029342 193500 1029591 sw
rect 181500 1028756 193500 1029342
tri 142100 1024530 142242 1024661 sw
tri 132100 1020756 133160 1021816 sw
tri 139040 1020756 140100 1021816 se
rect 140100 1020756 142242 1024530
rect 130100 1020170 142242 1020756
tri 130100 1019822 130448 1020170 ne
rect 130448 1019822 142242 1020170
rect 79057 1019813 96470 1019822
tri 79057 1018756 80114 1019813 ne
rect 80114 1018756 96470 1019813
tri 96470 1018756 97696 1019822 sw
tri 130448 1018756 131514 1019822 ne
rect 131514 1018756 142242 1019822
tri 142242 1018756 148496 1024530 sw
rect 181500 1020756 183500 1028756
tri 183500 1027696 184560 1028756 nw
tri 190440 1027696 191500 1028756 ne
tri 183500 1020756 184560 1021816 sw
tri 190440 1020756 191500 1021816 se
rect 191500 1020756 193500 1028756
tri 232900 1029342 233245 1029687 se
rect 233245 1029342 244278 1029687
tri 244278 1029342 244900 1029964 sw
tri 284856 1029698 285558 1030400 se
rect 285558 1030364 295442 1030400
tri 295442 1030364 295478 1030400 sw
tri 335953 1030395 336314 1030756 se
rect 336314 1030395 345486 1030756
tri 345486 1030395 345847 1030756 sw
rect 285558 1029698 295478 1030364
rect 232900 1028756 244900 1029342
rect 181500 1020170 193500 1020756
tri 181500 1019827 181843 1020170 ne
rect 181843 1019921 193500 1020170
tri 193500 1019921 198118 1024465 sw
rect 232900 1020756 234900 1028756
tri 234900 1027696 235960 1028756 nw
tri 241840 1027696 242900 1028756 ne
tri 234900 1020756 235960 1021816 sw
tri 241840 1020756 242900 1021816 se
rect 242900 1020756 244900 1028756
tri 284500 1029342 284856 1029698 se
rect 284856 1029342 295478 1029698
tri 295478 1029342 296500 1030364 sw
tri 335261 1029703 335953 1030395 se
rect 335953 1029703 345847 1030395
rect 284500 1028756 296500 1029342
rect 232900 1020170 244900 1020756
rect 181843 1019827 198118 1019921
tri 181843 1018756 182914 1019827 ne
rect 182914 1019825 198118 1019827
tri 198118 1019825 198216 1019921 sw
tri 232900 1019825 233245 1020170 ne
rect 233245 1019825 244900 1020170
rect 182914 1018756 198216 1019825
tri 198216 1018756 199302 1019825 sw
tri 233245 1018756 234314 1019825 ne
rect 234314 1019548 244900 1019825
tri 244900 1019548 249361 1024246 sw
rect 284500 1020756 286500 1028756
tri 286500 1027696 287560 1028756 nw
tri 293440 1027696 294500 1028756 ne
tri 286500 1020756 287560 1021816 sw
tri 293440 1020756 294500 1021816 se
rect 294500 1020756 296500 1028756
tri 334900 1029342 335261 1029703 se
rect 335261 1029342 345847 1029703
tri 345847 1029342 346900 1030395 sw
tri 387331 1030373 387714 1030756 se
rect 387714 1030373 396886 1030756
tri 386683 1029725 387331 1030373 se
rect 387331 1029725 396886 1030373
rect 334900 1028756 346900 1029342
rect 284500 1020170 296500 1020756
tri 284500 1019814 284856 1020170 ne
rect 284856 1019814 296500 1020170
rect 234314 1018757 249361 1019548
tri 249361 1018757 250113 1019548 sw
rect 234314 1018756 250113 1018757
tri 284856 1018756 285914 1019814 ne
rect 285914 1019809 296500 1019814
tri 296500 1019809 300131 1023967 sw
rect 334900 1020756 336900 1028756
tri 336900 1027696 337960 1028756 nw
tri 343840 1027696 344900 1028756 ne
tri 336900 1020756 337960 1021816 sw
tri 343840 1020756 344900 1021816 se
rect 344900 1020756 346900 1028756
tri 386300 1029342 386683 1029725 se
rect 386683 1029342 396886 1029725
tri 396886 1029342 398300 1030756 sw
tri 476367 1030409 476714 1030756 se
rect 476714 1030409 485886 1030756
tri 485886 1030409 486233 1030756 sw
rect 386300 1028756 398300 1029342
rect 334900 1020170 346900 1020756
tri 334900 1019809 335261 1020170 ne
rect 335261 1019809 346900 1020170
rect 285914 1019148 300131 1019809
tri 300131 1019148 300708 1019809 sw
rect 285914 1018756 300708 1019148
tri 300708 1018756 301050 1019148 sw
tri 335261 1018756 336314 1019809 ne
rect 336314 1019052 346900 1019809
tri 346900 1019052 351033 1023891 sw
rect 386300 1020756 388300 1028756
tri 388300 1027696 389360 1028756 nw
tri 395240 1027696 396300 1028756 ne
tri 388300 1020756 389360 1021816 sw
tri 395240 1020756 396300 1021816 se
rect 396300 1020756 398300 1028756
tri 475300 1029342 476367 1030409 se
rect 476367 1029689 486233 1030409
tri 486233 1029689 486953 1030409 sw
rect 476367 1029342 486953 1029689
tri 486953 1029342 487300 1029689 sw
tri 526774 1029416 528114 1030756 se
rect 528114 1029416 537286 1030756
tri 537286 1029416 538626 1030756 sw
tri 578130 1030372 578514 1030756 se
rect 578514 1030372 587686 1030756
tri 587686 1030372 588070 1030756 sw
tri 629542 1030384 629914 1030756 se
rect 629914 1030384 639086 1030756
tri 639086 1030384 639458 1030756 sw
rect 475300 1028756 487300 1029342
rect 386300 1020170 398300 1020756
tri 386300 1019787 386683 1020170 ne
rect 386683 1019787 398300 1020170
rect 336314 1018756 351033 1019052
tri 351033 1018756 351286 1019052 sw
tri 386683 1018756 387714 1019787 ne
rect 387714 1019477 398300 1019787
tri 398300 1019477 401547 1023601 sw
tri 469764 1019477 475300 1024633 se
rect 475300 1020756 477300 1028756
tri 477300 1027696 478360 1028756 nw
tri 484240 1027696 485300 1028756 ne
tri 477300 1020756 478360 1021816 sw
tri 484240 1020756 485300 1021816 se
rect 485300 1020756 487300 1028756
rect 475300 1020170 487300 1020756
rect 475300 1019823 486953 1020170
tri 486953 1019823 487300 1020170 nw
tri 526700 1029342 526774 1029416 se
rect 526774 1029342 538626 1029416
tri 538626 1029342 538700 1029416 sw
rect 526700 1028756 538700 1029342
rect 526700 1020756 528700 1028756
tri 528700 1027696 529760 1028756 nw
tri 535640 1027696 536700 1028756 ne
tri 528700 1020756 529760 1021816 sw
tri 535640 1020756 536700 1021816 se
rect 536700 1020756 538700 1028756
tri 577100 1029342 578130 1030372 se
rect 578130 1029726 588070 1030372
tri 588070 1029726 588716 1030372 sw
rect 578130 1029342 588716 1029726
tri 588716 1029342 589100 1029726 sw
rect 577100 1028756 589100 1029342
rect 526700 1020170 538700 1020756
rect 475300 1019477 486607 1019823
tri 486607 1019477 486953 1019823 nw
rect 387714 1018756 401547 1019477
tri 401547 1018756 402115 1019477 sw
tri 468990 1018756 469764 1019477 se
rect 469764 1018756 485886 1019477
tri 485886 1018756 486607 1019477 nw
tri 526700 1018830 528040 1020170 ne
rect 528040 1019270 537800 1020170
tri 537800 1019270 538700 1020170 nw
rect 528040 1019254 537784 1019270
tri 537784 1019254 537800 1019270 nw
rect 528040 1019166 537783 1019254
tri 537783 1019253 537784 1019254 nw
tri 537783 1019166 537800 1019250 sw
rect 528040 1018830 537800 1019166
tri 528040 1018756 528114 1018830 ne
rect 528114 1018756 537800 1018830
tri 573305 1018756 577100 1023591 se
rect 577100 1020756 579100 1028756
tri 579100 1027696 580160 1028756 nw
tri 586040 1027696 587100 1028756 ne
tri 579100 1020756 580160 1021816 sw
tri 586040 1020756 587100 1021816 se
rect 587100 1020756 589100 1028756
tri 628500 1029342 629542 1030384 se
rect 629542 1029714 639458 1030384
tri 639458 1029714 640128 1030384 sw
rect 629542 1029342 640128 1029714
tri 640128 1029342 640500 1029714 sw
rect 628500 1028756 640500 1029342
rect 577100 1020170 589100 1020756
rect 577100 1019786 588716 1020170
tri 588716 1019786 589100 1020170 nw
tri 622413 1020061 628500 1025025 se
rect 628500 1020756 630500 1028756
tri 630500 1027696 631560 1028756 nw
tri 637440 1027696 638500 1028756 ne
tri 630500 1020756 631560 1021816 sw
tri 637440 1020756 638500 1021816 se
rect 638500 1020756 640500 1028756
rect 628500 1020170 640500 1020756
rect 628500 1020061 640391 1020170
tri 640391 1020061 640500 1020170 nw
tri 622076 1019786 622413 1020061 se
rect 622413 1019786 639086 1020061
rect 577100 1018756 587686 1019786
tri 587686 1018756 588716 1019786 nw
tri 620813 1018756 622076 1019786 se
rect 622076 1018756 639086 1019786
tri 639086 1018756 640391 1020061 nw
tri 85504 1013761 91249 1018756 ne
rect 91249 1013761 97696 1018756
tri 97696 1013761 103441 1018756 sw
tri 91249 1013643 91384 1013761 ne
rect 91384 1013643 103441 1013761
tri 103441 1013643 103576 1013761 sw
tri 136703 1013643 142242 1018756 ne
rect 142242 1013643 148496 1018756
tri 148496 1013643 154035 1018756 sw
tri 187895 1013643 193092 1018756 ne
rect 193092 1013643 199302 1018756
tri 199302 1013643 204499 1018756 sw
tri 239081 1013643 243937 1018756 ne
rect 243937 1013821 250113 1018756
tri 250113 1013821 254800 1018756 sw
tri 290429 1013821 294739 1018756 ne
rect 294739 1014462 301050 1018756
tri 301050 1014462 304800 1018756 sw
rect 294739 1013821 304800 1014462
rect 243937 1013643 254800 1013821
tri 91384 1012883 92258 1013643 ne
rect 92258 1012883 103576 1013643
tri 103576 1012883 104450 1013643 sw
tri 142242 1012883 143065 1013643 ne
rect 143065 1012883 154035 1013643
tri 154035 1012883 154858 1013643 sw
tri 193092 1013487 193251 1013643 ne
rect 193251 1013487 204499 1013643
tri 204499 1013487 204658 1013643 sw
tri 193251 1013284 193457 1013487 ne
rect 193457 1013284 204658 1013487
tri 204658 1013284 204864 1013487 sw
tri 243937 1013284 244278 1013643 ne
rect 244278 1013285 254800 1013643
tri 254800 1013285 255309 1013821 sw
rect 244278 1013284 255309 1013285
tri 294739 1013284 295208 1013821 ne
rect 295208 1013284 304800 1013821
tri 193457 1012883 193864 1013284 ne
rect 193864 1012883 204864 1013284
tri 204864 1012883 205271 1013284 sw
tri 244278 1012883 244658 1013284 ne
rect 244658 1012883 255309 1013284
tri 255309 1012883 255690 1013284 sw
tri 295208 1012975 295478 1013284 ne
rect 295478 1012975 304800 1013284
tri 304800 1012975 306098 1014462 sw
tri 295478 1012883 295558 1012975 ne
rect 295558 1012884 306098 1012975
tri 306098 1012884 306178 1012975 sw
rect 295558 1012883 306178 1012884
tri 340765 1012883 345782 1018756 ne
rect 345782 1014642 351286 1018756
tri 351286 1014642 354800 1018756 sw
tri 391933 1017416 392988 1018756 ne
rect 392988 1017416 402115 1018756
tri 402115 1017416 403170 1018756 sw
tri 467551 1017416 468990 1018756 se
rect 468990 1017416 479288 1018756
tri 479288 1017416 480727 1018756 nw
tri 529740 1018434 529800 1018756 ne
tri 392988 1014643 395172 1017416 ne
rect 395172 1015346 403170 1017416
tri 403170 1015346 404800 1017416 sw
rect 395172 1014642 404800 1015346
tri 404800 1014642 405354 1015346 sw
tri 464573 1014642 467551 1017416 se
rect 467551 1014642 476310 1017416
tri 476310 1014642 479288 1017416 nw
rect 345782 1012883 354800 1014642
tri 354800 1012883 356302 1014642 sw
tri 395172 1012884 396557 1014642 ne
rect 396557 1012883 405354 1014642
tri 405354 1012883 406739 1014642 sw
tri 462684 1012883 464573 1014642 se
rect 464573 1012883 474421 1014642
tri 474421 1012883 476310 1014642 nw
tri 92258 1003159 103441 1012883 ne
rect 103441 1005623 104450 1012883
tri 104450 1005623 112800 1012883 sw
rect 103441 1003159 112800 1005623
tri 103441 1002756 103904 1003159 ne
rect 103904 1002756 112800 1003159
tri 143065 1002756 154035 1012883 ne
rect 154035 1005551 154858 1012883
tri 154858 1005551 162800 1012883 sw
rect 154035 1002756 162800 1005551
tri 103904 1002324 104401 1002756 ne
rect 104401 1002324 112800 1002756
tri 154035 1002324 154502 1002756 ne
rect 154502 1002324 162800 1002756
tri 193864 1002324 204597 1012883 ne
rect 204597 1005476 205271 1012883
tri 205271 1005476 212800 1012883 sw
rect 204597 1002324 212800 1005476
tri 244658 1002324 254685 1012883 ne
rect 254685 1005397 255690 1012883
tri 255690 1005397 262800 1012883 sw
rect 254685 1002324 262800 1005397
tri 295558 1002324 304778 1012883 ne
rect 304778 1005301 306178 1012883
tri 306178 1005301 312800 1012883 sw
rect 304778 1002324 312800 1005301
tri 345782 1002324 354800 1012883 ne
rect 354800 1005276 356302 1012883
tri 356302 1005276 362800 1012883 sw
tri 396557 1012493 396865 1012883 ne
rect 396865 1012493 406739 1012883
tri 406739 1012493 407046 1012883 sw
tri 396865 1008545 399973 1012493 ne
rect 399973 1008545 407046 1012493
tri 407046 1008545 410155 1012493 sw
tri 458026 1008545 462684 1012883 se
rect 462684 1008545 469764 1012883
tri 469764 1008545 474421 1012883 nw
tri 104401 1002049 104717 1002324 ne
rect 104717 1002049 112800 1002324
tri 154502 1002049 154800 1002324 ne
tri 104717 1001977 104800 1002049 ne
tri 7989 968355 8334 968700 se
rect 8334 968355 17506 968700
tri 17506 968355 17851 968700 sw
tri 7265 967631 7989 968355 se
rect 7989 967631 17851 968355
tri 6920 967286 7265 967631 se
rect 7265 967370 17851 967631
tri 17851 967370 18836 968355 sw
rect 7265 967286 18836 967370
tri 18836 967286 18920 967370 sw
rect 6920 966700 18920 967286
rect 6920 958700 8920 966700
tri 8920 965640 9980 966700 nw
tri 15860 965640 16920 966700 ne
tri 8920 958700 9980 959760 sw
tri 15860 958700 16920 959760 se
rect 16920 958700 18920 966700
rect 104800 964800 112800 1002049
rect 6920 958114 18920 958700
tri 6920 957769 7265 958114 ne
rect 7265 958030 18920 958114
tri 18920 958030 23586 962494 sw
rect 7265 957769 23586 958030
tri 7265 956700 8334 957769 ne
rect 8334 956700 23586 957769
tri 13405 951504 18836 956700 ne
rect 18836 951504 23586 956700
tri 23586 951504 30407 958030 sw
tri 18836 940433 30407 951504 ne
tri 30407 940433 41978 951504 sw
tri 30407 929361 41978 940433 ne
tri 41978 929361 53549 940433 sw
tri 41978 925500 46013 929361 ne
rect 46013 925500 53549 929361
tri 7991 925157 8334 925500 se
rect 8334 925157 17506 925500
tri 17506 925157 17849 925500 sw
tri 7263 924429 7991 925157 se
rect 7991 924429 17849 925157
tri 6920 924086 7263 924429 se
rect 7263 924389 17849 924429
tri 17849 924389 18617 925157 sw
rect 7263 924086 18617 924389
tri 18617 924086 18920 924389 sw
rect 6920 923500 18920 924086
rect 6920 915500 8920 923500
tri 8920 922440 9980 923500 nw
tri 15860 922440 16920 923500 ne
rect 16920 918289 18920 923500
tri 18920 918289 19816 919179 sw
tri 46013 918289 53549 925500 ne
tri 53549 922800 60405 929361 sw
rect 53549 918289 135457 922800
tri 135457 918289 139968 922800 sw
rect 154800 918289 162800 1002324
tri 204597 1002264 204658 1002324 ne
rect 204658 1002264 212800 1002324
tri 204658 1002203 204719 1002264 ne
rect 204719 1002203 212800 1002264
tri 254685 1002203 254800 1002324 ne
tri 204719 1002124 204800 1002203 ne
rect 204800 964800 212800 1002203
tri 162800 918289 164968 920457 sw
rect 254800 918289 262800 1002324
tri 304778 1002299 304800 1002324 ne
rect 304800 964800 312800 1002324
tri 262800 918289 264968 920457 sw
tri 8920 915500 9980 916560 sw
tri 15860 915500 16920 916560 se
rect 16920 915500 19816 918289
rect 6920 914914 19816 915500
tri 6920 914571 7263 914914 ne
rect 7263 914800 19816 914914
tri 19816 914800 23330 918289 sw
tri 53549 914800 57195 918289 ne
rect 57195 914800 139968 918289
tri 139968 914800 143457 918289 sw
rect 154800 917143 164968 918289
tri 164968 917143 166114 918289 sw
rect 254800 917143 264968 918289
tri 264968 917143 266114 918289 sw
tri 154800 914800 157143 917143 ne
rect 157143 914800 166114 917143
rect 7263 914611 23330 914800
tri 23330 914611 23520 914800 sw
rect 7263 914571 23520 914611
tri 7263 913500 8334 914571 ne
rect 8334 913500 23520 914571
tri 23520 913500 24639 914611 sw
tri 132143 913500 133443 914800 ne
rect 133443 913500 143457 914800
tri 13285 908206 18617 913500 ne
rect 18617 908206 24639 913500
tri 24639 908206 29971 913500 sw
tri 18617 903486 23370 908206 ne
rect 23370 903486 29971 908206
tri 29971 903486 34723 908206 sw
tri 133443 903486 143457 913500 ne
tri 143457 903486 154771 914800 sw
tri 157143 905829 166114 914800 ne
tri 166114 905829 177428 917143 sw
tri 254800 905829 266114 917143 ne
tri 266114 905829 277428 917143 sw
tri 166114 903486 168457 905829 ne
rect 168457 903486 177428 905829
tri 23370 896931 29971 903486 ne
rect 29971 897800 34723 903486
tri 34723 897800 40449 903486 sw
rect 29971 896931 85457 897800
tri 85457 896931 86326 897800 sw
tri 29971 892172 34762 896931 ne
rect 34762 892172 86326 896931
tri 86326 892172 91085 896931 sw
tri 143457 892172 154771 903486 ne
tri 154771 895457 162800 903486 sw
rect 154771 892172 162800 895457
tri 168457 894515 177428 903486 ne
tri 177428 894515 188742 905829 sw
tri 266114 894515 277428 905829 ne
tri 277428 894515 288742 905829 sw
tri 34762 892143 34791 892172 ne
rect 34791 892143 91085 892172
tri 91085 892143 91114 892172 sw
tri 154771 892143 154800 892172 ne
tri 34791 889800 37151 892143 ne
rect 37151 889800 91114 892143
tri 91114 889800 93457 892143 sw
tri 82143 883300 88643 889800 ne
rect 88643 883300 93457 889800
tri 7989 882955 8334 883300 se
rect 8334 882955 17506 883300
tri 17506 882955 17851 883300 sw
tri 88643 882955 88988 883300 ne
rect 88988 882955 93457 883300
tri 7265 882231 7989 882955 se
rect 7989 882231 17851 882955
tri 6920 881886 7265 882231 se
rect 7265 881946 17851 882231
tri 17851 881946 18860 882955 sw
tri 88988 881946 89997 882955 ne
rect 89997 881946 93457 882955
rect 7265 881886 18860 881946
tri 18860 881886 18920 881946 sw
rect 6920 881300 18920 881886
rect 6920 873300 8920 881300
tri 8920 880240 9980 881300 nw
tri 15860 880240 16920 881300 ne
tri 8920 873300 9980 874360 sw
tri 15860 873300 16920 874360 se
rect 16920 873300 18920 881300
tri 89997 878486 93457 881946 ne
tri 93457 878486 104771 889800 sw
tri 93457 877107 94836 878486 ne
rect 94836 877107 104771 878486
rect 6920 872714 18920 873300
tri 6920 872369 7265 872714 ne
rect 7265 872654 18920 872714
tri 18920 872654 23592 877107 sw
tri 94836 872654 99289 877107 ne
rect 99289 872654 104771 877107
rect 7265 872369 23592 872654
tri 7265 871300 8334 872369 ne
rect 8334 871300 23592 872369
tri 13418 866113 18860 871300 ne
rect 18860 866113 23592 871300
tri 23592 866113 30455 872654 sw
tri 99289 867172 104771 872654 ne
tri 104771 868800 114457 878486 sw
rect 104771 867172 112829 868800
tri 112829 867172 114457 868800 nw
tri 104771 866113 105830 867172 ne
rect 105830 866113 108800 867172
tri 18860 855061 30455 866113 ne
tri 30455 855061 42049 866113 sw
tri 105830 863143 108800 866113 ne
tri 108800 863143 112829 867172 nw
tri 30455 844009 42049 855061 ne
tri 42049 844009 53643 855061 sw
rect 154800 844009 162800 892172
tri 177428 883201 188742 894515 ne
tri 188742 883201 200056 894515 sw
tri 277428 883201 288742 894515 ne
tri 288742 883201 300056 894515 sw
tri 188742 871887 200056 883201 ne
tri 200056 874457 208800 883201 sw
tri 288742 874457 297486 883201 ne
rect 297486 874457 300056 883201
tri 300056 874457 308800 883201 sw
rect 200056 871887 208800 874457
tri 208800 871887 211370 874457 sw
tri 297486 871887 300056 874457 ne
rect 300056 871887 308800 874457
tri 308800 871887 311370 874457 sw
tri 200056 863143 208800 871887 ne
rect 208800 868800 211370 871887
tri 211370 868800 214457 871887 sw
tri 208800 863143 214457 868800 nw
tri 300056 863143 308800 871887 ne
rect 308800 868800 311370 871887
tri 311370 868800 314457 871887 sw
tri 308800 863143 314457 868800 nw
tri 162800 844009 164248 845457 sw
tri 42049 841100 45100 844009 ne
rect 45100 841100 53643 844009
tri 7991 840757 8334 841100 se
rect 8334 840757 17506 841100
tri 17506 840757 17849 841100 sw
tri 7263 840029 7991 840757 se
rect 7991 840118 17849 840757
tri 17849 840118 18488 840757 sw
rect 7991 840029 18488 840118
tri 6920 839686 7263 840029 se
rect 7263 839686 18488 840029
tri 18488 839686 18920 840118 sw
rect 6920 839100 18920 839686
rect 6920 831100 8920 839100
tri 8920 838040 9980 839100 nw
tri 15860 838040 16920 839100 ne
rect 16920 832957 18920 839100
tri 18920 832957 20642 834706 sw
tri 45100 832957 53643 841100 ne
tri 53643 835852 62199 844009 sw
rect 154800 842143 164248 844009
tri 164248 842143 166114 844009 sw
tri 154800 835852 161091 842143 ne
rect 161091 835852 166114 842143
rect 53643 832957 62199 835852
tri 62199 832957 65236 835852 sw
tri 161091 832957 163986 835852 ne
rect 163986 832957 166114 835852
tri 8920 831100 9980 832160 sw
tri 15860 831100 16920 832160 se
rect 16920 831100 20642 832957
rect 6920 830514 20642 831100
tri 6920 830171 7263 830514 ne
rect 7263 830171 20642 830514
tri 7263 829100 8334 830171 ne
rect 8334 830082 20642 830171
tri 20642 830082 23471 832957 sw
rect 8334 829100 23471 830082
tri 23471 829100 24437 830082 sw
tri 53643 829100 57688 832957 ne
rect 57688 832800 65236 832957
tri 65236 832800 65401 832957 sw
tri 163986 832800 164143 832957 ne
rect 164143 832800 166114 832957
tri 166114 832800 175457 842143 sw
rect 57688 829100 140457 832800
tri 13212 824800 17443 829100 ne
rect 17443 824800 24437 829100
tri 24437 824800 28668 829100 sw
tri 57688 824800 62199 829100 ne
rect 62199 824800 140457 829100
tri 140457 824800 148457 832800 sw
tri 164143 830829 166114 832800 ne
rect 166114 830829 250457 832800
tri 250457 830829 252428 832800 sw
tri 166114 824800 172143 830829 ne
rect 172143 824800 252428 830829
tri 252428 824800 258457 830829 sw
tri 17443 823739 18488 824800 ne
rect 18488 823739 28668 824800
tri 28668 823739 29713 824800 sw
tri 18488 820457 21717 823739 ne
rect 21717 820457 29713 823739
tri 29713 820457 32942 823739 sw
tri 137143 820457 141486 824800 ne
rect 141486 820457 148457 824800
tri 148457 820457 152800 824800 sw
tri 247143 820457 251486 824800 ne
rect 251486 820457 258457 824800
tri 258457 820457 262800 824800 sw
tri 21717 819900 22265 820457 ne
rect 22265 819900 32942 820457
tri 32942 819900 33490 820457 sw
tri 141486 819900 142043 820457 ne
rect 142043 819900 152800 820457
tri 152800 819900 153357 820457 sw
tri 251486 819900 252043 820457 ne
rect 252043 819900 262800 820457
tri 262800 819900 263357 820457 sw
tri 354243 819900 354800 820457 se
rect 354800 819900 362800 1005276
tri 399973 1002414 404800 1008545 ne
rect 404800 1005186 410155 1008545
tri 410155 1005186 412800 1008545 sw
rect 404800 964800 412800 1005186
tri 454800 1005541 458026 1008545 se
rect 458026 1005541 466539 1008545
tri 466539 1005541 469764 1008545 nw
rect 454800 1004460 465378 1005541
tri 465378 1004460 466539 1005541 nw
tri 445829 911486 454800 920457 se
rect 454800 917143 462800 1004460
tri 462800 1002059 465378 1004460 nw
tri 518486 984143 529800 995457 se
rect 529800 992143 537800 1018756
tri 572253 1017416 573305 1018756 se
rect 573305 1017416 582423 1018756
tri 582423 1017416 583475 1018756 nw
tri 619169 1017416 620813 1018756 se
rect 620813 1017416 622413 1018756
tri 570076 1014643 572253 1017416 se
tri 568695 1012883 570076 1014642 se
rect 570076 1012883 572253 1014643
tri 562083 1004460 568695 1012883 se
rect 568695 1004460 572253 1012883
tri 572253 1004460 582423 1017416 nw
tri 609753 1009738 619169 1017416 se
rect 619169 1009738 622413 1017416
tri 622413 1009738 633472 1018756 nw
tri 604800 1005700 609753 1009738 se
rect 609753 1005700 617461 1009738
tri 617461 1005700 622413 1009738 nw
rect 604800 1004460 615940 1005700
tri 615940 1004460 617461 1005700 nw
tri 529800 984143 537800 992143 nw
tri 554800 995182 562083 1004460 se
rect 562083 995182 564970 1004460
tri 564970 995182 572253 1004460 nw
tri 507172 972829 518486 984143 se
tri 518486 972829 529800 984143 nw
tri 503143 968800 507172 972829 se
rect 507172 968800 514457 972829
tri 514457 968800 518486 972829 nw
tri 503143 963143 508800 968800 ne
tri 508800 963143 514457 968800 nw
tri 543486 934143 554800 945457 se
rect 554800 942143 562800 995182
tri 562800 992418 564970 995182 nw
rect 604800 964800 612800 1004460
tri 612800 1001900 615940 1004460 nw
tri 699826 964756 700170 965100 se
rect 700170 964756 709342 965100
tri 709342 964756 709686 965100 sw
tri 698756 963686 699826 964756 se
rect 699826 964030 709686 964756
tri 709686 964030 710412 964756 sw
rect 699826 963686 710412 964030
tri 710412 963686 710756 964030 sw
rect 698756 963100 710756 963686
tri 693315 953671 698756 958888 se
rect 698756 955100 700756 963100
tri 700756 962040 701816 963100 nw
tri 707696 962040 708756 963100 ne
tri 700756 955100 701816 956160 sw
tri 707696 955100 708756 956160 se
rect 708756 955100 710756 963100
rect 698756 954514 710756 955100
rect 698756 954170 710412 954514
tri 710412 954170 710756 954514 nw
rect 698756 953671 709913 954170
tri 709913 953671 710412 954170 nw
tri 692719 953100 693315 953671 se
rect 693315 953100 709342 953671
tri 709342 953100 709913 953671 nw
tri 687192 947800 692719 953100 se
rect 692719 947800 698751 953100
tri 698751 947800 704279 953100 nw
tri 554800 934143 562800 942143 nw
tri 645829 936486 657143 947800 se
rect 657143 939800 690408 947800
tri 690408 939800 698751 947800 nw
tri 657143 936486 660457 939800 nw
tri 643486 934143 645829 936486 se
tri 532172 922829 543486 934143 se
tri 543486 922829 554800 934143 nw
tri 634515 925172 643486 934143 se
rect 643486 925172 645829 934143
tri 645829 925172 657143 936486 nw
tri 632172 922829 634515 925172 se
rect 634515 922829 643457 925172
tri 532143 922800 532172 922829 se
rect 532172 922800 543457 922829
tri 543457 922800 543486 922829 nw
tri 632143 922800 632172 922829 se
rect 632172 922800 643457 922829
tri 643457 922800 645829 925172 nw
tri 480443 921100 482143 922800 se
rect 482143 921100 541757 922800
tri 541757 921100 543457 922800 nw
tri 555443 921100 557143 922800 se
rect 557143 921100 641757 922800
tri 641757 921100 643457 922800 nw
rect 454800 911486 457143 917143
tri 457143 911486 462800 917143 nw
tri 470829 911486 480443 921100 se
rect 480443 914800 535457 921100
tri 535457 914800 541757 921100 nw
tri 549143 914800 555443 921100 se
rect 555443 914800 635457 921100
tri 635457 914800 641757 921100 nw
tri 699827 920757 700170 921100 se
rect 700170 920757 709342 921100
tri 709342 920757 709685 921100 sw
tri 698756 919686 699827 920757 se
rect 699827 920029 709685 920757
tri 709685 920029 710413 920757 sw
rect 699827 919686 710413 920029
tri 710413 919686 710756 920029 sw
rect 698756 919100 710756 919686
rect 480443 911486 482143 914800
tri 482143 911486 485457 914800 nw
tri 545829 911486 549143 914800 se
rect 549143 911486 557143 914800
tri 557143 911486 560457 914800 nw
tri 695589 911486 698756 914705 se
rect 698756 911486 700756 919100
tri 700756 918040 701816 919100 nw
tri 707696 918040 708756 919100 ne
tri 443486 909143 445829 911486 se
rect 445829 909143 454800 911486
tri 454800 909143 457143 911486 nw
tri 443443 909100 443486 909143 se
rect 443486 909100 454757 909143
tri 454757 909100 454800 909143 nw
tri 468443 909100 470829 911486 se
rect 470829 909100 479757 911486
tri 479757 909100 482143 911486 nw
tri 543443 909100 545829 911486 se
rect 545829 909100 554757 911486
tri 554757 909100 557143 911486 nw
tri 693487 909349 695589 911486 se
rect 695589 911100 700756 911486
tri 700756 911100 701816 912160 sw
tri 707696 911100 708756 912160 se
rect 708756 911100 710756 919100
rect 695589 910514 710756 911100
rect 695589 910171 710413 910514
tri 710413 910171 710756 910514 nw
rect 695589 909349 709591 910171
tri 709591 909349 710413 910171 nw
tri 693242 909100 693487 909349 se
rect 693487 909100 709342 909349
tri 709342 909100 709591 909349 nw
tri 434515 900172 443443 909100 se
rect 443443 900172 445829 909100
tri 445829 900172 454757 909100 nw
tri 459515 900172 468443 909100 se
rect 468443 900172 470829 909100
tri 470829 900172 479757 909100 nw
tri 534515 900172 543443 909100 se
rect 543443 900172 545829 909100
tri 545829 900172 554757 909100 nw
tri 684458 900172 693242 909100 se
rect 693242 900172 693487 909100
tri 432172 897829 434515 900172 se
rect 434515 897829 443486 900172
tri 443486 897829 445829 900172 nw
tri 420858 886515 432172 897829 se
tri 432172 886515 443486 897829 nw
tri 454800 895457 459515 900172 se
rect 459515 895457 466114 900172
tri 466114 895457 470829 900172 nw
tri 529800 895457 534515 900172 se
tri 409544 875201 420858 886515 se
tri 420858 875201 432172 886515 nw
tri 403143 868800 409544 875201 se
rect 409544 868800 414457 875201
tri 414457 868800 420858 875201 nw
tri 403143 863143 408800 868800 ne
tri 408800 863143 414457 868800 nw
tri 443486 834143 454800 845457 se
rect 454800 842143 462800 895457
tri 462800 892143 466114 895457 nw
tri 526486 892143 529800 895457 se
rect 529800 892143 534515 895457
tri 523201 888858 526486 892143 se
rect 526486 888858 534515 892143
tri 534515 888858 545829 900172 nw
tri 682264 897942 684458 900172 se
rect 684458 897942 693487 900172
tri 693487 897942 704465 909100 nw
tri 682124 897800 682264 897942 se
rect 682264 897800 693347 897942
tri 693347 897800 693487 897942 nw
tri 623201 888858 632143 897800 se
rect 632143 889800 685476 897800
tri 685476 889800 693347 897800 nw
tri 511887 877544 523201 888858 se
tri 523201 877544 534515 888858 nw
tri 620829 886486 623201 888858 se
rect 623201 886486 632143 888858
tri 632143 886486 635457 889800 nw
tri 611887 877544 620829 886486 se
rect 620829 877544 621557 886486
tri 510243 875900 511887 877544 se
rect 511887 875900 521557 877544
tri 521557 875900 523201 877544 nw
tri 610243 875900 611887 877544 se
rect 611887 875900 621557 877544
tri 621557 875900 632143 886486 nw
tri 509891 875548 510243 875900 se
rect 510243 875548 521205 875900
tri 521205 875548 521557 875900 nw
tri 609891 875548 610243 875900 se
rect 610243 875548 621205 875900
tri 621205 875548 621557 875900 nw
tri 699818 875548 700170 875900 se
rect 700170 875548 709342 875900
tri 709342 875548 709694 875900 sw
tri 504243 869900 509891 875548 se
rect 509891 869900 515557 875548
tri 515557 869900 521205 875548 nw
tri 609515 875172 609891 875548 se
rect 609891 875172 620829 875548
tri 620829 875172 621205 875548 nw
tri 604243 869900 609515 875172 se
rect 609515 869900 615557 875172
tri 615557 869900 620829 875172 nw
tri 698756 874486 699818 875548 se
rect 699818 874838 709694 875548
tri 709694 874838 710404 875548 sw
rect 699818 874486 710404 874838
tri 710404 874486 710756 874838 sw
rect 698756 873900 710756 874486
tri 503143 868800 504243 869900 se
rect 504243 868800 514457 869900
tri 514457 868800 515557 869900 nw
tri 603143 868800 604243 869900 se
rect 604243 868800 614457 869900
tri 614457 868800 615557 869900 nw
tri 503143 864815 507128 868800 ne
rect 507128 864815 510472 868800
tri 510472 864815 514457 868800 nw
tri 603143 864815 607128 868800 ne
rect 607128 864815 610472 868800
tri 610472 864815 614457 868800 nw
tri 693070 864815 698756 869900 se
rect 698756 865900 700756 873900
tri 700756 872840 701816 873900 nw
tri 707696 872840 708756 873900 ne
tri 700756 865900 701816 866960 sw
tri 707696 865900 708756 866960 se
rect 708756 865900 710756 873900
rect 698756 865314 710756 865900
rect 698756 864962 710404 865314
tri 710404 864962 710756 865314 nw
rect 698756 864815 710257 864962
tri 710257 864815 710404 864962 nw
tri 507128 863900 508043 864815 ne
rect 508043 863900 509557 864815
tri 509557 863900 510472 864815 nw
tri 607128 863900 608043 864815 ne
rect 608043 863900 609557 864815
tri 609557 863900 610472 864815 nw
tri 692047 863900 693070 864815 se
rect 693070 863900 709342 864815
tri 709342 863900 710257 864815 nw
tri 508043 863143 508800 863900 ne
tri 508800 863143 509557 863900 nw
tri 608043 863143 608800 863900 ne
tri 608800 863143 609557 863900 nw
tri 681069 854082 692047 863900 se
rect 692047 854082 693070 863900
tri 693070 854082 704048 863900 nw
tri 669068 843349 681069 854082 se
tri 681069 843349 693070 854082 nw
tri 454800 834143 462800 842143 nw
tri 658774 834143 669068 843349 se
rect 669068 834143 669273 843349
tri 441243 831900 443486 834143 se
rect 443486 831900 452557 834143
tri 452557 831900 454800 834143 nw
tri 657272 832800 658774 834143 se
rect 658774 832800 669273 834143
tri 669273 832800 681069 843349 nw
tri 466243 831900 467143 832800 se
rect 467143 831900 668267 832800
tri 668267 831900 669273 832800 nw
tri 432172 822829 441243 831900 se
rect 441243 822829 443486 831900
tri 443486 822829 452557 831900 nw
tri 465896 831553 466243 831900 se
rect 466243 831553 667879 831900
tri 667879 831553 668267 831900 nw
tri 699823 831553 700170 831900 se
rect 700170 831553 709342 831900
tri 709342 831553 709689 831900 sw
tri 459676 825333 465896 831553 se
rect 465896 825333 660924 831553
tri 660924 825333 667879 831553 nw
tri 698756 830486 699823 831553 se
rect 699823 830833 709689 831553
tri 709689 830833 710409 831553 sw
rect 699823 830486 710409 830833
tri 710409 830486 710756 830833 sw
rect 698756 829900 710756 830486
tri 457172 822829 459676 825333 se
rect 459676 824800 660328 825333
tri 660328 824800 660924 825333 nw
rect 459676 822829 468486 824800
tri 468486 822829 470457 824800 nw
tri 696420 822829 698756 825333 se
rect 698756 822829 700756 829900
tri 700756 828840 701816 829900 nw
tri 707696 828840 708756 829900 ne
tri 432143 822800 432172 822829 se
rect 432172 822800 443457 822829
tri 443457 822800 443486 822829 nw
tri 457143 822800 457172 822829 se
rect 457172 822800 468457 822829
tri 468457 822800 468486 822829 nw
tri 696393 822800 696420 822829 se
rect 696420 822800 700756 822829
tri 389243 819900 392143 822800 se
rect 392143 819900 440557 822800
tri 440557 819900 443457 822800 nw
tri 455829 821486 457143 822800 se
rect 457143 821486 467143 822800
tri 467143 821486 468457 822800 nw
tri 454243 819900 455829 821486 se
rect 455829 819900 465557 821486
tri 465557 819900 467143 821486 nw
tri 693687 819900 696393 822800 se
rect 696393 821900 700756 822800
tri 700756 821900 701816 822960 sw
tri 707696 821900 708756 822960 se
rect 708756 821900 710756 829900
rect 696393 821314 710756 821900
rect 696393 820967 710409 821314
tri 710409 820967 710756 821314 nw
rect 696393 819900 709342 820967
tri 709342 819900 710409 820967 nw
tri 22265 813486 28577 819900 ne
rect 28577 813486 33490 819900
tri 33490 813486 39801 819900 sw
tri 142043 813486 148457 819900 ne
rect 148457 816114 153357 819900
tri 153357 816114 157143 819900 sw
tri 252043 816114 255829 819900 ne
rect 255829 816114 263357 819900
rect 148457 813486 157143 816114
tri 157143 813486 159771 816114 sw
tri 255829 813486 258457 816114 ne
rect 258457 813486 263357 816114
tri 263357 813486 269771 819900 sw
tri 28577 812332 29713 813486 ne
rect 29713 812800 39801 813486
tri 39801 812800 40476 813486 sw
rect 29713 812332 125321 812800
tri 125321 812332 125847 812800 sw
tri 29713 804800 37124 812332 ne
rect 37124 804800 125847 812332
tri 125847 804800 134321 812332 sw
tri 148457 804800 157143 813486 ne
rect 157143 812800 159771 813486
tri 159771 812800 160457 813486 sw
tri 258457 812800 259143 813486 ne
rect 259143 812800 269771 813486
rect 157143 804800 230457 812800
tri 230457 804800 238457 812800 sw
tri 259143 804800 267143 812800 ne
rect 267143 804800 269771 812800
tri 122279 798900 128916 804800 ne
rect 128916 798900 134321 804800
tri 134321 798900 140958 804800 sw
tri 227143 798900 233043 804800 ne
rect 233043 798900 238457 804800
tri 7987 798553 8334 798900 se
rect 8334 798553 17506 798900
tri 17506 798553 17853 798900 sw
tri 128916 798553 129306 798900 ne
rect 129306 798553 140958 798900
tri 7267 797833 7987 798553 se
rect 7987 797833 17853 798553
tri 6920 797486 7267 797833 se
rect 7267 797486 17853 797833
tri 17853 797486 18920 798553 sw
rect 6920 796900 18920 797486
rect 6920 788900 8920 796900
tri 8920 795840 9980 796900 nw
tri 15860 795840 16920 796900 ne
rect 16920 792699 18920 796900
tri 129306 794096 134321 798553 ne
rect 134321 794096 140958 798553
tri 140958 794096 146363 798900 sw
tri 134321 793486 135007 794096 ne
rect 135007 793486 146363 794096
tri 146363 793486 147049 794096 sw
tri 233043 793486 238457 798900 ne
tri 238457 793486 249771 804800 sw
tri 267143 802172 269771 804800 ne
tri 269771 802172 281085 813486 sw
tri 344800 810457 354243 819900 se
rect 354243 817143 362800 819900
rect 354243 810457 356114 817143
tri 356114 810457 362800 817143 nw
tri 380829 811486 389243 819900 se
rect 389243 814800 435457 819900
tri 435457 814800 440557 819900 nw
tri 454170 819827 454243 819900 se
rect 454243 819827 465484 819900
tri 465484 819827 465557 819900 nw
tri 693619 819827 693687 819900 se
rect 693687 819827 704560 819900
tri 704560 819827 704628 819900 nw
tri 449143 814800 454170 819827 se
rect 454170 814800 460457 819827
tri 460457 814800 465484 819827 nw
tri 688928 814800 693619 819827 se
rect 693619 814800 698002 819827
rect 389243 811486 392143 814800
tri 392143 811486 395457 814800 nw
tri 447143 812800 449143 814800 se
rect 449143 812800 458457 814800
tri 458457 812800 460457 814800 nw
tri 687062 812800 688928 814800 se
rect 688928 812800 698002 814800
tri 698002 812800 704560 819827 nw
tri 445829 811486 447143 812800 se
rect 447143 811486 457143 812800
tri 457143 811486 458457 812800 nw
tri 475829 811486 477143 812800 se
rect 477143 811486 690538 812800
tri 379800 810457 380829 811486 se
tri 269771 793486 278457 802172 ne
rect 278457 793486 281085 802172
tri 135007 792779 135802 793486 ne
rect 135802 792779 147049 793486
tri 18920 792699 19006 792779 sw
tri 135802 792699 135892 792779 ne
rect 135892 792699 147049 792779
tri 8920 788900 9980 789960 sw
tri 15860 788900 16920 789960 se
rect 16920 788900 19006 792699
rect 6920 788314 19006 788900
tri 6920 787967 7267 788314 ne
rect 7267 787967 19006 788314
tri 7267 786900 8334 787967 ne
rect 8334 786900 19006 787967
tri 19006 786900 25233 792699 sw
tri 135892 786900 142416 792699 ne
rect 142416 786900 147049 792699
tri 147049 786900 154458 793486 sw
tri 238457 786900 245043 793486 ne
rect 245043 788457 249771 793486
tri 249771 788457 254800 793486 sw
tri 278457 790858 281085 793486 ne
tri 281085 790858 292399 802172 sw
tri 281085 788457 283486 790858 ne
rect 283486 788457 292399 790858
rect 245043 786900 254800 788457
tri 13494 782172 18572 786900 ne
rect 18572 782172 25233 786900
tri 25233 782172 30310 786900 sw
tri 142416 783392 146363 786900 ne
rect 146363 783392 154458 786900
tri 154458 783392 158405 786900 sw
tri 146363 782172 147735 783392 ne
rect 147735 782172 158405 783392
tri 158405 782172 159777 783392 sw
tri 245043 782172 249771 786900 ne
rect 249771 782172 254800 786900
tri 254800 782172 261085 788457 sw
tri 283486 782172 289771 788457 ne
rect 289771 782172 292399 788457
tri 18572 781768 19006 782172 ne
rect 19006 781768 30310 782172
tri 30310 781768 30744 782172 sw
tri 147735 781768 148190 782172 ne
rect 148190 781768 159777 782172
tri 19006 777143 23972 781768 ne
rect 23972 777143 30744 781768
tri 30744 777143 35710 781768 sw
tri 148190 777143 153393 781768 ne
rect 153393 777143 159777 781768
tri 159777 777143 165435 782172 sw
tri 249771 777143 254800 782172 ne
rect 254800 780457 261085 782172
tri 261085 780457 262800 782172 sw
tri 23972 770837 30744 777143 ne
rect 30744 772800 35710 777143
tri 35710 772800 40374 777143 sw
tri 153393 772800 158279 777143 ne
rect 158279 772800 165435 777143
tri 165435 772800 170321 777143 sw
rect 30744 770837 112800 772800
tri 158279 772688 158405 772800 ne
rect 158405 772688 212800 772800
tri 30744 764800 37226 770837 ne
rect 37226 764800 112800 770837
tri 158405 764800 167279 772688 ne
rect 167279 764800 212800 772688
tri 7975 755341 8334 755700 se
rect 8334 755341 17506 755700
tri 17506 755341 17865 755700 sw
tri 7279 754645 7975 755341 se
rect 7975 754645 17865 755341
tri 6920 754286 7279 754645 se
rect 7279 754286 17865 754645
tri 17865 754286 18920 755341 sw
rect 6920 753700 18920 754286
rect 6920 745700 8920 753700
tri 8920 752640 9980 753700 nw
tri 15860 752640 16920 753700 ne
rect 16920 749279 18920 753700
tri 18920 749279 19539 749812 sw
tri 8920 745700 9980 746760 sw
tri 15860 745700 16920 746760 se
rect 16920 745700 19539 749279
rect 6920 745114 19539 745700
tri 6920 744755 7279 745114 ne
rect 7279 744755 19539 745114
tri 7279 743700 8334 744755 ne
rect 8334 743700 19539 744755
tri 13757 738721 19539 743700 ne
tri 19539 738721 31799 749279 sw
tri 19539 728163 31799 738721 ne
tri 31799 728163 44058 738721 sw
tri 31799 717606 44058 728163 ne
tri 44058 722800 50285 728163 sw
rect 44058 717606 160457 722800
tri 160457 717606 165651 722800 sw
tri 44058 714800 47315 717606 ne
rect 47315 714800 165651 717606
tri 165651 714800 168457 717606 sw
tri 157143 712500 159443 714800 ne
rect 159443 712500 168457 714800
tri 7986 712152 8334 712500 se
rect 8334 712152 17506 712500
tri 17506 712152 17854 712500 sw
tri 159443 712152 159791 712500 ne
rect 159791 712152 168457 712500
tri 7268 711434 7986 712152 se
rect 7986 711434 17854 712152
tri 6920 711086 7268 711434 se
rect 7268 711086 17854 711434
tri 17854 711086 18920 712152 sw
rect 6920 710500 18920 711086
rect 6920 702500 8920 710500
tri 8920 709440 9980 710500 nw
tri 15860 709440 16920 710500 ne
rect 16920 706271 18920 710500
tri 159791 706408 165535 712152 ne
rect 165535 706408 168457 712152
tri 18920 706271 19069 706408 sw
tri 165535 706271 165672 706408 ne
rect 165672 706271 168457 706408
tri 8920 702500 9980 703560 sw
tri 15860 702500 16920 703560 se
rect 16920 702500 19069 706271
rect 6920 701914 19069 702500
tri 6920 701566 7268 701914 ne
rect 7268 701566 19069 701914
tri 7268 700500 8334 701566 ne
rect 8334 700500 19069 701566
tri 13525 695388 19069 700500 ne
tri 19069 695388 30870 706271 sw
tri 165672 703486 168457 706271 ne
tri 168457 703486 179771 714800 sw
tri 168457 695388 176555 703486 ne
rect 176555 695388 179771 703486
tri 19069 684505 30870 695388 ne
tri 30870 684505 42671 695388 sw
tri 176555 692172 179771 695388 ne
tri 179771 692172 191085 703486 sw
tri 179771 684505 187438 692172 ne
rect 187438 684505 191085 692172
tri 30870 673622 42671 684505 ne
tri 42671 675682 52237 684505 sw
tri 187438 680858 191085 684505 ne
tri 191085 680858 202399 692172 sw
tri 191085 675682 196261 680858 ne
rect 196261 675682 202399 680858
rect 42671 673622 52237 675682
tri 52237 673622 54471 675682 sw
tri 196261 673622 198321 675682 ne
rect 198321 674457 202399 675682
tri 202399 674457 208800 680858 sw
rect 198321 673622 208800 674457
tri 42671 669300 47357 673622 ne
rect 47357 672800 54471 673622
tri 54471 672800 55363 673622 sw
tri 198321 672800 199143 673622 ne
rect 199143 672800 208800 673622
rect 47357 669300 112800 672800
tri 199143 669544 202399 672800 ne
rect 202399 669544 208800 672800
tri 208800 669544 213713 674457 sw
rect 254800 672800 262800 780457
tri 289771 779544 292399 782172 ne
tri 292399 779544 303713 790858 sw
tri 292399 768230 303713 779544 ne
tri 303713 768800 314457 779544 sw
rect 303713 768230 313887 768800
tri 313887 768230 314457 768800 nw
tri 303713 763143 308800 768230 ne
tri 308800 763143 313887 768230 nw
tri 7990 668956 8334 669300 se
rect 8334 668956 17506 669300
tri 17506 668956 17850 669300 sw
tri 47357 668956 47730 669300 ne
rect 47730 668956 112800 669300
tri 7264 668230 7990 668956 se
rect 7990 668230 17850 668956
tri 6920 667886 7264 668230 se
rect 7264 668051 17850 668230
tri 17850 668051 18755 668956 sw
tri 47730 668051 48711 668956 ne
rect 48711 668051 112800 668956
rect 7264 667886 18755 668051
tri 18755 667886 18920 668051 sw
rect 6920 667300 18920 667886
rect 6920 659300 8920 667300
tri 8920 666240 9980 667300 nw
tri 15860 666240 16920 667300 ne
tri 8920 659300 9980 660360 sw
tri 15860 659300 16920 660360 se
rect 16920 659300 18920 667300
tri 48711 664800 52237 668051 ne
rect 52237 664800 112800 668051
tri 202399 664800 207143 669544 ne
rect 207143 668800 213713 669544
tri 213713 668800 214457 669544 sw
rect 207143 664800 208800 668800
tri 207143 663143 208800 664800 ne
tri 208800 663143 214457 668800 nw
rect 254800 664800 312800 672800
rect 6920 658714 18920 659300
tri 6920 658370 7264 658714 ne
rect 7264 658549 18920 658714
tri 18920 658549 23564 663053 sw
rect 7264 658370 23564 658549
tri 7264 657300 8334 658370 ne
rect 8334 657300 23564 658370
tri 13361 652069 18755 657300 ne
rect 18755 652069 23564 657300
tri 23564 652069 30246 658549 sw
tri 18755 640924 30246 652069 ne
tri 30246 640924 41736 652069 sw
tri 30246 629780 41736 640924 ne
tri 41736 629780 53225 640924 sw
tri 41736 626100 45529 629780 ne
rect 45529 626100 53225 629780
tri 53225 626100 57018 629780 sw
tri 7986 625752 8334 626100 se
rect 8334 625752 17506 626100
tri 17506 625752 17854 626100 sw
tri 45529 625752 45888 626100 ne
rect 45888 625752 57018 626100
tri 7268 625034 7986 625752 se
rect 7986 625034 17854 625752
tri 6920 624686 7268 625034 se
rect 7268 624686 17854 625034
tri 17854 624686 18920 625752 sw
rect 6920 624100 18920 624686
rect 6920 616100 8920 624100
tri 8920 623040 9980 624100 nw
tri 15860 623040 16920 624100 ne
rect 16920 619859 18920 624100
tri 45888 620023 51795 625752 ne
rect 51795 622800 57018 625752
tri 57018 622800 60421 626100 sw
rect 51795 620023 160457 622800
tri 18920 619859 19099 620023 sw
tri 51795 619859 51964 620023 ne
rect 51964 619859 160457 620023
tri 8920 616100 9980 617160 sw
tri 15860 616100 16920 617160 se
rect 16920 617143 19099 619859
tri 19099 617143 22057 619859 sw
tri 51964 618636 53225 619859 ne
rect 53225 618636 160457 619859
tri 160457 618636 164621 622800 sw
tri 53225 617143 54763 618636 ne
rect 54763 617143 164621 618636
tri 164621 617143 166114 618636 sw
rect 16920 616100 22057 617143
rect 6920 615514 22057 616100
tri 6920 615166 7268 615514 ne
rect 7268 615166 22057 615514
tri 7268 614100 8334 615166 ne
rect 8334 614100 22057 615166
tri 13541 608998 19099 614100 ne
rect 19099 608998 22057 614100
tri 22057 608998 30930 617143 sw
tri 54763 614800 57179 617143 ne
rect 57179 614800 166114 617143
tri 166114 614800 168457 617143 sw
tri 157143 608998 162945 614800 ne
rect 162945 608998 168457 614800
tri 19099 598137 30930 608998 ne
tri 30930 598137 42761 608998 sw
tri 162945 603486 168457 608998 ne
tri 168457 603486 179771 614800 sw
tri 168457 598137 173806 603486 ne
rect 173806 598137 179771 603486
tri 30930 587276 42761 598137 ne
tri 42761 587276 54591 598137 sw
tri 173806 592172 179771 598137 ne
tri 179771 592172 191085 603486 sw
tri 179771 587276 184667 592172 ne
rect 184667 587276 191085 592172
tri 42761 582900 47527 587276 ne
rect 47527 582900 54591 587276
tri 7977 582543 8334 582900 se
rect 8334 582543 17506 582900
tri 17506 582543 17863 582900 sw
tri 47527 582543 47916 582900 ne
rect 47916 582543 54591 582900
tri 7277 581843 7977 582543 se
rect 7977 581843 17863 582543
tri 6920 581486 7277 581843 se
rect 7277 581486 17863 581843
tri 17863 581486 18920 582543 sw
rect 6920 580900 18920 581486
rect 6920 572900 8920 580900
tri 8920 579840 9980 580900 nw
tri 15860 579840 16920 580900 ne
rect 16920 576498 18920 580900
tri 47916 576993 53961 582543 ne
rect 53961 576993 54591 582543
tri 18920 576498 19492 576993 sw
tri 53961 576498 54500 576993 ne
rect 54500 576498 54591 576993
tri 8920 572900 9980 573960 sw
tri 15860 572900 16920 573960 se
rect 16920 572900 19492 576498
rect 6920 572314 19492 572900
tri 6920 571957 7277 572314 ne
rect 7277 571957 19492 572314
tri 7277 570900 8334 571957 ne
rect 8334 570900 19492 571957
tri 13735 565910 19492 570900 ne
tri 19492 565910 31705 576498 sw
tri 54500 576415 54591 576498 ne
tri 54591 576415 66421 587276 sw
tri 184667 580858 191085 587276 ne
tri 191085 580858 202399 592172 sw
tri 191085 576415 195528 580858 ne
rect 195528 576415 202399 580858
tri 54591 565910 66033 576415 ne
rect 66033 572800 66421 576415
tri 66421 572800 70358 576415 sw
tri 195528 572800 199143 576415 ne
rect 199143 574457 202399 576415
tri 202399 574457 208800 580858 sw
rect 199143 572800 208800 574457
rect 66033 565910 112800 572800
tri 199143 569544 202399 572800 ne
rect 202399 569544 208800 572800
tri 208800 569544 213713 574457 sw
tri 19492 561300 24810 565910 ne
rect 24810 562800 31705 565910
tri 31705 562800 35292 565910 sw
tri 66033 565554 66421 565910 ne
rect 66421 565554 112800 565910
tri 66421 564800 67242 565554 ne
rect 67242 564800 112800 565554
tri 202399 564800 207143 569544 ne
rect 207143 568800 213713 569544
tri 213713 568800 214457 569544 sw
rect 207143 564800 208800 568800
tri 207143 563143 208800 564800 ne
tri 208800 563143 214457 568800 nw
rect 24810 561300 45457 562800
tri 45457 561300 46957 562800 sw
tri 24810 555323 31705 561300 ne
rect 31705 555323 46957 561300
tri 46957 555323 52934 561300 sw
tri 31705 554800 32308 555323 ne
rect 32308 554800 52934 555323
tri 52934 554800 53457 555323 sw
tri 42143 549300 47643 554800 ne
rect 47643 549300 53457 554800
tri 53457 549300 58957 554800 sw
tri 47643 543486 53457 549300 ne
rect 53457 543486 58957 549300
tri 58957 543486 64771 549300 sw
tri 53457 539700 57243 543486 ne
rect 57243 539700 64771 543486
tri 6920 538286 8334 539700 se
rect 8334 538286 17506 539700
tri 17506 538286 18920 539700 sw
rect 6920 537719 18920 538286
tri 57243 537805 59138 539700 ne
rect 59138 537805 64771 539700
tri 18920 537719 45451 537805 se
rect 6920 537700 45451 537719
rect 6920 529700 8920 537700
tri 8920 536640 9980 537700 nw
tri 15860 536640 16920 537700 ne
rect 16920 532172 45451 537700
tri 45451 532172 51085 537805 sw
tri 59138 532172 64771 537805 ne
tri 64771 532172 76085 543486 sw
tri 8920 529700 9980 530760 sw
tri 15860 529700 16920 530760 se
rect 16920 529795 51085 532172
tri 51085 529795 53462 532172 sw
tri 64771 529795 67148 532172 ne
rect 67148 529795 76085 532172
rect 16920 529700 18920 529795
tri 18920 529719 42149 529795 nw
tri 42149 529719 42225 529795 ne
rect 42225 529719 53462 529795
rect 6920 529114 18920 529700
tri 6920 527700 8334 529114 ne
rect 8334 527700 17506 529114
tri 17506 527700 18920 529114 nw
tri 42225 527700 44244 529719 ne
rect 44244 527700 53462 529719
tri 44244 518482 53462 527700 ne
tri 53462 520858 62399 529795 sw
tri 67148 520858 76085 529795 ne
tri 76085 522800 85457 532172 sw
rect 76085 520858 160457 522800
tri 160457 520858 162399 522800 sw
rect 53462 518482 62399 520858
tri 62399 518482 64775 520858 sw
tri 76085 518482 78461 520858 ne
rect 78461 518482 162399 520858
tri 53462 517300 54644 518482 ne
rect 54644 517300 64775 518482
tri 64775 517300 65957 518482 sw
tri 78461 517300 79643 518482 ne
rect 79643 517300 162399 518482
tri 162399 517300 165957 520858 sw
tri 54644 507169 64775 517300 ne
rect 64775 514800 65957 517300
tri 65957 514800 68457 517300 sw
tri 79643 514800 82143 517300 ne
rect 82143 514800 165957 517300
tri 165957 514800 168457 517300 sw
rect 64775 507169 68457 514800
tri 68457 507169 76088 514800 sw
tri 157143 507169 164774 514800 ne
rect 164774 507169 168457 514800
tri 64775 505300 66644 507169 ne
rect 66644 505300 76088 507169
tri 76088 505300 77957 507169 sw
tri 164774 505300 166643 507169 ne
rect 166643 505300 168457 507169
tri 168457 505300 177957 514800 sw
tri 66644 496500 75444 505300 ne
rect 75444 496500 77957 505300
tri 7991 496157 8334 496500 se
rect 8334 496157 17506 496500
tri 17506 496157 17849 496500 sw
tri 75444 496157 75787 496500 ne
rect 75787 496157 77957 496500
tri 7263 495429 7991 496157 se
rect 7991 495503 17849 496157
tri 17849 495503 18503 496157 sw
tri 75787 495856 76088 496157 ne
rect 76088 495856 77957 496157
tri 77957 495856 87401 505300 sw
tri 166643 503486 168457 505300 ne
rect 168457 503486 177957 505300
tri 177957 503486 179771 505300 sw
tri 168457 495856 176087 503486 ne
rect 176087 495856 179771 503486
tri 76088 495503 76441 495856 ne
rect 76441 495503 87401 495856
rect 7991 495429 18503 495503
tri 6920 495086 7263 495429 se
rect 7263 495086 18503 495429
tri 18503 495086 18920 495503 sw
rect 6920 494500 18920 495086
rect 6920 486500 8920 494500
tri 8920 493440 9980 494500 nw
tri 15860 493440 16920 494500 ne
tri 8920 486500 9980 487560 sw
tri 15860 486500 16920 487560 se
rect 16920 486500 18920 494500
tri 76441 490115 81829 495503 ne
rect 81829 490115 87401 495503
rect 6920 485914 18920 486500
tri 6920 485571 7263 485914 ne
rect 7263 485571 18920 485914
tri 7263 484500 8334 485571 ne
rect 8334 485497 18920 485571
tri 18920 485497 23477 490115 sw
tri 81829 485497 86447 490115 ne
rect 86447 485497 87401 490115
rect 8334 484500 23477 485497
tri 13220 479147 18503 484500 ne
rect 18503 479147 23477 484500
tri 23477 479147 29743 485497 sw
tri 86447 484543 87401 485497 ne
tri 87401 484543 98714 495856 sw
tri 176087 492172 179771 495856 ne
tri 179771 492172 191085 503486 sw
tri 179771 484543 187400 492172 ne
rect 187400 484543 191085 492172
tri 87401 479147 92797 484543 ne
rect 92797 479147 98714 484543
tri 18503 473300 24272 479147 ne
rect 24272 473300 29743 479147
tri 29743 473300 35512 479147 sw
tri 92797 473300 98644 479147 ne
rect 98644 474457 98714 479147
tri 98714 474457 108800 484543 sw
tri 187400 480858 191085 484543 ne
tri 191085 480858 202399 492172 sw
tri 191085 474457 197486 480858 ne
rect 197486 474457 202399 480858
tri 202399 474457 208800 480858 sw
rect 98644 473300 108800 474457
tri 108800 473300 109957 474457 sw
tri 197486 473300 198643 474457 ne
rect 198643 473300 208800 474457
tri 208800 473300 209957 474457 sw
tri 24272 467756 29743 473300 ne
rect 29743 467756 35512 473300
tri 35512 467756 40983 473300 sw
tri 98644 473230 98714 473300 ne
rect 98714 473230 109957 473300
tri 109957 473230 110027 473300 sw
tri 198643 473230 198713 473300 ne
rect 198713 473230 209957 473300
tri 98714 467756 104187 473230 ne
rect 104187 468800 110027 473230
tri 110027 468800 114457 473230 sw
tri 198713 469544 202399 473230 ne
rect 202399 469544 209957 473230
tri 209957 469544 213713 473300 sw
rect 104187 467756 108800 468800
tri 29743 461300 36113 467756 ne
rect 36113 461300 40983 467756
tri 40983 461300 47353 467756 sw
tri 104187 463143 108800 467756 ne
tri 108800 463143 114457 468800 nw
tri 202399 463143 208800 469544 ne
rect 208800 468800 213713 469544
tri 213713 468800 214457 469544 sw
tri 208800 463143 214457 468800 nw
tri 36113 456365 40983 461300 ne
rect 40983 456365 47353 461300
tri 47353 456365 52223 461300 sw
tri 40983 454300 43020 456365 ne
rect 43020 454300 52223 456365
tri 7990 453956 8334 454300 se
rect 8334 453956 17506 454300
tri 17506 453956 17850 454300 sw
tri 43020 453956 43360 454300 ne
rect 43360 453956 52223 454300
tri 7264 453230 7990 453956 se
rect 7990 453230 17850 453956
tri 6920 452886 7264 453230 se
rect 7264 453028 17850 453230
tri 17850 453028 18778 453956 sw
tri 43360 453028 44275 453956 ne
rect 44275 453028 52223 453956
rect 7264 452886 18778 453028
tri 18778 452886 18920 453028 sw
rect 6920 452300 18920 452886
rect 6920 444300 8920 452300
tri 8920 451240 9980 452300 nw
tri 15860 451240 16920 452300 ne
tri 8920 444300 9980 445360 sw
tri 15860 444300 16920 445360 se
rect 16920 444300 18920 452300
tri 44275 448065 49172 453028 ne
rect 49172 448065 52223 453028
rect 6920 443714 18920 444300
tri 6920 443370 7264 443714 ne
rect 7264 443572 18920 443714
tri 18920 443572 23570 448065 sw
tri 49172 444974 52223 448065 ne
tri 52223 444974 63462 456365 sw
rect 254800 452143 262800 664800
rect 344800 628457 352800 810457
tri 352800 807143 356114 810457 nw
tri 376486 807143 379800 810457 se
rect 379800 807143 380829 810457
tri 369515 800172 376486 807143 se
rect 376486 800172 380829 807143
tri 380829 800172 392143 811486 nw
tri 444515 810172 445829 811486 se
rect 445829 810172 455829 811486
tri 455829 810172 457143 811486 nw
tri 474515 810172 475829 811486 se
rect 475829 810172 690538 811486
tri 435829 801486 444515 810172 se
rect 444515 801486 447143 810172
tri 447143 801486 455829 810172 nw
tri 465829 801486 474515 810172 se
rect 474515 804800 690538 810172
tri 690538 804800 698002 812800 nw
rect 474515 801486 477143 804800
tri 477143 801486 480457 804800 nw
tri 434515 800172 435829 801486 se
rect 435829 800172 445829 801486
tri 445829 800172 447143 801486 nw
tri 464515 800172 465829 801486 se
rect 465829 800172 466114 801486
tri 364800 795457 369515 800172 se
rect 369515 795457 376114 800172
tri 376114 795457 380829 800172 nw
tri 433201 798858 434515 800172 se
rect 434515 798858 444515 800172
tri 444515 798858 445829 800172 nw
tri 429800 795457 433201 798858 se
rect 433201 795457 441114 798858
tri 441114 795457 444515 798858 nw
tri 459800 795457 464515 800172 se
rect 464515 795457 466114 800172
rect 364800 647352 372800 795457
tri 372800 792143 376114 795457 nw
tri 426486 792143 429800 795457 se
rect 429800 792143 437800 795457
tri 437800 792143 441114 795457 nw
tri 456486 792143 459800 795457 se
rect 459800 792143 466114 795457
tri 421887 787544 426486 792143 se
rect 426486 787544 433201 792143
tri 433201 787544 437800 792143 nw
tri 454800 790457 456486 792143 se
rect 456486 790457 466114 792143
tri 466114 790457 477143 801486 nw
tri 410573 776230 421887 787544 se
tri 421887 776230 433201 787544 nw
tri 403143 768800 410573 776230 se
rect 410573 768800 414457 776230
tri 414457 768800 421887 776230 nw
tri 403143 763143 408800 768800 ne
tri 408800 763143 414457 768800 nw
tri 403143 668800 408800 674457 se
tri 403143 667027 404916 668800 ne
rect 404916 667027 408800 668800
tri 408800 667027 416230 674457 sw
tri 404916 663143 408800 667027 ne
rect 408800 663143 416230 667027
tri 408800 655713 416230 663143 ne
tri 416230 655713 427544 667027 sw
tri 416230 650248 421695 655713 ne
rect 421695 651500 427544 655713
tri 427544 651500 431757 655713 sw
rect 421695 650248 431757 651500
tri 431757 650248 433009 651500 sw
tri 372800 647352 375214 650248 sw
tri 421695 647352 424591 650248 ne
rect 424591 647352 433009 650248
tri 433009 647352 435905 650248 sw
tri 364800 639500 371343 647352 ne
rect 371343 639501 375214 647352
tri 375214 639501 381757 647352 sw
tri 424591 644399 427544 647352 ne
rect 427544 644399 435905 647352
tri 435905 644399 438858 647352 sw
rect 371343 639500 381757 639501
tri 427544 639500 432443 644399 ne
rect 432443 640457 438858 644399
tri 438858 640457 442800 644399 sw
rect 432443 639771 442800 640457
tri 442800 639771 443486 640457 sw
tri 454114 639771 454800 640457 se
rect 454800 639771 462800 790457
tri 462800 787143 466114 790457 nw
tri 699822 786352 700170 786700 se
rect 700170 786352 709342 786700
tri 709342 786352 709690 786700 sw
tri 698756 785286 699822 786352 se
rect 699822 785634 709690 786352
tri 709690 785634 710408 786352 sw
rect 699822 785286 710408 785634
tri 710408 785286 710756 785634 sw
rect 698756 784700 710756 785286
tri 693795 774700 698756 780088 se
rect 698756 776700 700756 784700
tri 700756 783640 701816 784700 nw
tri 707696 783640 708756 784700 ne
tri 700756 776700 701816 777760 sw
tri 707696 776700 708756 777760 se
rect 708756 776700 710756 784700
rect 698756 776114 710756 776700
rect 698756 775766 710408 776114
tri 710408 775766 710756 776114 nw
rect 698756 774700 709342 775766
tri 709342 774700 710408 775766 nw
tri 693649 774541 693795 774700 se
rect 693795 774541 704523 774700
tri 704523 774541 704669 774700 nw
tri 693572 774457 693649 774541 se
rect 693649 774457 702920 774541
tri 503143 768800 508800 774457 se
tri 503143 768056 503887 768800 ne
rect 503887 768056 508800 768800
tri 508800 768056 515201 774457 sw
tri 692046 772800 693572 774457 se
rect 693572 772800 702920 774457
tri 702920 772800 704523 774541 nw
rect 604800 768056 698552 772800
tri 698552 768056 702920 772800 nw
tri 503887 763143 508800 768056 ne
rect 508800 763143 515201 768056
tri 508800 756742 515201 763143 ne
tri 515201 756742 526515 768056 sw
rect 604800 764800 695554 768056
tri 695554 764800 698552 768056 nw
tri 515201 745428 526515 756742 ne
tri 526515 745428 537829 756742 sw
tri 526515 734114 537829 745428 ne
tri 537829 741700 541557 745428 sw
rect 537829 741355 541557 741700
tri 541557 741355 541902 741700 sw
tri 699825 741355 700170 741700 se
rect 700170 741355 709342 741700
tri 709342 741355 709687 741700 sw
rect 537829 735172 541902 741355
tri 541902 735172 548085 741355 sw
tri 698756 740286 699825 741355 se
rect 699825 740631 709687 741355
tri 709687 740631 710411 741355 sw
rect 699825 740286 710411 740631
tri 710411 740286 710756 740631 sw
rect 698756 739700 710756 740286
rect 537829 734114 548085 735172
tri 548085 734114 549143 735172 sw
tri 537829 722800 549143 734114 ne
tri 549143 729700 553557 734114 sw
tri 693590 729700 698756 735172 se
rect 698756 731700 700756 739700
tri 700756 738640 701816 739700 nw
tri 707696 738640 708756 739700 ne
tri 700756 731700 701816 732760 sw
tri 707696 731700 708756 732760 se
rect 708756 731700 710756 739700
rect 698756 731114 710756 731700
rect 698756 730769 710411 731114
tri 710411 730769 710756 731114 nw
rect 698756 729700 709342 730769
tri 709342 729700 710411 730769 nw
rect 549143 722800 553557 729700
tri 553557 722800 560457 729700 sw
tri 687075 722800 693590 729700 se
rect 693590 722800 698078 729700
tri 698078 722800 704594 729700 nw
tri 549143 714800 557143 722800 ne
rect 557143 714800 690525 722800
tri 690525 714800 698078 722800 nw
tri 699825 696355 700170 696700 se
rect 700170 696355 709342 696700
tri 709342 696355 709687 696700 sw
tri 698756 695286 699825 696355 se
rect 699825 695631 709687 696355
tri 709687 695631 710411 696355 sw
rect 699825 695286 710411 695631
tri 710411 695286 710756 695631 sw
rect 698756 694700 710756 695286
tri 693559 684784 698756 690215 se
rect 698756 686700 700756 694700
tri 700756 693640 701816 694700 nw
tri 707696 693640 708756 694700 ne
tri 700756 686700 701816 687760 sw
tri 707696 686700 708756 687760 se
rect 708756 686700 710756 694700
rect 698756 686114 710756 686700
rect 698756 685769 710411 686114
tri 710411 685769 710756 686114 nw
rect 698756 684784 709426 685769
tri 709426 684784 710411 685769 nw
tri 693479 684700 693559 684784 se
rect 693559 684700 709342 684784
tri 709342 684700 709426 684784 nw
tri 683677 674457 693479 684700 se
rect 693479 674457 693559 684700
tri 503143 668800 508800 674457 se
tri 503143 668056 503887 668800 ne
rect 503887 668056 508800 668800
tri 508800 668056 515201 674457 sw
tri 682486 673212 683677 674457 se
rect 683677 673212 693559 674457
tri 693559 673212 704551 684700 nw
tri 682091 672800 682486 673212 se
rect 682486 672800 693165 673212
tri 693165 672800 693559 673212 nw
rect 604800 668056 688625 672800
tri 688625 668056 693165 672800 nw
tri 503887 663143 508800 668056 ne
rect 508800 663143 515201 668056
tri 508800 656742 515201 663143 ne
tri 515201 656742 526515 668056 sw
rect 604800 664800 685509 668056
tri 685509 664800 688625 668056 nw
tri 515201 645428 526515 656742 ne
tri 526515 651500 531757 656742 sw
rect 526515 651156 531757 651500
tri 531757 651156 532101 651500 sw
tri 699826 651156 700170 651500 se
rect 700170 651156 709342 651500
tri 709342 651156 709686 651500 sw
rect 526515 645428 532101 651156
tri 532101 645428 537829 651156 sw
tri 698756 650086 699826 651156 se
rect 699826 650430 709686 651156
tri 709686 650430 710412 651156 sw
rect 699826 650086 710412 650430
tri 710412 650086 710756 650430 sw
rect 698756 649500 710756 650086
rect 432443 639500 443486 639771
tri 443486 639500 443757 639771 sw
tri 453843 639500 454114 639771 se
rect 454114 639500 462800 639771
tri 371343 634855 375214 639500 ne
rect 375214 634855 381757 639500
tri 381757 634855 385629 639500 sw
tri 432443 634855 437088 639500 ne
rect 437088 634855 443757 639500
tri 443757 634855 448402 639500 sw
tri 449198 634855 453843 639500 se
rect 453843 637143 462800 639500
rect 453843 634855 454800 637143
tri 375214 630457 378879 634855 ne
rect 378879 630457 385629 634855
tri 352800 628457 354800 630457 sw
tri 378879 628457 380545 630457 ne
rect 380545 628457 385629 630457
rect 344800 627143 354800 628457
tri 354800 627143 356114 628457 sw
tri 380545 627143 381640 628457 ne
rect 381640 627143 385629 628457
tri 344800 626100 345843 627143 ne
rect 345843 626100 356114 627143
tri 345843 617143 354800 626100 ne
rect 354800 620457 356114 626100
tri 356114 620457 362800 627143 sw
tri 381640 622357 385629 627143 ne
tri 385629 622800 395674 634855 sw
tri 437088 633085 438858 634855 ne
rect 438858 634457 448402 634855
tri 448402 634457 448800 634855 sw
tri 448800 634457 449198 634855 se
rect 449198 634457 454800 634855
rect 438858 633085 454800 634457
tri 438858 629143 442800 633085 ne
rect 442800 629143 454800 633085
tri 454800 629143 462800 637143 nw
tri 526515 634114 537829 645428 ne
tri 537829 645066 538191 645428 sw
rect 537829 639679 538191 645066
tri 538191 639679 543578 645066 sw
tri 693519 639679 698756 645066 se
rect 698756 641500 700756 649500
tri 700756 648440 701816 649500 nw
tri 707696 648440 708756 649500 ne
tri 700756 641500 701816 642560 sw
tri 707696 641500 708756 642560 se
rect 708756 641500 710756 649500
rect 698756 640914 710756 641500
rect 698756 640570 710412 640914
tri 710412 640570 710756 640914 nw
rect 698756 639679 709521 640570
tri 709521 639679 710412 640570 nw
rect 537829 639500 543578 639679
tri 543578 639500 543757 639679 sw
tri 693345 639500 693519 639679 se
rect 693519 639500 709342 639679
tri 709342 639500 709521 639679 nw
rect 537829 634114 543757 639500
tri 543757 634114 549143 639500 sw
tri 537829 629143 542800 634114 ne
rect 542800 629143 549143 634114
tri 549143 629143 554114 634114 sw
tri 683277 629143 693345 639500 se
rect 693345 629143 693519 639500
tri 442800 628800 443143 629143 ne
rect 443143 628800 454457 629143
tri 454457 628800 454800 629143 nw
tri 443143 623143 448800 628800 ne
rect 448800 628457 454457 628800
tri 454457 628457 454800 628800 sw
tri 542800 628457 543486 629143 ne
rect 543486 628457 554114 629143
tri 554114 628457 554800 629143 sw
tri 682610 628457 683277 629143 se
rect 683277 628457 693519 629143
rect 448800 623143 454800 628457
tri 454800 623143 460114 628457 sw
tri 543486 623143 548800 628457 ne
rect 548800 628202 554800 628457
tri 554800 628202 555055 628457 sw
tri 682362 628202 682610 628457 se
rect 682610 628202 693519 628457
tri 693519 628202 704502 639500 nw
rect 548800 623143 555055 628202
tri 555055 623143 560114 628202 sw
tri 677443 623143 682362 628202 se
rect 682362 623143 688267 628202
tri 448800 622800 449143 623143 ne
rect 449143 622800 460114 623143
tri 460114 622800 460457 623143 sw
tri 548800 622800 549143 623143 ne
rect 549143 622800 560114 623143
tri 560114 622800 560457 623143 sw
tri 677110 622800 677443 623143 se
rect 677443 622800 688267 623143
tri 688267 622800 693519 628202 nw
rect 385629 622357 425457 622800
tri 425457 622357 425900 622800 sw
tri 449143 622357 449586 622800 ne
rect 449586 622357 460457 622800
tri 460457 622357 460900 622800 sw
tri 549143 622357 549586 622800 ne
rect 549586 622357 680490 622800
rect 354800 582800 362800 620457
tri 385629 614800 391926 622357 ne
rect 391926 614800 425900 622357
tri 425900 614800 433457 622357 sw
tri 449586 621771 450172 622357 ne
rect 450172 621771 460900 622357
tri 460900 621771 461486 622357 sw
tri 549586 621771 550172 622357 ne
rect 550172 621771 680490 622357
tri 450172 614800 457143 621771 ne
rect 457143 614800 461486 621771
tri 461486 614800 468457 621771 sw
tri 550172 614800 557143 621771 ne
rect 557143 614800 680490 621771
tri 680490 614800 688267 622800 nw
tri 422143 606500 430443 614800 ne
rect 430443 606500 433457 614800
tri 433457 606500 441757 614800 sw
tri 457143 610457 461486 614800 ne
rect 461486 610457 468457 614800
tri 468457 610457 472800 614800 sw
tri 461486 607143 464800 610457 ne
tri 430443 603486 433457 606500 ne
rect 433457 603486 441757 606500
tri 441757 603486 444771 606500 sw
tri 433457 594500 442443 603486 ne
rect 442443 595457 444771 603486
tri 444771 595457 452800 603486 sw
rect 442443 594500 452800 595457
tri 442443 592172 444771 594500 ne
rect 444771 592172 452800 594500
tri 444771 592143 444800 592172 ne
tri 347701 580858 349643 582800 se
rect 349643 580858 362800 582800
tri 341643 574800 347701 580858 se
rect 347701 574800 362800 580858
tri 341300 574457 341643 574800 se
rect 341643 574457 352614 574800
tri 352614 574457 352957 574800 nw
tri 339643 572800 341300 574457 se
rect 341300 572800 347701 574457
rect 304800 569544 347701 572800
tri 347701 569544 352614 574457 nw
rect 304800 564800 342957 569544
tri 342957 564800 347701 569544 nw
rect 354800 562800 362800 574800
tri 364643 562800 374643 572800 se
rect 374643 564800 412800 572800
rect 374643 562800 375957 564800
tri 375957 562800 377957 564800 nw
rect 354800 554800 367957 562800
tri 367957 554800 375957 562800 nw
rect 354800 482800 362800 554800
rect 444800 528457 452800 592172
rect 464800 547143 472800 610457
tri 699826 606156 700170 606500 se
rect 700170 606156 709342 606500
tri 709342 606156 709686 606500 sw
tri 698756 605086 699826 606156 se
rect 699826 605430 709686 606156
tri 709686 605430 710412 606156 sw
rect 699826 605086 710412 605430
tri 710412 605086 710756 605430 sw
rect 698756 604500 710756 605086
tri 693508 594706 698756 600080 se
rect 698756 596500 700756 604500
tri 700756 603440 701816 604500 nw
tri 707696 603440 708756 604500 ne
tri 700756 596500 701816 597560 sw
tri 707696 596500 708756 597560 se
rect 708756 596500 710756 604500
rect 698756 595914 710756 596500
rect 698756 595570 710412 595914
tri 710412 595570 710756 595914 nw
rect 698756 594706 709548 595570
tri 709548 594706 710412 595570 nw
tri 693307 594500 693508 594706 se
rect 693508 594500 709342 594706
tri 709342 594500 709548 594706 nw
tri 682327 583256 693307 594500 se
rect 693307 583256 693508 594500
tri 693508 583256 704488 594500 nw
tri 673733 574457 682327 583256 se
rect 682327 574457 683297 583256
tri 503143 568800 508800 574457 se
tri 503143 566742 505201 568800 ne
rect 505201 566742 508800 568800
tri 508800 566742 516515 574457 sw
tri 672115 572800 673733 574457 se
rect 673733 572800 683297 574457
tri 683297 572800 693508 583256 nw
rect 604800 566742 677381 572800
tri 677381 566742 683297 572800 nw
tri 505201 563143 508800 566742 ne
rect 508800 563143 516515 566742
tri 508800 555428 516515 563143 ne
tri 516515 561300 521957 566742 sw
rect 604800 564800 675485 566742
tri 675485 564800 677381 566742 nw
rect 516515 560957 521957 561300
tri 521957 560957 522300 561300 sw
tri 699827 560957 700170 561300 se
rect 700170 560957 709342 561300
tri 709342 560957 709685 561300 sw
rect 516515 555428 522300 560957
tri 522300 555428 527829 560957 sw
tri 698756 559886 699827 560957 se
rect 699827 560229 709685 560957
tri 709685 560229 710413 560957 sw
rect 699827 559886 710413 560229
tri 710413 559886 710756 560229 sw
rect 698756 559300 710756 559886
tri 464800 545428 466515 547143 ne
rect 466515 545428 472800 547143
tri 472800 545428 477829 550457 sw
tri 466515 539143 472800 545428 ne
rect 472800 544114 477829 545428
tri 477829 544114 479143 545428 sw
tri 516515 544114 527829 555428 ne
tri 527829 554891 528366 555428 sw
rect 527829 549523 528366 554891
tri 528366 549523 533734 554891 sw
tri 693499 549523 698756 554891 se
rect 698756 551300 700756 559300
tri 700756 558240 701816 559300 nw
tri 707696 558240 708756 559300 ne
tri 700756 551300 701816 552360 sw
tri 707696 551300 708756 552360 se
rect 708756 551300 710756 559300
rect 698756 550714 710756 551300
rect 698756 550371 710413 550714
tri 710413 550371 710756 550714 nw
rect 698756 549523 709565 550371
tri 709565 549523 710413 550371 nw
rect 527829 549300 533734 549523
tri 533734 549300 533957 549523 sw
tri 693281 549300 693499 549523 se
rect 693499 549300 709342 549523
tri 709342 549300 709565 549523 nw
rect 527829 544114 533957 549300
tri 533957 544114 539143 549300 sw
rect 472800 539143 479143 544114
tri 472800 534114 477829 539143 ne
rect 477829 534114 479143 539143
tri 479143 534114 489143 544114 sw
tri 477829 530457 481486 534114 ne
rect 481486 532800 489143 534114
tri 489143 532800 490457 534114 sw
tri 527829 532800 539143 544114 ne
tri 539143 538090 545167 544114 sw
tri 682301 538090 693281 549300 se
rect 693281 538090 693499 549300
tri 693499 538090 704479 549300 nw
rect 539143 532800 545167 538090
tri 545167 532800 550457 538090 sw
tri 677119 532800 682301 538090 se
rect 682301 532800 688317 538090
tri 688317 532800 693499 538090 nw
rect 481486 530457 490457 532800
tri 490457 530457 492800 532800 sw
tri 539143 530457 541486 532800 ne
rect 541486 530457 680481 532800
tri 452800 528457 454800 530457 sw
tri 481486 528457 483486 530457 ne
rect 483486 528457 492800 530457
tri 492800 528457 494800 530457 sw
tri 541486 528457 543486 530457 ne
rect 543486 528457 680481 530457
rect 444800 527143 454800 528457
tri 454800 527143 456114 528457 sw
tri 483486 527143 484800 528457 ne
rect 484800 527143 494800 528457
tri 494800 527143 496114 528457 sw
tri 543486 527143 544800 528457 ne
rect 544800 527143 680481 528457
tri 444800 517300 454643 527143 ne
rect 454643 520457 456114 527143
tri 456114 520457 462800 527143 sw
tri 484800 522800 489143 527143 ne
rect 489143 524800 496114 527143
tri 496114 524800 498457 527143 sw
tri 544800 524800 547143 527143 ne
rect 547143 524800 680481 527143
tri 680481 524800 688317 532800 nw
rect 489143 522800 498457 524800
tri 498457 522800 500457 524800 sw
rect 454643 517300 462800 520457
tri 454643 517143 454800 517300 ne
tri 347701 480858 349643 482800 se
rect 349643 480858 362800 482800
tri 341643 474800 347701 480858 se
rect 347701 474800 362800 480858
tri 341300 474457 341643 474800 se
rect 341643 474457 352614 474800
tri 352614 474457 352957 474800 nw
tri 340143 473300 341300 474457 se
rect 341300 473300 351457 474457
tri 351457 473300 352614 474457 nw
tri 339643 472800 340143 473300 se
rect 340143 472800 347701 473300
rect 304800 469544 347701 472800
tri 347701 469544 351457 473300 nw
rect 304800 464800 342957 469544
tri 342957 464800 347701 469544 nw
rect 354800 462800 362800 474800
rect 454800 482143 462800 517300
tri 489143 514800 497143 522800 ne
rect 497143 517300 535457 522800
tri 535457 517300 540957 522800 sw
rect 497143 516536 540957 517300
tri 540957 516536 541721 517300 sw
tri 699406 516536 700170 517300 se
rect 700170 516536 709342 517300
tri 709342 516536 710106 517300 sw
rect 497143 514800 541721 516536
tri 532143 512800 534143 514800 ne
rect 534143 513119 541721 514800
tri 541721 513119 545138 516536 sw
tri 698756 515886 699406 516536 se
rect 699406 515886 710106 516536
tri 710106 515886 710756 516536 sw
rect 698756 515300 710756 515886
rect 698756 513119 700756 515300
tri 700756 514240 701816 515300 nw
tri 707696 514240 708756 515300 ne
rect 534143 512800 545138 513119
tri 545138 512800 545457 513119 sw
tri 697995 512800 698755 513119 se
rect 698755 512800 700756 513119
tri 534143 511486 535457 512800 ne
rect 535457 511486 700756 512800
tri 535457 505300 541643 511486 ne
rect 541643 507300 700756 511486
tri 700756 507300 701816 508360 sw
tri 707696 507300 708756 508360 se
rect 708756 507300 710756 515300
rect 541643 506714 710756 507300
rect 541643 505950 709992 506714
tri 709992 505950 710756 506714 nw
rect 541643 505300 709342 505950
tri 709342 505300 709992 505950 nw
tri 541643 504800 542143 505300 ne
rect 542143 504800 699605 505300
tri 699605 504800 700796 505300 nw
tri 462800 482143 466114 485457 sw
tri 454800 474457 462486 482143 ne
rect 462486 474457 466114 482143
tri 466114 474457 473800 482143 sw
tri 462486 472800 464143 474457 ne
rect 464143 472800 473800 474457
tri 473800 472800 475457 474457 sw
tri 507143 472800 508800 474457 se
tri 508800 473300 509957 474457 sw
rect 508800 472800 509957 473300
tri 509957 472800 510457 473300 sw
tri 699670 472800 700170 473300 se
rect 700170 472800 709342 473300
tri 709342 472800 709842 473300 sw
tri 371387 469544 374643 472800 se
rect 374643 469544 412800 472800
tri 464143 470829 466114 472800 ne
rect 466114 470829 512800 472800
tri 366643 464800 371387 469544 se
rect 371387 464800 412800 469544
tri 466114 468056 468887 470829 ne
rect 468887 468056 512800 470829
rect 604800 472363 709842 472800
tri 709842 472363 710279 472800 sw
rect 604800 471886 710279 472363
tri 710279 471886 710756 472363 sw
rect 604800 471300 710756 471886
tri 512800 468056 515201 470457 sw
tri 468887 464800 472143 468056 ne
rect 472143 464800 515201 468056
tri 515201 464800 518457 468056 sw
rect 604800 464800 700756 471300
tri 700756 470240 701816 471300 nw
tri 707696 470240 708756 471300 ne
tri 364986 463143 366643 464800 se
rect 366643 463143 375957 464800
tri 364643 462800 364986 463143 se
rect 364986 462800 375957 463143
tri 375957 462800 377957 464800 nw
tri 507143 463143 508800 464800 ne
rect 508800 463143 518457 464800
tri 508800 462800 509143 463143 ne
rect 509143 462800 518457 463143
tri 518457 462800 520457 464800 sw
rect 698756 463300 700756 464800
tri 700756 463300 701816 464360 sw
tri 707696 463300 708756 464360 se
rect 708756 463300 710756 471300
rect 354800 461300 374457 462800
tri 374457 461300 375957 462800 nw
tri 509143 461300 510643 462800 ne
rect 510643 461300 520457 462800
tri 520457 461300 521957 462800 sw
rect 698756 462714 710756 463300
tri 698756 461300 700170 462714 ne
rect 700170 462237 710279 462714
tri 710279 462237 710756 462714 nw
rect 700170 461777 709819 462237
tri 709819 461777 710279 462237 nw
rect 700170 461300 709342 461777
tri 709342 461300 709819 461777 nw
rect 354800 456365 369522 461300
tri 369522 456365 374457 461300 nw
tri 510643 456742 515201 461300 ne
rect 515201 456742 521957 461300
tri 521957 456742 526515 461300 sw
tri 515201 456365 515578 456742 ne
rect 515578 456365 526515 456742
tri 526515 456365 526892 456742 sw
tri 254800 445428 261515 452143 ne
rect 261515 445428 262800 452143
tri 262800 445428 272829 455457 sw
rect 354800 454800 367957 456365
tri 367957 454800 369522 456365 nw
tri 515578 454800 517143 456365 ne
rect 517143 454800 526892 456365
tri 526892 454800 528457 456365 sw
tri 261515 444974 261969 445428 ne
rect 261969 444974 272829 445428
tri 272829 444974 273283 445428 sw
tri 52223 443572 53606 444974 ne
rect 53606 443572 63462 444974
rect 7264 443370 23570 443572
tri 7264 442300 8334 443370 ne
rect 8334 442300 23570 443370
tri 13373 437078 18778 442300 ne
rect 18778 437078 23570 442300
tri 23570 437078 30292 443572 sw
tri 53606 437078 60013 443572 ne
rect 60013 437078 63462 443572
tri 18778 429100 27034 437078 ne
rect 27034 429100 30292 437078
tri 30292 429100 38548 437078 sw
tri 60013 433583 63462 437078 ne
tri 63462 436191 72127 444974 sw
tri 261969 444143 262800 444974 ne
rect 262800 444143 273283 444974
tri 262800 436191 270752 444143 ne
rect 270752 436191 273283 444143
tri 273283 436191 282066 444974 sw
rect 63462 433583 72127 436191
tri 72127 433583 74700 436191 sw
tri 270752 434114 272829 436191 ne
rect 272829 434114 282066 436191
tri 282066 434114 284143 436191 sw
tri 272829 433583 273360 434114 ne
rect 273360 433583 284143 434114
tri 284143 433583 284674 434114 sw
tri 63462 429100 67884 433583 ne
rect 67884 432800 74700 433583
tri 74700 432800 75473 433583 sw
tri 273360 432800 274143 433583 ne
rect 274143 432800 284674 433583
tri 284674 432800 285457 433583 sw
rect 67884 429100 175457 432800
tri 175457 429100 179157 432800 sw
tri 274143 429100 277843 432800 ne
rect 277843 429100 285457 432800
tri 285457 429100 289157 432800 sw
tri 27034 425953 30292 429100 ne
rect 30292 425953 38548 429100
tri 38548 425953 41806 429100 sw
tri 67884 425953 70989 429100 ne
rect 70989 426114 179157 429100
tri 179157 426114 182143 429100 sw
tri 277843 426114 280829 429100 ne
rect 280829 426114 289157 429100
tri 289157 426114 292143 429100 sw
rect 70989 425953 182143 426114
tri 30292 417100 39454 425953 ne
rect 39454 417100 41806 425953
tri 41806 417100 50967 425953 sw
tri 70989 424800 72127 425953 ne
rect 72127 424800 182143 425953
tri 182143 424800 183457 426114 sw
tri 280829 424800 282143 426114 ne
rect 282143 424800 292143 426114
tri 292143 424800 293457 426114 sw
tri 172143 417100 179843 424800 ne
rect 179843 422800 183457 424800
tri 183457 422800 185457 424800 sw
tri 282143 422800 284143 424800 ne
rect 284143 422800 293457 424800
tri 293457 422800 295457 424800 sw
rect 179843 417100 260457 422800
tri 260457 417100 266157 422800 sw
tri 284143 417100 289843 422800 ne
rect 289843 417100 320457 422800
tri 320457 417100 326157 422800 sw
rect 354800 418457 362800 454800
tri 517143 445428 526515 454800 ne
rect 526515 445428 528457 454800
tri 528457 445428 537829 454800 sw
tri 526515 434114 537829 445428 ne
tri 537829 434114 549143 445428 sw
tri 537829 422800 549143 434114 ne
tri 549143 429100 554157 434114 sw
rect 549143 428685 554157 429100
tri 554157 428685 554572 429100 sw
tri 699755 428685 700170 429100 se
rect 700170 428685 709342 429100
tri 709342 428685 709757 429100 sw
rect 549143 423702 554572 428685
tri 554572 423702 559555 428685 sw
tri 698756 427686 699755 428685 se
rect 699755 428101 709757 428685
tri 709757 428101 710341 428685 sw
rect 699755 427686 710341 428101
tri 710341 427686 710756 428101 sw
rect 698756 427100 710756 427686
rect 549143 422800 559555 423702
tri 559555 422800 560457 423702 sw
tri 697507 422800 698756 423702 se
rect 698756 422800 700756 427100
tri 700756 426040 701816 427100 nw
tri 707696 426040 708756 427100 ne
tri 549143 420457 551486 422800 ne
rect 551486 420457 700756 422800
tri 362800 418457 364800 420457 sw
tri 551486 418457 553486 420457 ne
rect 553486 419100 700756 420457
tri 700756 419100 701816 420160 sw
tri 707696 419100 708756 420160 se
rect 708756 419100 710756 427100
rect 553486 418514 710756 419100
rect 553486 418457 710341 418514
rect 354800 417143 364800 418457
tri 364800 417143 366114 418457 sw
tri 553486 417143 554800 418457 ne
rect 554800 418099 710341 418457
tri 710341 418099 710756 418514 nw
rect 554800 417143 709342 418099
tri 354800 417100 354843 417143 ne
rect 354843 417100 366114 417143
tri 366114 417100 366157 417143 sw
tri 554800 417100 554843 417143 ne
rect 554843 417100 709342 417143
tri 709342 417100 710341 418099 nw
tri 39454 414828 41806 417100 ne
rect 41806 415925 50967 417100
tri 50967 415925 52183 417100 sw
tri 179843 415925 181018 417100 ne
rect 181018 415925 266157 417100
rect 41806 414828 52183 415925
tri 52183 414828 53318 415925 sw
tri 181018 414828 182115 415925 ne
rect 182115 414828 266157 415925
tri 41806 412100 44628 414828 ne
rect 44628 412800 53318 414828
tri 53318 412800 55417 414828 sw
tri 182115 414800 182143 414828 ne
rect 182143 414800 266157 414828
tri 266157 414800 268457 417100 sw
tri 289843 414800 292143 417100 ne
rect 292143 414800 326157 417100
tri 326157 414800 328457 417100 sw
tri 354843 414800 357143 417100 ne
rect 357143 414800 366157 417100
tri 257143 412800 259143 414800 ne
rect 259143 412800 268457 414800
rect 44628 412100 170457 412800
tri 7990 411756 8334 412100 se
rect 8334 411756 17506 412100
tri 17506 411756 17850 412100 sw
tri 44628 411756 44984 412100 ne
rect 44984 411756 170457 412100
tri 7264 411030 7990 411756 se
rect 7990 411241 17850 411756
tri 17850 411241 18365 411756 sw
tri 44984 411241 45517 411756 ne
rect 45517 411241 170457 411756
rect 7990 411030 18365 411241
tri 6920 410686 7264 411030 se
rect 7264 410686 18365 411030
tri 18365 410686 18920 411241 sw
rect 6920 410100 18920 410686
rect 6920 402100 8920 410100
tri 8920 409040 9980 410100 nw
tri 15860 409040 16920 410100 ne
tri 8920 402100 9980 403160 sw
tri 15860 402100 16920 403160 se
rect 16920 402100 18920 410100
tri 45517 405633 51321 411241 ne
rect 51321 405633 170457 411241
rect 6920 401514 18920 402100
tri 6920 401170 7264 401514 ne
rect 7264 401170 18920 401514
tri 7264 400100 8334 401170 ne
rect 8334 400959 18920 401170
tri 18920 400959 23416 405633 sw
tri 51321 404800 52183 405633 ne
rect 52183 404800 170457 405633
tri 170457 404800 178457 412800 sw
tri 259143 404800 267143 412800 ne
rect 267143 404800 268457 412800
tri 167143 400959 170984 404800 ne
rect 170984 400959 178457 404800
rect 8334 400100 23416 400959
tri 13141 394670 18365 400100 ne
rect 18365 394670 23416 400100
tri 23416 394670 29466 400959 sw
tri 170984 394670 177273 400959 ne
rect 177273 394670 178457 400959
tri 18365 384100 28532 394670 ne
rect 28532 384100 29466 394670
tri 29466 384100 39633 394670 sw
tri 177273 393486 178457 394670 ne
tri 178457 393486 189771 404800 sw
tri 267143 403486 268457 404800 ne
tri 268457 403486 279771 414800 sw
tri 317143 413085 318858 414800 ne
rect 318858 413085 328457 414800
tri 328457 413085 330172 414800 sw
tri 318858 411486 320457 413085 ne
rect 320457 411486 330172 413085
tri 320457 403486 328457 411486 ne
rect 328457 407143 330172 411486
tri 330172 407143 336114 413085 sw
tri 357143 407143 364800 414800 ne
rect 364800 410457 366157 414800
tri 366157 410457 372800 417100 sw
tri 554843 414800 557143 417100 ne
rect 557143 414800 700093 417100
tri 700093 414800 703279 417100 nw
rect 328457 403486 336114 407143
tri 336114 403486 339771 407143 sw
tri 268457 393486 278457 403486 ne
rect 278457 393486 279771 403486
tri 178457 384100 187843 393486 ne
rect 187843 384100 189771 393486
tri 189771 384100 199157 393486 sw
tri 278457 392172 279771 393486 ne
tri 279771 392172 291085 403486 sw
tri 328457 401771 330172 403486 ne
rect 330172 401771 339771 403486
tri 339771 401771 341486 403486 sw
tri 330172 392172 339771 401771 ne
rect 339771 392172 341486 401771
tri 341486 392172 351085 401771 sw
tri 279771 384100 287843 392172 ne
rect 287843 384100 291085 392172
tri 291085 384100 299157 392172 sw
tri 339771 390457 341486 392172 ne
rect 341486 390457 351085 392172
tri 351085 390457 352800 392172 sw
tri 341486 387143 344800 390457 ne
tri 28532 383130 29466 384100 ne
rect 29466 383130 39633 384100
tri 39633 383130 40567 384100 sw
tri 187843 383130 188813 384100 ne
rect 188813 383130 199157 384100
tri 29466 372100 40075 383130 ne
rect 40075 372800 40567 383130
tri 40567 372800 50503 383130 sw
tri 188813 382172 189771 383130 ne
rect 189771 382172 199157 383130
tri 199157 382172 201085 384100 sw
tri 287843 382172 289771 384100 ne
rect 289771 382172 299157 384100
tri 189771 372800 199143 382172 ne
rect 199143 374457 201085 382172
tri 201085 374457 208800 382172 sw
tri 289771 380858 291085 382172 ne
rect 291085 380858 299157 382172
tri 299157 380858 302399 384100 sw
tri 291085 374457 297486 380858 ne
rect 297486 374457 302399 380858
tri 302399 374457 308800 380858 sw
rect 199143 372800 208800 374457
rect 40075 372100 112800 372800
tri 199143 372100 199843 372800 ne
rect 199843 372100 208800 372800
tri 208800 372100 211157 374457 sw
tri 297486 372100 299843 374457 ne
rect 299843 372100 308800 374457
tri 308800 372100 311157 374457 sw
tri 40075 371589 40567 372100 ne
rect 40567 371589 112800 372100
tri 40567 368900 43153 371589 ne
rect 43153 368900 112800 371589
tri 199843 370858 201085 372100 ne
rect 201085 370858 211157 372100
tri 211157 370858 212399 372100 sw
tri 299843 370858 301085 372100 ne
rect 301085 370858 311157 372100
tri 7984 368550 8334 368900 se
rect 8334 368550 17506 368900
tri 17506 368550 17856 368900 sw
tri 43153 368550 43490 368900 ne
rect 43490 368550 112800 368900
tri 7270 367836 7984 368550 se
rect 7984 368343 17856 368550
tri 17856 368343 18063 368550 sw
tri 43490 368343 43689 368550 ne
rect 43689 368343 112800 368550
rect 7984 367836 18063 368343
tri 6920 367486 7270 367836 se
rect 7270 367486 18063 367836
tri 18063 367486 18920 368343 sw
rect 6920 366900 18920 367486
rect 6920 358900 8920 366900
tri 8920 365840 9980 366900 nw
tri 15860 365840 16920 366900 ne
tri 8920 358900 9980 359960 sw
tri 15860 358900 16920 359960 se
rect 16920 358900 18920 366900
tri 43689 364800 47097 368343 ne
rect 47097 364800 112800 368343
tri 201085 364800 207143 370858 ne
rect 207143 368800 212399 370858
tri 212399 368800 214457 370858 sw
tri 301085 369544 302399 370858 ne
rect 302399 369544 311157 370858
tri 311157 369544 313713 372100 sw
rect 207143 364800 208800 368800
tri 207143 363143 208800 364800 ne
tri 208800 363143 214457 368800 nw
tri 302399 363143 308800 369544 ne
rect 308800 368800 313713 369544
tri 313713 368800 314457 369544 sw
tri 308800 363143 314457 368800 nw
rect 6920 358314 18920 358900
tri 6920 357964 7270 358314 ne
rect 7270 357964 18920 358314
tri 7270 356900 8334 357964 ne
rect 8334 357457 18920 357964
tri 18920 357457 23245 362233 sw
rect 8334 356900 23245 357457
tri 12957 351262 18063 356900 ne
rect 18063 351262 23245 356900
tri 23245 351262 28856 357457 sw
tri 18063 339344 28856 351262 ne
tri 28856 339344 39649 351262 sw
tri 28856 338900 29258 339344 ne
rect 29258 338900 39649 339344
tri 39649 338900 40051 339344 sw
tri 29258 327425 39649 338900 ne
rect 39649 332800 40051 338900
tri 40051 332800 45574 338900 sw
rect 39649 327425 250457 332800
tri 250457 327425 255832 332800 sw
tri 39649 326900 40124 327425 ne
rect 40124 326900 255832 327425
tri 255832 326900 256357 327425 sw
tri 40124 325700 41211 326900 ne
rect 41211 325700 256357 326900
tri 7991 325357 8334 325700 se
rect 8334 325357 17506 325700
tri 17506 325357 17849 325700 sw
tri 41211 325357 41521 325700 ne
rect 41521 325357 256357 325700
tri 7263 324629 7991 325357 se
rect 7991 324639 17849 325357
tri 17849 324639 18567 325357 sw
tri 41521 324800 42026 325357 ne
rect 42026 324800 256357 325357
tri 256357 324800 258457 326900 sw
tri 247143 324639 247304 324800 ne
rect 247304 324639 258457 324800
rect 7991 324629 18567 324639
tri 6920 324286 7263 324629 se
rect 7263 324286 18567 324629
tri 18567 324286 18920 324639 sw
rect 6920 323700 18920 324286
rect 6920 315700 8920 323700
tri 8920 322640 9980 323700 nw
tri 15860 322640 16920 323700 ne
tri 8920 315700 9980 316760 sw
tri 15860 315700 16920 316760 se
rect 16920 315700 18920 323700
tri 247304 319351 252592 324639 ne
rect 252592 319351 258457 324639
rect 6920 315114 18920 315700
tri 6920 314771 7263 315114 ne
rect 7263 314771 18920 315114
tri 7263 313700 8334 314771 ne
rect 8334 314761 18920 314771
tri 18920 314761 23501 319351 sw
tri 252592 314761 257182 319351 ne
rect 257182 314761 258457 319351
rect 8334 313700 23501 314761
tri 13257 308381 18567 313700 ne
rect 18567 312800 23501 313700
tri 23501 312800 25459 314761 sw
tri 257182 313486 258457 314761 ne
tri 258457 313486 269771 324800 sw
tri 258457 312800 259143 313486 ne
rect 259143 312800 269771 313486
rect 18567 308381 170457 312800
tri 170457 308381 174876 312800 sw
tri 259143 308381 263562 312800 ne
rect 263562 308381 269771 312800
tri 18567 304800 22141 308381 ne
rect 22141 304800 174876 308381
tri 174876 304800 178457 308381 sw
tri 263562 304800 267143 308381 ne
rect 267143 304800 269771 308381
tri 167143 293900 178043 304800 ne
rect 178043 293900 178457 304800
tri 178457 293900 189357 304800 sw
tri 267143 302172 269771 304800 ne
tri 269771 302172 281085 313486 sw
tri 269771 293900 278043 302172 ne
rect 278043 293900 281085 302172
tri 281085 293900 289357 302172 sw
tri 178043 293486 178457 293900 ne
rect 178457 293486 189357 293900
tri 189357 293486 189771 293900 sw
tri 278043 293486 278457 293900 ne
rect 278457 293486 289357 293900
tri 178457 282500 189443 293486 ne
rect 189443 282500 189771 293486
tri 7910 282076 8334 282500 se
rect 8334 282076 17506 282500
tri 17506 282076 17930 282500 sw
tri 189443 282172 189771 282500 ne
tri 189771 282172 201085 293486 sw
tri 278457 290858 281085 293486 ne
rect 281085 290858 289357 293486
tri 289357 290858 292399 293900 sw
tri 281085 282172 289771 290858 ne
rect 289771 282172 292399 290858
tri 189771 282076 189867 282172 ne
rect 189867 282076 201085 282172
tri 7344 281510 7910 282076 se
rect 7910 281510 17930 282076
tri 6920 281086 7344 281510 se
rect 7344 281086 17930 281510
tri 17930 281086 18920 282076 sw
tri 189867 281900 190043 282076 ne
rect 190043 281900 201085 282076
tri 201085 281900 201357 282172 sw
tri 289771 281900 290043 282172 ne
rect 290043 281900 292399 282172
tri 292399 281900 301357 290858 sw
rect 6920 280500 18920 281086
rect 6920 272500 8920 280500
tri 8920 279440 9980 280500 nw
tri 15860 279440 16920 280500 ne
rect 16920 275546 18920 280500
tri 190043 277154 194789 281900 ne
rect 194789 277154 201357 281900
tri 18920 275546 21193 277154 sw
tri 194789 275546 196397 277154 ne
rect 196397 275546 201357 277154
tri 8920 272500 9980 273560 sw
tri 15860 272500 16920 273560 se
rect 16920 272800 21193 275546
tri 21193 272800 25072 275546 sw
tri 196397 272800 199143 275546 ne
rect 199143 274457 201357 275546
tri 201357 274457 208800 281900 sw
tri 290043 279544 292399 281900 ne
rect 292399 279544 301357 281900
tri 301357 279544 303713 281900 sw
tri 292399 274457 297486 279544 ne
rect 297486 274457 303713 279544
rect 199143 272800 208800 274457
rect 16920 272500 112800 272800
rect 6920 271914 112800 272500
tri 6920 271490 7344 271914 ne
rect 7344 271490 112800 271914
tri 7344 270500 8334 271490 ne
rect 8334 270500 112800 271490
tri 199143 270858 201085 272800 ne
rect 201085 270858 208800 272800
tri 208800 270858 212399 274457 sw
tri 297486 270858 301085 274457 ne
rect 301085 270858 303713 274457
tri 14474 265745 21193 270500 ne
rect 21193 265745 112800 270500
tri 21193 264800 22528 265745 ne
rect 22528 264800 112800 265745
tri 201085 264800 207143 270858 ne
rect 207143 268800 212399 270858
tri 212399 268800 214457 270858 sw
rect 207143 264800 208800 268800
tri 207143 263143 208800 264800 ne
tri 208800 263143 214457 268800 nw
tri 301085 268230 303713 270858 ne
tri 303713 268800 314457 279544 sw
rect 303713 268230 313887 268800
tri 313887 268230 314457 268800 nw
tri 303713 263143 308800 268230 ne
tri 308800 263143 313887 268230 nw
tri 341486 252143 344800 255457 se
rect 344800 252143 352800 390457
tri 336771 247428 341486 252143 se
rect 341486 247428 348085 252143
tri 348085 247428 352800 252143 nw
rect 364800 322800 372800 410457
tri 699808 383738 700170 384100 se
rect 700170 383738 709342 384100
tri 709342 383738 709704 384100 sw
tri 698756 382686 699808 383738 se
rect 699808 383048 709704 383738
tri 709704 383048 710394 383738 sw
rect 699808 382686 710394 383048
tri 710394 382686 710756 383048 sw
rect 698756 382100 710756 382686
tri 694284 374457 698756 378253 se
rect 698756 374457 700756 382100
tri 700756 381040 701816 382100 nw
tri 707696 381040 708756 382100 ne
tri 406443 372100 408800 374457 se
tri 408800 372100 411157 374457 sw
tri 506443 372100 508800 374457 se
tri 508800 372100 511157 374457 sw
tri 692855 373244 694284 374457 se
rect 694284 374100 700756 374457
tri 700756 374100 701816 375160 sw
tri 707696 374100 708756 375160 se
rect 708756 374100 710756 382100
rect 694284 373514 710756 374100
rect 694284 373244 710486 373514
tri 710486 373244 710756 373514 nw
tri 692331 372800 692855 373244 se
rect 692855 372800 709342 373244
rect 604800 372100 709342 372800
tri 709342 372100 710486 373244 nw
tri 403887 369544 406443 372100 se
rect 406443 369544 411157 372100
tri 411157 369544 413713 372100 sw
tri 503887 369544 506443 372100 se
rect 506443 369544 511157 372100
tri 511157 369544 513713 372100 sw
rect 604800 369544 700858 372100
tri 700858 369544 703869 372100 nw
tri 403143 368800 403887 369544 se
rect 403887 368800 413713 369544
tri 403143 367027 404916 368800 ne
rect 404916 367027 413713 368800
tri 413713 367027 416230 369544 sw
tri 503143 368800 503887 369544 se
tri 503143 368056 503887 368800 ne
rect 503887 368056 513713 369544
tri 513713 368056 515201 369544 sw
rect 604800 368056 699105 369544
tri 699105 368056 700858 369544 nw
tri 503887 367027 504916 368056 ne
rect 504916 367027 515201 368056
tri 515201 367027 516230 368056 sw
rect 604800 367027 697893 368056
tri 697893 367027 699105 368056 nw
tri 404916 363143 408800 367027 ne
rect 408800 363143 416230 367027
tri 416230 363143 420114 367027 sw
tri 504916 363143 508800 367027 ne
rect 508800 363143 516230 367027
tri 516230 363143 520114 367027 sw
rect 604800 364800 695269 367027
tri 695269 364800 697893 367027 nw
tri 408800 362233 409710 363143 ne
rect 409710 362233 420114 363143
tri 420114 362233 421024 363143 sw
tri 508800 362233 509710 363143 ne
rect 509710 362233 520114 363143
tri 520114 362233 521024 363143 sw
tri 409710 357457 414486 362233 ne
rect 414486 357457 421024 362233
tri 421024 357457 425800 362233 sw
tri 509710 357457 514486 362233 ne
rect 514486 357457 521024 362233
tri 521024 357457 525800 362233 sw
tri 414486 355713 416230 357457 ne
rect 416230 355713 425800 357457
tri 425800 355713 427544 357457 sw
tri 514486 356742 515201 357457 ne
rect 515201 356742 525800 357457
tri 525800 356742 526515 357457 sw
tri 515201 355713 516230 356742 ne
rect 516230 355713 526515 356742
tri 526515 355713 527544 356742 sw
tri 416230 351262 420681 355713 ne
rect 420681 351262 427544 355713
tri 427544 351262 431995 355713 sw
tri 516230 351262 520681 355713 ne
rect 520681 351262 527544 355713
tri 527544 351262 531995 355713 sw
tri 420681 344399 427544 351262 ne
rect 427544 344399 431995 351262
tri 431995 344399 438858 351262 sw
tri 520681 345428 526515 351262 ne
rect 526515 345428 531995 351262
tri 531995 345428 537829 351262 sw
tri 526515 344399 527544 345428 ne
rect 527544 344399 537829 345428
tri 537829 344399 538858 345428 sw
tri 427544 339344 432599 344399 ne
rect 432599 339344 438858 344399
tri 438858 339344 443913 344399 sw
tri 527544 339344 532599 344399 ne
rect 532599 339344 538858 344399
tri 538858 339344 543913 344399 sw
tri 432599 338900 433043 339344 ne
rect 433043 338900 443913 339344
tri 443913 338900 444357 339344 sw
tri 532599 338900 533043 339344 ne
rect 533043 338900 543913 339344
tri 543913 338900 544357 339344 sw
tri 433043 333085 438858 338900 ne
rect 438858 333085 444357 338900
tri 444357 333085 450172 338900 sw
tri 533043 334114 537829 338900 ne
rect 537829 338546 544357 338900
tri 544357 338546 544711 338900 sw
tri 699816 338546 700170 338900 se
rect 700170 338546 709342 338900
tri 709342 338546 709696 338900 sw
rect 537829 334114 544711 338546
tri 544711 334114 549143 338546 sw
tri 698756 337486 699816 338546 se
rect 699816 337840 709696 338546
tri 709696 337840 710402 338546 sw
rect 699816 337486 710402 337840
tri 710402 337486 710756 337840 sw
rect 698756 336900 710756 337486
tri 537829 333085 538858 334114 ne
rect 538858 333085 549143 334114
tri 549143 333085 550172 334114 sw
tri 438858 332800 439143 333085 ne
rect 439143 332800 450172 333085
tri 450172 332800 450457 333085 sw
tri 538858 332800 539143 333085 ne
rect 539143 332935 550172 333085
tri 550172 332935 550322 333085 sw
rect 539143 332800 550322 332935
tri 550322 332800 550457 332935 sw
tri 698603 332800 698756 332935 se
rect 698756 332800 700756 336900
tri 700756 335840 701816 336900 nw
tri 707696 335840 708756 336900 ne
tri 439143 327425 444518 332800 ne
rect 444518 327425 450457 332800
tri 450457 327425 455832 332800 sw
tri 539143 327425 544518 332800 ne
rect 544518 327870 550457 332800
tri 550457 327870 555387 332800 sw
tri 693024 327870 698603 332800 se
rect 698603 328900 700756 332800
tri 700756 328900 701816 329960 sw
tri 707696 328900 708756 329960 se
rect 708756 328900 710756 336900
rect 698603 328314 710756 328900
rect 698603 327960 710402 328314
tri 710402 327960 710756 328314 nw
rect 698603 327870 710312 327960
tri 710312 327870 710402 327960 nw
rect 544518 327425 555387 327870
tri 555387 327425 555832 327870 sw
tri 692520 327425 693024 327870 se
rect 693024 327425 709342 327870
tri 444518 326900 445043 327425 ne
rect 445043 326900 455832 327425
tri 455832 326900 456357 327425 sw
tri 544518 326900 545043 327425 ne
rect 545043 326900 555832 327425
tri 555832 326900 556357 327425 sw
tri 691926 326900 692520 327425 se
rect 692520 326900 709342 327425
tri 709342 326900 710312 327870 nw
tri 445043 324800 447143 326900 ne
rect 447143 324800 456357 326900
tri 456357 324800 458457 326900 sw
tri 545043 324800 547143 326900 ne
rect 547143 324800 556357 326900
tri 556357 324800 558457 326900 sw
tri 689550 324800 691926 326900 se
rect 691926 324800 699367 326900
rect 364800 321771 425457 322800
tri 425457 321771 426486 322800 sw
tri 447143 321771 450172 324800 ne
rect 450172 321771 458457 324800
tri 458457 321771 461486 324800 sw
tri 547143 322800 549143 324800 ne
rect 549143 322800 558457 324800
tri 558457 322800 560457 324800 sw
tri 687286 322800 689550 324800 se
rect 689550 322800 699367 324800
tri 699367 322800 704007 326900 nw
tri 549143 321771 550172 322800 ne
rect 550172 321771 690314 322800
rect 364800 318085 426486 321771
tri 426486 318085 430172 321771 sw
rect 364800 314800 430172 318085
tri 328643 239300 336771 247428 se
rect 336771 239300 339957 247428
tri 339957 239300 348085 247428 nw
tri 7985 238951 8334 239300 se
rect 8334 238951 17506 239300
tri 17506 238951 17855 239300 sw
tri 328294 238951 328643 239300 se
rect 328643 238951 339608 239300
tri 339608 238951 339957 239300 nw
tri 7269 238235 7985 238951 se
rect 7985 238235 17855 238951
tri 6920 237886 7269 238235 se
rect 7269 237886 17855 238235
tri 17855 237886 18920 238951 sw
rect 6920 237300 18920 237886
rect 6920 229300 8920 237300
tri 8920 236240 9980 237300 nw
tri 15860 236240 16920 237300 ne
rect 16920 233043 18920 237300
tri 325457 236114 328294 238951 se
rect 328294 236114 336771 238951
tri 336771 236114 339608 238951 nw
tri 322581 233238 325457 236114 se
rect 325457 235457 336114 236114
tri 336114 235457 336771 236114 nw
rect 325457 233238 333895 235457
tri 333895 233238 336114 235457 nw
tri 362581 233238 364800 235457 se
rect 364800 233238 372800 314800
tri 422143 313486 423457 314800 ne
rect 423457 313486 430172 314800
tri 430172 313486 434771 318085 sw
tri 450172 313486 458457 321771 ne
rect 458457 313486 461486 321771
tri 461486 313486 469771 321771 sw
tri 550172 314800 557143 321771 ne
rect 557143 314800 690314 321771
tri 690314 314800 699367 322800 nw
tri 423457 306771 430172 313486 ne
rect 430172 310457 434771 313486
tri 434771 310457 437800 313486 sw
tri 458457 310457 461486 313486 ne
rect 461486 310457 469771 313486
tri 469771 310457 472800 313486 sw
rect 430172 307143 437800 310457
tri 437800 307143 441114 310457 sw
tri 461486 307143 464800 310457 ne
rect 430172 306771 441114 307143
tri 441114 306771 441486 307143 sw
tri 430172 302172 434771 306771 ne
rect 434771 302172 441486 306771
tri 441486 302172 446085 306771 sw
tri 434771 295457 441486 302172 ne
rect 441486 295457 446085 302172
tri 446085 295457 452800 302172 sw
tri 441486 293900 443043 295457 ne
rect 443043 293900 452800 295457
tri 443043 292143 444800 293900 ne
tri 402581 233238 404800 235457 se
rect 404800 233238 412800 272800
tri 18920 233043 19134 233238 sw
tri 322386 233043 322581 233238 se
rect 322581 233043 333700 233238
tri 333700 233043 333895 233238 nw
tri 362386 233043 362581 233238 se
rect 362581 233043 372800 233238
tri 402386 233043 402581 233238 se
rect 402581 233043 412800 233238
tri 8920 229300 9980 230360 sw
tri 15860 229300 16920 230360 se
rect 16920 229300 19134 233043
rect 6920 228714 19134 229300
tri 6920 228365 7269 228714 ne
rect 7269 228365 19134 228714
tri 7269 227300 8334 228365 ne
rect 8334 227300 19134 228365
tri 13559 222210 19134 227300 ne
tri 19134 222800 30351 233043 sw
tri 322143 232800 322386 233043 se
rect 322386 232800 332800 233043
tri 264143 224800 272143 232800 se
rect 272143 232143 332800 232800
tri 332800 232143 333700 233043 nw
tri 361486 232143 362386 233043 se
rect 362386 232143 372800 233043
tri 401486 232143 402386 233043 se
rect 402386 232143 412800 233043
rect 272143 226085 326742 232143
tri 326742 226085 332800 232143 nw
tri 355428 226085 361486 232143 se
rect 361486 226085 366742 232143
tri 366742 226085 372800 232143 nw
tri 395428 226085 401486 232143 se
rect 401486 226085 406742 232143
tri 406742 226085 412800 232143 nw
rect 272143 224800 325457 226085
tri 325457 224800 326742 226085 nw
tri 264114 224771 264143 224800 se
rect 264143 224771 275428 224800
tri 275428 224771 275457 224800 nw
tri 262143 222800 264114 224771 se
rect 264114 224143 274800 224771
tri 274800 224143 275428 224771 nw
tri 353486 224143 355428 226085 se
rect 355428 224143 364800 226085
tri 364800 224143 366742 226085 nw
rect 264114 222800 273457 224143
tri 273457 222800 274800 224143 nw
tri 352143 222800 353486 224143 se
rect 353486 222800 363457 224143
tri 363457 222800 364800 224143 nw
tri 392143 222800 395428 226085 se
rect 395428 222800 403457 226085
tri 403457 222800 406742 226085 nw
rect 19134 222210 160457 222800
tri 160457 222210 161047 222800 sw
tri 261553 222210 262143 222800 se
rect 262143 222210 272867 222800
tri 272867 222210 273457 222800 nw
tri 351553 222210 352143 222800 se
rect 352143 222210 362867 222800
tri 362867 222210 363457 222800 nw
tri 391553 222210 392143 222800 se
rect 392143 222210 402867 222800
tri 402867 222210 403457 222800 nw
tri 19134 214800 27249 222210 ne
rect 27249 214800 161047 222210
tri 161047 214800 168457 222210 sw
tri 254143 214800 261553 222210 se
rect 261553 214800 265457 222210
tri 265457 214800 272867 222210 nw
tri 344143 214800 351553 222210 se
rect 351553 214800 355457 222210
tri 355457 214800 362867 222210 nw
tri 384143 214800 391553 222210 se
rect 391553 214800 395457 222210
tri 395457 214800 402867 222210 nw
tri 157143 203700 168243 214800 ne
rect 168243 203700 168457 214800
tri 168457 203700 179557 214800 sw
tri 252800 213457 254143 214800 se
rect 254143 214771 265428 214800
tri 265428 214771 265457 214800 nw
tri 344114 214771 344143 214800 se
rect 344143 214771 355428 214800
tri 355428 214771 355457 214800 nw
tri 384114 214771 384143 214800 se
rect 384143 214771 395428 214800
tri 395428 214771 395457 214800 nw
rect 254143 213457 264114 214771
tri 264114 213457 265428 214771 nw
tri 244800 205457 252800 213457 se
rect 252800 212829 263486 213457
tri 263486 212829 264114 213457 nw
tri 342172 212829 344114 214771 se
rect 344114 212829 353486 214771
tri 353486 212829 355428 214771 nw
rect 252800 212800 263457 212829
tri 263457 212800 263486 212829 nw
tri 342143 212800 342172 212829 se
rect 342172 212800 344357 212829
rect 252800 205457 255457 212800
rect 244800 204800 255457 205457
tri 255457 204800 263457 212800 nw
tri 274143 204800 282143 212800 se
rect 282143 207399 325457 212800
tri 325457 207399 330858 212800 sw
tri 336742 207399 342143 212800 se
rect 342143 207399 344357 212800
rect 282143 204800 330858 207399
tri 330858 204800 333457 207399 sw
tri 334143 204800 336742 207399 se
rect 336742 204800 344357 207399
rect 244800 203700 254357 204800
tri 254357 203700 255457 204800 nw
tri 273043 203700 274143 204800 se
rect 274143 203700 284357 204800
tri 284357 203700 285457 204800 nw
tri 322143 203700 323243 204800 ne
rect 323243 204457 333457 204800
tri 333457 204457 333800 204800 sw
tri 333800 204457 334143 204800 se
rect 334143 204457 344357 204800
rect 323243 203700 344357 204457
tri 344357 203700 353486 212829 nw
tri 373043 203700 384114 214771 se
rect 384114 203700 384357 214771
tri 384357 203700 395428 214771 nw
tri 168243 203486 168457 203700 ne
rect 168457 203486 179557 203700
tri 179557 203486 179771 203700 sw
rect 244800 203486 254143 203700
tri 254143 203486 254357 203700 nw
tri 272829 203486 273043 203700 se
rect 273043 203486 284143 203700
tri 284143 203486 284357 203700 nw
tri 323243 203486 323457 203700 ne
rect 323457 203486 344143 203700
tri 344143 203486 344357 203700 nw
tri 372829 203486 373043 203700 se
rect 373043 203486 384143 203700
tri 384143 203486 384357 203700 nw
tri 168457 196100 175843 203486 ne
rect 175843 196100 179771 203486
tri 7991 195757 8334 196100 se
rect 8334 195757 17506 196100
tri 17506 195757 17849 196100 sw
tri 175843 195757 176186 196100 ne
rect 176186 195757 179771 196100
tri 7263 195029 7991 195757 se
rect 7991 195139 17849 195757
tri 17849 195139 18467 195757 sw
tri 176186 195139 176804 195757 ne
rect 176804 195139 179771 195757
rect 7991 195029 18467 195139
tri 6920 194686 7263 195029 se
rect 7263 194686 18467 195029
tri 18467 194686 18920 195139 sw
rect 6920 194100 18920 194686
rect 6920 186100 8920 194100
tri 8920 193040 9980 194100 nw
tri 15860 193040 16920 194100 ne
tri 8920 186100 9980 187160 sw
tri 15860 186100 16920 187160 se
rect 16920 186100 18920 194100
tri 176804 192172 179771 195139 ne
tri 179771 192172 191085 203486 sw
rect 244800 203457 254114 203486
tri 254114 203457 254143 203486 nw
tri 272800 203457 272829 203486 se
rect 272829 203457 284114 203486
tri 284114 203457 284143 203486 nw
tri 323457 203457 323486 203486 ne
rect 323486 203457 344114 203486
tri 344114 203457 344143 203486 nw
tri 372800 203457 372829 203486 se
rect 372829 203457 384114 203486
tri 384114 203457 384143 203486 nw
tri 179771 191700 180243 192172 ne
rect 180243 191700 191085 192172
tri 191085 191700 191557 192172 sw
tri 180243 189693 182250 191700 ne
rect 182250 189693 191557 191700
rect 6920 185514 18920 186100
tri 6920 185171 7263 185514 ne
rect 7263 185171 18920 185514
tri 7263 184100 8334 185171 ne
rect 8334 185061 18920 185171
tri 18920 185061 23461 189693 sw
tri 182250 185061 186882 189693 ne
rect 186882 185061 191557 189693
rect 8334 184100 23461 185061
tri 13200 178728 18467 184100 ne
rect 18467 178728 23461 184100
tri 23461 178728 29670 185061 sw
tri 186882 180858 191085 185061 ne
rect 191085 180858 191557 185061
tri 191557 180858 202399 191700 sw
tri 191085 178728 193215 180858 ne
rect 193215 178728 202399 180858
tri 18467 167300 29670 178728 ne
tri 29670 172800 35480 178728 sw
tri 193215 172800 199143 178728 ne
rect 199143 174457 202399 178728
tri 202399 174457 208800 180858 sw
rect 199143 172800 208800 174457
rect 29670 167300 112800 172800
tri 199143 169544 202399 172800 ne
rect 202399 169544 208800 172800
tri 208800 169544 213713 174457 sw
tri 29670 164800 32120 167300 ne
rect 32120 164800 112800 167300
tri 202399 164800 207143 169544 ne
rect 207143 168800 213713 169544
tri 213713 168800 214457 169544 sw
rect 207143 164800 208800 168800
tri 207143 163143 208800 164800 ne
tri 208800 163143 214457 168800 nw
tri 241486 152143 244800 155457 se
rect 244800 152143 252800 203457
tri 252800 202143 254114 203457 nw
tri 236771 147428 241486 152143 se
rect 241486 147428 248085 152143
tri 248085 147428 252800 152143 nw
tri 264800 195457 272800 203457 se
rect 272800 195457 272829 203457
rect 264800 192172 272829 195457
tri 272829 192172 284114 203457 nw
tri 323486 201515 325428 203457 ne
rect 325428 201515 342172 203457
tri 342172 201515 344114 203457 nw
tri 325428 198800 328143 201515 ne
rect 328143 198800 339457 201515
tri 339457 198800 342172 201515 nw
tri 328143 193486 333457 198800 ne
rect 333457 196085 339457 198800
tri 339457 196085 342172 198800 sw
rect 333457 193486 342172 196085
tri 342172 193486 344771 196085 sw
tri 364800 195457 372800 203457 se
rect 372800 203354 384011 203457
tri 384011 203354 384114 203457 nw
rect 372800 197571 378228 203354
tri 378228 197571 384011 203354 nw
rect 372800 195457 373065 197571
tri 333457 193143 333800 193486 ne
rect 333800 193143 344771 193486
tri 333800 192172 334771 193143 ne
rect 334771 192172 344771 193143
tri 225457 136114 236771 147428 se
rect 236771 145457 246114 147428
tri 246114 145457 248085 147428 nw
rect 236771 142143 242800 145457
tri 242800 142143 246114 145457 nw
tri 261486 142143 264800 145457 se
rect 264800 142143 272800 192172
tri 272800 192143 272829 192172 nw
tri 334771 192143 334800 192172 ne
rect 334800 192143 344771 192172
tri 334800 191700 335243 192143 ne
rect 335243 191700 344771 192143
tri 335243 182172 344771 191700 ne
tri 344771 185457 352800 193486 sw
rect 344771 182172 352800 185457
tri 344771 182143 344800 182172 ne
tri 303887 169544 308800 174457 se
tri 308800 169544 313713 174457 sw
tri 303143 168800 303887 169544 se
rect 303887 168800 313713 169544
tri 313713 168800 314457 169544 sw
tri 299114 164771 303143 168800 se
rect 303143 164771 310428 168800
tri 310428 164771 314457 168800 nw
tri 297486 163143 299114 164771 se
rect 299114 163143 308800 164771
tri 308800 163143 310428 164771 nw
tri 287800 153457 297486 163143 se
rect 297486 158700 304357 163143
tri 304357 158700 308800 163143 nw
rect 297486 153457 299114 158700
tri 299114 153457 304357 158700 nw
rect 236771 138742 239399 142143
tri 239399 138742 242800 142143 nw
tri 258085 138742 261486 142143 se
rect 261486 138742 269399 142143
tri 269399 138742 272800 142143 nw
tri 279800 145457 287800 153457 se
rect 287800 146700 292357 153457
tri 292357 146700 299114 153457 nw
tri 236771 136114 239399 138742 nw
tri 255457 136114 258085 138742 se
rect 258085 136114 266114 138742
tri 222143 132800 225457 136114 se
rect 225457 132800 228085 136114
tri 149143 124800 157143 132800 se
rect 157143 127428 228085 132800
tri 228085 127428 236771 136114 nw
tri 246771 127428 255457 136114 se
rect 255457 135457 266114 136114
tri 266114 135457 269399 138742 nw
rect 255457 132143 262800 135457
tri 262800 132143 266114 135457 nw
tri 276486 132143 279800 135457 se
rect 279800 132143 287800 145457
tri 287800 142143 292357 146700 nw
tri 341486 142143 344800 145457 se
rect 344800 142143 352800 182172
tri 333486 134143 341486 142143 se
rect 341486 134143 344800 142143
tri 344800 134143 352800 142143 nw
rect 364800 192408 373065 195457
tri 373065 192408 378228 197571 nw
rect 364800 192172 372829 192408
tri 372829 192172 373065 192408 nw
rect 255457 131085 261742 132143
tri 261742 131085 262800 132143 nw
tri 275428 131085 276486 132143 se
rect 276486 131085 286742 132143
tri 286742 131085 287800 132143 nw
tri 330428 131085 333486 134143 se
rect 255457 127428 258085 131085
tri 258085 127428 261742 131085 nw
tri 271771 127428 275428 131085 se
rect 275428 127428 279357 131085
rect 157143 124800 225457 127428
tri 225457 124800 228085 127428 nw
tri 148043 123700 149143 124800 se
rect 149143 123700 159357 124800
tri 159357 123700 160457 124800 nw
tri 243043 123700 246771 127428 se
rect 246771 123700 254357 127428
tri 254357 123700 258085 127428 nw
tri 268043 123700 271771 127428 se
rect 271771 123700 279357 127428
tri 279357 123700 286742 131085 nw
tri 323043 123700 330428 131085 se
rect 330428 123700 333486 131085
tri 7434 122800 8334 123700 se
rect 8334 122800 17506 123700
tri 17506 122800 18406 123700 sw
tri 147143 122800 148043 123700 se
rect 148043 122800 151771 123700
tri 6920 122286 7434 122800 se
rect 7434 122798 18406 122800
tri 18406 122798 18408 122800 sw
tri 18419 122798 18429 122800 se
rect 18429 122798 151771 122800
rect 7434 122796 18408 122798
tri 18408 122796 18410 122798 sw
tri 18410 122796 18419 122798 se
rect 18419 122796 151771 122798
rect 7434 122286 151771 122796
rect 6920 121700 151771 122286
rect 6920 113700 8920 121700
tri 8920 120640 9980 121700 nw
tri 15860 120640 16920 121700 ne
rect 16920 116114 151771 121700
tri 151771 116114 159357 123700 nw
tri 235457 116114 243043 123700 se
rect 243043 119771 250428 123700
tri 250428 119771 254357 123700 nw
tri 264114 119771 268043 123700 se
rect 268043 119771 275428 123700
tri 275428 119771 279357 123700 nw
tri 322172 122829 323043 123700 se
rect 323043 122829 333486 123700
tri 333486 122829 344800 134143 nw
tri 322143 122800 322172 122829 se
rect 322172 122800 333457 122829
tri 333457 122800 333486 122829 nw
tri 294114 119771 297143 122800 se
rect 297143 119771 325457 122800
rect 243043 116114 246771 119771
tri 246771 116114 250428 119771 nw
tri 260457 116114 264114 119771 se
rect 264114 116114 269157 119771
rect 16920 114800 150457 116114
tri 150457 114800 151771 116114 nw
tri 8920 113700 9980 114760 sw
tri 15860 113700 16920 114760 se
rect 16920 113700 18920 114800
tri 18920 114753 19171 114800 nw
rect 6920 113114 18920 113700
tri 6920 113033 7001 113114 ne
rect 7001 113033 18839 113114
tri 18839 113033 18920 113114 nw
tri 7001 111700 8334 113033 ne
rect 8334 111700 17506 113033
tri 17506 111700 18839 113033 nw
tri 232143 112800 235457 116114 se
rect 235457 112800 242357 116114
tri 171043 111700 172143 112800 se
rect 172143 111700 242357 112800
tri 242357 111700 246771 116114 nw
tri 256043 111700 260457 116114 se
rect 260457 113500 269157 116114
tri 269157 113500 275428 119771 nw
tri 287843 113500 294114 119771 se
rect 294114 114800 325457 119771
tri 325457 114800 333457 122800 nw
rect 294114 113500 297143 114800
rect 260457 111700 267357 113500
tri 267357 111700 269157 113500 nw
tri 286043 111700 287843 113500 se
rect 287843 111700 297143 113500
tri 164143 104800 171043 111700 se
rect 171043 108457 239114 111700
tri 239114 108457 242357 111700 nw
tri 252800 108457 256043 111700 se
rect 256043 108457 264114 111700
tri 264114 108457 267357 111700 nw
tri 285829 111486 286043 111700 se
rect 286043 111486 297143 111700
tri 297143 111486 300457 114800 nw
tri 282800 108457 285829 111486 se
rect 171043 104800 235457 108457
tri 235457 104800 239114 108457 nw
tri 249143 104800 252800 108457 se
rect 252800 104800 257157 108457
tri 162800 103457 164143 104800 se
rect 164143 103457 174114 104800
tri 174114 103457 175457 104800 nw
tri 154800 95457 162800 103457 se
tri 7979 81145 8334 81500 se
rect 8334 81145 17506 81500
tri 7275 80441 7979 81145 se
rect 7979 80441 17506 81145
tri 6920 80086 7275 80441 se
rect 7275 80086 17506 80441
tri 17506 80086 18920 81500 sw
rect 6920 79500 18920 80086
rect 6920 71500 8920 79500
tri 8920 78440 9980 79500 nw
tri 15860 78440 16920 79500 ne
rect 16920 72800 18920 79500
tri 18920 72800 20612 74727 sw
tri 8920 71500 9980 72560 sw
tri 15860 71500 16920 72560 se
rect 16920 71500 112800 72800
rect 6920 70914 112800 71500
tri 6920 70559 7275 70914 ne
rect 7275 70559 112800 70914
tri 7275 69500 8334 70559 ne
rect 8334 69500 112800 70559
tri 12863 64800 16988 69500 ne
rect 16988 64800 112800 69500
tri 154143 64800 154800 65457 se
rect 154800 64800 162800 95457
tri 162800 92143 174114 103457 nw
tri 244800 100457 249143 104800 se
rect 249143 101500 257157 104800
tri 257157 101500 264114 108457 nw
tri 275843 101500 282800 108457 se
rect 282800 101500 285829 108457
rect 249143 100457 252800 101500
tri 207143 72800 208800 74457 se
tri 208800 72800 210457 74457 sw
tri 203143 68800 207143 72800 se
rect 207143 68800 210457 72800
tri 210457 68800 214457 72800 sw
tri 199143 64800 203143 68800 se
rect 203143 64800 210457 68800
tri 210457 64800 214457 68800 nw
tri 151486 62143 154143 64800 se
rect 154143 62143 162800 64800
tri 148085 58742 151486 62143 se
rect 151486 58742 159399 62143
tri 159399 58742 162800 62143 nw
tri 193085 58742 199143 64800 se
rect 199143 58742 204399 64800
tri 204399 58742 210457 64800 nw
tri 136771 47428 148085 58742 se
tri 148085 47428 159399 58742 nw
tri 181771 47428 193085 58742 se
tri 193085 47428 204399 58742 nw
tri 241771 47428 244800 50457 se
rect 244800 47428 252800 100457
tri 252800 97143 257157 101500 nw
tri 274515 100172 275843 101500 se
rect 275843 100172 285829 101500
tri 285829 100172 297143 111486 nw
tri 271486 97143 274515 100172 se
rect 274515 97143 276114 100172
tri 125457 36114 136771 47428 se
tri 136771 36114 148085 47428 nw
tri 170457 36114 181771 47428 se
tri 181771 36114 193085 47428 nw
tri 241486 47143 241771 47428 se
rect 241771 47143 252800 47428
tri 230457 36114 241486 47143 se
rect 241486 36114 241771 47143
tri 241771 36114 252800 47143 nw
tri 264800 90457 271486 97143 se
rect 271486 90457 276114 97143
tri 276114 90457 285829 100172 nw
tri 122143 32800 125457 36114 se
rect 125457 32800 133457 36114
tri 133457 32800 136771 36114 nw
tri 167143 32800 170457 36114 se
tri 93440 24800 102256 32800 se
rect 102256 24800 125457 32800
tri 125457 24800 133457 32800 nw
tri 145067 24800 151968 32800 se
rect 151968 24800 170457 32800
tri 170457 24800 181771 36114 nw
tri 227143 32800 230457 36114 se
tri 199562 24800 207068 32800 se
rect 207068 24800 230457 32800
tri 230457 24800 241771 36114 nw
tri 254585 24801 264800 35412 se
rect 264800 32188 272800 90457
tri 272800 87143 276114 90457 nw
tri 361486 77143 364800 80457 se
rect 364800 77143 372800 192172
tri 372800 192143 372829 192172 nw
rect 404800 132143 412800 172800
rect 444800 144114 452800 293900
rect 464800 147143 472800 310457
tri 699821 293551 700170 293900 se
rect 700170 293551 709342 293900
tri 709342 293551 709691 293900 sw
tri 698756 292486 699821 293551 se
rect 699821 292835 709691 293551
tri 709691 292835 710407 293551 sw
rect 699821 292486 710407 292835
tri 710407 292486 710756 292835 sw
rect 698756 291900 710756 292486
tri 693142 282726 698756 287843 se
rect 698756 283900 700756 291900
tri 700756 290840 701816 291900 nw
tri 707696 290840 708756 291900 ne
tri 700756 283900 701816 284960 sw
tri 707696 283900 708756 284960 se
rect 708756 283900 710756 291900
rect 698756 283314 710756 283900
rect 698756 282965 710407 283314
tri 710407 282965 710756 283314 nw
rect 698756 282726 710168 282965
tri 710168 282726 710407 282965 nw
tri 692236 281900 693142 282726 se
rect 693142 281900 709342 282726
tri 709342 281900 710168 282726 nw
tri 689651 279544 692236 281900 se
rect 692236 279544 694126 281900
tri 684069 274457 689651 279544 se
rect 689651 274457 694126 279544
tri 507143 272800 508800 274457 se
tri 508800 272800 510457 274457 sw
tri 682251 272800 684069 274457 se
rect 684069 272800 694126 274457
tri 694126 272800 704112 281900 nw
tri 503143 268800 507143 272800 se
rect 507143 268800 510457 272800
tri 503143 268056 503887 268800 ne
rect 503887 268056 510457 268800
tri 510457 268056 515201 272800 sw
rect 604800 268056 688921 272800
tri 688921 268056 694126 272800 nw
tri 503887 263143 508800 268056 ne
rect 508800 263143 515201 268056
tri 508800 256742 515201 263143 ne
tri 515201 256742 526515 268056 sw
rect 604800 264800 685349 268056
tri 685349 264800 688921 268056 nw
tri 515201 245428 526515 256742 ne
tri 526515 248900 534357 256742 sw
rect 526515 248553 534357 248900
tri 534357 248553 534704 248900 sw
tri 699823 248553 700170 248900 se
rect 700170 248553 709342 248900
tri 709342 248553 709689 248900 sw
rect 526515 245428 534704 248553
tri 534704 245428 537829 248553 sw
tri 698756 247486 699823 248553 se
rect 699823 247833 709689 248553
tri 709689 247833 710409 248553 sw
rect 699823 247486 710409 247833
tri 710409 247486 710756 247833 sw
rect 698756 246900 710756 247486
tri 526515 234114 537829 245428 ne
tri 537829 242787 540470 245428 sw
rect 537829 237636 540470 242787
tri 540470 237636 545621 242787 sw
tri 693208 237636 698756 242787 se
rect 698756 238900 700756 246900
tri 700756 245840 701816 246900 nw
tri 707696 245840 708756 246900 ne
tri 700756 238900 701816 239960 sw
tri 707696 238900 708756 239960 se
rect 708756 238900 710756 246900
rect 698756 238314 710756 238900
rect 698756 237967 710409 238314
tri 710409 237967 710756 238314 nw
rect 698756 237636 710078 237967
tri 710078 237636 710409 237967 nw
rect 537829 236900 545621 237636
tri 545621 236900 546357 237636 sw
tri 692415 236900 693208 237636 se
rect 693208 236900 709342 237636
tri 709342 236900 710078 237636 nw
rect 537829 234114 546357 236900
tri 546357 234114 549143 236900 sw
tri 537829 226085 545858 234114 ne
rect 545858 226718 549143 234114
tri 549143 226718 556539 234114 sw
tri 681449 226718 692415 236900 se
rect 692415 226718 693208 236900
tri 693208 226718 704173 236900 nw
rect 545858 226085 556539 226718
tri 556539 226085 557172 226718 sw
tri 680767 226085 681449 226718 se
rect 681449 226085 688987 226718
tri 545858 222800 549143 226085 ne
rect 549143 222800 557172 226085
tri 557172 222800 560457 226085 sw
tri 677229 222800 680767 226085 se
rect 680767 222800 688987 226085
tri 688987 222800 693208 226718 nw
tri 549143 222210 549733 222800 ne
rect 549733 222210 680371 222800
tri 549733 214800 557143 222210 ne
rect 557143 214800 680371 222210
tri 680371 214800 688987 222800 nw
tri 699824 203354 700170 203700 se
rect 700170 203354 709342 203700
tri 709342 203354 709688 203700 sw
tri 698756 202286 699824 203354 se
rect 699824 202632 709688 203354
tri 709688 202632 710410 203354 sw
rect 699824 202286 710410 202632
tri 710410 202286 710756 202632 sw
rect 698756 201700 710756 202286
tri 693226 192408 698756 197571 se
rect 698756 193700 700756 201700
tri 700756 200640 701816 201700 nw
tri 707696 200640 708756 201700 ne
tri 700756 193700 701816 194760 sw
tri 707696 193700 708756 194760 se
rect 708756 193700 710756 201700
rect 698756 193114 710756 193700
rect 698756 192768 710410 193114
tri 710410 192768 710756 193114 nw
rect 698756 192408 710050 192768
tri 710050 192408 710410 192768 nw
tri 692973 192172 693226 192408 se
rect 693226 192172 709342 192408
tri 692468 191700 692973 192172 se
rect 692973 191700 709342 192172
tri 709342 191700 710050 192408 nw
tri 681503 181463 692468 191700 se
rect 692468 181463 693226 191700
tri 693226 181463 704192 191700 nw
tri 680855 180858 681503 181463 se
rect 681503 180858 683946 181463
tri 673998 174457 680855 180858 se
rect 680855 174457 683946 180858
tri 672223 172800 673998 174457 se
rect 673998 172800 683946 174457
tri 683946 172800 693226 181463 nw
rect 504800 166742 545457 172800
tri 545457 166742 551515 172800 sw
rect 604800 166742 677457 172800
tri 677457 166742 683946 172800 nw
rect 504800 164800 551515 166742
tri 542143 155428 551515 164800 ne
tri 551515 158700 559557 166742 sw
rect 604800 164800 675377 166742
tri 675377 164800 677457 166742 nw
rect 551515 158352 559557 158700
tri 559557 158352 559905 158700 sw
tri 699822 158352 700170 158700 se
rect 700170 158352 709342 158700
tri 709342 158352 709690 158700 sw
rect 551515 155428 559905 158352
tri 559905 155428 562829 158352 sw
tri 698756 157286 699822 158352 se
rect 699822 157634 709690 158352
tri 709690 157634 710408 158352 sw
rect 699822 157286 710408 157634
tri 710408 157286 710756 157634 sw
rect 698756 156700 710756 157286
tri 452800 144114 454143 145457 sw
tri 464800 144114 467829 147143 ne
rect 467829 144114 472800 147143
tri 472800 144114 479143 150457 sw
tri 551515 144114 562829 155428 ne
tri 562829 152612 565645 155428 sw
rect 698756 152612 700756 156700
tri 700756 155640 701816 156700 nw
tri 707696 155640 708756 156700 ne
rect 562829 147477 565645 152612
tri 565645 147477 570780 152612 sw
tri 693179 147477 698755 152612 se
rect 698755 148700 700756 152612
tri 700756 148700 701816 149760 sw
tri 707696 148700 708756 149760 se
rect 708756 148700 710756 156700
rect 698755 148114 710756 148700
rect 698755 147766 710408 148114
tri 710408 147766 710756 148114 nw
rect 698755 147477 710119 147766
tri 710119 147477 710408 147766 nw
rect 562829 146700 570780 147477
tri 570780 146700 571557 147477 sw
tri 692335 146700 693179 147477 se
rect 693179 146700 709342 147477
tri 709342 146700 710119 147477 nw
rect 562829 144114 571557 146700
tri 571557 144114 574143 146700 sw
rect 444800 142143 454143 144114
tri 444800 135457 451486 142143 ne
rect 451486 139143 454143 142143
tri 454143 139143 459114 144114 sw
tri 467829 139143 472800 144114 ne
rect 472800 139143 479143 144114
rect 451486 135457 459114 139143
tri 459114 135457 462800 139143 sw
tri 472800 135457 476486 139143 ne
rect 476486 135457 479143 139143
tri 479143 135457 487800 144114 sw
tri 562829 135457 571486 144114 ne
rect 571486 136602 574143 144114
tri 574143 136602 581655 144114 sw
tri 681369 136602 692335 146700 se
rect 692335 136602 693179 146700
tri 693179 136602 704145 146700 nw
rect 571486 135457 581655 136602
tri 581655 135457 582800 136602 sw
tri 680125 135457 681369 136602 se
rect 681369 135457 689049 136602
tri 404800 131085 405858 132143 ne
rect 405858 131085 412800 132143
tri 412800 131085 417172 135457 sw
tri 451486 135428 451515 135457 ne
rect 451515 135428 462800 135457
tri 462800 135428 462829 135457 sw
tri 451515 134143 452800 135428 ne
rect 452800 134143 462829 135428
tri 452800 131085 455858 134143 ne
rect 455858 132800 462829 134143
tri 462829 132800 465457 135428 sw
tri 476486 132800 479143 135457 ne
rect 479143 132800 487800 135457
tri 487800 132800 490457 135457 sw
tri 571486 132800 574143 135457 ne
rect 574143 132800 582800 135457
tri 582800 132800 585457 135457 sw
tri 677239 132800 680125 135457 se
rect 680125 132800 689049 135457
tri 689049 132800 693179 136602 nw
rect 455858 131085 465457 132800
tri 465457 131085 467172 132800 sw
tri 479143 131085 480858 132800 ne
rect 480858 131085 550457 132800
tri 550457 131085 552172 132800 sw
tri 574143 131085 575858 132800 ne
rect 575858 131085 680361 132800
tri 405858 130713 406230 131085 ne
rect 406230 130713 417172 131085
tri 417172 130713 417544 131085 sw
tri 455858 130713 456230 131085 ne
rect 456230 130713 467172 131085
tri 467172 130713 467544 131085 sw
tri 480858 130713 481230 131085 ne
rect 481230 130713 552172 131085
tri 552172 130713 552544 131085 sw
tri 575858 130713 576230 131085 ne
rect 576230 130713 680361 131085
tri 406230 124143 412800 130713 ne
rect 412800 124143 417544 130713
tri 412800 123700 413243 124143 ne
rect 413243 123700 417544 124143
tri 417544 123700 424557 130713 sw
tri 456230 124114 462829 130713 ne
rect 462829 124800 467544 130713
tri 467544 124800 473457 130713 sw
tri 481230 124800 487143 130713 ne
rect 487143 124800 552544 130713
tri 552544 124800 558457 130713 sw
tri 576230 124800 582143 130713 ne
rect 582143 124800 680361 130713
tri 680361 124800 689049 132800 nw
rect 462829 124114 473457 124800
tri 473457 124114 474143 124800 sw
tri 547143 124114 547829 124800 ne
rect 547829 124114 558457 124800
tri 558457 124114 559143 124800 sw
tri 462829 123700 463243 124114 ne
rect 463243 123700 474143 124114
tri 474143 123700 474557 124114 sw
tri 547829 123700 548243 124114 ne
rect 548243 123700 559143 124114
tri 559143 123700 559557 124114 sw
tri 413243 119771 417172 123700 ne
rect 417172 119771 424557 123700
tri 424557 119771 428486 123700 sw
tri 463243 119771 467172 123700 ne
rect 467172 121486 474557 123700
tri 474557 121486 476771 123700 sw
tri 548243 121486 550457 123700 ne
rect 550457 121486 559557 123700
rect 467172 119771 476771 121486
tri 476771 119771 478486 121486 sw
tri 550457 119771 552172 121486 ne
rect 552172 119771 559557 121486
tri 559557 119771 563486 123700 sw
tri 417172 119399 417544 119771 ne
rect 417544 119399 428486 119771
tri 428486 119399 428858 119771 sw
tri 467172 119399 467544 119771 ne
rect 467544 119399 478486 119771
tri 478486 119399 478858 119771 sw
tri 552172 119399 552544 119771 ne
rect 552544 119399 563486 119771
tri 563486 119399 563858 119771 sw
tri 417544 113500 423443 119399 ne
rect 423443 113500 428858 119399
tri 428858 113500 434757 119399 sw
tri 467544 113500 473443 119399 ne
rect 473443 113500 478858 119399
tri 478858 113500 484757 119399 sw
tri 552544 113500 558443 119399 ne
rect 558443 113500 563858 119399
tri 563858 113500 569757 119399 sw
tri 423443 111700 425243 113500 ne
rect 425243 111700 434757 113500
tri 434757 111700 436557 113500 sw
tri 473443 112800 474143 113500 ne
rect 474143 112800 484757 113500
tri 484757 112800 485457 113500 sw
tri 558443 112800 559143 113500 ne
rect 559143 112800 569757 113500
tri 569757 112800 570457 113500 sw
tri 699470 112800 700170 113500 se
rect 700170 112800 709342 113500
tri 709342 112800 710042 113500 sw
tri 474143 111700 475243 112800 ne
rect 475243 112561 540457 112800
tri 540457 112561 540696 112800 sw
tri 559143 112561 559382 112800 ne
rect 559382 112758 699231 112800
tri 699231 112758 699417 112800 sw
tri 699428 112758 699470 112800 se
rect 699470 112758 710042 112800
rect 559382 112756 699420 112758
tri 699420 112756 699426 112758 sw
tri 699426 112756 699428 112758 se
rect 699428 112756 710042 112758
rect 559382 112561 710042 112756
rect 475243 111700 540696 112561
tri 540696 111700 541557 112561 sw
tri 559382 111700 560243 112561 ne
rect 560243 112086 710042 112561
tri 710042 112086 710756 112800 sw
rect 560243 111700 710756 112086
tri 425243 108457 428486 111700 ne
rect 428486 108457 436557 111700
tri 436557 108457 439800 111700 sw
tri 475243 108457 478486 111700 ne
rect 478486 108457 541557 111700
tri 541557 108457 544800 111700 sw
tri 560243 108457 563486 111700 ne
rect 563486 111500 710756 111700
rect 563486 108457 700756 111500
tri 700756 110440 701816 111500 nw
tri 707696 110440 708756 111500 ne
tri 428486 108085 428858 108457 ne
rect 428858 108085 439800 108457
tri 439800 108085 440172 108457 sw
tri 478486 108085 478858 108457 ne
rect 478858 108085 544800 108457
tri 544800 108085 545172 108457 sw
tri 563486 108085 563858 108457 ne
rect 563858 108085 700756 108457
tri 428858 101500 435443 108085 ne
rect 435443 101500 440172 108085
tri 440172 101500 446757 108085 sw
tri 478858 104800 482143 108085 ne
rect 482143 104800 545172 108085
tri 545172 104800 548457 108085 sw
tri 563858 104800 567143 108085 ne
rect 567143 104800 700756 108085
tri 537143 101771 540172 104800 ne
rect 540172 104715 548457 104800
tri 548457 104715 548542 104800 sw
tri 698369 104715 698756 104800 ne
rect 540172 102739 548542 104715
tri 548542 102739 550518 104715 sw
rect 698756 103500 700756 104800
tri 700756 103500 701816 104560 sw
tri 707696 103500 708756 104560 se
rect 708756 103500 710756 111500
rect 698756 102914 710756 103500
tri 698756 102739 698931 102914 ne
rect 698931 102739 710581 102914
tri 710581 102739 710756 102914 nw
rect 540172 101771 550518 102739
tri 550518 101771 551486 102739 sw
tri 540172 101500 540443 101771 ne
rect 540443 101500 551486 101771
tri 551486 101500 551757 101771 sw
tri 698931 101500 700170 102739 ne
rect 700170 101500 709342 102739
tri 709342 101500 710581 102739 nw
tri 435443 97143 439800 101500 ne
rect 439800 97143 446757 101500
tri 446757 97143 451114 101500 sw
tri 540443 101486 540457 101500 ne
rect 540457 101486 551757 101500
tri 540457 97143 544800 101486 ne
rect 544800 97143 551757 101486
tri 551757 97143 556114 101500 sw
tri 439800 96771 440172 97143 ne
rect 440172 96771 451114 97143
tri 451114 96771 451486 97143 sw
tri 544800 96771 545172 97143 ne
rect 545172 96771 556114 97143
tri 556114 96771 556486 97143 sw
tri 440172 85457 451486 96771 ne
tri 451486 85457 462800 96771 sw
tri 545172 90457 551486 96771 ne
rect 551486 90457 556486 96771
tri 556486 90457 562800 96771 sw
tri 551486 87143 554800 90457 ne
tri 451486 82143 454800 85457 ne
tri 357143 72800 361486 77143 se
rect 361486 72800 368457 77143
tri 368457 72800 372800 77143 nw
tri 86960 18920 93440 24800 se
rect 93440 19526 99531 24800
tri 99531 19526 105344 24800 nw
tri 140516 19526 145067 24800 se
rect 145067 19526 151082 24800
tri 151082 19526 155632 24800 nw
tri 194613 19526 199562 24800 se
rect 199562 20538 206533 24800
tri 206533 20538 210532 24800 nw
tri 253696 23877 254585 24800 se
rect 254585 23877 264800 24801
tri 264800 23877 272800 32188 nw
tri 250482 20538 253696 23877 se
rect 253696 20538 261586 23877
tri 261586 20538 264800 23877 nw
rect 199562 19526 205583 20538
tri 205583 19526 206533 20538 nw
tri 249507 19526 250482 20538 se
rect 250482 19526 260611 20538
tri 260611 19526 261586 20538 nw
tri 303716 19526 304800 20538 se
rect 304800 19526 312800 72800
rect 93440 18920 98864 19526
tri 98864 18920 99531 19526 nw
tri 139993 18920 140516 19526 se
rect 140516 18920 150559 19526
tri 150559 18920 151082 19526 nw
tri 194080 18958 194613 19526 se
rect 194613 18958 205050 19526
tri 205050 18958 205583 19526 nw
tri 248961 18958 249507 19526 se
rect 249507 18958 260028 19526
tri 194044 18920 194080 18958 se
rect 194080 18920 205014 18958
tri 205014 18920 205050 18958 nw
tri 248924 18920 248961 18958 se
rect 248961 18920 260028 18958
tri 260028 18920 260611 19526 nw
tri 303067 18920 303716 19526 se
rect 303716 18920 312800 19526
tri 354800 70457 357143 72800 se
rect 357143 70457 362800 72800
tri 354703 18922 354800 19302 se
rect 354800 18922 362800 70457
tri 362800 67143 368457 72800 nw
rect 354703 18920 362800 18922
tri 80867 18073 81714 18920 se
rect 81714 18073 97930 18920
tri 97930 18073 98864 18920 nw
tri 80650 17856 80867 18073 se
rect 80867 17864 97700 18073
tri 97700 17864 97930 18073 nw
tri 134458 17864 135514 18920 se
rect 135514 17864 146100 18920
rect 80867 17856 92300 17864
tri 80300 17506 80650 17856 se
rect 80650 17506 92300 17856
rect 80300 16920 92300 17506
rect 80300 8920 82300 16920
tri 82300 15860 83360 16920 nw
tri 89240 15860 90300 16920 ne
tri 82300 8920 83360 9980 sw
tri 89240 8920 90300 9980 se
rect 90300 8920 92300 16920
tri 92300 12964 97700 17864 nw
tri 134100 17506 134458 17864 se
rect 134458 17506 146100 17864
rect 134100 16920 146100 17506
rect 80300 8334 92300 8920
tri 80300 7984 80650 8334 ne
rect 80650 7984 91236 8334
tri 80650 7270 81364 7984 ne
rect 81364 7270 91236 7984
tri 91236 7270 92300 8334 nw
rect 134100 8920 136100 16920
tri 136100 15860 137160 16920 nw
tri 143040 15860 144100 16920 ne
tri 136100 8920 137160 9980 sw
tri 143040 8920 144100 9980 se
rect 144100 8920 146100 16920
tri 146100 13751 150559 18920 nw
tri 188246 17852 189314 18920 se
rect 189314 17852 199900 18920
tri 187900 17506 188246 17852 se
rect 188246 17506 199900 17852
rect 187900 16920 199900 17506
rect 134100 8334 146100 8920
tri 134100 7976 134458 8334 ne
rect 134458 7976 145044 8334
tri 134458 7278 135156 7976 ne
rect 135156 7278 145044 7976
tri 145044 7278 146100 8334 nw
rect 187900 8920 189900 16920
tri 189900 15860 190960 16920 nw
tri 196840 15860 197900 16920 ne
tri 189900 8920 190960 9980 sw
tri 196840 8920 197900 9980 se
rect 197900 8920 199900 16920
tri 199900 13469 205014 18920 nw
tri 243044 17850 244114 18920 se
rect 244114 18510 259633 18920
tri 259633 18510 260028 18920 nw
rect 244114 18058 259198 18510
tri 259198 18058 259633 18510 nw
rect 244114 17850 254700 18058
tri 242700 17506 243044 17850 se
rect 243044 17506 254700 17850
rect 242700 16920 254700 17506
rect 187900 8334 199900 8920
tri 187900 7988 188246 8334 ne
rect 188246 7988 198832 8334
tri 81364 6920 81714 7270 ne
rect 81714 6920 90886 7270
tri 90886 6920 91236 7270 nw
tri 135156 6920 135514 7278 ne
rect 135514 6920 144686 7278
tri 144686 6920 145044 7278 nw
tri 188246 7266 188968 7988 ne
rect 188968 7266 198832 7988
tri 198832 7266 199900 8334 nw
rect 242700 8920 244700 16920
tri 244700 15860 245760 16920 nw
tri 251640 15860 252700 16920 ne
tri 244700 8920 245760 9980 sw
tri 251640 8920 252700 9980 se
rect 252700 8920 254700 16920
tri 254700 13385 259198 18058 nw
tri 296500 17506 297914 18920 se
rect 297914 17506 312800 18920
tri 352435 18641 352714 18920 se
rect 352714 18641 362800 18920
rect 296500 17062 312800 17506
rect 296500 16920 308500 17062
rect 242700 8334 254700 8920
tri 242700 7990 243044 8334 ne
rect 243044 7990 254148 8334
tri 188968 6920 189314 7266 ne
rect 189314 6920 198486 7266
tri 198486 6920 198832 7266 nw
tri 243044 7264 243770 7990 ne
rect 243770 7782 254148 7990
tri 254148 7782 254700 8334 nw
rect 296500 8920 298500 16920
tri 298500 15860 299560 16920 nw
tri 305440 15860 306500 16920 ne
tri 298500 8920 299560 9980 sw
tri 305440 8920 306500 9980 se
rect 306500 8920 308500 16920
tri 308500 13048 312800 17062 nw
tri 351300 17506 352435 18641 se
rect 352435 18298 362800 18641
rect 352435 18079 362744 18298
tri 362744 18080 362800 18298 nw
rect 404800 18921 412800 72800
rect 454800 25026 462800 85457
rect 504800 27380 512800 72800
rect 554800 32333 562800 90457
rect 604800 35305 612800 72800
tri 612800 35305 612991 35491 sw
tri 554800 30220 556591 32333 ne
rect 556591 30220 562800 32333
tri 562800 30220 567078 35267 sw
rect 604800 32109 612991 35305
tri 604800 30220 606745 32109 ne
rect 606745 30220 612991 32109
tri 612991 30220 618226 35305 sw
tri 462800 25026 462873 25125 sw
tri 504800 25026 506712 27380 ne
rect 506712 25026 512800 27380
tri 512800 25026 517019 30220 sw
tri 556591 25026 560993 30220 ne
rect 560993 25026 567078 30220
tri 567078 25026 571481 30220 sw
tri 606745 25026 612093 30220 ne
rect 612093 25026 618226 30220
tri 618226 25026 623575 30220 sw
rect 454800 22475 462873 25026
tri 454800 19846 456757 22475 ne
rect 456757 19846 462873 22475
tri 462873 19846 466730 25026 sw
tri 506712 19846 510920 25026 ne
rect 510920 19846 517019 25026
tri 517019 19846 521227 25026 sw
tri 560993 24828 561161 25026 ne
rect 561161 24828 571481 25026
tri 571481 24828 571649 25026 sw
tri 561161 22895 562800 24828 ne
rect 562800 24154 571649 24828
tri 571649 24154 572220 24828 sw
tri 612093 24154 612991 25026 ne
rect 612991 24154 623575 25026
tri 623575 24154 624473 25026 sw
rect 562800 22895 572220 24154
tri 562800 19846 565384 22895 ne
rect 565384 19846 572220 22895
tri 572220 19846 575872 24154 sw
tri 612991 19846 617426 24154 ne
rect 617426 19846 624473 24154
tri 624473 19846 628909 24154 sw
tri 412800 18921 413319 19846 sw
rect 404800 18920 413319 18921
tri 456757 18920 457446 19846 ne
rect 457446 18920 466730 19846
tri 466730 18920 467419 19846 sw
tri 510920 18920 511672 19846 ne
rect 511672 18920 521227 19846
tri 521227 18920 521979 19846 sw
tri 565384 18920 566169 19846 ne
rect 566169 18920 575872 19846
tri 575872 18920 576657 19846 sw
tri 617426 18920 618380 19846 ne
rect 618380 18920 628909 19846
tri 628909 18920 629862 19846 sw
rect 352435 18063 362741 18079
tri 362741 18067 362744 18079 nw
tri 362741 18063 362743 18065 sw
rect 352435 18062 362743 18063
tri 362743 18062 362744 18063 sw
rect 352435 18008 362744 18062
tri 362744 18008 362798 18062 sw
rect 404800 18060 416686 18920
tri 416686 18060 417546 18920 sw
tri 457446 18061 458086 18920 ne
rect 458086 18060 471486 18920
rect 352435 18006 362798 18008
tri 362798 18006 362800 18008 sw
rect 352435 17506 362800 18006
tri 362800 17506 363300 18006 sw
rect 351300 16920 363300 17506
rect 296500 8334 308500 8920
tri 296500 7987 296847 8334 ne
rect 296847 7987 307432 8334
rect 243770 7264 253630 7782
tri 253630 7264 254148 7782 nw
tri 296847 7266 297568 7987 ne
rect 297568 7266 307432 7987
tri 307432 7266 308500 8334 nw
rect 351300 8920 353300 16920
tri 353300 15860 354360 16920 nw
tri 360240 15860 361300 16920 ne
tri 353300 8920 354360 9980 sw
tri 360240 8920 361300 9980 se
rect 361300 8920 363300 16920
rect 404800 17754 417546 18060
tri 404800 15437 406100 17754 ne
rect 406100 17506 417546 17754
tri 417546 17506 418100 18060 sw
rect 406100 16920 418100 17506
rect 351300 8334 363300 8920
tri 351300 8055 351579 8334 ne
rect 351579 8055 363021 8334
tri 363021 8055 363300 8334 nw
rect 406100 8920 408100 16920
tri 408100 15860 409160 16920 nw
tri 415040 15860 416100 16920 ne
tri 408100 8920 409160 9980 sw
tri 415040 8920 416100 9980 se
rect 416100 8920 418100 16920
tri 458086 14281 460900 18060 ne
rect 460900 17909 471486 18060
tri 471486 17909 472497 18920 sw
tri 511672 18825 511749 18920 ne
rect 511749 18825 526286 18920
rect 460900 17506 472497 17909
tri 472497 17506 472900 17909 sw
tri 511749 17532 512800 18825 ne
rect 512800 17879 526286 18825
tri 526286 17879 527327 18920 sw
tri 566169 18655 566393 18920 ne
rect 566393 18655 581086 18920
tri 566393 17879 567051 18655 ne
rect 567051 17879 581086 18655
rect 512800 17532 527327 17879
rect 460900 16920 472900 17506
rect 406100 8334 418100 8920
tri 243770 6920 244114 7264 ne
rect 244114 6920 253286 7264
tri 253286 6920 253630 7264 nw
tri 297568 6920 297914 7266 ne
rect 297914 6920 307086 7266
tri 307086 6920 307432 7266 nw
tri 351579 6920 352714 8055 ne
rect 352714 6920 361886 8055
tri 361886 6920 363021 8055 nw
tri 406100 7474 406960 8334 ne
rect 406960 7780 417546 8334
tri 417546 7780 418100 8334 nw
rect 460900 8920 462900 16920
tri 462900 15860 463960 16920 nw
tri 469840 15860 470900 16920 ne
tri 462900 8920 463960 9980 sw
tri 469840 8920 470900 9980 se
rect 470900 8920 472900 16920
tri 512800 13961 515700 17532 ne
rect 515700 17506 527327 17532
tri 527327 17506 527700 17879 sw
rect 515700 16920 527700 17506
rect 460900 8334 472900 8920
rect 406960 7474 417240 7780
tri 417240 7474 417546 7780 nw
tri 406960 6920 407514 7474 ne
rect 407514 6920 416686 7474
tri 416686 6920 417240 7474 nw
tri 460900 6920 462314 8334 ne
rect 462314 7931 472497 8334
tri 472497 7931 472900 8334 nw
rect 515700 8920 517700 16920
tri 517700 15860 518760 16920 nw
tri 524640 15860 525700 16920 ne
tri 517700 8920 518760 9980 sw
tri 524640 8920 525700 9980 se
rect 525700 8920 527700 16920
tri 567051 13810 570500 17879 ne
rect 570500 17868 581086 17879
tri 581086 17868 582138 18920 sw
rect 570500 17506 582138 17868
tri 582138 17506 582500 17868 sw
tri 618380 17679 619658 18920 ne
rect 619658 17850 634886 18920
tri 634886 17850 635956 18920 sw
rect 619658 17679 635956 17850
rect 570500 16920 582500 17506
rect 515700 8334 527700 8920
rect 462314 7323 471889 7931
tri 471889 7323 472497 7931 nw
rect 462314 6920 471486 7323
tri 471486 6920 471889 7323 nw
tri 515700 7293 516741 8334 ne
rect 516741 7961 527327 8334
tri 527327 7961 527700 8334 nw
rect 570500 8920 572500 16920
tri 572500 15860 573560 16920 nw
tri 579440 15860 580500 16920 ne
tri 572500 8920 573560 9980 sw
tri 579440 8920 580500 9980 se
rect 580500 8920 582500 16920
tri 619658 13171 624300 17679 ne
rect 624300 17506 635956 17679
tri 635956 17506 636300 17850 sw
rect 624300 16920 636300 17506
rect 570500 8334 582500 8920
rect 516741 7293 526659 7961
tri 526659 7293 527327 7961 nw
tri 516741 6920 517114 7293 ne
rect 517114 6920 526286 7293
tri 526286 6920 526659 7293 nw
tri 570500 7282 571552 8334 ne
rect 571552 7972 582138 8334
tri 582138 7972 582500 8334 nw
rect 624300 8920 626300 16920
tri 626300 15860 627360 16920 nw
tri 633240 15860 634300 16920 ne
tri 626300 8920 627360 9980 sw
tri 633240 8920 634300 9980 se
rect 634300 8920 636300 16920
rect 624300 8334 636300 8920
tri 624300 8161 624473 8334 ne
rect 624473 8161 635956 8334
rect 571552 7282 581448 7972
tri 581448 7282 582138 7972 nw
tri 571552 6920 571914 7282 ne
rect 571914 6920 581086 7282
tri 581086 6920 581448 7282 nw
tri 624473 7264 625370 8161 ne
rect 625370 7990 635956 8161
tri 635956 7990 636300 8334 nw
rect 625370 7264 635230 7990
tri 635230 7264 635956 7990 nw
tri 625370 6920 625714 7264 ne
rect 625714 6920 634886 7264
tri 634886 6920 635230 7264 nw
use bump_bond0  bump_bond0_0
timestamp 1611856895
transform -1 0 108800 0 -1 68800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_0
timestamp 1611856895
transform -1 0 208800 0 -1 68800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_1
timestamp 1611856895
transform 0 1 308800 -1 0 68800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_2
timestamp 1611856895
transform 0 1 408800 -1 0 68800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_3
timestamp 1611856895
transform 0 1 508800 -1 0 68800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_4
timestamp 1611856895
transform 0 1 608800 -1 0 68800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_5
timestamp 1611856895
transform -1 0 108800 0 -1 168800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_9
timestamp 1611856895
transform -1 0 108800 0 -1 268800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_1
timestamp 1611856895
transform 0 -1 208800 1 0 168800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_3
timestamp 1611856895
transform 0 -1 208800 1 0 268800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_2
timestamp 1611856895
transform -1 0 308800 0 -1 168800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_4
timestamp 1611856895
transform 0 -1 308800 1 0 268800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_6
timestamp 1611856895
transform 0 1 408800 -1 0 168800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_10
timestamp 1611856895
transform 0 1 408800 -1 0 268800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_7
timestamp 1611856895
transform 1 0 508800 0 1 168800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_5
timestamp 1611856895
transform 0 1 508800 -1 0 268800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_11
timestamp 1611856895
transform 1 0 608800 0 1 268800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_8
timestamp 1611856895
transform 1 0 608800 0 1 168800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_10
timestamp 1611856895
transform 0 -1 108800 1 0 468800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_12
timestamp 1611856895
transform -1 0 108800 0 -1 368800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_11
timestamp 1611856895
transform 0 -1 208800 1 0 468800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_6
timestamp 1611856895
transform 0 -1 208800 1 0 368800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_14
timestamp 1611856895
transform 1 0 308800 0 1 468800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_7
timestamp 1611856895
transform 0 -1 308800 1 0 368800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_32
timestamp 1611856895
transform -1 0 508800 0 -1 468800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_15
timestamp 1611856895
transform -1 0 408800 0 -1 468800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_8
timestamp 1611856895
transform 0 1 408800 -1 0 368800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_12
timestamp 1611856895
transform 0 1 508800 -1 0 468800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_9
timestamp 1611856895
transform 0 1 508800 -1 0 368800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_16
timestamp 1611856895
transform 1 0 608800 0 1 468800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_13
timestamp 1611856895
transform 1 0 608800 0 1 368800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_21
timestamp 1611856895
transform -1 0 108800 0 -1 668800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_17
timestamp 1611856895
transform -1 0 108800 0 -1 568800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_22
timestamp 1611856895
transform -1 0 308800 0 -1 668800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_15
timestamp 1611856895
transform 0 -1 208800 1 0 668800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_18
timestamp 1611856895
transform 1 0 308800 0 1 568800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_13
timestamp 1611856895
transform 0 -1 208800 1 0 568800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_17
timestamp 1611856895
transform 0 1 508800 -1 0 668800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_16
timestamp 1611856895
transform 0 1 408800 -1 0 668800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_14
timestamp 1611856895
transform 0 1 508800 -1 0 568800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_19
timestamp 1611856895
transform -1 0 408800 0 -1 568800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_23
timestamp 1611856895
transform 1 0 608800 0 1 668800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_20
timestamp 1611856895
transform 1 0 608800 0 1 568800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_21
timestamp 1611856895
transform 0 -1 108800 1 0 868800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_25
timestamp 1611856895
transform -1 0 208800 0 -1 768800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_24
timestamp 1611856895
transform -1 0 108800 0 -1 768800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_23
timestamp 1611856895
transform 0 -1 308800 1 0 868800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_22
timestamp 1611856895
transform 0 -1 208800 1 0 868800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_18
timestamp 1611856895
transform 0 -1 308800 1 0 768800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_25
timestamp 1611856895
transform 1 0 508800 0 1 868800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_24
timestamp 1611856895
transform 1 0 408800 0 1 868800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_20
timestamp 1611856895
transform 0 1 508800 -1 0 768800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_19
timestamp 1611856895
transform 1 0 408800 0 1 768800
box -27000 -27000 27000 27000
use bump_bond45  bump_bond45_26
timestamp 1611856895
transform 1 0 608800 0 1 868800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_26
timestamp 1611856895
transform 1 0 608800 0 1 768800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_27
timestamp 1611856895
transform 0 -1 108800 1 0 968800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_29
timestamp 1611856895
transform 0 -1 308800 1 0 968800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_28
timestamp 1611856895
transform 0 -1 208800 1 0 968800
box -26897 -26897 38184 26897
use bump_bond45  bump_bond45_27
timestamp 1611856895
transform 1 0 508800 0 1 968800
box -27000 -27000 27000 27000
use bump_bond0  bump_bond0_30
timestamp 1611856895
transform 0 -1 408800 1 0 968800
box -26897 -26897 38184 26897
use bump_bond0  bump_bond0_31
timestamp 1611856895
transform 0 -1 608800 1 0 968800
box -26897 -26897 38184 26897
<< end >>
