magic
tech sky130A
magscale 1 2
timestamp 1625156099
<< metal1 >>
rect 80560 1002267 80566 1002319
rect 80618 1002307 80624 1002319
rect 82288 1002307 82294 1002319
rect 80618 1002279 82294 1002307
rect 80618 1002267 80624 1002279
rect 82288 1002267 82294 1002279
rect 82346 1002267 82352 1002319
rect 483664 1002267 483670 1002319
rect 483722 1002307 483728 1002319
rect 486736 1002307 486742 1002319
rect 483722 1002279 486742 1002307
rect 483722 1002267 483728 1002279
rect 486736 1002267 486742 1002279
rect 486794 1002267 486800 1002319
rect 535696 991463 535702 991515
rect 535754 991503 535760 991515
rect 538576 991503 538582 991515
rect 535754 991475 538582 991503
rect 535754 991463 535760 991475
rect 538576 991463 538582 991475
rect 538634 991463 538640 991515
rect 388624 990723 388630 990775
rect 388682 990763 388688 990775
rect 389584 990763 389590 990775
rect 388682 990735 389590 990763
rect 388682 990723 388688 990735
rect 389584 990723 389590 990735
rect 389642 990723 389648 990775
rect 240880 982953 240886 983005
rect 240938 982993 240944 983005
rect 241936 982993 241942 983005
rect 240938 982965 241942 982993
rect 240938 982953 240944 982965
rect 241936 982953 241942 982965
rect 241994 982953 242000 983005
rect 292528 982953 292534 983005
rect 292586 982993 292592 983005
rect 296656 982993 296662 983005
rect 292586 982965 296662 982993
rect 292586 982953 292592 982965
rect 296656 982953 296662 982965
rect 296714 982953 296720 983005
rect 40144 961863 40150 961915
rect 40202 961903 40208 961915
rect 60016 961903 60022 961915
rect 40202 961875 60022 961903
rect 40202 961863 40208 961875
rect 60016 961863 60022 961875
rect 60074 961863 60080 961915
rect 653776 960457 653782 960509
rect 653834 960497 653840 960509
rect 679696 960497 679702 960509
rect 653834 960469 679702 960497
rect 653834 960457 653840 960469
rect 679696 960457 679702 960469
rect 679754 960457 679760 960509
rect 655408 892969 655414 893021
rect 655466 893009 655472 893021
rect 676240 893009 676246 893021
rect 655466 892981 676246 893009
rect 655466 892969 655472 892981
rect 676240 892969 676246 892981
rect 676298 892969 676304 893021
rect 655216 892895 655222 892947
rect 655274 892935 655280 892947
rect 676144 892935 676150 892947
rect 655274 892907 676150 892935
rect 655274 892895 655280 892907
rect 676144 892895 676150 892907
rect 676202 892895 676208 892947
rect 655120 892821 655126 892873
rect 655178 892861 655184 892873
rect 676048 892861 676054 892873
rect 655178 892833 676054 892861
rect 655178 892821 655184 892833
rect 676048 892821 676054 892833
rect 676106 892821 676112 892873
rect 673360 892377 673366 892429
rect 673418 892417 673424 892429
rect 676048 892417 676054 892429
rect 673418 892389 676054 892417
rect 673418 892377 673424 892389
rect 676048 892377 676054 892389
rect 676106 892377 676112 892429
rect 670960 891415 670966 891467
rect 671018 891455 671024 891467
rect 676048 891455 676054 891467
rect 671018 891427 676054 891455
rect 671018 891415 671024 891427
rect 676048 891415 676054 891427
rect 676106 891415 676112 891467
rect 670864 890379 670870 890431
rect 670922 890419 670928 890431
rect 676048 890419 676054 890431
rect 670922 890391 676054 890419
rect 670922 890379 670928 890391
rect 676048 890379 676054 890391
rect 676106 890379 676112 890431
rect 674224 887493 674230 887545
rect 674282 887533 674288 887545
rect 676048 887533 676054 887545
rect 674282 887505 676054 887533
rect 674282 887493 674288 887505
rect 676048 887493 676054 887505
rect 676106 887493 676112 887545
rect 675088 887123 675094 887175
rect 675146 887163 675152 887175
rect 676240 887163 676246 887175
rect 675146 887135 676246 887163
rect 675146 887123 675152 887135
rect 676240 887123 676246 887135
rect 676298 887123 676304 887175
rect 675184 887049 675190 887101
rect 675242 887089 675248 887101
rect 676048 887089 676054 887101
rect 675242 887061 676054 887089
rect 675242 887049 675248 887061
rect 676048 887049 676054 887061
rect 676106 887049 676112 887101
rect 674032 885051 674038 885103
rect 674090 885091 674096 885103
rect 676048 885091 676054 885103
rect 674090 885063 676054 885091
rect 674090 885051 674096 885063
rect 676048 885051 676054 885063
rect 676106 885051 676112 885103
rect 674896 884385 674902 884437
rect 674954 884425 674960 884437
rect 676048 884425 676054 884437
rect 674954 884397 676054 884425
rect 674954 884385 674960 884397
rect 676048 884385 676054 884397
rect 676106 884385 676112 884437
rect 674896 884163 674902 884215
rect 674954 884203 674960 884215
rect 676240 884203 676246 884215
rect 674954 884175 676246 884203
rect 674954 884163 674960 884175
rect 676240 884163 676246 884175
rect 676298 884163 676304 884215
rect 674608 883571 674614 883623
rect 674666 883611 674672 883623
rect 676048 883611 676054 883623
rect 674666 883583 676054 883611
rect 674666 883571 674672 883583
rect 676048 883571 676054 883583
rect 676106 883571 676112 883623
rect 675280 882831 675286 882883
rect 675338 882871 675344 882883
rect 679696 882871 679702 882883
rect 675338 882843 679702 882871
rect 675338 882831 675344 882843
rect 679696 882831 679702 882843
rect 679754 882831 679760 882883
rect 675760 882239 675766 882291
rect 675818 882279 675824 882291
rect 680080 882279 680086 882291
rect 675818 882251 680086 882279
rect 675818 882239 675824 882251
rect 680080 882239 680086 882251
rect 680138 882239 680144 882291
rect 674416 881943 674422 881995
rect 674474 881983 674480 881995
rect 676048 881983 676054 881995
rect 674474 881955 676054 881983
rect 674474 881943 674480 881955
rect 676048 881943 676054 881955
rect 676106 881943 676112 881995
rect 674320 881647 674326 881699
rect 674378 881687 674384 881699
rect 680272 881687 680278 881699
rect 674378 881659 680278 881687
rect 674378 881647 674384 881659
rect 680272 881647 680278 881659
rect 680330 881647 680336 881699
rect 649456 881425 649462 881477
rect 649514 881465 649520 881477
rect 679792 881465 679798 881477
rect 649514 881437 679798 881465
rect 649514 881425 649520 881437
rect 679792 881425 679798 881437
rect 679850 881425 679856 881477
rect 655312 881351 655318 881403
rect 655370 881391 655376 881403
rect 675472 881391 675478 881403
rect 655370 881363 675478 881391
rect 655370 881351 655376 881363
rect 675472 881351 675478 881363
rect 675530 881351 675536 881403
rect 674128 880981 674134 881033
rect 674186 881021 674192 881033
rect 674416 881021 674422 881033
rect 674186 880993 674422 881021
rect 674186 880981 674192 880993
rect 674416 880981 674422 880993
rect 674474 880981 674480 881033
rect 674416 880833 674422 880885
rect 674474 880873 674480 880885
rect 675088 880873 675094 880885
rect 674474 880845 675094 880873
rect 674474 880833 674480 880845
rect 675088 880833 675094 880845
rect 675146 880833 675152 880885
rect 675088 880685 675094 880737
rect 675146 880725 675152 880737
rect 680176 880725 680182 880737
rect 675146 880697 680182 880725
rect 675146 880685 675152 880697
rect 680176 880685 680182 880697
rect 680234 880685 680240 880737
rect 674992 879501 674998 879553
rect 675050 879541 675056 879553
rect 679984 879541 679990 879553
rect 675050 879513 679990 879541
rect 675050 879501 675056 879513
rect 679984 879501 679990 879513
rect 680042 879501 680048 879553
rect 674512 878613 674518 878665
rect 674570 878653 674576 878665
rect 675184 878653 675190 878665
rect 674570 878625 675190 878653
rect 674570 878613 674576 878625
rect 675184 878613 675190 878625
rect 675242 878613 675248 878665
rect 675184 878465 675190 878517
rect 675242 878505 675248 878517
rect 679888 878505 679894 878517
rect 675242 878477 679894 878505
rect 675242 878465 675248 878477
rect 679888 878465 679894 878477
rect 679946 878465 679952 878517
rect 675760 878317 675766 878369
rect 675818 878317 675824 878369
rect 675778 877851 675806 878317
rect 675760 877799 675766 877851
rect 675818 877799 675824 877851
rect 674320 876689 674326 876741
rect 674378 876729 674384 876741
rect 675280 876729 675286 876741
rect 674378 876701 675286 876729
rect 674378 876689 674384 876701
rect 675280 876689 675286 876701
rect 675338 876689 675344 876741
rect 675088 874913 675094 874965
rect 675146 874953 675152 874965
rect 675472 874953 675478 874965
rect 675146 874925 675478 874953
rect 675146 874913 675152 874925
rect 675472 874913 675478 874925
rect 675530 874913 675536 874965
rect 675184 874247 675190 874299
rect 675242 874287 675248 874299
rect 675472 874287 675478 874299
rect 675242 874259 675478 874287
rect 675242 874247 675248 874259
rect 675472 874247 675478 874259
rect 675530 874247 675536 874299
rect 674992 873507 674998 873559
rect 675050 873547 675056 873559
rect 675376 873547 675382 873559
rect 675050 873519 675382 873547
rect 675050 873507 675056 873519
rect 675376 873507 675382 873519
rect 675434 873507 675440 873559
rect 674896 872915 674902 872967
rect 674954 872955 674960 872967
rect 675376 872955 675382 872967
rect 674954 872927 675382 872955
rect 674954 872915 674960 872927
rect 675376 872915 675382 872927
rect 675434 872915 675440 872967
rect 674032 872693 674038 872745
rect 674090 872733 674096 872745
rect 674896 872733 674902 872745
rect 674090 872705 674902 872733
rect 674090 872693 674096 872705
rect 674896 872693 674902 872705
rect 674954 872693 674960 872745
rect 654160 872619 654166 872671
rect 654218 872659 654224 872671
rect 675088 872659 675094 872671
rect 654218 872631 675094 872659
rect 654218 872619 654224 872631
rect 675088 872619 675094 872631
rect 675146 872619 675152 872671
rect 674224 870547 674230 870599
rect 674282 870587 674288 870599
rect 675472 870587 675478 870599
rect 674282 870559 675478 870587
rect 674282 870547 674288 870559
rect 675472 870547 675478 870559
rect 675530 870547 675536 870599
rect 674608 869955 674614 870007
rect 674666 869995 674672 870007
rect 675376 869995 675382 870007
rect 674666 869967 675382 869995
rect 674666 869955 674672 869967
rect 675376 869955 675382 869967
rect 675434 869955 675440 870007
rect 674512 869733 674518 869785
rect 674570 869773 674576 869785
rect 674992 869773 674998 869785
rect 674570 869745 674998 869773
rect 674570 869733 674576 869745
rect 674992 869733 674998 869745
rect 675050 869733 675056 869785
rect 674128 868771 674134 868823
rect 674186 868811 674192 868823
rect 675184 868811 675190 868823
rect 674186 868783 675190 868811
rect 674186 868771 674192 868783
rect 675184 868771 675190 868783
rect 675242 868771 675248 868823
rect 674896 867365 674902 867417
rect 674954 867405 674960 867417
rect 675472 867405 675478 867417
rect 674954 867377 675478 867405
rect 674954 867365 674960 867377
rect 675472 867365 675478 867377
rect 675530 867365 675536 867417
rect 674416 865737 674422 865789
rect 674474 865777 674480 865789
rect 675184 865777 675190 865789
rect 674474 865749 675190 865777
rect 674474 865737 674480 865749
rect 675184 865737 675190 865749
rect 675242 865737 675248 865789
rect 653776 863961 653782 864013
rect 653834 864001 653840 864013
rect 675088 864001 675094 864013
rect 653834 863973 675094 864001
rect 653834 863961 653840 863973
rect 675088 863961 675094 863973
rect 675146 863961 675152 864013
rect 41776 816601 41782 816653
rect 41834 816641 41840 816653
rect 47440 816641 47446 816653
rect 41834 816613 47446 816641
rect 41834 816601 41840 816613
rect 47440 816601 47446 816613
rect 47498 816601 47504 816653
rect 41776 816083 41782 816135
rect 41834 816123 41840 816135
rect 44848 816123 44854 816135
rect 41834 816095 44854 816123
rect 41834 816083 41840 816095
rect 44848 816083 44854 816095
rect 44906 816083 44912 816135
rect 41584 815343 41590 815395
rect 41642 815383 41648 815395
rect 44944 815383 44950 815395
rect 41642 815355 44950 815383
rect 41642 815343 41648 815355
rect 44944 815343 44950 815355
rect 45002 815343 45008 815395
rect 41776 814603 41782 814655
rect 41834 814643 41840 814655
rect 43216 814643 43222 814655
rect 41834 814615 43222 814643
rect 41834 814603 41840 814615
rect 43216 814603 43222 814615
rect 43274 814603 43280 814655
rect 41584 813419 41590 813471
rect 41642 813459 41648 813471
rect 44656 813459 44662 813471
rect 41642 813431 44662 813459
rect 41642 813419 41648 813431
rect 44656 813419 44662 813431
rect 44714 813419 44720 813471
rect 41776 812531 41782 812583
rect 41834 812571 41840 812583
rect 44752 812571 44758 812583
rect 41834 812543 44758 812571
rect 41834 812531 41840 812543
rect 44752 812531 44758 812543
rect 44810 812531 44816 812583
rect 41584 810089 41590 810141
rect 41642 810129 41648 810141
rect 42736 810129 42742 810141
rect 41642 810101 42742 810129
rect 41642 810089 41648 810101
rect 42736 810089 42742 810101
rect 42794 810089 42800 810141
rect 41584 808387 41590 808439
rect 41642 808427 41648 808439
rect 42832 808427 42838 808439
rect 41642 808399 42838 808427
rect 41642 808387 41648 808399
rect 42832 808387 42838 808399
rect 42890 808387 42896 808439
rect 41776 807203 41782 807255
rect 41834 807243 41840 807255
rect 43024 807243 43030 807255
rect 41834 807215 43030 807243
rect 41834 807203 41840 807215
rect 43024 807203 43030 807215
rect 43082 807203 43088 807255
rect 41584 806907 41590 806959
rect 41642 806947 41648 806959
rect 42640 806947 42646 806959
rect 41642 806919 42646 806947
rect 41642 806907 41648 806919
rect 42640 806907 42646 806919
rect 42698 806907 42704 806959
rect 41776 803799 41782 803851
rect 41834 803839 41840 803851
rect 43120 803839 43126 803851
rect 41834 803811 43126 803839
rect 41834 803799 41840 803811
rect 43120 803799 43126 803811
rect 43178 803799 43184 803851
rect 41488 803725 41494 803777
rect 41546 803765 41552 803777
rect 44560 803765 44566 803777
rect 41546 803737 44566 803765
rect 41546 803725 41552 803737
rect 44560 803725 44566 803737
rect 44618 803725 44624 803777
rect 41584 803651 41590 803703
rect 41642 803691 41648 803703
rect 42928 803691 42934 803703
rect 41642 803663 42934 803691
rect 41642 803651 41648 803663
rect 42928 803651 42934 803663
rect 42986 803651 42992 803703
rect 42736 800839 42742 800891
rect 42794 800879 42800 800891
rect 43504 800879 43510 800891
rect 42794 800851 43510 800879
rect 42794 800839 42800 800851
rect 43504 800839 43510 800851
rect 43562 800839 43568 800891
rect 42832 800765 42838 800817
rect 42890 800805 42896 800817
rect 43408 800805 43414 800817
rect 42890 800777 43414 800805
rect 42890 800765 42896 800777
rect 43408 800765 43414 800777
rect 43466 800765 43472 800817
rect 42736 800691 42742 800743
rect 42794 800731 42800 800743
rect 57712 800731 57718 800743
rect 42794 800703 57718 800731
rect 42794 800691 42800 800703
rect 57712 800691 57718 800703
rect 57770 800691 57776 800743
rect 42832 800617 42838 800669
rect 42890 800657 42896 800669
rect 57616 800657 57622 800669
rect 42890 800629 57622 800657
rect 42890 800617 42896 800629
rect 57616 800617 57622 800629
rect 57674 800617 57680 800669
rect 41392 800469 41398 800521
rect 41450 800509 41456 800521
rect 43696 800509 43702 800521
rect 41450 800481 43702 800509
rect 41450 800469 41456 800481
rect 43696 800469 43702 800481
rect 43754 800469 43760 800521
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 42064 800173 42070 800225
rect 42122 800213 42128 800225
rect 43312 800213 43318 800225
rect 42122 800185 43318 800213
rect 42122 800173 42128 800185
rect 43312 800173 43318 800185
rect 43370 800173 43376 800225
rect 41890 800003 41918 800173
rect 41872 799951 41878 800003
rect 41930 799951 41936 800003
rect 42640 797879 42646 797931
rect 42698 797919 42704 797931
rect 42698 797891 42878 797919
rect 42698 797879 42704 797891
rect 42064 797435 42070 797487
rect 42122 797475 42128 797487
rect 42736 797475 42742 797487
rect 42122 797447 42742 797475
rect 42122 797435 42128 797447
rect 42736 797435 42742 797447
rect 42794 797435 42800 797487
rect 42850 797401 42878 797891
rect 42754 797373 42878 797401
rect 42754 797339 42782 797373
rect 42736 797287 42742 797339
rect 42794 797287 42800 797339
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 43024 796291 43030 796303
rect 42218 796263 43030 796291
rect 42218 796251 42224 796263
rect 43024 796251 43030 796263
rect 43082 796251 43088 796303
rect 43024 796103 43030 796155
rect 43082 796143 43088 796155
rect 43312 796143 43318 796155
rect 43082 796115 43318 796143
rect 43082 796103 43088 796115
rect 43312 796103 43318 796115
rect 43370 796103 43376 796155
rect 42064 795585 42070 795637
rect 42122 795625 42128 795637
rect 42832 795625 42838 795637
rect 42122 795597 42838 795625
rect 42122 795585 42128 795597
rect 42832 795585 42838 795597
rect 42890 795585 42896 795637
rect 42160 794771 42166 794823
rect 42218 794811 42224 794823
rect 42928 794811 42934 794823
rect 42218 794783 42934 794811
rect 42218 794771 42224 794783
rect 42928 794771 42934 794783
rect 42986 794771 42992 794823
rect 42928 794623 42934 794675
rect 42986 794663 42992 794675
rect 43408 794663 43414 794675
rect 42986 794635 43414 794663
rect 42986 794623 42992 794635
rect 43408 794623 43414 794635
rect 43466 794623 43472 794675
rect 42064 794253 42070 794305
rect 42122 794293 42128 794305
rect 42736 794293 42742 794305
rect 42122 794265 42742 794293
rect 42122 794253 42128 794265
rect 42736 794253 42742 794265
rect 42794 794253 42800 794305
rect 42160 793809 42166 793861
rect 42218 793849 42224 793861
rect 43120 793849 43126 793861
rect 42218 793821 43126 793849
rect 42218 793809 42224 793821
rect 43120 793809 43126 793821
rect 43178 793809 43184 793861
rect 43120 793661 43126 793713
rect 43178 793701 43184 793713
rect 43504 793701 43510 793713
rect 43178 793673 43510 793701
rect 43178 793661 43184 793673
rect 43504 793661 43510 793673
rect 43562 793661 43568 793713
rect 42256 792107 42262 792159
rect 42314 792147 42320 792159
rect 43024 792147 43030 792159
rect 42314 792119 43030 792147
rect 42314 792107 42320 792119
rect 43024 792107 43030 792119
rect 43082 792107 43088 792159
rect 655216 792033 655222 792085
rect 655274 792073 655280 792085
rect 675376 792073 675382 792085
rect 655274 792045 675382 792073
rect 655274 792033 655280 792045
rect 675376 792033 675382 792045
rect 675434 792033 675440 792085
rect 42256 790109 42262 790161
rect 42314 790149 42320 790161
rect 43120 790149 43126 790161
rect 42314 790121 43126 790149
rect 42314 790109 42320 790121
rect 43120 790109 43126 790121
rect 43178 790109 43184 790161
rect 43120 789961 43126 790013
rect 43178 790001 43184 790013
rect 43696 790001 43702 790013
rect 43178 789973 43702 790001
rect 43178 789961 43184 789973
rect 43696 789961 43702 789973
rect 43754 789961 43760 790013
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 42736 789927 42742 789939
rect 42218 789899 42742 789927
rect 42218 789887 42224 789899
rect 42736 789887 42742 789899
rect 42794 789887 42800 789939
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 43024 789483 43030 789495
rect 42218 789455 43030 789483
rect 42218 789443 42224 789455
rect 43024 789443 43030 789455
rect 43082 789443 43088 789495
rect 42736 789147 42742 789199
rect 42794 789187 42800 789199
rect 58192 789187 58198 789199
rect 42794 789159 58198 789187
rect 42794 789147 42800 789159
rect 58192 789147 58198 789159
rect 58250 789147 58256 789199
rect 44944 789073 44950 789125
rect 45002 789113 45008 789125
rect 58384 789113 58390 789125
rect 45002 789085 58390 789113
rect 45002 789073 45008 789085
rect 58384 789073 58390 789085
rect 58442 789073 58448 789125
rect 42160 786853 42166 786905
rect 42218 786893 42224 786905
rect 43120 786893 43126 786905
rect 42218 786865 43126 786893
rect 42218 786853 42224 786865
rect 43120 786853 43126 786865
rect 43178 786853 43184 786905
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42832 786449 42838 786461
rect 42218 786421 42838 786449
rect 42218 786409 42224 786421
rect 42832 786409 42838 786421
rect 42890 786409 42896 786461
rect 42064 785595 42070 785647
rect 42122 785635 42128 785647
rect 42928 785635 42934 785647
rect 42122 785607 42934 785635
rect 42122 785595 42128 785607
rect 42928 785595 42934 785607
rect 42986 785595 42992 785647
rect 44848 785521 44854 785573
rect 44906 785561 44912 785573
rect 59152 785561 59158 785573
rect 44906 785533 59158 785561
rect 44906 785521 44912 785533
rect 59152 785521 59158 785533
rect 59210 785521 59216 785573
rect 47440 785373 47446 785425
rect 47498 785413 47504 785425
rect 59632 785413 59638 785425
rect 47498 785385 59638 785413
rect 47498 785373 47504 785385
rect 59632 785373 59638 785385
rect 59690 785373 59696 785425
rect 42160 785151 42166 785203
rect 42218 785191 42224 785203
rect 42736 785191 42742 785203
rect 42218 785163 42742 785191
rect 42218 785151 42224 785163
rect 42736 785151 42742 785163
rect 42794 785151 42800 785203
rect 655024 783449 655030 783501
rect 655082 783489 655088 783501
rect 674992 783489 674998 783501
rect 655082 783461 674998 783489
rect 655082 783449 655088 783461
rect 674992 783449 674998 783461
rect 675050 783449 675056 783501
rect 673264 782931 673270 782983
rect 673322 782971 673328 782983
rect 675376 782971 675382 782983
rect 673322 782943 675382 782971
rect 673322 782931 673328 782943
rect 675376 782931 675382 782943
rect 675434 782931 675440 782983
rect 654352 780489 654358 780541
rect 654410 780529 654416 780541
rect 675280 780529 675286 780541
rect 654410 780501 675286 780529
rect 654410 780489 654416 780501
rect 675280 780489 675286 780501
rect 675338 780489 675344 780541
rect 674992 778861 674998 778913
rect 675050 778901 675056 778913
rect 675376 778901 675382 778913
rect 675050 778873 675382 778901
rect 675050 778861 675056 778873
rect 675376 778861 675382 778873
rect 675434 778861 675440 778913
rect 673168 778713 673174 778765
rect 673226 778753 673232 778765
rect 675472 778753 675478 778765
rect 673226 778725 675478 778753
rect 673226 778713 673232 778725
rect 675472 778713 675478 778725
rect 675530 778713 675536 778765
rect 674608 773607 674614 773659
rect 674666 773647 674672 773659
rect 675280 773647 675286 773659
rect 674666 773619 675286 773647
rect 674666 773607 674672 773619
rect 675280 773607 675286 773619
rect 675338 773607 675344 773659
rect 41776 773459 41782 773511
rect 41834 773499 41840 773511
rect 47440 773499 47446 773511
rect 41834 773471 47446 773499
rect 41834 773459 41840 773471
rect 47440 773459 47446 773471
rect 47498 773459 47504 773511
rect 41776 772867 41782 772919
rect 41834 772907 41840 772919
rect 44944 772907 44950 772919
rect 41834 772879 44950 772907
rect 41834 772867 41840 772879
rect 44944 772867 44950 772879
rect 45002 772867 45008 772919
rect 41776 772275 41782 772327
rect 41834 772315 41840 772327
rect 45040 772315 45046 772327
rect 41834 772287 45046 772315
rect 41834 772275 41840 772287
rect 45040 772275 45046 772287
rect 45098 772275 45104 772327
rect 41584 772127 41590 772179
rect 41642 772167 41648 772179
rect 61840 772167 61846 772179
rect 41642 772139 61846 772167
rect 41642 772127 41648 772139
rect 61840 772127 61846 772139
rect 61898 772127 61904 772179
rect 41776 771979 41782 772031
rect 41834 772019 41840 772031
rect 43216 772019 43222 772031
rect 41834 771991 43222 772019
rect 41834 771979 41840 771991
rect 43216 771979 43222 771991
rect 43274 771979 43280 772031
rect 41488 771905 41494 771957
rect 41546 771945 41552 771957
rect 62032 771945 62038 771957
rect 41546 771917 62038 771945
rect 41546 771905 41552 771917
rect 62032 771905 62038 771917
rect 62090 771905 62096 771957
rect 41776 771387 41782 771439
rect 41834 771427 41840 771439
rect 43216 771427 43222 771439
rect 41834 771399 43222 771427
rect 41834 771387 41840 771399
rect 43216 771387 43222 771399
rect 43274 771387 43280 771439
rect 41584 767391 41590 767443
rect 41642 767431 41648 767443
rect 43024 767431 43030 767443
rect 41642 767403 43030 767431
rect 41642 767391 41648 767403
rect 43024 767391 43030 767403
rect 43082 767391 43088 767443
rect 41584 766281 41590 766333
rect 41642 766321 41648 766333
rect 42928 766321 42934 766333
rect 41642 766293 42934 766321
rect 41642 766281 41648 766293
rect 42928 766281 42934 766293
rect 42986 766281 42992 766333
rect 41776 765393 41782 765445
rect 41834 765433 41840 765445
rect 43120 765433 43126 765445
rect 41834 765405 43126 765433
rect 41834 765393 41840 765405
rect 43120 765393 43126 765405
rect 43178 765393 43184 765445
rect 41776 763395 41782 763447
rect 41834 763435 41840 763447
rect 42832 763435 42838 763447
rect 41834 763407 42838 763435
rect 41834 763395 41840 763407
rect 42832 763395 42838 763407
rect 42890 763395 42896 763447
rect 41584 760731 41590 760783
rect 41642 760771 41648 760783
rect 44848 760771 44854 760783
rect 41642 760743 44854 760771
rect 41642 760731 41648 760743
rect 44848 760731 44854 760743
rect 44906 760731 44912 760783
rect 42832 757475 42838 757527
rect 42890 757515 42896 757527
rect 58672 757515 58678 757527
rect 42890 757487 58678 757515
rect 42890 757475 42896 757487
rect 58672 757475 58678 757487
rect 58730 757475 58736 757527
rect 41296 757401 41302 757453
rect 41354 757441 41360 757453
rect 43408 757441 43414 757453
rect 41354 757413 43414 757441
rect 41354 757401 41360 757413
rect 43408 757401 43414 757413
rect 43466 757401 43472 757453
rect 40336 757327 40342 757379
rect 40394 757367 40400 757379
rect 40394 757339 41438 757367
rect 40394 757327 40400 757339
rect 41410 756775 41438 757339
rect 41680 757327 41686 757379
rect 41738 757367 41744 757379
rect 42736 757367 42742 757379
rect 41738 757339 42742 757367
rect 41738 757327 41744 757339
rect 42736 757327 42742 757339
rect 42794 757327 42800 757379
rect 43024 757327 43030 757379
rect 43082 757367 43088 757379
rect 43600 757367 43606 757379
rect 43082 757339 43606 757367
rect 43082 757327 43088 757339
rect 43600 757327 43606 757339
rect 43658 757327 43664 757379
rect 42928 757253 42934 757305
rect 42986 757293 42992 757305
rect 43504 757293 43510 757305
rect 42986 757265 43510 757293
rect 42986 757253 42992 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 42160 757179 42166 757231
rect 42218 757219 42224 757231
rect 43312 757219 43318 757231
rect 42218 757191 43318 757219
rect 42218 757179 42224 757191
rect 43312 757179 43318 757191
rect 43370 757179 43376 757231
rect 42064 757105 42070 757157
rect 42122 757145 42128 757157
rect 43120 757145 43126 757157
rect 42122 757117 43126 757145
rect 42122 757105 42128 757117
rect 43120 757105 43126 757117
rect 43178 757105 43184 757157
rect 41776 757031 41782 757083
rect 41834 757071 41840 757083
rect 43024 757071 43030 757083
rect 41834 757043 43030 757071
rect 41834 757031 41840 757043
rect 43024 757031 43030 757043
rect 43082 757031 43088 757083
rect 41872 756957 41878 757009
rect 41930 756997 41936 757009
rect 42928 756997 42934 757009
rect 41930 756969 42934 756997
rect 41930 756957 41936 756969
rect 42928 756957 42934 756969
rect 42986 756957 42992 757009
rect 41776 756775 41782 756787
rect 41410 756747 41782 756775
rect 41776 756735 41782 756747
rect 41834 756735 41840 756787
rect 42064 754885 42070 754937
rect 42122 754925 42128 754937
rect 42736 754925 42742 754937
rect 42122 754897 42742 754925
rect 42122 754885 42128 754897
rect 42736 754885 42742 754897
rect 42794 754885 42800 754937
rect 42160 754071 42166 754123
rect 42218 754111 42224 754123
rect 42832 754111 42838 754123
rect 42218 754083 42838 754111
rect 42218 754071 42224 754083
rect 42832 754071 42838 754083
rect 42890 754071 42896 754123
rect 42832 753923 42838 753975
rect 42890 753963 42896 753975
rect 43312 753963 43318 753975
rect 42890 753935 43318 753963
rect 42890 753923 42896 753935
rect 43312 753923 43318 753935
rect 43370 753923 43376 753975
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 42928 753075 42934 753087
rect 42122 753047 42934 753075
rect 42122 753035 42128 753047
rect 42928 753035 42934 753047
rect 42986 753035 42992 753087
rect 42928 752887 42934 752939
rect 42986 752927 42992 752939
rect 43408 752927 43414 752939
rect 42986 752899 43414 752927
rect 42986 752887 42992 752899
rect 43408 752887 43414 752899
rect 43466 752887 43472 752939
rect 42160 751999 42166 752051
rect 42218 752039 42224 752051
rect 43312 752039 43318 752051
rect 42218 752011 43318 752039
rect 42218 751999 42224 752011
rect 43312 751999 43318 752011
rect 43370 751999 43376 752051
rect 42064 751777 42070 751829
rect 42122 751817 42128 751829
rect 43024 751817 43030 751829
rect 42122 751789 43030 751817
rect 42122 751777 42128 751789
rect 43024 751777 43030 751789
rect 43082 751777 43088 751829
rect 42064 751111 42070 751163
rect 42122 751151 42128 751163
rect 43120 751151 43126 751163
rect 42122 751123 43126 751151
rect 42122 751111 42128 751123
rect 43120 751111 43126 751123
rect 43178 751111 43184 751163
rect 43120 750963 43126 751015
rect 43178 751003 43184 751015
rect 43504 751003 43510 751015
rect 43178 750975 43510 751003
rect 43178 750963 43184 750975
rect 43504 750963 43510 750975
rect 43562 750963 43568 751015
rect 42160 750593 42166 750645
rect 42218 750633 42224 750645
rect 42832 750633 42838 750645
rect 42218 750605 42838 750633
rect 42218 750593 42224 750605
rect 42832 750593 42838 750605
rect 42890 750593 42896 750645
rect 42064 749779 42070 749831
rect 42122 749819 42128 749831
rect 42736 749819 42742 749831
rect 42122 749791 42742 749819
rect 42122 749779 42128 749791
rect 42736 749779 42742 749791
rect 42794 749779 42800 749831
rect 655696 748817 655702 748869
rect 655754 748857 655760 748869
rect 675376 748857 675382 748869
rect 655754 748829 675382 748857
rect 655754 748817 655760 748829
rect 675376 748817 675382 748829
rect 675434 748817 675440 748869
rect 42160 747411 42166 747463
rect 42218 747451 42224 747463
rect 43120 747451 43126 747463
rect 42218 747423 43126 747451
rect 42218 747411 42224 747423
rect 43120 747411 43126 747423
rect 43178 747411 43184 747463
rect 42832 747263 42838 747315
rect 42890 747303 42896 747315
rect 43120 747303 43126 747315
rect 42890 747275 43126 747303
rect 42890 747263 42896 747275
rect 43120 747263 43126 747275
rect 43178 747263 43184 747315
rect 42160 746893 42166 746945
rect 42218 746933 42224 746945
rect 42928 746933 42934 746945
rect 42218 746905 42934 746933
rect 42218 746893 42224 746905
rect 42928 746893 42934 746905
rect 42986 746893 42992 746945
rect 42928 746745 42934 746797
rect 42986 746785 42992 746797
rect 43600 746785 43606 746797
rect 42986 746757 43606 746785
rect 42986 746745 42992 746757
rect 43600 746745 43606 746757
rect 43658 746745 43664 746797
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 43024 746119 43030 746131
rect 42122 746091 43030 746119
rect 42122 746079 42128 746091
rect 43024 746079 43030 746091
rect 43082 746079 43088 746131
rect 42352 745931 42358 745983
rect 42410 745971 42416 745983
rect 54640 745971 54646 745983
rect 42410 745943 54646 745971
rect 42410 745931 42416 745943
rect 54640 745931 54646 745943
rect 54698 745931 54704 745983
rect 54736 745931 54742 745983
rect 54794 745971 54800 745983
rect 57616 745971 57622 745983
rect 54794 745943 57622 745971
rect 54794 745931 54800 745943
rect 57616 745931 57622 745943
rect 57674 745931 57680 745983
rect 43312 745561 43318 745613
rect 43370 745601 43376 745613
rect 59632 745601 59638 745613
rect 43370 745573 59638 745601
rect 43370 745561 43376 745573
rect 59632 745561 59638 745573
rect 59690 745561 59696 745613
rect 42160 745487 42166 745539
rect 42218 745527 42224 745539
rect 42928 745527 42934 745539
rect 42218 745499 42934 745527
rect 42218 745487 42224 745499
rect 42928 745487 42934 745499
rect 42986 745487 42992 745539
rect 45040 745339 45046 745391
rect 45098 745379 45104 745391
rect 58480 745379 58486 745391
rect 45098 745351 58486 745379
rect 45098 745339 45104 745351
rect 58480 745339 58486 745351
rect 58538 745339 58544 745391
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 43120 743825 43126 743837
rect 42218 743797 43126 743825
rect 42218 743785 42224 743797
rect 43120 743785 43126 743797
rect 43178 743785 43184 743837
rect 42064 743193 42070 743245
rect 42122 743233 42128 743245
rect 42832 743233 42838 743245
rect 42122 743205 42838 743233
rect 42122 743193 42128 743205
rect 42832 743193 42838 743205
rect 42890 743193 42896 743245
rect 47440 742971 47446 743023
rect 47498 743011 47504 743023
rect 59632 743011 59638 743023
rect 47498 742983 59638 743011
rect 47498 742971 47504 742983
rect 59632 742971 59638 742983
rect 59690 742971 59696 743023
rect 44944 742897 44950 742949
rect 45002 742937 45008 742949
rect 59728 742937 59734 742949
rect 45002 742909 59734 742937
rect 45002 742897 45008 742909
rect 59728 742897 59734 742909
rect 59786 742897 59792 742949
rect 674416 742749 674422 742801
rect 674474 742789 674480 742801
rect 675184 742789 675190 742801
rect 674474 742761 675190 742789
rect 674474 742749 674480 742761
rect 675184 742749 675190 742761
rect 675242 742749 675248 742801
rect 42160 742601 42166 742653
rect 42218 742641 42224 742653
rect 42736 742641 42742 742653
rect 42218 742613 42742 742641
rect 42218 742601 42224 742613
rect 42736 742601 42742 742613
rect 42794 742601 42800 742653
rect 42160 741935 42166 741987
rect 42218 741975 42224 741987
rect 42352 741975 42358 741987
rect 42218 741947 42358 741975
rect 42218 741935 42224 741947
rect 42352 741935 42358 741947
rect 42410 741935 42416 741987
rect 674896 741417 674902 741469
rect 674954 741457 674960 741469
rect 675184 741457 675190 741469
rect 674954 741429 675190 741457
rect 674954 741417 674960 741429
rect 675184 741417 675190 741429
rect 675242 741417 675248 741469
rect 670768 737495 670774 737547
rect 670826 737535 670832 737547
rect 675280 737535 675286 737547
rect 670826 737507 675286 737535
rect 670826 737495 670832 737507
rect 675280 737495 675286 737507
rect 675338 737495 675344 737547
rect 654064 737421 654070 737473
rect 654122 737461 654128 737473
rect 674512 737461 674518 737473
rect 654122 737433 674518 737461
rect 654122 737421 654128 737433
rect 674512 737421 674518 737433
rect 674570 737421 674576 737473
rect 654160 737347 654166 737399
rect 654218 737387 654224 737399
rect 675280 737387 675286 737399
rect 654218 737359 675286 737387
rect 654218 737347 654224 737359
rect 675280 737347 675286 737359
rect 675338 737347 675344 737399
rect 672592 734905 672598 734957
rect 672650 734945 672656 734957
rect 675376 734945 675382 734957
rect 672650 734917 675382 734945
rect 672650 734905 672656 734917
rect 675376 734905 675382 734917
rect 675434 734905 675440 734957
rect 672976 734387 672982 734439
rect 673034 734427 673040 734439
rect 675376 734427 675382 734439
rect 673034 734399 675382 734427
rect 673034 734387 673040 734399
rect 675376 734387 675382 734399
rect 675434 734387 675440 734439
rect 673072 734165 673078 734217
rect 673130 734205 673136 734217
rect 675376 734205 675382 734217
rect 673130 734177 675382 734205
rect 673130 734165 673136 734177
rect 675376 734165 675382 734177
rect 675434 734165 675440 734217
rect 675184 733869 675190 733921
rect 675242 733909 675248 733921
rect 675472 733909 675478 733921
rect 675242 733881 675478 733909
rect 675242 733869 675248 733881
rect 675472 733869 675478 733881
rect 675530 733869 675536 733921
rect 672880 732315 672886 732367
rect 672938 732355 672944 732367
rect 675472 732355 675478 732367
rect 672938 732327 675478 732355
rect 672938 732315 672944 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 674512 732019 674518 732071
rect 674570 732059 674576 732071
rect 675376 732059 675382 732071
rect 674570 732031 675382 732059
rect 674570 732019 674576 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 674416 730465 674422 730517
rect 674474 730505 674480 730517
rect 675472 730505 675478 730517
rect 674474 730477 675478 730505
rect 674474 730465 674480 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 41776 730391 41782 730443
rect 41834 730431 41840 730443
rect 47536 730431 47542 730443
rect 41834 730403 47542 730431
rect 41834 730391 41840 730403
rect 47536 730391 47542 730403
rect 47594 730391 47600 730443
rect 41776 729873 41782 729925
rect 41834 729913 41840 729925
rect 44944 729913 44950 729925
rect 41834 729885 44950 729913
rect 41834 729873 41840 729885
rect 44944 729873 44950 729885
rect 45002 729873 45008 729925
rect 41776 729355 41782 729407
rect 41834 729395 41840 729407
rect 45040 729395 45046 729407
rect 41834 729367 45046 729395
rect 41834 729355 41840 729367
rect 45040 729355 45046 729367
rect 45098 729355 45104 729407
rect 41776 728985 41782 729037
rect 41834 729025 41840 729037
rect 43216 729025 43222 729037
rect 41834 728997 43222 729025
rect 41834 728985 41840 728997
rect 43216 728985 43222 728997
rect 43274 728985 43280 729037
rect 41584 728911 41590 728963
rect 41642 728951 41648 728963
rect 62224 728951 62230 728963
rect 41642 728923 62230 728951
rect 41642 728911 41648 728923
rect 62224 728911 62230 728923
rect 62282 728911 62288 728963
rect 41680 728689 41686 728741
rect 41738 728729 41744 728741
rect 62416 728729 62422 728741
rect 41738 728701 62422 728729
rect 41738 728689 41744 728701
rect 62416 728689 62422 728701
rect 62474 728689 62480 728741
rect 674128 728615 674134 728667
rect 674186 728655 674192 728667
rect 675472 728655 675478 728667
rect 674186 728627 675478 728655
rect 674186 728615 674192 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 41776 728319 41782 728371
rect 41834 728359 41840 728371
rect 43312 728359 43318 728371
rect 41834 728331 43318 728359
rect 41834 728319 41840 728331
rect 43312 728319 43318 728331
rect 43370 728319 43376 728371
rect 41776 727875 41782 727927
rect 41834 727915 41840 727927
rect 43408 727915 43414 727927
rect 41834 727887 43414 727915
rect 41834 727875 41840 727887
rect 43408 727875 43414 727887
rect 43466 727875 43472 727927
rect 41776 726839 41782 726891
rect 41834 726879 41840 726891
rect 43216 726879 43222 726891
rect 41834 726851 43222 726879
rect 41834 726839 41840 726851
rect 43216 726839 43222 726851
rect 43274 726839 43280 726891
rect 41776 725951 41782 726003
rect 41834 725991 41840 726003
rect 42928 725991 42934 726003
rect 41834 725963 42934 725991
rect 41834 725951 41840 725963
rect 42928 725951 42934 725963
rect 42986 725951 42992 726003
rect 41584 720993 41590 721045
rect 41642 721033 41648 721045
rect 43024 721033 43030 721045
rect 41642 721005 43030 721033
rect 41642 720993 41648 721005
rect 43024 720993 43030 721005
rect 43082 720993 43088 721045
rect 41584 720623 41590 720675
rect 41642 720663 41648 720675
rect 43120 720663 43126 720675
rect 41642 720635 43126 720663
rect 41642 720623 41648 720635
rect 43120 720623 43126 720635
rect 43178 720623 43184 720675
rect 42256 719735 42262 719787
rect 42314 719775 42320 719787
rect 42832 719775 42838 719787
rect 42314 719747 42838 719775
rect 42314 719735 42320 719747
rect 42832 719735 42838 719747
rect 42890 719735 42896 719787
rect 42160 719439 42166 719491
rect 42218 719479 42224 719491
rect 43120 719479 43126 719491
rect 42218 719451 43126 719479
rect 42218 719439 42224 719451
rect 43120 719439 43126 719451
rect 43178 719439 43184 719491
rect 41584 719291 41590 719343
rect 41642 719331 41648 719343
rect 43120 719331 43126 719343
rect 41642 719303 43126 719331
rect 41642 719291 41648 719303
rect 43120 719291 43126 719303
rect 43178 719291 43184 719343
rect 41488 717663 41494 717715
rect 41546 717703 41552 717715
rect 47440 717703 47446 717715
rect 41546 717675 47446 717703
rect 41546 717663 41552 717675
rect 47440 717663 47446 717675
rect 47498 717663 47504 717715
rect 41584 717515 41590 717567
rect 41642 717555 41648 717567
rect 42928 717555 42934 717567
rect 41642 717527 42934 717555
rect 41642 717515 41648 717527
rect 42928 717515 42934 717527
rect 42986 717515 42992 717567
rect 41872 715591 41878 715643
rect 41930 715631 41936 715643
rect 42736 715631 42742 715643
rect 41930 715603 42742 715631
rect 41930 715591 41936 715603
rect 42736 715591 42742 715603
rect 42794 715591 42800 715643
rect 655600 714703 655606 714755
rect 655658 714743 655664 714755
rect 676240 714743 676246 714755
rect 655658 714715 676246 714743
rect 655658 714703 655664 714715
rect 676240 714703 676246 714715
rect 676298 714703 676304 714755
rect 655408 714555 655414 714607
rect 655466 714595 655472 714607
rect 676144 714595 676150 714607
rect 655466 714567 676150 714595
rect 655466 714555 655472 714567
rect 676144 714555 676150 714567
rect 676202 714555 676208 714607
rect 655120 714407 655126 714459
rect 655178 714447 655184 714459
rect 676336 714447 676342 714459
rect 655178 714419 676342 714447
rect 655178 714407 655184 714419
rect 676336 714407 676342 714419
rect 676394 714407 676400 714459
rect 42832 714259 42838 714311
rect 42890 714299 42896 714311
rect 59632 714299 59638 714311
rect 42890 714271 59638 714299
rect 42890 714259 42896 714271
rect 59632 714259 59638 714271
rect 59690 714259 59696 714311
rect 43024 714185 43030 714237
rect 43082 714225 43088 714237
rect 43504 714225 43510 714237
rect 43082 714197 43510 714225
rect 43082 714185 43088 714197
rect 43504 714185 43510 714197
rect 43562 714185 43568 714237
rect 673360 714185 673366 714237
rect 673418 714225 673424 714237
rect 676048 714225 676054 714237
rect 673418 714197 676054 714225
rect 673418 714185 673424 714197
rect 676048 714185 676054 714197
rect 676106 714185 676112 714237
rect 41680 714037 41686 714089
rect 41738 714077 41744 714089
rect 43024 714077 43030 714089
rect 41738 714049 43030 714077
rect 41738 714037 41744 714049
rect 43024 714037 43030 714049
rect 43082 714037 43088 714089
rect 41776 713815 41782 713867
rect 41834 713815 41840 713867
rect 41794 713571 41822 713815
rect 42256 713741 42262 713793
rect 42314 713781 42320 713793
rect 43600 713781 43606 713793
rect 42314 713753 43606 713781
rect 42314 713741 42320 713753
rect 43600 713741 43606 713753
rect 43658 713741 43664 713793
rect 41776 713519 41782 713571
rect 41834 713519 41840 713571
rect 672784 713371 672790 713423
rect 672842 713411 672848 713423
rect 676240 713411 676246 713423
rect 672842 713383 676246 713411
rect 672842 713371 672848 713383
rect 676240 713371 676246 713383
rect 676298 713371 676304 713423
rect 669712 713075 669718 713127
rect 669770 713115 669776 713127
rect 670960 713115 670966 713127
rect 669770 713087 670966 713115
rect 669770 713075 669776 713087
rect 670960 713075 670966 713087
rect 671018 713115 671024 713127
rect 676048 713115 676054 713127
rect 671018 713087 676054 713115
rect 671018 713075 671024 713087
rect 676048 713075 676054 713087
rect 676106 713075 676112 713127
rect 670672 712631 670678 712683
rect 670730 712671 670736 712683
rect 676048 712671 676054 712683
rect 670730 712643 676054 712671
rect 670730 712631 670736 712643
rect 676048 712631 676054 712643
rect 676106 712631 676112 712683
rect 669520 711891 669526 711943
rect 669578 711931 669584 711943
rect 670864 711931 670870 711943
rect 669578 711903 670870 711931
rect 669578 711891 669584 711903
rect 670864 711891 670870 711903
rect 670922 711931 670928 711943
rect 676240 711931 676246 711943
rect 670922 711903 676246 711931
rect 670922 711891 670928 711903
rect 676240 711891 676246 711903
rect 676298 711891 676304 711943
rect 42064 711669 42070 711721
rect 42122 711709 42128 711721
rect 42736 711709 42742 711721
rect 42122 711681 42742 711709
rect 42122 711669 42128 711681
rect 42736 711669 42742 711681
rect 42794 711669 42800 711721
rect 42736 711521 42742 711573
rect 42794 711561 42800 711573
rect 43504 711561 43510 711573
rect 42794 711533 43510 711561
rect 42794 711521 42800 711533
rect 43504 711521 43510 711533
rect 43562 711521 43568 711573
rect 670576 711521 670582 711573
rect 670634 711561 670640 711573
rect 676048 711561 676054 711573
rect 670634 711533 676054 711561
rect 670634 711521 670640 711533
rect 676048 711521 676054 711533
rect 676106 711521 676112 711573
rect 43024 711299 43030 711351
rect 43082 711299 43088 711351
rect 674608 711299 674614 711351
rect 674666 711339 674672 711351
rect 676048 711339 676054 711351
rect 674666 711311 676054 711339
rect 674666 711299 674672 711311
rect 676048 711299 676054 711311
rect 676106 711299 676112 711351
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 42832 710895 42838 710907
rect 42218 710867 42838 710895
rect 42218 710855 42224 710867
rect 42832 710855 42838 710867
rect 42890 710855 42896 710907
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 42736 709933 42742 709945
rect 42218 709905 42742 709933
rect 42218 709893 42224 709905
rect 42736 709893 42742 709905
rect 42794 709893 42800 709945
rect 42736 709745 42742 709797
rect 42794 709785 42800 709797
rect 43042 709785 43070 711299
rect 42794 709757 43070 709785
rect 42794 709745 42800 709757
rect 42064 708487 42070 708539
rect 42122 708527 42128 708539
rect 43504 708527 43510 708539
rect 42122 708499 43510 708527
rect 42122 708487 42128 708499
rect 43504 708487 43510 708499
rect 43562 708487 43568 708539
rect 674992 708413 674998 708465
rect 675050 708453 675056 708465
rect 676048 708453 676054 708465
rect 675050 708425 676054 708453
rect 675050 708413 675056 708425
rect 676048 708413 676054 708425
rect 676106 708413 676112 708465
rect 42064 708339 42070 708391
rect 42122 708379 42128 708391
rect 43024 708379 43030 708391
rect 42122 708351 43030 708379
rect 42122 708339 42128 708351
rect 43024 708339 43030 708351
rect 43082 708339 43088 708391
rect 42160 707377 42166 707429
rect 42218 707417 42224 707429
rect 43120 707417 43126 707429
rect 42218 707389 43126 707417
rect 42218 707377 42224 707389
rect 43120 707377 43126 707389
rect 43178 707377 43184 707429
rect 42160 706563 42166 706615
rect 42218 706603 42224 706615
rect 42736 706603 42742 706615
rect 42218 706575 42742 706603
rect 42218 706563 42224 706575
rect 42736 706563 42742 706575
rect 42794 706563 42800 706615
rect 673264 705527 673270 705579
rect 673322 705567 673328 705579
rect 676048 705567 676054 705579
rect 673322 705539 676054 705567
rect 673322 705527 673328 705539
rect 676048 705527 676054 705539
rect 676106 705527 676112 705579
rect 673168 704861 673174 704913
rect 673226 704901 673232 704913
rect 676240 704901 676246 704913
rect 673226 704873 676246 704901
rect 673226 704861 673232 704873
rect 676240 704861 676246 704873
rect 676298 704861 676304 704913
rect 42352 704787 42358 704839
rect 42410 704827 42416 704839
rect 43600 704827 43606 704839
rect 42410 704799 43606 704827
rect 42410 704787 42416 704799
rect 43600 704787 43606 704799
rect 43658 704787 43664 704839
rect 42160 704269 42166 704321
rect 42218 704309 42224 704321
rect 42928 704309 42934 704321
rect 42218 704281 42934 704309
rect 42218 704269 42224 704281
rect 42928 704269 42934 704281
rect 42986 704269 42992 704321
rect 42064 703529 42070 703581
rect 42122 703569 42128 703581
rect 43024 703569 43030 703581
rect 42122 703541 43030 703569
rect 42122 703529 42128 703541
rect 43024 703529 43030 703541
rect 43082 703529 43088 703581
rect 42160 702863 42166 702915
rect 42218 702903 42224 702915
rect 42352 702903 42358 702915
rect 42218 702875 42358 702903
rect 42218 702863 42224 702875
rect 42352 702863 42358 702875
rect 42410 702863 42416 702915
rect 654352 702789 654358 702841
rect 654410 702829 654416 702841
rect 675376 702829 675382 702841
rect 654410 702801 675382 702829
rect 654410 702789 654416 702801
rect 675376 702789 675382 702801
rect 675434 702789 675440 702841
rect 649456 702715 649462 702767
rect 649514 702755 649520 702767
rect 679984 702755 679990 702767
rect 649514 702727 679990 702755
rect 649514 702715 649520 702727
rect 679984 702715 679990 702727
rect 680042 702715 680048 702767
rect 43504 702641 43510 702693
rect 43562 702681 43568 702693
rect 58768 702681 58774 702693
rect 43562 702653 58774 702681
rect 43562 702641 43568 702653
rect 58768 702641 58774 702653
rect 58826 702641 58832 702693
rect 45040 702567 45046 702619
rect 45098 702607 45104 702619
rect 58672 702607 58678 702619
rect 45098 702579 58678 702607
rect 45098 702567 45104 702579
rect 58672 702567 58678 702579
rect 58730 702567 58736 702619
rect 42160 702419 42166 702471
rect 42218 702459 42224 702471
rect 42832 702459 42838 702471
rect 42218 702431 42838 702459
rect 42218 702419 42224 702431
rect 42832 702419 42838 702431
rect 42890 702419 42896 702471
rect 42064 700495 42070 700547
rect 42122 700535 42128 700547
rect 43120 700535 43126 700547
rect 42122 700507 43126 700535
rect 42122 700495 42128 700507
rect 43120 700495 43126 700507
rect 43178 700495 43184 700547
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42928 700091 42934 700103
rect 42218 700063 42934 700091
rect 42218 700051 42224 700063
rect 42928 700051 42934 700063
rect 42986 700051 42992 700103
rect 47536 699755 47542 699807
rect 47594 699795 47600 699807
rect 59248 699795 59254 699807
rect 47594 699767 59254 699795
rect 47594 699755 47600 699767
rect 59248 699755 59254 699767
rect 59306 699755 59312 699807
rect 44944 699681 44950 699733
rect 45002 699721 45008 699733
rect 58864 699721 58870 699733
rect 45002 699693 58870 699721
rect 45002 699681 45008 699693
rect 58864 699681 58870 699693
rect 58922 699681 58928 699733
rect 42160 699385 42166 699437
rect 42218 699425 42224 699437
rect 42736 699425 42742 699437
rect 42218 699397 42742 699425
rect 42218 699385 42224 699397
rect 42736 699385 42742 699397
rect 42794 699385 42800 699437
rect 42064 698423 42070 698475
rect 42122 698463 42128 698475
rect 43792 698463 43798 698475
rect 42122 698435 43798 698463
rect 42122 698423 42128 698435
rect 43792 698423 43798 698435
rect 43850 698423 43856 698475
rect 654160 694279 654166 694331
rect 654218 694319 654224 694331
rect 674992 694319 674998 694331
rect 654218 694291 674998 694319
rect 654218 694279 654224 694291
rect 674992 694279 674998 694291
rect 675050 694279 675056 694331
rect 670960 693613 670966 693665
rect 671018 693653 671024 693665
rect 675472 693653 675478 693665
rect 671018 693625 675478 693653
rect 671018 693613 671024 693625
rect 675472 693613 675478 693625
rect 675530 693613 675536 693665
rect 674896 692873 674902 692925
rect 674954 692913 674960 692925
rect 675376 692913 675382 692925
rect 674954 692885 675382 692913
rect 674954 692873 674960 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 654064 691319 654070 691371
rect 654122 691359 654128 691371
rect 675184 691359 675190 691371
rect 654122 691331 675190 691359
rect 654122 691319 654128 691331
rect 675184 691319 675190 691331
rect 675242 691319 675248 691371
rect 674608 690431 674614 690483
rect 674666 690471 674672 690483
rect 675472 690471 675478 690483
rect 674666 690443 675478 690471
rect 674666 690431 674672 690443
rect 675472 690431 675478 690443
rect 675530 690431 675536 690483
rect 673168 689765 673174 689817
rect 673226 689805 673232 689817
rect 675376 689805 675382 689817
rect 673226 689777 675382 689805
rect 673226 689765 673232 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 673360 689321 673366 689373
rect 673418 689361 673424 689373
rect 675376 689361 675382 689373
rect 673418 689333 675382 689361
rect 673418 689321 673424 689333
rect 675376 689321 675382 689333
rect 675434 689321 675440 689373
rect 673264 689099 673270 689151
rect 673322 689139 673328 689151
rect 675376 689139 675382 689151
rect 673322 689111 675382 689139
rect 673322 689099 673328 689111
rect 675376 689099 675382 689111
rect 675434 689099 675440 689151
rect 674992 688877 674998 688929
rect 675050 688917 675056 688929
rect 675472 688917 675478 688929
rect 675050 688889 675478 688917
rect 675050 688877 675056 688889
rect 675472 688877 675478 688889
rect 675530 688877 675536 688929
rect 672688 687323 672694 687375
rect 672746 687363 672752 687375
rect 675472 687363 675478 687375
rect 672746 687335 675478 687363
rect 672746 687323 672752 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 675184 687027 675190 687079
rect 675242 687067 675248 687079
rect 675472 687067 675478 687079
rect 675242 687039 675478 687067
rect 675242 687027 675248 687039
rect 675472 687027 675478 687039
rect 675530 687027 675536 687079
rect 41776 686805 41782 686857
rect 41834 686845 41840 686857
rect 50320 686845 50326 686857
rect 41834 686817 50326 686845
rect 41834 686805 41840 686817
rect 50320 686805 50326 686817
rect 50378 686805 50384 686857
rect 41776 686287 41782 686339
rect 41834 686327 41840 686339
rect 47632 686327 47638 686339
rect 41834 686299 47638 686327
rect 41834 686287 41840 686299
rect 47632 686287 47638 686299
rect 47690 686287 47696 686339
rect 41584 685547 41590 685599
rect 41642 685587 41648 685599
rect 47728 685587 47734 685599
rect 41642 685559 47734 685587
rect 41642 685547 41648 685559
rect 47728 685547 47734 685559
rect 47786 685547 47792 685599
rect 674320 685473 674326 685525
rect 674378 685513 674384 685525
rect 675472 685513 675478 685525
rect 674378 685485 675478 685513
rect 674378 685473 674384 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 41776 685325 41782 685377
rect 41834 685365 41840 685377
rect 43312 685365 43318 685377
rect 41834 685337 43318 685365
rect 41834 685325 41840 685337
rect 43312 685325 43318 685337
rect 43370 685325 43376 685377
rect 41776 684807 41782 684859
rect 41834 684847 41840 684859
rect 43600 684847 43606 684859
rect 41834 684819 43606 684847
rect 41834 684807 41840 684819
rect 43600 684807 43606 684819
rect 43658 684807 43664 684859
rect 41776 683845 41782 683897
rect 41834 683885 41840 683897
rect 43408 683885 43414 683897
rect 41834 683857 43414 683885
rect 41834 683845 41840 683857
rect 43408 683845 43414 683857
rect 43466 683885 43472 683897
rect 44944 683885 44950 683897
rect 43466 683857 44950 683885
rect 43466 683845 43472 683857
rect 44944 683845 44950 683857
rect 45002 683845 45008 683897
rect 674224 683623 674230 683675
rect 674282 683663 674288 683675
rect 675472 683663 675478 683675
rect 674282 683635 675478 683663
rect 674282 683623 674288 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 41584 682957 41590 683009
rect 41642 682997 41648 683009
rect 43216 682997 43222 683009
rect 41642 682969 43222 682997
rect 41642 682957 41648 682969
rect 43216 682957 43222 682969
rect 43274 682997 43280 683009
rect 45136 682997 45142 683009
rect 43274 682969 45142 682997
rect 43274 682957 43280 682969
rect 45136 682957 45142 682969
rect 45194 682957 45200 683009
rect 41776 680663 41782 680715
rect 41834 680703 41840 680715
rect 43024 680703 43030 680715
rect 41834 680675 43030 680703
rect 41834 680663 41840 680675
rect 43024 680663 43030 680675
rect 43082 680663 43088 680715
rect 41584 676075 41590 676127
rect 41642 676115 41648 676127
rect 43120 676115 43126 676127
rect 41642 676087 43126 676115
rect 41642 676075 41648 676087
rect 43120 676075 43126 676087
rect 43178 676075 43184 676127
rect 41584 674299 41590 674351
rect 41642 674339 41648 674351
rect 42928 674339 42934 674351
rect 41642 674311 42934 674339
rect 41642 674299 41648 674311
rect 42928 674299 42934 674311
rect 42986 674299 42992 674351
rect 41584 674003 41590 674055
rect 41642 674043 41648 674055
rect 47536 674043 47542 674055
rect 41642 674015 47542 674043
rect 41642 674003 41648 674015
rect 47536 674003 47542 674015
rect 47594 674003 47600 674055
rect 39760 673855 39766 673907
rect 39818 673895 39824 673907
rect 41488 673895 41494 673907
rect 39818 673867 41494 673895
rect 39818 673855 39824 673867
rect 41488 673855 41494 673867
rect 41546 673855 41552 673907
rect 34480 672523 34486 672575
rect 34538 672563 34544 672575
rect 42160 672563 42166 672575
rect 34538 672535 42166 672563
rect 34538 672523 34544 672535
rect 42160 672523 42166 672535
rect 42218 672523 42224 672575
rect 41968 671339 41974 671391
rect 42026 671379 42032 671391
rect 43120 671379 43126 671391
rect 42026 671351 43126 671379
rect 42026 671339 42032 671351
rect 43120 671339 43126 671351
rect 43178 671339 43184 671391
rect 37360 671265 37366 671317
rect 37418 671305 37424 671317
rect 43696 671305 43702 671317
rect 37418 671277 43702 671305
rect 37418 671265 37424 671277
rect 43696 671265 43702 671277
rect 43754 671265 43760 671317
rect 41488 671191 41494 671243
rect 41546 671231 41552 671243
rect 43504 671231 43510 671243
rect 41546 671203 43510 671231
rect 41546 671191 41552 671203
rect 43504 671191 43510 671203
rect 43562 671191 43568 671243
rect 42160 671117 42166 671169
rect 42218 671157 42224 671169
rect 43312 671157 43318 671169
rect 42218 671129 43318 671157
rect 42218 671117 42224 671129
rect 43312 671117 43318 671129
rect 43370 671117 43376 671169
rect 42832 671043 42838 671095
rect 42890 671083 42896 671095
rect 59632 671083 59638 671095
rect 42890 671055 59638 671083
rect 42890 671043 42896 671055
rect 59632 671043 59638 671055
rect 59690 671043 59696 671095
rect 41776 670599 41782 670651
rect 41834 670599 41840 670651
rect 42256 670599 42262 670651
rect 42314 670639 42320 670651
rect 43408 670639 43414 670651
rect 42314 670611 43414 670639
rect 42314 670599 42320 670611
rect 43408 670599 43414 670611
rect 43466 670599 43472 670651
rect 41794 670355 41822 670599
rect 41776 670303 41782 670355
rect 41834 670303 41840 670355
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 43024 668567 43030 668579
rect 42218 668539 43030 668567
rect 42218 668527 42224 668539
rect 43024 668527 43030 668539
rect 43082 668527 43088 668579
rect 43120 668453 43126 668505
rect 43178 668453 43184 668505
rect 43138 668209 43166 668453
rect 655504 668379 655510 668431
rect 655562 668419 655568 668431
rect 676240 668419 676246 668431
rect 655562 668391 676246 668419
rect 655562 668379 655568 668391
rect 676240 668379 676246 668391
rect 676298 668379 676304 668431
rect 43120 668157 43126 668209
rect 43178 668157 43184 668209
rect 655312 668157 655318 668209
rect 655370 668197 655376 668209
rect 676240 668197 676246 668209
rect 655370 668169 676246 668197
rect 655370 668157 655376 668169
rect 676240 668157 676246 668169
rect 676298 668157 676304 668209
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 42832 667901 42838 667913
rect 42218 667873 42838 667901
rect 42218 667861 42224 667873
rect 42832 667861 42838 667873
rect 42890 667861 42896 667913
rect 42832 667713 42838 667765
rect 42890 667753 42896 667765
rect 43312 667753 43318 667765
rect 42890 667725 43318 667753
rect 42890 667713 42896 667725
rect 43312 667713 43318 667725
rect 43370 667713 43376 667765
rect 672784 667565 672790 667617
rect 672842 667605 672848 667617
rect 675952 667605 675958 667617
rect 672842 667577 675958 667605
rect 672842 667565 672848 667577
rect 675952 667565 675958 667577
rect 676010 667565 676016 667617
rect 652240 666751 652246 666803
rect 652298 666791 652304 666803
rect 668752 666791 668758 666803
rect 652298 666763 668758 666791
rect 652298 666751 652304 666763
rect 668752 666751 668758 666763
rect 668810 666751 668816 666803
rect 672784 666751 672790 666803
rect 672842 666791 672848 666803
rect 676240 666791 676246 666803
rect 672842 666763 676246 666791
rect 672842 666751 672848 666763
rect 676240 666751 676246 666763
rect 676298 666751 676304 666803
rect 649744 666677 649750 666729
rect 649802 666717 649808 666729
rect 670672 666717 670678 666729
rect 649802 666689 670678 666717
rect 649802 666677 649808 666689
rect 670672 666677 670678 666689
rect 670730 666717 670736 666729
rect 676144 666717 676150 666729
rect 670730 666689 676150 666717
rect 670730 666677 670736 666689
rect 676144 666677 676150 666689
rect 676202 666677 676208 666729
rect 670384 666011 670390 666063
rect 670442 666051 670448 666063
rect 675952 666051 675958 666063
rect 670442 666023 675958 666051
rect 670442 666011 670448 666023
rect 675952 666011 675958 666023
rect 676010 666011 676016 666063
rect 668752 665493 668758 665545
rect 668810 665533 668816 665545
rect 670576 665533 670582 665545
rect 668810 665505 670582 665533
rect 668810 665493 668816 665505
rect 670576 665493 670582 665505
rect 670634 665533 670640 665545
rect 675952 665533 675958 665545
rect 670634 665505 675958 665533
rect 670634 665493 670640 665505
rect 675952 665493 675958 665505
rect 676010 665493 676016 665545
rect 655216 665419 655222 665471
rect 655274 665459 655280 665471
rect 676048 665459 676054 665471
rect 655274 665431 676054 665459
rect 655274 665419 655280 665431
rect 676048 665419 676054 665431
rect 676106 665419 676112 665471
rect 42160 665345 42166 665397
rect 42218 665385 42224 665397
rect 42928 665385 42934 665397
rect 42218 665357 42934 665385
rect 42218 665345 42224 665357
rect 42928 665345 42934 665357
rect 42986 665345 42992 665397
rect 42064 665271 42070 665323
rect 42122 665311 42128 665323
rect 45040 665311 45046 665323
rect 42122 665283 45046 665311
rect 42122 665271 42128 665283
rect 45040 665271 45046 665283
rect 45098 665271 45104 665323
rect 42928 665197 42934 665249
rect 42986 665237 42992 665249
rect 43408 665237 43414 665249
rect 42986 665209 43414 665237
rect 42986 665197 42992 665209
rect 43408 665197 43414 665209
rect 43466 665197 43472 665249
rect 674416 665197 674422 665249
rect 674474 665237 674480 665249
rect 676048 665237 676054 665249
rect 674474 665209 676054 665237
rect 674474 665197 674480 665209
rect 676048 665197 676054 665209
rect 676106 665197 676112 665249
rect 670672 664975 670678 665027
rect 670730 665015 670736 665027
rect 675952 665015 675958 665027
rect 670730 664987 675958 665015
rect 670730 664975 670736 664987
rect 675952 664975 675958 664987
rect 676010 664975 676016 665027
rect 42064 663939 42070 663991
rect 42122 663979 42128 663991
rect 43024 663979 43030 663991
rect 42122 663951 43030 663979
rect 42122 663939 42128 663951
rect 43024 663939 43030 663951
rect 43082 663939 43088 663991
rect 43120 663495 43126 663547
rect 43178 663495 43184 663547
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 43138 663387 43166 663495
rect 42218 663359 43166 663387
rect 42218 663347 42224 663359
rect 43120 663273 43126 663325
rect 43178 663313 43184 663325
rect 43696 663313 43702 663325
rect 43178 663285 43702 663313
rect 43178 663273 43184 663285
rect 43696 663273 43702 663285
rect 43754 663273 43760 663325
rect 674128 662311 674134 662363
rect 674186 662351 674192 662363
rect 676048 662351 676054 662363
rect 674186 662323 676054 662351
rect 674186 662311 674192 662323
rect 676048 662311 676054 662323
rect 676106 662311 676112 662363
rect 670768 660461 670774 660513
rect 670826 660501 670832 660513
rect 676048 660501 676054 660513
rect 670826 660473 676054 660501
rect 670826 660461 670832 660473
rect 676048 660461 676054 660473
rect 676106 660461 676112 660513
rect 42064 660387 42070 660439
rect 42122 660427 42128 660439
rect 42928 660427 42934 660439
rect 42122 660399 42934 660427
rect 42122 660387 42128 660399
rect 42928 660387 42934 660399
rect 42986 660387 42992 660439
rect 672880 660091 672886 660143
rect 672938 660131 672944 660143
rect 676048 660131 676054 660143
rect 672938 660103 676054 660131
rect 672938 660091 672944 660103
rect 676048 660091 676054 660103
rect 676106 660091 676112 660143
rect 42160 659869 42166 659921
rect 42218 659909 42224 659921
rect 42832 659909 42838 659921
rect 42218 659881 42838 659909
rect 42218 659869 42224 659881
rect 42832 659869 42838 659881
rect 42890 659869 42896 659921
rect 672976 659721 672982 659773
rect 673034 659761 673040 659773
rect 676240 659761 676246 659773
rect 673034 659733 676246 659761
rect 673034 659721 673040 659733
rect 676240 659721 676246 659733
rect 676298 659721 676304 659773
rect 47728 659425 47734 659477
rect 47786 659465 47792 659477
rect 59152 659465 59158 659477
rect 47786 659437 59158 659465
rect 47786 659425 47792 659437
rect 59152 659425 59158 659437
rect 59210 659425 59216 659477
rect 45040 659351 45046 659403
rect 45098 659391 45104 659403
rect 58768 659391 58774 659403
rect 45098 659363 58774 659391
rect 45098 659351 45104 659363
rect 58768 659351 58774 659363
rect 58826 659351 58832 659403
rect 42064 659055 42070 659107
rect 42122 659095 42128 659107
rect 43120 659095 43126 659107
rect 42122 659067 43126 659095
rect 42122 659055 42128 659067
rect 43120 659055 43126 659067
rect 43178 659055 43184 659107
rect 672592 658611 672598 658663
rect 672650 658651 672656 658663
rect 676048 658651 676054 658663
rect 672650 658623 676054 658651
rect 672650 658611 672656 658623
rect 676048 658611 676054 658623
rect 676106 658611 676112 658663
rect 673072 658241 673078 658293
rect 673130 658281 673136 658293
rect 676240 658281 676246 658293
rect 673130 658253 676246 658281
rect 673130 658241 673136 658253
rect 676240 658241 676246 658253
rect 676298 658241 676304 658293
rect 42064 657353 42070 657405
rect 42122 657393 42128 657405
rect 43024 657393 43030 657405
rect 42122 657365 43030 657393
rect 42122 657353 42128 657365
rect 43024 657353 43030 657365
rect 43082 657353 43088 657405
rect 42160 656835 42166 656887
rect 42218 656875 42224 656887
rect 42832 656875 42838 656887
rect 42218 656847 42838 656875
rect 42218 656835 42224 656847
rect 42832 656835 42838 656847
rect 42890 656835 42896 656887
rect 654160 656687 654166 656739
rect 654218 656727 654224 656739
rect 675376 656727 675382 656739
rect 654218 656699 675382 656727
rect 654218 656687 654224 656699
rect 675376 656687 675382 656699
rect 675434 656687 675440 656739
rect 50320 656613 50326 656665
rect 50378 656653 50384 656665
rect 58192 656653 58198 656665
rect 50378 656625 58198 656653
rect 50378 656613 50384 656625
rect 58192 656613 58198 656625
rect 58250 656613 58256 656665
rect 47632 656539 47638 656591
rect 47690 656579 47696 656591
rect 58384 656579 58390 656591
rect 47690 656551 58390 656579
rect 47690 656539 47696 656551
rect 58384 656539 58390 656551
rect 58442 656539 58448 656591
rect 42160 656169 42166 656221
rect 42218 656209 42224 656221
rect 42928 656209 42934 656221
rect 42218 656181 42934 656209
rect 42218 656169 42224 656181
rect 42928 656169 42934 656181
rect 42986 656169 42992 656221
rect 42160 655503 42166 655555
rect 42218 655543 42224 655555
rect 45904 655543 45910 655555
rect 42218 655515 45910 655543
rect 42218 655503 42224 655515
rect 45904 655503 45910 655515
rect 45962 655503 45968 655555
rect 679984 654137 679990 654149
rect 659506 654109 679990 654137
rect 649552 654023 649558 654075
rect 649610 654063 649616 654075
rect 659506 654063 659534 654109
rect 679984 654097 679990 654109
rect 680042 654097 680048 654149
rect 649610 654035 659534 654063
rect 649610 654023 649616 654035
rect 670864 648917 670870 648969
rect 670922 648957 670928 648969
rect 675184 648957 675190 648969
rect 670922 648929 675190 648957
rect 670922 648917 670928 648929
rect 675184 648917 675190 648929
rect 675242 648917 675248 648969
rect 670768 648325 670774 648377
rect 670826 648365 670832 648377
rect 675184 648365 675190 648377
rect 670826 648337 675190 648365
rect 670826 648325 670832 648337
rect 675184 648325 675190 648337
rect 675242 648325 675248 648377
rect 655792 648251 655798 648303
rect 655850 648291 655856 648303
rect 674992 648291 674998 648303
rect 655850 648263 674998 648291
rect 655850 648251 655856 648263
rect 674992 648251 674998 648263
rect 675050 648251 675056 648303
rect 673840 648029 673846 648081
rect 673898 648069 673904 648081
rect 675184 648069 675190 648081
rect 673898 648041 675190 648069
rect 673898 648029 673904 648041
rect 675184 648029 675190 648041
rect 675242 648029 675248 648081
rect 655984 645143 655990 645195
rect 656042 645183 656048 645195
rect 675280 645183 675286 645195
rect 656042 645155 675286 645183
rect 656042 645143 656048 645155
rect 675280 645143 675286 645155
rect 675338 645143 675344 645195
rect 672976 644551 672982 644603
rect 673034 644591 673040 644603
rect 675376 644591 675382 644603
rect 673034 644563 675382 644591
rect 673034 644551 673040 644563
rect 675376 644551 675382 644563
rect 675434 644551 675440 644603
rect 670576 644033 670582 644085
rect 670634 644073 670640 644085
rect 675472 644073 675478 644085
rect 670634 644045 675478 644073
rect 670634 644033 670640 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 41776 643663 41782 643715
rect 41834 643703 41840 643715
rect 50320 643703 50326 643715
rect 41834 643675 50326 643703
rect 41834 643663 41840 643675
rect 50320 643663 50326 643675
rect 50378 643663 50384 643715
rect 674992 643663 674998 643715
rect 675050 643703 675056 643715
rect 675376 643703 675382 643715
rect 675050 643675 675382 643703
rect 675050 643663 675056 643675
rect 675376 643663 675382 643675
rect 675434 643663 675440 643715
rect 672880 643589 672886 643641
rect 672938 643629 672944 643641
rect 675472 643629 675478 643641
rect 672938 643601 675478 643629
rect 672938 643589 672944 643601
rect 675472 643589 675478 643601
rect 675530 643589 675536 643641
rect 41776 643071 41782 643123
rect 41834 643111 41840 643123
rect 47728 643111 47734 643123
rect 41834 643083 47734 643111
rect 41834 643071 41840 643083
rect 47728 643071 47734 643083
rect 47786 643071 47792 643123
rect 41488 642553 41494 642605
rect 41546 642593 41552 642605
rect 61936 642593 61942 642605
rect 41546 642565 61942 642593
rect 41546 642553 41552 642565
rect 61936 642553 61942 642565
rect 61994 642553 62000 642605
rect 41680 642479 41686 642531
rect 41738 642519 41744 642531
rect 62128 642519 62134 642531
rect 41738 642491 62134 642519
rect 41738 642479 41744 642491
rect 62128 642479 62134 642491
rect 62186 642479 62192 642531
rect 41584 642331 41590 642383
rect 41642 642371 41648 642383
rect 47824 642371 47830 642383
rect 41642 642343 47830 642371
rect 41642 642331 41648 642343
rect 47824 642331 47830 642343
rect 47882 642331 47888 642383
rect 670480 642257 670486 642309
rect 670538 642297 670544 642309
rect 675472 642297 675478 642309
rect 670538 642269 675478 642297
rect 670538 642257 670544 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 41776 642183 41782 642235
rect 41834 642223 41840 642235
rect 43504 642223 43510 642235
rect 41834 642195 43510 642223
rect 41834 642183 41840 642195
rect 43504 642183 43510 642195
rect 43562 642183 43568 642235
rect 41776 641591 41782 641643
rect 41834 641631 41840 641643
rect 43600 641631 43606 641643
rect 41834 641603 43606 641631
rect 41834 641591 41840 641603
rect 43600 641591 43606 641603
rect 43658 641591 43664 641643
rect 41776 640111 41782 640163
rect 41834 640151 41840 640163
rect 43408 640151 43414 640163
rect 41834 640123 43414 640151
rect 41834 640111 41840 640123
rect 43408 640111 43414 640123
rect 43466 640111 43472 640163
rect 41584 633895 41590 633947
rect 41642 633935 41648 633947
rect 43120 633935 43126 633947
rect 41642 633907 43126 633935
rect 41642 633895 41648 633907
rect 43120 633895 43126 633907
rect 43178 633895 43184 633947
rect 41872 631083 41878 631135
rect 41930 631123 41936 631135
rect 43024 631123 43030 631135
rect 41930 631095 43030 631123
rect 41930 631083 41936 631095
rect 43024 631083 43030 631095
rect 43082 631083 43088 631135
rect 41584 630787 41590 630839
rect 41642 630827 41648 630839
rect 47632 630827 47638 630839
rect 41642 630799 47638 630827
rect 41642 630787 41648 630799
rect 47632 630787 47638 630799
rect 47690 630787 47696 630839
rect 43120 628123 43126 628175
rect 43178 628163 43184 628175
rect 43504 628163 43510 628175
rect 43178 628135 43510 628163
rect 43178 628123 43184 628135
rect 43504 628123 43510 628135
rect 43562 628123 43568 628175
rect 37360 627975 37366 628027
rect 37418 628015 37424 628027
rect 43888 628015 43894 628027
rect 37418 627987 43894 628015
rect 37418 627975 37424 627987
rect 43888 627975 43894 627987
rect 43946 627975 43952 628027
rect 34480 627901 34486 627953
rect 34538 627941 34544 627953
rect 43792 627941 43798 627953
rect 34538 627913 43798 627941
rect 34538 627901 34544 627913
rect 43792 627901 43798 627913
rect 43850 627901 43856 627953
rect 40144 627827 40150 627879
rect 40202 627867 40208 627879
rect 43696 627867 43702 627879
rect 40202 627839 43702 627867
rect 40202 627827 40208 627839
rect 43696 627827 43702 627839
rect 43754 627827 43760 627879
rect 41488 627679 41494 627731
rect 41546 627719 41552 627731
rect 43120 627719 43126 627731
rect 41546 627691 43126 627719
rect 41546 627679 41552 627691
rect 43120 627679 43126 627691
rect 43178 627679 43184 627731
rect 43216 627679 43222 627731
rect 43274 627719 43280 627731
rect 43274 627691 43358 627719
rect 43274 627679 43280 627691
rect 42256 627605 42262 627657
rect 42314 627645 42320 627657
rect 43024 627645 43030 627657
rect 42314 627617 43030 627645
rect 42314 627605 42320 627617
rect 43024 627605 43030 627617
rect 43082 627605 43088 627657
rect 42160 627531 42166 627583
rect 42218 627571 42224 627583
rect 43216 627571 43222 627583
rect 42218 627543 43222 627571
rect 42218 627531 42224 627543
rect 43216 627531 43222 627543
rect 43274 627531 43280 627583
rect 43330 627571 43358 627691
rect 43330 627543 43454 627571
rect 43426 627509 43454 627543
rect 43408 627457 43414 627509
rect 43466 627457 43472 627509
rect 41776 627383 41782 627435
rect 41834 627383 41840 627435
rect 41794 627213 41822 627383
rect 41776 627161 41782 627213
rect 41834 627161 41840 627213
rect 42832 625163 42838 625215
rect 42890 625203 42896 625215
rect 43216 625203 43222 625215
rect 42890 625175 43222 625203
rect 42890 625163 42896 625175
rect 43216 625163 43222 625175
rect 43274 625163 43280 625215
rect 655408 624941 655414 624993
rect 655466 624981 655472 624993
rect 676240 624981 676246 624993
rect 655466 624953 676246 624981
rect 655466 624941 655472 624953
rect 676240 624941 676246 624953
rect 676298 624941 676304 624993
rect 42160 624275 42166 624327
rect 42218 624315 42224 624327
rect 58960 624315 58966 624327
rect 42218 624287 58966 624315
rect 42218 624275 42224 624287
rect 58960 624275 58966 624287
rect 59018 624275 59024 624327
rect 672784 623979 672790 624031
rect 672842 624019 672848 624031
rect 676048 624019 676054 624031
rect 672842 623991 676054 624019
rect 672842 623979 672848 623991
rect 676048 623979 676054 623991
rect 676106 623979 676112 624031
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 42928 623501 42934 623513
rect 42218 623473 42934 623501
rect 42218 623461 42224 623473
rect 42928 623461 42934 623473
rect 42986 623461 42992 623513
rect 672592 623387 672598 623439
rect 672650 623427 672656 623439
rect 676048 623427 676054 623439
rect 672650 623399 676054 623427
rect 672650 623387 672656 623399
rect 676048 623387 676054 623399
rect 676106 623387 676112 623439
rect 42928 623313 42934 623365
rect 42986 623353 42992 623365
rect 43408 623353 43414 623365
rect 42986 623325 43414 623353
rect 42986 623313 42992 623325
rect 43408 623313 43414 623325
rect 43466 623313 43472 623365
rect 669616 623165 669622 623217
rect 669674 623205 669680 623217
rect 670384 623205 670390 623217
rect 669674 623177 670390 623205
rect 669674 623165 669680 623177
rect 670384 623165 670390 623177
rect 670442 623205 670448 623217
rect 676336 623205 676342 623217
rect 670442 623177 676342 623205
rect 670442 623165 670448 623177
rect 676336 623165 676342 623177
rect 676394 623165 676400 623217
rect 670192 622425 670198 622477
rect 670250 622465 670256 622477
rect 676048 622465 676054 622477
rect 670250 622437 676054 622465
rect 670250 622425 670256 622437
rect 676048 622425 676054 622437
rect 676106 622425 676112 622477
rect 655600 622351 655606 622403
rect 655658 622391 655664 622403
rect 676240 622391 676246 622403
rect 655658 622363 676246 622391
rect 655658 622351 655664 622363
rect 676240 622351 676246 622363
rect 676298 622351 676304 622403
rect 655120 622203 655126 622255
rect 655178 622243 655184 622255
rect 676144 622243 676150 622255
rect 655178 622215 676150 622243
rect 655178 622203 655184 622215
rect 676144 622203 676150 622215
rect 676202 622203 676208 622255
rect 42160 622055 42166 622107
rect 42218 622095 42224 622107
rect 47920 622095 47926 622107
rect 42218 622067 47926 622095
rect 42218 622055 42224 622067
rect 47920 622055 47926 622067
rect 47978 622055 47984 622107
rect 674320 621981 674326 622033
rect 674378 622021 674384 622033
rect 676240 622021 676246 622033
rect 674378 621993 676246 622021
rect 674378 621981 674384 621993
rect 676240 621981 676246 621993
rect 676298 621981 676304 622033
rect 42160 621907 42166 621959
rect 42218 621947 42224 621959
rect 43024 621947 43030 621959
rect 42218 621919 43030 621947
rect 42218 621907 42224 621919
rect 43024 621907 43030 621919
rect 43082 621907 43088 621959
rect 670672 621907 670678 621959
rect 670730 621947 670736 621959
rect 676048 621947 676054 621959
rect 670730 621919 676054 621947
rect 670730 621907 670736 621919
rect 676048 621907 676054 621919
rect 676106 621907 676112 621959
rect 43024 621759 43030 621811
rect 43082 621799 43088 621811
rect 43696 621799 43702 621811
rect 43082 621771 43702 621799
rect 43082 621759 43088 621771
rect 43696 621759 43702 621771
rect 43754 621759 43760 621811
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 43504 621651 43510 621663
rect 42218 621623 43510 621651
rect 42218 621611 42224 621623
rect 43504 621611 43510 621623
rect 43562 621611 43568 621663
rect 670288 621315 670294 621367
rect 670346 621355 670352 621367
rect 676048 621355 676054 621367
rect 670346 621327 676054 621355
rect 670346 621315 670352 621327
rect 676048 621315 676054 621327
rect 676106 621315 676112 621367
rect 42928 620985 42934 620997
rect 42082 620957 42934 620985
rect 42082 620923 42110 620957
rect 42928 620945 42934 620957
rect 42986 620945 42992 620997
rect 42064 620871 42070 620923
rect 42122 620871 42128 620923
rect 42928 620797 42934 620849
rect 42986 620837 42992 620849
rect 43792 620837 43798 620849
rect 42986 620809 43798 620837
rect 42986 620797 42992 620809
rect 43792 620797 43798 620809
rect 43850 620797 43856 620849
rect 43216 620649 43222 620701
rect 43274 620689 43280 620701
rect 43600 620689 43606 620701
rect 43274 620661 43606 620689
rect 43274 620649 43280 620661
rect 43600 620649 43606 620661
rect 43658 620649 43664 620701
rect 42160 620353 42166 620405
rect 42218 620393 42224 620405
rect 43120 620393 43126 620405
rect 42218 620365 43126 620393
rect 42218 620353 42224 620365
rect 43120 620353 43126 620365
rect 43178 620353 43184 620405
rect 43120 620205 43126 620257
rect 43178 620245 43184 620257
rect 43888 620245 43894 620257
rect 43178 620217 43894 620245
rect 43178 620205 43184 620217
rect 43888 620205 43894 620217
rect 43946 620205 43952 620257
rect 669808 619835 669814 619887
rect 669866 619875 669872 619887
rect 670672 619875 670678 619887
rect 669866 619847 670678 619875
rect 669866 619835 669872 619847
rect 670672 619835 670678 619847
rect 670730 619835 670736 619887
rect 674608 619021 674614 619073
rect 674666 619061 674672 619073
rect 676048 619061 676054 619073
rect 674666 619033 676054 619061
rect 674666 619021 674672 619033
rect 676048 619021 676054 619033
rect 676106 619021 676112 619073
rect 674224 618799 674230 618851
rect 674282 618839 674288 618851
rect 676240 618839 676246 618851
rect 674282 618811 676246 618839
rect 674282 618799 674288 618811
rect 676240 618799 676246 618811
rect 676298 618799 676304 618851
rect 42064 617837 42070 617889
rect 42122 617877 42128 617889
rect 42832 617877 42838 617889
rect 42122 617849 42838 617877
rect 42122 617837 42128 617849
rect 42832 617837 42838 617849
rect 42890 617837 42896 617889
rect 42736 617319 42742 617371
rect 42794 617319 42800 617371
rect 42160 617171 42166 617223
rect 42218 617211 42224 617223
rect 42754 617211 42782 617319
rect 42218 617183 42782 617211
rect 42218 617171 42224 617183
rect 670960 617097 670966 617149
rect 671018 617137 671024 617149
rect 676240 617137 676246 617149
rect 671018 617109 676246 617137
rect 671018 617097 671024 617109
rect 676240 617097 676246 617109
rect 676298 617097 676304 617149
rect 42160 616653 42166 616705
rect 42218 616693 42224 616705
rect 42928 616693 42934 616705
rect 42218 616665 42934 616693
rect 42218 616653 42224 616665
rect 42928 616653 42934 616665
rect 42986 616653 42992 616705
rect 672688 616505 672694 616557
rect 672746 616545 672752 616557
rect 676048 616545 676054 616557
rect 672746 616517 676054 616545
rect 672746 616505 672752 616517
rect 676048 616505 676054 616517
rect 676106 616505 676112 616557
rect 47824 616283 47830 616335
rect 47882 616323 47888 616335
rect 58960 616323 58966 616335
rect 47882 616295 58966 616323
rect 47882 616283 47888 616295
rect 58960 616283 58966 616295
rect 59018 616283 59024 616335
rect 47920 616209 47926 616261
rect 47978 616249 47984 616261
rect 59632 616249 59638 616261
rect 47978 616221 59638 616249
rect 47978 616209 47984 616221
rect 59632 616209 59638 616221
rect 59690 616209 59696 616261
rect 42160 615987 42166 616039
rect 42218 616027 42224 616039
rect 43024 616027 43030 616039
rect 42218 615999 43030 616027
rect 42218 615987 42224 615999
rect 43024 615987 43030 615999
rect 43082 615987 43088 616039
rect 673360 615913 673366 615965
rect 673418 615953 673424 615965
rect 676048 615953 676054 615965
rect 673418 615925 676054 615953
rect 673418 615913 673424 615925
rect 676048 615913 676054 615925
rect 676106 615913 676112 615965
rect 673168 615173 673174 615225
rect 673226 615213 673232 615225
rect 676240 615213 676246 615225
rect 673226 615185 676246 615213
rect 673226 615173 673232 615185
rect 676240 615173 676246 615185
rect 676298 615173 676304 615225
rect 673264 614433 673270 614485
rect 673322 614473 673328 614485
rect 676048 614473 676054 614485
rect 673322 614445 676054 614473
rect 673322 614433 673328 614445
rect 676048 614433 676054 614445
rect 676106 614433 676112 614485
rect 42160 614137 42166 614189
rect 42218 614177 42224 614189
rect 43120 614177 43126 614189
rect 42218 614149 43126 614177
rect 42218 614137 42224 614149
rect 43120 614137 43126 614149
rect 43178 614137 43184 614189
rect 42160 613619 42166 613671
rect 42218 613659 42224 613671
rect 42832 613659 42838 613671
rect 42218 613631 42838 613659
rect 42218 613619 42224 613631
rect 42832 613619 42838 613631
rect 42890 613619 42896 613671
rect 655120 613471 655126 613523
rect 655178 613511 655184 613523
rect 675376 613511 675382 613523
rect 655178 613483 675382 613511
rect 655178 613471 655184 613483
rect 675376 613471 675382 613483
rect 675434 613471 675440 613523
rect 50320 613397 50326 613449
rect 50378 613437 50384 613449
rect 59632 613437 59638 613449
rect 50378 613409 59638 613437
rect 50378 613397 50384 613409
rect 59632 613397 59638 613409
rect 59690 613397 59696 613449
rect 47728 613323 47734 613375
rect 47786 613363 47792 613375
rect 59536 613363 59542 613375
rect 47786 613335 59542 613363
rect 47786 613323 47792 613335
rect 59536 613323 59542 613335
rect 59594 613323 59600 613375
rect 42064 612953 42070 613005
rect 42122 612993 42128 613005
rect 42736 612993 42742 613005
rect 42122 612965 42742 612993
rect 42122 612953 42128 612965
rect 42736 612953 42742 612965
rect 42794 612953 42800 613005
rect 42160 612361 42166 612413
rect 42218 612401 42224 612413
rect 45904 612401 45910 612413
rect 42218 612373 45910 612401
rect 42218 612361 42224 612373
rect 45904 612361 45910 612373
rect 45962 612361 45968 612413
rect 649648 610659 649654 610711
rect 649706 610699 649712 610711
rect 679984 610699 679990 610711
rect 649706 610671 679990 610699
rect 649706 610659 649712 610671
rect 679984 610659 679990 610671
rect 680042 610659 680048 610711
rect 673264 606885 673270 606937
rect 673322 606925 673328 606937
rect 675184 606925 675190 606937
rect 673322 606897 675190 606925
rect 673322 606885 673328 606897
rect 675184 606885 675190 606897
rect 675242 606885 675248 606937
rect 670960 603259 670966 603311
rect 671018 603299 671024 603311
rect 675376 603299 675382 603311
rect 671018 603271 675382 603299
rect 671018 603259 671024 603271
rect 675376 603259 675382 603271
rect 675434 603259 675440 603311
rect 673360 603037 673366 603089
rect 673418 603077 673424 603089
rect 675376 603077 675382 603089
rect 673418 603049 675382 603077
rect 673418 603037 673424 603049
rect 675376 603037 675382 603049
rect 675434 603037 675440 603089
rect 655792 602075 655798 602127
rect 655850 602115 655856 602127
rect 674992 602115 674998 602127
rect 655850 602087 674998 602115
rect 655850 602075 655856 602087
rect 674992 602075 674998 602087
rect 675050 602075 675056 602127
rect 653776 602001 653782 602053
rect 653834 602041 653840 602053
rect 674896 602041 674902 602053
rect 653834 602013 674902 602041
rect 653834 602001 653840 602013
rect 674896 602001 674902 602013
rect 674954 602001 674960 602053
rect 673072 601927 673078 601979
rect 673130 601967 673136 601979
rect 675280 601967 675286 601979
rect 673130 601939 675286 601967
rect 673130 601927 673136 601939
rect 675280 601927 675286 601939
rect 675338 601927 675344 601979
rect 41776 600447 41782 600499
rect 41834 600487 41840 600499
rect 50320 600487 50326 600499
rect 41834 600459 50326 600487
rect 41834 600447 41840 600459
rect 50320 600447 50326 600459
rect 50378 600447 50384 600499
rect 41584 599707 41590 599759
rect 41642 599747 41648 599759
rect 47824 599747 47830 599759
rect 41642 599719 47830 599747
rect 41642 599707 41648 599719
rect 47824 599707 47830 599719
rect 47882 599707 47888 599759
rect 673168 599559 673174 599611
rect 673226 599599 673232 599611
rect 675376 599599 675382 599611
rect 673226 599571 675382 599599
rect 673226 599559 673232 599571
rect 675376 599559 675382 599571
rect 675434 599559 675440 599611
rect 41776 599337 41782 599389
rect 41834 599377 41840 599389
rect 47920 599377 47926 599389
rect 41834 599349 47926 599377
rect 41834 599337 41840 599349
rect 47920 599337 47926 599349
rect 47978 599337 47984 599389
rect 670672 599263 670678 599315
rect 670730 599303 670736 599315
rect 675376 599303 675382 599315
rect 670730 599275 675382 599303
rect 670730 599263 670736 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 41776 598967 41782 599019
rect 41834 599007 41840 599019
rect 43216 599007 43222 599019
rect 41834 598979 43222 599007
rect 41834 598967 41840 598979
rect 43216 598967 43222 598979
rect 43274 598967 43280 599019
rect 672784 598893 672790 598945
rect 672842 598933 672848 598945
rect 675376 598933 675382 598945
rect 672842 598905 675382 598933
rect 672842 598893 672848 598905
rect 675376 598893 675382 598905
rect 675434 598893 675440 598945
rect 674992 598671 674998 598723
rect 675050 598711 675056 598723
rect 675472 598711 675478 598723
rect 675050 598683 675478 598711
rect 675050 598671 675056 598683
rect 675472 598671 675478 598683
rect 675530 598671 675536 598723
rect 41584 598227 41590 598279
rect 41642 598267 41648 598279
rect 43504 598267 43510 598279
rect 41642 598239 43510 598267
rect 41642 598227 41648 598239
rect 43504 598227 43510 598239
rect 43562 598227 43568 598279
rect 672688 597117 672694 597169
rect 672746 597157 672752 597169
rect 675472 597157 675478 597169
rect 672746 597129 675478 597157
rect 672746 597117 672752 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 674896 596821 674902 596873
rect 674954 596861 674960 596873
rect 675376 596861 675382 596873
rect 674954 596833 675382 596861
rect 674954 596821 674960 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 41584 596155 41590 596207
rect 41642 596195 41648 596207
rect 43312 596195 43318 596207
rect 41642 596167 43318 596195
rect 41642 596155 41648 596167
rect 43312 596155 43318 596167
rect 43370 596195 43376 596207
rect 45040 596195 45046 596207
rect 43370 596167 45046 596195
rect 43370 596155 43376 596167
rect 45040 596155 45046 596167
rect 45098 596155 45104 596207
rect 41776 593491 41782 593543
rect 41834 593531 41840 593543
rect 43024 593531 43030 593543
rect 41834 593503 43030 593531
rect 41834 593491 41840 593503
rect 43024 593491 43030 593503
rect 43082 593491 43088 593543
rect 41872 590901 41878 590953
rect 41930 590941 41936 590953
rect 43120 590941 43126 590953
rect 41930 590913 43126 590941
rect 41930 590901 41936 590913
rect 43120 590901 43126 590913
rect 43178 590901 43184 590953
rect 41584 590531 41590 590583
rect 41642 590571 41648 590583
rect 42832 590571 42838 590583
rect 41642 590543 42838 590571
rect 41642 590531 41648 590543
rect 42832 590531 42838 590543
rect 42890 590531 42896 590583
rect 41968 589495 41974 589547
rect 42026 589535 42032 589547
rect 43120 589535 43126 589547
rect 42026 589507 43126 589535
rect 42026 589495 42032 589507
rect 43120 589495 43126 589507
rect 43178 589495 43184 589547
rect 41584 589347 41590 589399
rect 41642 589387 41648 589399
rect 43120 589387 43126 589399
rect 41642 589359 43126 589387
rect 41642 589347 41648 589359
rect 43120 589347 43126 589359
rect 43178 589347 43184 589399
rect 41584 587867 41590 587919
rect 41642 587907 41648 587919
rect 42832 587907 42838 587919
rect 41642 587879 42838 587907
rect 41642 587867 41648 587879
rect 42832 587867 42838 587879
rect 42890 587867 42896 587919
rect 41584 587571 41590 587623
rect 41642 587611 41648 587623
rect 47728 587611 47734 587623
rect 41642 587583 47734 587611
rect 41642 587571 41648 587583
rect 47728 587571 47734 587583
rect 47786 587571 47792 587623
rect 42352 584611 42358 584663
rect 42410 584651 42416 584663
rect 43408 584651 43414 584663
rect 42410 584623 43414 584651
rect 42410 584611 42416 584623
rect 43408 584611 43414 584623
rect 43466 584611 43472 584663
rect 42064 584537 42070 584589
rect 42122 584577 42128 584589
rect 43312 584577 43318 584589
rect 42122 584549 43318 584577
rect 42122 584537 42128 584549
rect 43312 584537 43318 584549
rect 43370 584537 43376 584589
rect 42160 584463 42166 584515
rect 42218 584503 42224 584515
rect 43216 584503 43222 584515
rect 42218 584475 43222 584503
rect 42218 584463 42224 584475
rect 43216 584463 43222 584475
rect 43274 584463 43280 584515
rect 41776 584167 41782 584219
rect 41834 584167 41840 584219
rect 41794 583997 41822 584167
rect 41776 583945 41782 583997
rect 41834 583945 41840 583997
rect 42160 582095 42166 582147
rect 42218 582135 42224 582147
rect 43024 582135 43030 582147
rect 42218 582107 43030 582135
rect 42218 582095 42224 582107
rect 43024 582095 43030 582107
rect 43082 582095 43088 582147
rect 43024 581947 43030 581999
rect 43082 581987 43088 581999
rect 43216 581987 43222 581999
rect 43082 581959 43222 581987
rect 43082 581947 43088 581959
rect 43216 581947 43222 581959
rect 43274 581947 43280 581999
rect 42160 580837 42166 580889
rect 42218 580877 42224 580889
rect 58960 580877 58966 580889
rect 42218 580849 58966 580877
rect 42218 580837 42224 580849
rect 58960 580837 58966 580849
rect 59018 580837 59024 580889
rect 42064 580245 42070 580297
rect 42122 580285 42128 580297
rect 42928 580285 42934 580297
rect 42122 580257 42934 580285
rect 42122 580245 42128 580257
rect 42928 580245 42934 580257
rect 42986 580245 42992 580297
rect 42928 580097 42934 580149
rect 42986 580137 42992 580149
rect 43312 580137 43318 580149
rect 42986 580109 43318 580137
rect 42986 580097 42992 580109
rect 43312 580097 43318 580109
rect 43370 580097 43376 580149
rect 655696 579283 655702 579335
rect 655754 579323 655760 579335
rect 676240 579323 676246 579335
rect 655754 579295 676246 579323
rect 655754 579283 655760 579295
rect 676240 579283 676246 579295
rect 676298 579283 676304 579335
rect 655504 579135 655510 579187
rect 655562 579175 655568 579187
rect 676336 579175 676342 579187
rect 655562 579147 676342 579175
rect 655562 579135 655568 579147
rect 676336 579135 676342 579147
rect 676394 579135 676400 579187
rect 655312 578987 655318 579039
rect 655370 579027 655376 579039
rect 676144 579027 676150 579039
rect 655370 578999 676150 579027
rect 655370 578987 655376 578999
rect 676144 578987 676150 578999
rect 676202 578987 676208 579039
rect 42160 578913 42166 578965
rect 42218 578953 42224 578965
rect 48016 578953 48022 578965
rect 42218 578925 48022 578953
rect 42218 578913 42224 578925
rect 48016 578913 48022 578925
rect 48074 578913 48080 578965
rect 42160 578765 42166 578817
rect 42218 578805 42224 578817
rect 42832 578805 42838 578817
rect 42218 578777 42838 578805
rect 42218 578765 42224 578777
rect 42832 578765 42838 578777
rect 42890 578765 42896 578817
rect 672592 578765 672598 578817
rect 672650 578805 672656 578817
rect 676240 578805 676246 578817
rect 672650 578777 676246 578805
rect 672650 578765 672656 578777
rect 676240 578765 676246 578777
rect 676298 578765 676304 578817
rect 42160 577803 42166 577855
rect 42218 577843 42224 577855
rect 43120 577843 43126 577855
rect 42218 577815 43126 577843
rect 42218 577803 42224 577815
rect 43120 577803 43126 577815
rect 43178 577803 43184 577855
rect 672496 577803 672502 577855
rect 672554 577843 672560 577855
rect 676240 577843 676246 577855
rect 672554 577815 676246 577843
rect 672554 577803 672560 577815
rect 676240 577803 676246 577815
rect 676298 577803 676304 577855
rect 670096 577433 670102 577485
rect 670154 577473 670160 577485
rect 676048 577473 676054 577485
rect 670154 577445 676054 577473
rect 670154 577433 670160 577445
rect 676048 577433 676054 577445
rect 676106 577433 676112 577485
rect 672592 577063 672598 577115
rect 672650 577103 672656 577115
rect 676048 577103 676054 577115
rect 672650 577075 676054 577103
rect 672650 577063 672656 577075
rect 676048 577063 676054 577075
rect 676106 577063 676112 577115
rect 42064 576915 42070 576967
rect 42122 576955 42128 576967
rect 43024 576955 43030 576967
rect 42122 576927 43030 576955
rect 42122 576915 42128 576927
rect 43024 576915 43030 576927
rect 43082 576915 43088 576967
rect 670288 576545 670294 576597
rect 670346 576585 670352 576597
rect 676048 576585 676054 576597
rect 670346 576557 676054 576585
rect 670346 576545 670352 576557
rect 676048 576545 676054 576557
rect 676106 576545 676112 576597
rect 669904 576027 669910 576079
rect 669962 576067 669968 576079
rect 670288 576067 670294 576079
rect 669962 576039 670294 576067
rect 669962 576027 669968 576039
rect 670288 576027 670294 576039
rect 670346 576027 670352 576079
rect 670384 575879 670390 575931
rect 670442 575919 670448 575931
rect 676048 575919 676054 575931
rect 670442 575891 676054 575919
rect 670442 575879 670448 575891
rect 676048 575879 676054 575891
rect 676106 575879 676112 575931
rect 42160 574547 42166 574599
rect 42218 574587 42224 574599
rect 43120 574587 43126 574599
rect 42218 574559 43126 574587
rect 42218 574547 42224 574559
rect 43120 574547 43126 574559
rect 43178 574547 43184 574599
rect 42160 574103 42166 574155
rect 42218 574143 42224 574155
rect 42928 574143 42934 574155
rect 42218 574115 42934 574143
rect 42218 574103 42224 574115
rect 42928 574103 42934 574115
rect 42986 574103 42992 574155
rect 47920 573067 47926 573119
rect 47978 573107 47984 573119
rect 58960 573107 58966 573119
rect 47978 573079 58966 573107
rect 47978 573067 47984 573079
rect 58960 573067 58966 573079
rect 59018 573067 59024 573119
rect 48016 572993 48022 573045
rect 48074 573033 48080 573045
rect 59632 573033 59638 573045
rect 48074 573005 59638 573033
rect 48074 572993 48080 573005
rect 59632 572993 59638 573005
rect 59690 572993 59696 573045
rect 42160 572623 42166 572675
rect 42218 572663 42224 572675
rect 42832 572663 42838 572675
rect 42218 572635 42838 572663
rect 42218 572623 42224 572635
rect 42832 572623 42838 572635
rect 42890 572623 42896 572675
rect 670864 572253 670870 572305
rect 670922 572293 670928 572305
rect 676240 572293 676246 572305
rect 670922 572265 676246 572293
rect 670922 572253 670928 572265
rect 676240 572253 676246 572265
rect 676298 572253 676304 572305
rect 670768 571513 670774 571565
rect 670826 571553 670832 571565
rect 676048 571553 676054 571565
rect 670826 571525 676054 571553
rect 670826 571513 670832 571525
rect 676048 571513 676054 571525
rect 676106 571513 676112 571565
rect 670480 571069 670486 571121
rect 670538 571109 670544 571121
rect 676048 571109 676054 571121
rect 670538 571081 676054 571109
rect 670538 571069 670544 571081
rect 676048 571069 676054 571081
rect 676106 571069 676112 571121
rect 670576 570551 670582 570603
rect 670634 570591 670640 570603
rect 676048 570591 676054 570603
rect 670634 570563 676054 570591
rect 670634 570551 670640 570563
rect 676048 570551 676054 570563
rect 676106 570551 676112 570603
rect 42064 570403 42070 570455
rect 42122 570443 42128 570455
rect 43024 570443 43030 570455
rect 42122 570415 43030 570443
rect 42122 570403 42128 570415
rect 43024 570403 43030 570415
rect 43082 570403 43088 570455
rect 42160 570329 42166 570381
rect 42218 570369 42224 570381
rect 42928 570369 42934 570381
rect 42218 570341 42934 570369
rect 42218 570329 42224 570341
rect 42928 570329 42934 570341
rect 42986 570329 42992 570381
rect 50320 570181 50326 570233
rect 50378 570221 50384 570233
rect 59344 570221 59350 570233
rect 50378 570193 59350 570221
rect 50378 570181 50384 570193
rect 59344 570181 59350 570193
rect 59402 570181 59408 570233
rect 673840 570181 673846 570233
rect 673898 570221 673904 570233
rect 676240 570221 676246 570233
rect 673898 570193 676246 570221
rect 673898 570181 673904 570193
rect 676240 570181 676246 570193
rect 676298 570181 676304 570233
rect 47824 570107 47830 570159
rect 47882 570147 47888 570159
rect 59536 570147 59542 570159
rect 47882 570119 59542 570147
rect 47882 570107 47888 570119
rect 59536 570107 59542 570119
rect 59594 570107 59600 570159
rect 42064 569663 42070 569715
rect 42122 569703 42128 569715
rect 42928 569703 42934 569715
rect 42122 569675 42934 569703
rect 42122 569663 42128 569675
rect 42928 569663 42934 569675
rect 42986 569663 42992 569715
rect 672976 569589 672982 569641
rect 673034 569629 673040 569641
rect 676048 569629 676054 569641
rect 673034 569601 676054 569629
rect 673034 569589 673040 569601
rect 676048 569589 676054 569601
rect 676106 569589 676112 569641
rect 42160 569145 42166 569197
rect 42218 569185 42224 569197
rect 46192 569185 46198 569197
rect 42218 569157 46198 569185
rect 42218 569145 42224 569157
rect 46192 569145 46198 569157
rect 46250 569145 46256 569197
rect 672880 569071 672886 569123
rect 672938 569111 672944 569123
rect 676048 569111 676054 569123
rect 672938 569083 676054 569111
rect 672938 569071 672944 569083
rect 676048 569071 676054 569083
rect 676106 569071 676112 569123
rect 655696 567443 655702 567495
rect 655754 567483 655760 567495
rect 675376 567483 675382 567495
rect 655754 567455 675382 567483
rect 655754 567443 655760 567455
rect 675376 567443 675382 567455
rect 675434 567443 675440 567495
rect 649840 567369 649846 567421
rect 649898 567409 649904 567421
rect 679984 567409 679990 567421
rect 649898 567381 679990 567409
rect 649898 567369 649904 567381
rect 679984 567369 679990 567381
rect 680042 567369 680048 567421
rect 674416 559525 674422 559577
rect 674474 559565 674480 559577
rect 675376 559565 675382 559577
rect 674474 559537 675382 559565
rect 674474 559525 674480 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 656560 558785 656566 558837
rect 656618 558825 656624 558837
rect 674992 558825 674998 558837
rect 656618 558797 674998 558825
rect 656618 558785 656624 558797
rect 674992 558785 674998 558797
rect 675050 558785 675056 558837
rect 674608 558045 674614 558097
rect 674666 558085 674672 558097
rect 675376 558085 675382 558097
rect 674666 558057 675382 558085
rect 674666 558045 674672 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 673840 555973 673846 556025
rect 673898 556013 673904 556025
rect 675280 556013 675286 556025
rect 673898 555985 675286 556013
rect 673898 555973 673904 555985
rect 675280 555973 675286 555985
rect 675338 555973 675344 556025
rect 654160 555825 654166 555877
rect 654218 555865 654224 555877
rect 675280 555865 675286 555877
rect 654218 555837 675286 555865
rect 654218 555825 654224 555837
rect 675280 555825 675286 555837
rect 675338 555825 675344 555877
rect 674896 555011 674902 555063
rect 674954 555051 674960 555063
rect 675472 555051 675478 555063
rect 674954 555023 675478 555051
rect 674954 555011 674960 555023
rect 675472 555011 675478 555023
rect 675530 555011 675536 555063
rect 673744 554345 673750 554397
rect 673802 554385 673808 554397
rect 675376 554385 675382 554397
rect 673802 554357 675382 554385
rect 673802 554345 673808 554357
rect 675376 554345 675382 554357
rect 675434 554345 675440 554397
rect 672880 553901 672886 553953
rect 672938 553941 672944 553953
rect 675472 553941 675478 553953
rect 672938 553913 675478 553941
rect 672938 553901 672944 553913
rect 675472 553901 675478 553913
rect 675530 553901 675536 553953
rect 674992 553457 674998 553509
rect 675050 553497 675056 553509
rect 675376 553497 675382 553509
rect 675050 553469 675382 553497
rect 675050 553457 675056 553469
rect 675376 553457 675382 553469
rect 675434 553457 675440 553509
rect 673648 553309 673654 553361
rect 673706 553349 673712 553361
rect 675472 553349 675478 553361
rect 673706 553321 675478 553349
rect 673706 553309 673712 553321
rect 675472 553309 675478 553321
rect 675530 553309 675536 553361
rect 670864 551903 670870 551955
rect 670922 551943 670928 551955
rect 675472 551943 675478 551955
rect 670922 551915 675478 551943
rect 670922 551903 670928 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 674320 548869 674326 548921
rect 674378 548909 674384 548921
rect 675280 548909 675286 548921
rect 674378 548881 675286 548909
rect 674378 548869 674384 548881
rect 675280 548869 675286 548881
rect 675338 548869 675344 548921
rect 674224 548203 674230 548255
rect 674282 548243 674288 548255
rect 675280 548243 675286 548255
rect 674282 548215 675286 548243
rect 674282 548203 674288 548215
rect 675280 548203 675286 548215
rect 675338 548203 675344 548255
rect 41584 543023 41590 543075
rect 41642 543063 41648 543075
rect 50512 543063 50518 543075
rect 41642 543035 50518 543063
rect 41642 543023 41648 543035
rect 50512 543023 50518 543035
rect 50570 543023 50576 543075
rect 41776 542653 41782 542705
rect 41834 542693 41840 542705
rect 48784 542693 48790 542705
rect 41834 542665 48790 542693
rect 41834 542653 41840 542665
rect 48784 542653 48790 542665
rect 48842 542653 48848 542705
rect 41776 542135 41782 542187
rect 41834 542175 41840 542187
rect 48880 542175 48886 542187
rect 41834 542147 48886 542175
rect 41834 542135 41840 542147
rect 48880 542135 48886 542147
rect 48938 542135 48944 542187
rect 41776 541765 41782 541817
rect 41834 541805 41840 541817
rect 43216 541805 43222 541817
rect 41834 541777 43222 541805
rect 41834 541765 41840 541777
rect 43216 541765 43222 541777
rect 43274 541765 43280 541817
rect 42736 541543 42742 541595
rect 42794 541583 42800 541595
rect 57712 541583 57718 541595
rect 42794 541555 57718 541583
rect 42794 541543 42800 541555
rect 57712 541543 57718 541555
rect 57770 541543 57776 541595
rect 42832 541469 42838 541521
rect 42890 541509 42896 541521
rect 57616 541509 57622 541521
rect 42890 541481 57622 541509
rect 42890 541469 42896 541481
rect 57616 541469 57622 541481
rect 57674 541469 57680 541521
rect 42160 539693 42166 539745
rect 42218 539733 42224 539745
rect 42928 539733 42934 539745
rect 42218 539705 42934 539733
rect 42218 539693 42224 539705
rect 42928 539693 42934 539705
rect 42986 539693 42992 539745
rect 42160 538139 42166 538191
rect 42218 538179 42224 538191
rect 42736 538179 42742 538191
rect 42218 538151 42742 538179
rect 42218 538139 42224 538151
rect 42736 538139 42742 538151
rect 42794 538139 42800 538191
rect 42160 536437 42166 536489
rect 42218 536477 42224 536489
rect 42832 536477 42838 536489
rect 42218 536449 42838 536477
rect 42218 536437 42224 536449
rect 42832 536437 42838 536449
rect 42890 536437 42896 536489
rect 672496 533773 672502 533825
rect 672554 533813 672560 533825
rect 675952 533813 675958 533825
rect 672554 533785 675958 533813
rect 672554 533773 672560 533785
rect 675952 533773 675958 533785
rect 676010 533773 676016 533825
rect 42064 533699 42070 533751
rect 42122 533739 42128 533751
rect 42736 533739 42742 533751
rect 42122 533711 42742 533739
rect 42122 533699 42128 533711
rect 42736 533699 42742 533711
rect 42794 533699 42800 533751
rect 655600 533255 655606 533307
rect 655658 533295 655664 533307
rect 676048 533295 676054 533307
rect 655658 533267 676054 533295
rect 655658 533255 655664 533267
rect 676048 533255 676054 533267
rect 676106 533255 676112 533307
rect 655408 533107 655414 533159
rect 655466 533147 655472 533159
rect 676144 533147 676150 533159
rect 655466 533119 676150 533147
rect 655466 533107 655472 533119
rect 676144 533107 676150 533119
rect 676202 533107 676208 533159
rect 655216 532959 655222 533011
rect 655274 532999 655280 533011
rect 676240 532999 676246 533011
rect 655274 532971 676246 532999
rect 655274 532959 655280 532971
rect 676240 532959 676246 532971
rect 676298 532959 676304 533011
rect 672400 532663 672406 532715
rect 672458 532703 672464 532715
rect 672592 532703 672598 532715
rect 672458 532675 672598 532703
rect 672458 532663 672464 532675
rect 672592 532663 672598 532675
rect 672650 532703 672656 532715
rect 676048 532703 676054 532715
rect 672650 532675 676054 532703
rect 672650 532663 672656 532675
rect 676048 532663 676054 532675
rect 676106 532663 676112 532715
rect 42160 531479 42166 531531
rect 42218 531519 42224 531531
rect 42736 531519 42742 531531
rect 42218 531491 42742 531519
rect 42218 531479 42224 531491
rect 42736 531479 42742 531491
rect 42794 531479 42800 531531
rect 670288 531479 670294 531531
rect 670346 531519 670352 531531
rect 676240 531519 676246 531531
rect 670346 531491 676246 531519
rect 670346 531479 670352 531491
rect 676240 531479 676246 531491
rect 676298 531479 676304 531531
rect 42160 530887 42166 530939
rect 42218 530927 42224 530939
rect 42832 530927 42838 530939
rect 42218 530899 42838 530927
rect 42218 530887 42224 530899
rect 42832 530887 42838 530899
rect 42890 530887 42896 530939
rect 42160 529407 42166 529459
rect 42218 529447 42224 529459
rect 43024 529447 43030 529459
rect 42218 529419 43030 529447
rect 42218 529407 42224 529419
rect 43024 529407 43030 529419
rect 43082 529407 43088 529459
rect 673264 528001 673270 528053
rect 673322 528041 673328 528053
rect 676240 528041 676246 528053
rect 673322 528013 676246 528041
rect 673322 528001 673328 528013
rect 676240 528001 676246 528013
rect 676298 528001 676304 528053
rect 42160 527779 42166 527831
rect 42218 527819 42224 527831
rect 43120 527819 43126 527831
rect 42218 527791 43126 527819
rect 42218 527779 42224 527791
rect 43120 527779 43126 527791
rect 43178 527779 43184 527831
rect 48880 527483 48886 527535
rect 48938 527523 48944 527535
rect 59632 527523 59638 527535
rect 48938 527495 59638 527523
rect 48938 527483 48944 527495
rect 59632 527483 59638 527495
rect 59690 527483 59696 527535
rect 673072 527409 673078 527461
rect 673130 527449 673136 527461
rect 676240 527449 676246 527461
rect 673130 527421 676246 527449
rect 673130 527409 673136 527421
rect 676240 527409 676246 527421
rect 676298 527409 676304 527461
rect 42064 527187 42070 527239
rect 42122 527227 42128 527239
rect 42832 527227 42838 527239
rect 42122 527199 42838 527227
rect 42122 527187 42128 527199
rect 42832 527187 42838 527199
rect 42890 527187 42896 527239
rect 670960 526669 670966 526721
rect 671018 526709 671024 526721
rect 676048 526709 676054 526721
rect 671018 526681 676054 526709
rect 671018 526669 671024 526681
rect 676048 526669 676054 526681
rect 676106 526669 676112 526721
rect 42160 526447 42166 526499
rect 42218 526487 42224 526499
rect 42928 526487 42934 526499
rect 42218 526459 42934 526487
rect 42218 526447 42224 526459
rect 42928 526447 42934 526459
rect 42986 526447 42992 526499
rect 672688 526299 672694 526351
rect 672746 526339 672752 526351
rect 676048 526339 676054 526351
rect 672746 526311 676054 526339
rect 672746 526299 672752 526311
rect 676048 526299 676054 526311
rect 676106 526299 676112 526351
rect 42064 525929 42070 525981
rect 42122 525969 42128 525981
rect 46672 525969 46678 525981
rect 42122 525941 46678 525969
rect 42122 525929 42128 525941
rect 46672 525929 46678 525941
rect 46730 525929 46736 525981
rect 670672 525929 670678 525981
rect 670730 525969 670736 525981
rect 676240 525969 676246 525981
rect 670730 525941 676246 525969
rect 670730 525929 670736 525941
rect 676240 525929 676246 525941
rect 676298 525929 676304 525981
rect 673360 525189 673366 525241
rect 673418 525229 673424 525241
rect 676048 525229 676054 525241
rect 673418 525201 676054 525229
rect 673418 525189 673424 525201
rect 676048 525189 676054 525201
rect 676106 525189 676112 525241
rect 48784 524967 48790 525019
rect 48842 525007 48848 525019
rect 59632 525007 59638 525019
rect 48842 524979 59638 525007
rect 48842 524967 48848 524979
rect 59632 524967 59638 524979
rect 59690 524967 59696 525019
rect 673168 524819 673174 524871
rect 673226 524859 673232 524871
rect 676048 524859 676054 524871
rect 673226 524831 676054 524859
rect 673226 524819 673232 524831
rect 676048 524819 676054 524831
rect 676106 524819 676112 524871
rect 50512 524671 50518 524723
rect 50570 524711 50576 524723
rect 59344 524711 59350 524723
rect 50570 524683 59350 524711
rect 50570 524671 50576 524683
rect 59344 524671 59350 524683
rect 59402 524671 59408 524723
rect 672784 524449 672790 524501
rect 672842 524489 672848 524501
rect 676240 524489 676246 524501
rect 672842 524461 676246 524489
rect 672842 524449 672848 524461
rect 676240 524449 676246 524461
rect 676298 524449 676304 524501
rect 42352 524227 42358 524279
rect 42410 524267 42416 524279
rect 47824 524267 47830 524279
rect 42410 524239 47830 524267
rect 42410 524227 42416 524239
rect 47824 524227 47830 524239
rect 47882 524227 47888 524279
rect 649936 521267 649942 521319
rect 649994 521307 650000 521319
rect 679792 521307 679798 521319
rect 649994 521279 679798 521307
rect 649994 521267 650000 521279
rect 679792 521267 679798 521279
rect 679850 521267 679856 521319
rect 43408 519935 43414 519987
rect 43466 519935 43472 519987
rect 43426 519765 43454 519935
rect 43408 519713 43414 519765
rect 43466 519713 43472 519765
rect 43312 514089 43318 514141
rect 43370 514129 43376 514141
rect 43504 514129 43510 514141
rect 43370 514101 43510 514129
rect 43370 514089 43376 514101
rect 43504 514089 43510 514101
rect 43562 514089 43568 514141
rect 655504 490039 655510 490091
rect 655562 490079 655568 490091
rect 676240 490079 676246 490091
rect 655562 490051 676246 490079
rect 655562 490039 655568 490051
rect 676240 490039 676246 490051
rect 676298 490039 676304 490091
rect 655312 489891 655318 489943
rect 655370 489931 655376 489943
rect 676144 489931 676150 489943
rect 655370 489903 676150 489931
rect 655370 489891 655376 489903
rect 676144 489891 676150 489903
rect 676202 489891 676208 489943
rect 655120 489743 655126 489795
rect 655178 489783 655184 489795
rect 676336 489783 676342 489795
rect 655178 489755 676342 489783
rect 655178 489743 655184 489755
rect 676336 489743 676342 489755
rect 676394 489743 676400 489795
rect 670000 488115 670006 488167
rect 670058 488155 670064 488167
rect 676048 488155 676054 488167
rect 670058 488127 676054 488155
rect 670058 488115 670064 488127
rect 676048 488115 676054 488127
rect 676106 488155 676112 488167
rect 676624 488155 676630 488167
rect 676106 488127 676630 488155
rect 676106 488115 676112 488127
rect 676624 488115 676630 488127
rect 676682 488115 676688 488167
rect 670192 487079 670198 487131
rect 670250 487119 670256 487131
rect 676240 487119 676246 487131
rect 670250 487091 676246 487119
rect 670250 487079 670256 487091
rect 676240 487079 676246 487091
rect 676298 487119 676304 487131
rect 676528 487119 676534 487131
rect 676298 487091 676534 487119
rect 676298 487079 676304 487091
rect 676528 487079 676534 487091
rect 676586 487079 676592 487131
rect 674896 486635 674902 486687
rect 674954 486675 674960 486687
rect 676048 486675 676054 486687
rect 674954 486647 676054 486675
rect 674954 486635 674960 486647
rect 676048 486635 676054 486647
rect 676106 486635 676112 486687
rect 674320 486561 674326 486613
rect 674378 486601 674384 486613
rect 675952 486601 675958 486613
rect 674378 486573 675958 486601
rect 674378 486561 674384 486573
rect 675952 486561 675958 486573
rect 676010 486561 676016 486613
rect 674416 486487 674422 486539
rect 674474 486527 674480 486539
rect 676240 486527 676246 486539
rect 674474 486499 676246 486527
rect 674474 486487 674480 486499
rect 676240 486487 676246 486499
rect 676298 486487 676304 486539
rect 674608 483749 674614 483801
rect 674666 483789 674672 483801
rect 676048 483789 676054 483801
rect 674666 483761 676054 483789
rect 674666 483749 674672 483761
rect 676048 483749 676054 483761
rect 676106 483749 676112 483801
rect 674224 483675 674230 483727
rect 674282 483715 674288 483727
rect 675952 483715 675958 483727
rect 674282 483687 675958 483715
rect 674282 483675 674288 483687
rect 675952 483675 675958 483687
rect 676010 483675 676016 483727
rect 670864 481899 670870 481951
rect 670922 481939 670928 481951
rect 676048 481939 676054 481951
rect 670922 481911 676054 481939
rect 670922 481899 670928 481911
rect 676048 481899 676054 481911
rect 676106 481899 676112 481951
rect 672880 481529 672886 481581
rect 672938 481569 672944 481581
rect 676240 481569 676246 481581
rect 672938 481541 676246 481569
rect 672938 481529 672944 481541
rect 676240 481529 676246 481541
rect 676298 481529 676304 481581
rect 673840 480789 673846 480841
rect 673898 480829 673904 480841
rect 676048 480829 676054 480841
rect 673898 480801 676054 480829
rect 673898 480789 673904 480801
rect 676048 480789 676054 480801
rect 676106 480789 676112 480841
rect 673744 480419 673750 480471
rect 673802 480459 673808 480471
rect 676048 480459 676054 480471
rect 673802 480431 676054 480459
rect 673802 480419 673808 480431
rect 676048 480419 676054 480431
rect 676106 480419 676112 480471
rect 673648 480049 673654 480101
rect 673706 480089 673712 480101
rect 676240 480089 676246 480101
rect 673706 480061 676246 480089
rect 673706 480049 673712 480061
rect 676240 480049 676246 480061
rect 676298 480049 676304 480101
rect 676624 479235 676630 479287
rect 676682 479275 676688 479287
rect 679696 479275 679702 479287
rect 676682 479247 679702 479275
rect 676682 479235 676688 479247
rect 679696 479235 679702 479247
rect 679754 479235 679760 479287
rect 650032 478125 650038 478177
rect 650090 478165 650096 478177
rect 679888 478165 679894 478177
rect 650090 478137 679894 478165
rect 650090 478125 650096 478137
rect 679888 478125 679894 478137
rect 679946 478125 679952 478177
rect 41584 429211 41590 429263
rect 41642 429251 41648 429263
rect 53200 429251 53206 429263
rect 41642 429223 53206 429251
rect 41642 429211 41648 429223
rect 53200 429211 53206 429223
rect 53258 429211 53264 429263
rect 673840 429137 673846 429189
rect 673898 429177 673904 429189
rect 675280 429177 675286 429189
rect 673898 429149 675286 429177
rect 673898 429137 673904 429149
rect 675280 429137 675286 429149
rect 675338 429137 675344 429189
rect 41776 428915 41782 428967
rect 41834 428955 41840 428967
rect 50320 428955 50326 428967
rect 41834 428927 50326 428955
rect 41834 428915 41840 428927
rect 50320 428915 50326 428927
rect 50378 428915 50384 428967
rect 41776 428323 41782 428375
rect 41834 428363 41840 428375
rect 48016 428363 48022 428375
rect 41834 428335 48022 428363
rect 41834 428323 41840 428335
rect 48016 428323 48022 428335
rect 48074 428323 48080 428375
rect 41776 427953 41782 428005
rect 41834 427993 41840 428005
rect 43312 427993 43318 428005
rect 41834 427965 43318 427993
rect 41834 427953 41840 427965
rect 43312 427953 43318 427965
rect 43370 427953 43376 428005
rect 41776 427361 41782 427413
rect 41834 427401 41840 427413
rect 43408 427401 43414 427413
rect 41834 427373 43414 427401
rect 41834 427361 41840 427373
rect 43408 427361 43414 427373
rect 43466 427361 43472 427413
rect 41680 427213 41686 427265
rect 41738 427253 41744 427265
rect 45328 427253 45334 427265
rect 41738 427225 45334 427253
rect 41738 427213 41744 427225
rect 45328 427213 45334 427225
rect 45386 427213 45392 427265
rect 41776 426843 41782 426895
rect 41834 426883 41840 426895
rect 43312 426883 43318 426895
rect 41834 426855 43318 426883
rect 41834 426843 41840 426855
rect 43312 426843 43318 426855
rect 43370 426843 43376 426895
rect 41776 420405 41782 420457
rect 41834 420445 41840 420457
rect 45520 420445 45526 420457
rect 41834 420417 45526 420445
rect 41834 420405 41840 420417
rect 45520 420405 45526 420417
rect 45578 420405 45584 420457
rect 41776 419073 41782 419125
rect 41834 419113 41840 419125
rect 42832 419113 42838 419125
rect 41834 419085 42838 419113
rect 41834 419073 41840 419085
rect 42832 419073 42838 419085
rect 42890 419073 42896 419125
rect 41776 418555 41782 418607
rect 41834 418595 41840 418607
rect 43120 418595 43126 418607
rect 41834 418567 43126 418595
rect 41834 418555 41840 418567
rect 43120 418555 43126 418567
rect 43178 418555 43184 418607
rect 41584 417815 41590 417867
rect 41642 417855 41648 417867
rect 42928 417855 42934 417867
rect 41642 417827 42934 417855
rect 41642 417815 41648 417827
rect 42928 417815 42934 417827
rect 42986 417815 42992 417867
rect 41776 417741 41782 417793
rect 41834 417781 41840 417793
rect 43024 417781 43030 417793
rect 41834 417753 43030 417781
rect 41834 417741 41840 417753
rect 43024 417741 43030 417753
rect 43082 417741 43088 417793
rect 41776 416927 41782 416979
rect 41834 416967 41840 416979
rect 47920 416967 47926 416979
rect 41834 416939 47926 416967
rect 41834 416927 41840 416939
rect 47920 416927 47926 416939
rect 47978 416927 47984 416979
rect 41776 413375 41782 413427
rect 41834 413375 41840 413427
rect 41794 413205 41822 413375
rect 41776 413153 41782 413205
rect 41834 413153 41840 413205
rect 42832 409823 42838 409875
rect 42890 409863 42896 409875
rect 43216 409863 43222 409875
rect 42890 409835 43222 409863
rect 42890 409823 42896 409835
rect 43216 409823 43222 409835
rect 43274 409823 43280 409875
rect 42160 409675 42166 409727
rect 42218 409715 42224 409727
rect 42832 409715 42838 409727
rect 42218 409687 42838 409715
rect 42218 409675 42224 409687
rect 42832 409675 42838 409687
rect 42890 409675 42896 409727
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42928 409493 42934 409505
rect 42218 409465 42934 409493
rect 42218 409453 42224 409465
rect 42928 409453 42934 409465
rect 42986 409453 42992 409505
rect 42928 409305 42934 409357
rect 42986 409345 42992 409357
rect 43120 409345 43126 409357
rect 42986 409317 43126 409345
rect 42986 409305 42992 409317
rect 43120 409305 43126 409317
rect 43178 409305 43184 409357
rect 43216 409009 43222 409061
rect 43274 409049 43280 409061
rect 43408 409049 43414 409061
rect 43274 409021 43414 409049
rect 43274 409009 43280 409021
rect 43408 409009 43414 409021
rect 43466 409009 43472 409061
rect 42064 408047 42070 408099
rect 42122 408087 42128 408099
rect 43024 408087 43030 408099
rect 42122 408059 43030 408087
rect 42122 408047 42128 408059
rect 43024 408047 43030 408059
rect 43082 408047 43088 408099
rect 42160 407973 42166 408025
rect 42218 407973 42224 408025
rect 42178 407865 42206 407973
rect 42928 407865 42934 407877
rect 42178 407837 42934 407865
rect 42928 407825 42934 407837
rect 42986 407825 42992 407877
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 43120 407495 43126 407507
rect 42122 407467 43126 407495
rect 42122 407455 42128 407467
rect 43120 407455 43126 407467
rect 43178 407455 43184 407507
rect 42160 406863 42166 406915
rect 42218 406903 42224 406915
rect 43024 406903 43030 406915
rect 42218 406875 43030 406903
rect 42218 406863 42224 406875
rect 43024 406863 43030 406875
rect 43082 406863 43088 406915
rect 42832 406049 42838 406101
rect 42890 406089 42896 406101
rect 58480 406089 58486 406101
rect 42890 406061 58486 406089
rect 42890 406049 42896 406061
rect 58480 406049 58486 406061
rect 58538 406049 58544 406101
rect 42928 402571 42934 402623
rect 42986 402611 42992 402623
rect 59344 402611 59350 402623
rect 42986 402583 59350 402611
rect 42986 402571 42992 402583
rect 59344 402571 59350 402583
rect 59402 402571 59408 402623
rect 655120 400573 655126 400625
rect 655178 400613 655184 400625
rect 676144 400613 676150 400625
rect 655178 400585 676150 400613
rect 655178 400573 655184 400585
rect 676144 400573 676150 400585
rect 676202 400573 676208 400625
rect 655504 400499 655510 400551
rect 655562 400539 655568 400551
rect 676240 400539 676246 400551
rect 655562 400511 676246 400539
rect 655562 400499 655568 400511
rect 676240 400499 676246 400511
rect 676298 400499 676304 400551
rect 655312 400425 655318 400477
rect 655370 400465 655376 400477
rect 676048 400465 676054 400477
rect 655370 400437 676054 400465
rect 655370 400425 655376 400437
rect 676048 400425 676054 400437
rect 676106 400425 676112 400477
rect 673360 400351 673366 400403
rect 673418 400391 673424 400403
rect 676240 400391 676246 400403
rect 673418 400363 676246 400391
rect 673418 400351 673424 400363
rect 676240 400351 676246 400363
rect 676298 400351 676304 400403
rect 53200 400277 53206 400329
rect 53258 400317 53264 400329
rect 59728 400317 59734 400329
rect 53258 400289 59734 400317
rect 53258 400277 53264 400289
rect 59728 400277 59734 400289
rect 59786 400277 59792 400329
rect 50320 400203 50326 400255
rect 50378 400243 50384 400255
rect 59536 400243 59542 400255
rect 50378 400215 59542 400243
rect 50378 400203 50384 400215
rect 59536 400203 59542 400215
rect 59594 400203 59600 400255
rect 48016 400129 48022 400181
rect 48074 400169 48080 400181
rect 59632 400169 59638 400181
rect 48074 400141 59638 400169
rect 48074 400129 48080 400141
rect 59632 400129 59638 400141
rect 59690 400129 59696 400181
rect 672496 400129 672502 400181
rect 672554 400169 672560 400181
rect 673840 400169 673846 400181
rect 672554 400141 673846 400169
rect 672554 400129 672560 400141
rect 673840 400129 673846 400141
rect 673898 400169 673904 400181
rect 676048 400169 676054 400181
rect 673898 400141 676054 400169
rect 673898 400129 673904 400141
rect 676048 400129 676054 400141
rect 676106 400129 676112 400181
rect 673072 397983 673078 398035
rect 673130 398023 673136 398035
rect 675952 398023 675958 398035
rect 673130 397995 675958 398023
rect 673130 397983 673136 397995
rect 675952 397983 675958 397995
rect 676010 397983 676016 398035
rect 675184 397909 675190 397961
rect 675242 397949 675248 397961
rect 676624 397949 676630 397961
rect 675242 397921 676630 397949
rect 675242 397909 675248 397921
rect 676624 397909 676630 397921
rect 676682 397909 676688 397961
rect 674512 397687 674518 397739
rect 674570 397727 674576 397739
rect 676048 397727 676054 397739
rect 674570 397699 676054 397727
rect 674570 397687 674576 397699
rect 676048 397687 676054 397699
rect 676106 397687 676112 397739
rect 673168 395541 673174 395593
rect 673226 395581 673232 395593
rect 676048 395581 676054 395593
rect 673226 395553 676054 395581
rect 673226 395541 673232 395553
rect 676048 395541 676054 395553
rect 676106 395541 676112 395593
rect 42064 394505 42070 394557
rect 42122 394545 42128 394557
rect 57712 394545 57718 394557
rect 42122 394517 57718 394545
rect 42122 394505 42128 394517
rect 57712 394505 57718 394517
rect 57770 394505 57776 394557
rect 650128 388807 650134 388859
rect 650186 388847 650192 388859
rect 679792 388847 679798 388859
rect 650186 388819 679798 388847
rect 650186 388807 650192 388819
rect 679792 388807 679798 388819
rect 679850 388807 679856 388859
rect 41776 386439 41782 386491
rect 41834 386479 41840 386491
rect 53200 386479 53206 386491
rect 41834 386451 53206 386479
rect 41834 386439 41840 386451
rect 53200 386439 53206 386451
rect 53258 386439 53264 386491
rect 673264 385847 673270 385899
rect 673322 385887 673328 385899
rect 674512 385887 674518 385899
rect 673322 385859 674518 385887
rect 673322 385847 673328 385859
rect 674512 385847 674518 385859
rect 674570 385847 674576 385899
rect 41584 385699 41590 385751
rect 41642 385739 41648 385751
rect 50320 385739 50326 385751
rect 41642 385711 50326 385739
rect 41642 385699 41648 385711
rect 50320 385699 50326 385711
rect 50378 385699 50384 385751
rect 41776 385329 41782 385381
rect 41834 385369 41840 385381
rect 48112 385369 48118 385381
rect 41834 385341 48118 385369
rect 41834 385329 41840 385341
rect 48112 385329 48118 385341
rect 48170 385329 48176 385381
rect 41584 385181 41590 385233
rect 41642 385221 41648 385233
rect 43216 385221 43222 385233
rect 41642 385193 43222 385221
rect 41642 385181 41648 385193
rect 43216 385181 43222 385193
rect 43274 385181 43280 385233
rect 41776 384367 41782 384419
rect 41834 384407 41840 384419
rect 43504 384407 43510 384419
rect 41834 384379 43510 384407
rect 41834 384367 41840 384379
rect 43504 384367 43510 384379
rect 43562 384367 43568 384419
rect 41776 383479 41782 383531
rect 41834 383519 41840 383531
rect 43312 383519 43318 383531
rect 41834 383491 43318 383519
rect 41834 383479 41840 383491
rect 43312 383479 43318 383491
rect 43370 383519 43376 383531
rect 45424 383519 45430 383531
rect 43370 383491 45430 383519
rect 43370 383479 43376 383491
rect 45424 383479 45430 383491
rect 45482 383479 45488 383531
rect 653776 381629 653782 381681
rect 653834 381669 653840 381681
rect 675088 381669 675094 381681
rect 653834 381641 675094 381669
rect 653834 381629 653840 381641
rect 675088 381629 675094 381641
rect 675146 381629 675152 381681
rect 34480 381555 34486 381607
rect 34538 381595 34544 381607
rect 43312 381595 43318 381607
rect 34538 381567 43318 381595
rect 34538 381555 34544 381567
rect 43312 381555 43318 381567
rect 43370 381555 43376 381607
rect 652336 381555 652342 381607
rect 652394 381595 652400 381607
rect 674992 381595 674998 381607
rect 652394 381567 674998 381595
rect 652394 381555 652400 381567
rect 674992 381555 674998 381567
rect 675050 381555 675056 381607
rect 40240 377189 40246 377241
rect 40298 377229 40304 377241
rect 45616 377229 45622 377241
rect 40298 377201 45622 377229
rect 40298 377189 40304 377201
rect 45616 377189 45622 377201
rect 45674 377189 45680 377241
rect 41776 376893 41782 376945
rect 41834 376933 41840 376945
rect 42928 376933 42934 376945
rect 41834 376905 42934 376933
rect 41834 376893 41840 376905
rect 42928 376893 42934 376905
rect 42986 376893 42992 376945
rect 41776 374747 41782 374799
rect 41834 374787 41840 374799
rect 43024 374787 43030 374799
rect 41834 374759 43030 374787
rect 41834 374747 41840 374759
rect 43024 374747 43030 374759
rect 43082 374747 43088 374799
rect 41584 374599 41590 374651
rect 41642 374639 41648 374651
rect 42832 374639 42838 374651
rect 41642 374611 42838 374639
rect 41642 374599 41648 374611
rect 42832 374599 42838 374611
rect 42890 374599 42896 374651
rect 39280 374303 39286 374355
rect 39338 374343 39344 374355
rect 41776 374343 41782 374355
rect 39338 374315 41782 374343
rect 39338 374303 39344 374315
rect 41776 374303 41782 374315
rect 41834 374303 41840 374355
rect 39664 374229 39670 374281
rect 39722 374269 39728 374281
rect 43120 374269 43126 374281
rect 39722 374241 43126 374269
rect 39722 374229 39728 374241
rect 43120 374229 43126 374241
rect 43178 374229 43184 374281
rect 41872 373859 41878 373911
rect 41930 373899 41936 373911
rect 48016 373899 48022 373911
rect 41930 373871 48022 373899
rect 41930 373859 41936 373871
rect 48016 373859 48022 373871
rect 48074 373859 48080 373911
rect 673168 372083 673174 372135
rect 673226 372123 673232 372135
rect 675376 372123 675382 372135
rect 673226 372095 675382 372123
rect 673226 372083 673232 372095
rect 675376 372083 675382 372095
rect 675434 372083 675440 372135
rect 41776 370159 41782 370211
rect 41834 370159 41840 370211
rect 41794 369989 41822 370159
rect 41776 369937 41782 369989
rect 41834 369937 41840 369989
rect 42928 366681 42934 366733
rect 42986 366721 42992 366733
rect 43216 366721 43222 366733
rect 42986 366693 43222 366721
rect 42986 366681 42992 366693
rect 43216 366681 43222 366693
rect 43274 366681 43280 366733
rect 42160 366533 42166 366585
rect 42218 366573 42224 366585
rect 42928 366573 42934 366585
rect 42218 366545 42934 366573
rect 42218 366533 42224 366545
rect 42928 366533 42934 366545
rect 42986 366533 42992 366585
rect 42064 366237 42070 366289
rect 42122 366277 42128 366289
rect 43120 366277 43126 366289
rect 42122 366249 43126 366277
rect 42122 366237 42128 366249
rect 43120 366237 43126 366249
rect 43178 366237 43184 366289
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 42832 365019 42838 365031
rect 42218 364991 42838 365019
rect 42218 364979 42224 364991
rect 42832 364979 42838 364991
rect 42890 364979 42896 365031
rect 42064 364683 42070 364735
rect 42122 364723 42128 364735
rect 42832 364723 42838 364735
rect 42122 364695 42838 364723
rect 42122 364683 42128 364695
rect 42832 364683 42838 364695
rect 42890 364683 42896 364735
rect 42064 364239 42070 364291
rect 42122 364279 42128 364291
rect 43120 364279 43126 364291
rect 42122 364251 43126 364279
rect 42122 364239 42128 364251
rect 43120 364239 43126 364251
rect 43178 364239 43184 364291
rect 42160 363795 42166 363847
rect 42218 363835 42224 363847
rect 43024 363835 43030 363847
rect 42218 363807 43030 363835
rect 42218 363795 42224 363807
rect 43024 363795 43030 363807
rect 43082 363795 43088 363847
rect 42928 361427 42934 361479
rect 42986 361467 42992 361479
rect 58480 361467 58486 361479
rect 42986 361439 58486 361467
rect 42986 361427 42992 361439
rect 58480 361427 58486 361439
rect 58538 361427 58544 361479
rect 42832 359947 42838 359999
rect 42890 359987 42896 359999
rect 59152 359987 59158 359999
rect 42890 359959 59158 359987
rect 42890 359947 42896 359959
rect 59152 359947 59158 359959
rect 59210 359947 59216 359999
rect 655120 357135 655126 357187
rect 655178 357175 655184 357187
rect 676240 357175 676246 357187
rect 655178 357147 676246 357175
rect 655178 357135 655184 357147
rect 676240 357135 676246 357147
rect 676298 357135 676304 357187
rect 53200 357061 53206 357113
rect 53258 357101 53264 357113
rect 58384 357101 58390 357113
rect 53258 357073 58390 357101
rect 53258 357061 53264 357073
rect 58384 357061 58390 357073
rect 58442 357061 58448 357113
rect 50320 356987 50326 357039
rect 50378 357027 50384 357039
rect 58480 357027 58486 357039
rect 50378 356999 58486 357027
rect 50378 356987 50384 356999
rect 58480 356987 58486 356999
rect 58538 356987 58544 357039
rect 48112 356913 48118 356965
rect 48170 356953 48176 356965
rect 59632 356953 59638 356965
rect 48170 356925 59638 356953
rect 48170 356913 48176 356925
rect 59632 356913 59638 356925
rect 59690 356913 59696 356965
rect 673360 356173 673366 356225
rect 673418 356213 673424 356225
rect 676240 356213 676246 356225
rect 673418 356185 676246 356213
rect 673418 356173 673424 356185
rect 676240 356173 676246 356185
rect 676298 356173 676304 356225
rect 673264 354767 673270 354819
rect 673322 354807 673328 354819
rect 675952 354807 675958 354819
rect 673322 354779 675958 354807
rect 673322 354767 673328 354779
rect 675952 354767 675958 354779
rect 676010 354767 676016 354819
rect 672592 354397 672598 354449
rect 672650 354437 672656 354449
rect 673264 354437 673270 354449
rect 672650 354409 673270 354437
rect 672650 354397 672656 354409
rect 673264 354397 673270 354409
rect 673322 354397 673328 354449
rect 655312 354323 655318 354375
rect 655370 354363 655376 354375
rect 676048 354363 676054 354375
rect 655370 354335 676054 354363
rect 655370 354323 655376 354335
rect 676048 354323 676054 354335
rect 676106 354323 676112 354375
rect 655216 354249 655222 354301
rect 655274 354289 655280 354301
rect 676144 354289 676150 354301
rect 655274 354261 676150 354289
rect 655274 354249 655280 354261
rect 676144 354249 676150 354261
rect 676202 354249 676208 354301
rect 672784 353879 672790 353931
rect 672842 353919 672848 353931
rect 676048 353919 676054 353931
rect 672842 353891 676054 353919
rect 672842 353879 672848 353891
rect 676048 353879 676054 353891
rect 676106 353879 676112 353931
rect 42160 351289 42166 351341
rect 42218 351329 42224 351341
rect 57712 351329 57718 351341
rect 42218 351301 57718 351329
rect 42218 351289 42224 351301
rect 57712 351289 57718 351301
rect 57770 351289 57776 351341
rect 674416 348625 674422 348677
rect 674474 348665 674480 348677
rect 675952 348665 675958 348677
rect 674474 348637 675958 348665
rect 674474 348625 674480 348637
rect 675952 348625 675958 348637
rect 676010 348625 676016 348677
rect 675280 348551 675286 348603
rect 675338 348591 675344 348603
rect 676240 348591 676246 348603
rect 675338 348563 676246 348591
rect 675338 348551 675344 348563
rect 676240 348551 676246 348563
rect 676298 348551 676304 348603
rect 675184 348477 675190 348529
rect 675242 348517 675248 348529
rect 676048 348517 676054 348529
rect 675242 348489 676054 348517
rect 675242 348477 675248 348489
rect 676048 348477 676054 348489
rect 676106 348477 676112 348529
rect 674800 347515 674806 347567
rect 674858 347555 674864 347567
rect 676048 347555 676054 347567
rect 674858 347527 676054 347555
rect 674858 347515 674864 347527
rect 676048 347515 676054 347527
rect 676106 347515 676112 347567
rect 674896 345739 674902 345791
rect 674954 345779 674960 345791
rect 676144 345779 676150 345791
rect 674954 345751 676150 345779
rect 674954 345739 674960 345751
rect 676144 345739 676150 345751
rect 676202 345739 676208 345791
rect 674992 345665 674998 345717
rect 675050 345705 675056 345717
rect 676240 345705 676246 345717
rect 675050 345677 676246 345705
rect 675050 345665 675056 345677
rect 676240 345665 676246 345677
rect 676298 345665 676304 345717
rect 675088 345591 675094 345643
rect 675146 345631 675152 345643
rect 676048 345631 676054 345643
rect 675146 345603 676054 345631
rect 675146 345591 675152 345603
rect 676048 345591 676054 345603
rect 676106 345591 676112 345643
rect 41584 343223 41590 343275
rect 41642 343263 41648 343275
rect 53200 343263 53206 343275
rect 41642 343235 53206 343263
rect 41642 343223 41648 343235
rect 53200 343223 53206 343235
rect 53258 343223 53264 343275
rect 41776 342853 41782 342905
rect 41834 342893 41840 342905
rect 50320 342893 50326 342905
rect 41834 342865 50326 342893
rect 41834 342853 41840 342865
rect 50320 342853 50326 342865
rect 50378 342853 50384 342905
rect 650224 342705 650230 342757
rect 650282 342745 650288 342757
rect 679696 342745 679702 342757
rect 650282 342717 679702 342745
rect 650282 342705 650288 342717
rect 679696 342705 679702 342717
rect 679754 342705 679760 342757
rect 41776 342335 41782 342387
rect 41834 342375 41840 342387
rect 48112 342375 48118 342387
rect 41834 342347 48118 342375
rect 41834 342335 41840 342347
rect 48112 342335 48118 342347
rect 48170 342335 48176 342387
rect 41776 341965 41782 342017
rect 41834 342005 41840 342017
rect 43504 342005 43510 342017
rect 41834 341977 43510 342005
rect 41834 341965 41840 341977
rect 43504 341965 43510 341977
rect 43562 341965 43568 342017
rect 41776 341373 41782 341425
rect 41834 341413 41840 341425
rect 43216 341413 43222 341425
rect 41834 341385 43222 341413
rect 41834 341373 41840 341385
rect 43216 341373 43222 341385
rect 43274 341373 43280 341425
rect 675760 341373 675766 341425
rect 675818 341373 675824 341425
rect 41776 340855 41782 340907
rect 41834 340895 41840 340907
rect 43408 340895 43414 340907
rect 41834 340867 43414 340895
rect 41834 340855 41840 340867
rect 43408 340855 43414 340867
rect 43466 340855 43472 340907
rect 675778 340759 675806 341373
rect 675760 340707 675766 340759
rect 675818 340707 675824 340759
rect 666640 340633 666646 340685
rect 666698 340673 666704 340685
rect 675472 340673 675478 340685
rect 666698 340645 675478 340673
rect 666698 340633 666704 340645
rect 675472 340633 675478 340645
rect 675530 340633 675536 340685
rect 41776 340485 41782 340537
rect 41834 340525 41840 340537
rect 43312 340525 43318 340537
rect 41834 340497 43318 340525
rect 41834 340485 41840 340497
rect 43312 340485 43318 340497
rect 43370 340525 43376 340537
rect 45712 340525 45718 340537
rect 43370 340497 45718 340525
rect 43370 340485 43376 340497
rect 45712 340485 45718 340497
rect 45770 340485 45776 340537
rect 45616 339933 45622 339945
rect 44962 339905 45622 339933
rect 41776 339819 41782 339871
rect 41834 339859 41840 339871
rect 43600 339859 43606 339871
rect 41834 339831 43606 339859
rect 41834 339819 41840 339831
rect 43600 339819 43606 339831
rect 43658 339819 43664 339871
rect 41584 339745 41590 339797
rect 41642 339785 41648 339797
rect 44962 339785 44990 339905
rect 45616 339893 45622 339905
rect 45674 339933 45680 339945
rect 62608 339933 62614 339945
rect 45674 339905 62614 339933
rect 45674 339893 45680 339905
rect 62608 339893 62614 339905
rect 62666 339893 62672 339945
rect 41642 339757 44990 339785
rect 41642 339745 41648 339757
rect 675184 337229 675190 337281
rect 675242 337269 675248 337281
rect 675472 337269 675478 337281
rect 675242 337241 675478 337269
rect 675242 337229 675248 337241
rect 675472 337229 675478 337241
rect 675530 337229 675536 337281
rect 674416 336563 674422 336615
rect 674474 336603 674480 336615
rect 675376 336603 675382 336615
rect 674474 336575 675382 336603
rect 674474 336563 674480 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 675088 336045 675094 336097
rect 675146 336085 675152 336097
rect 675376 336085 675382 336097
rect 675146 336057 675382 336085
rect 675146 336045 675152 336057
rect 675376 336045 675382 336057
rect 675434 336045 675440 336097
rect 41776 333085 41782 333137
rect 41834 333125 41840 333137
rect 42736 333125 42742 333137
rect 41834 333097 42742 333125
rect 41834 333085 41840 333097
rect 42736 333085 42742 333097
rect 42794 333085 42800 333137
rect 674992 332715 674998 332767
rect 675050 332755 675056 332767
rect 675376 332755 675382 332767
rect 675050 332727 675382 332755
rect 675050 332715 675056 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 674800 332197 674806 332249
rect 674858 332237 674864 332249
rect 675472 332237 675478 332249
rect 674858 332209 675478 332237
rect 674858 332197 674864 332209
rect 675472 332197 675478 332209
rect 675530 332197 675536 332249
rect 674896 331753 674902 331805
rect 674954 331793 674960 331805
rect 675376 331793 675382 331805
rect 674954 331765 675382 331793
rect 674954 331753 674960 331765
rect 675376 331753 675382 331765
rect 675434 331753 675440 331805
rect 41776 331531 41782 331583
rect 41834 331571 41840 331583
rect 42928 331571 42934 331583
rect 41834 331543 42934 331571
rect 41834 331531 41840 331543
rect 42928 331531 42934 331543
rect 42986 331531 42992 331583
rect 41872 330939 41878 330991
rect 41930 330979 41936 330991
rect 48208 330979 48214 330991
rect 41930 330951 48214 330979
rect 41930 330939 41936 330951
rect 48208 330939 48214 330951
rect 48266 330939 48272 330991
rect 41584 328719 41590 328771
rect 41642 328759 41648 328771
rect 43024 328759 43030 328771
rect 41642 328731 43030 328759
rect 41642 328719 41648 328731
rect 43024 328719 43030 328731
rect 43082 328719 43088 328771
rect 654160 328275 654166 328327
rect 654218 328315 654224 328327
rect 666640 328315 666646 328327
rect 654218 328287 666646 328315
rect 654218 328275 654224 328287
rect 666640 328275 666646 328287
rect 666698 328275 666704 328327
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326625 41822 327017
rect 41776 326573 41782 326625
rect 41834 326573 41840 326625
rect 42928 325759 42934 325811
rect 42986 325799 42992 325811
rect 43120 325799 43126 325811
rect 42986 325771 43126 325799
rect 42986 325759 42992 325771
rect 43120 325759 43126 325771
rect 43178 325759 43184 325811
rect 42064 323317 42070 323369
rect 42122 323357 42128 323369
rect 42448 323357 42454 323369
rect 42122 323329 42454 323357
rect 42122 323317 42128 323329
rect 42448 323317 42454 323329
rect 42506 323317 42512 323369
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 43024 323135 43030 323147
rect 42218 323107 43030 323135
rect 42218 323095 42224 323107
rect 43024 323095 43030 323107
rect 43082 323095 43088 323147
rect 41968 321615 41974 321667
rect 42026 321655 42032 321667
rect 43120 321655 43126 321667
rect 42026 321627 43126 321655
rect 42026 321615 42032 321627
rect 43120 321615 43126 321627
rect 43178 321615 43184 321667
rect 42160 321467 42166 321519
rect 42218 321507 42224 321519
rect 43120 321507 43126 321519
rect 42218 321479 43126 321507
rect 42218 321467 42224 321479
rect 43120 321467 43126 321479
rect 43178 321467 43184 321519
rect 42160 321245 42166 321297
rect 42218 321285 42224 321297
rect 43024 321285 43030 321297
rect 42218 321257 43030 321285
rect 42218 321245 42224 321257
rect 43024 321245 43030 321257
rect 43082 321245 43088 321297
rect 42448 319617 42454 319669
rect 42506 319657 42512 319669
rect 58480 319657 58486 319669
rect 42506 319629 58486 319657
rect 42506 319617 42512 319629
rect 58480 319617 58486 319629
rect 58538 319617 58544 319669
rect 43120 316731 43126 316783
rect 43178 316771 43184 316783
rect 59152 316771 59158 316783
rect 43178 316743 59158 316771
rect 43178 316731 43184 316743
rect 59152 316731 59158 316743
rect 59210 316731 59216 316783
rect 53200 313845 53206 313897
rect 53258 313885 53264 313897
rect 59728 313885 59734 313897
rect 53258 313857 59734 313885
rect 53258 313845 53264 313857
rect 59728 313845 59734 313857
rect 59786 313845 59792 313897
rect 50320 313771 50326 313823
rect 50378 313811 50384 313823
rect 59536 313811 59542 313823
rect 50378 313783 59542 313811
rect 50378 313771 50384 313783
rect 59536 313771 59542 313783
rect 59594 313771 59600 313823
rect 48112 313697 48118 313749
rect 48170 313737 48176 313749
rect 59632 313737 59638 313749
rect 48170 313709 59638 313737
rect 48170 313697 48176 313709
rect 59632 313697 59638 313709
rect 59690 313697 59696 313749
rect 654256 311181 654262 311233
rect 654314 311221 654320 311233
rect 676240 311221 676246 311233
rect 654314 311193 676246 311221
rect 654314 311181 654320 311193
rect 676240 311181 676246 311193
rect 676298 311181 676304 311233
rect 654160 311107 654166 311159
rect 654218 311147 654224 311159
rect 676144 311147 676150 311159
rect 654218 311119 676150 311147
rect 654218 311107 654224 311119
rect 676144 311107 676150 311119
rect 676202 311107 676208 311159
rect 654064 311033 654070 311085
rect 654122 311073 654128 311085
rect 676336 311073 676342 311085
rect 654122 311045 676342 311073
rect 654122 311033 654128 311045
rect 676336 311033 676342 311045
rect 676394 311033 676400 311085
rect 42160 308073 42166 308125
rect 42218 308113 42224 308125
rect 59056 308113 59062 308125
rect 42218 308085 59062 308113
rect 42218 308073 42224 308085
rect 59056 308073 59062 308085
rect 59114 308073 59120 308125
rect 45520 307777 45526 307829
rect 45578 307817 45584 307829
rect 46096 307817 46102 307829
rect 45578 307789 46102 307817
rect 45578 307777 45584 307789
rect 46096 307777 46102 307789
rect 46154 307777 46160 307829
rect 674608 305335 674614 305387
rect 674666 305375 674672 305387
rect 676048 305375 676054 305387
rect 674666 305347 676054 305375
rect 674666 305335 674672 305347
rect 676048 305335 676054 305347
rect 676106 305335 676112 305387
rect 675088 305261 675094 305313
rect 675146 305301 675152 305313
rect 676240 305301 676246 305313
rect 675146 305273 676246 305301
rect 675146 305261 675152 305273
rect 676240 305261 676246 305273
rect 676298 305261 676304 305313
rect 674224 302597 674230 302649
rect 674282 302637 674288 302649
rect 675952 302637 675958 302649
rect 674282 302609 675958 302637
rect 674282 302597 674288 302609
rect 675952 302597 675958 302609
rect 676010 302597 676016 302649
rect 674416 302523 674422 302575
rect 674474 302563 674480 302575
rect 676048 302563 676054 302575
rect 674474 302535 676054 302563
rect 674474 302523 674480 302535
rect 676048 302523 676054 302535
rect 676106 302523 676112 302575
rect 674704 302449 674710 302501
rect 674762 302489 674768 302501
rect 676240 302489 676246 302501
rect 674762 302461 676246 302489
rect 674762 302449 674768 302461
rect 676240 302449 676246 302461
rect 676298 302449 676304 302501
rect 674896 302375 674902 302427
rect 674954 302415 674960 302427
rect 676048 302415 676054 302427
rect 674954 302387 676054 302415
rect 674954 302375 674960 302387
rect 676048 302375 676054 302387
rect 676106 302375 676112 302427
rect 46096 302301 46102 302353
rect 46154 302341 46160 302353
rect 54640 302341 54646 302353
rect 46154 302313 54646 302341
rect 46154 302301 46160 302313
rect 54640 302301 54646 302313
rect 54698 302301 54704 302353
rect 43408 300895 43414 300947
rect 43466 300935 43472 300947
rect 44272 300935 44278 300947
rect 43466 300907 44278 300935
rect 43466 300895 43472 300907
rect 44272 300895 44278 300907
rect 44330 300935 44336 300947
rect 62896 300935 62902 300947
rect 44330 300907 62902 300935
rect 44330 300895 44336 300907
rect 62896 300895 62902 300907
rect 62954 300895 62960 300947
rect 41776 299711 41782 299763
rect 41834 299751 41840 299763
rect 50704 299751 50710 299763
rect 41834 299723 50710 299751
rect 41834 299711 41840 299723
rect 50704 299711 50710 299723
rect 50762 299711 50768 299763
rect 650320 299711 650326 299763
rect 650378 299751 650384 299763
rect 679984 299751 679990 299763
rect 650378 299723 679990 299751
rect 650378 299711 650384 299723
rect 679984 299711 679990 299723
rect 680042 299711 680048 299763
rect 41872 299637 41878 299689
rect 41930 299677 41936 299689
rect 44272 299677 44278 299689
rect 41930 299649 44278 299677
rect 41930 299637 41936 299649
rect 44272 299637 44278 299649
rect 44330 299637 44336 299689
rect 674320 299637 674326 299689
rect 674378 299677 674384 299689
rect 676048 299677 676054 299689
rect 674378 299649 676054 299677
rect 674378 299637 674384 299649
rect 676048 299637 676054 299649
rect 676106 299637 676112 299689
rect 41584 299563 41590 299615
rect 41642 299603 41648 299615
rect 60208 299603 60214 299615
rect 41642 299575 60214 299603
rect 41642 299563 41648 299575
rect 60208 299563 60214 299575
rect 60266 299563 60272 299615
rect 674992 299563 674998 299615
rect 675050 299603 675056 299615
rect 676240 299603 676246 299615
rect 675050 299575 676246 299603
rect 675050 299563 675056 299575
rect 676240 299563 676246 299575
rect 676298 299563 676304 299615
rect 41776 298749 41782 298801
rect 41834 298789 41840 298801
rect 43216 298789 43222 298801
rect 41834 298761 43222 298789
rect 41834 298749 41840 298761
rect 43216 298749 43222 298761
rect 43274 298749 43280 298801
rect 41776 298157 41782 298209
rect 41834 298197 41840 298209
rect 43408 298197 43414 298209
rect 41834 298169 43414 298197
rect 41834 298157 41840 298169
rect 43408 298157 43414 298169
rect 43466 298157 43472 298209
rect 43600 298083 43606 298135
rect 43658 298123 43664 298135
rect 62992 298123 62998 298135
rect 43658 298095 62998 298123
rect 43658 298083 43664 298095
rect 62992 298083 62998 298095
rect 63050 298083 63056 298135
rect 41776 297639 41782 297691
rect 41834 297679 41840 297691
rect 43216 297679 43222 297691
rect 41834 297651 43222 297679
rect 41834 297639 41840 297651
rect 43216 297639 43222 297651
rect 43274 297639 43280 297691
rect 39856 296751 39862 296803
rect 39914 296791 39920 296803
rect 43600 296791 43606 296803
rect 39914 296763 43606 296791
rect 39914 296751 39920 296763
rect 43600 296751 43606 296763
rect 43658 296751 43664 296803
rect 41776 296677 41782 296729
rect 41834 296717 41840 296729
rect 43312 296717 43318 296729
rect 41834 296689 43318 296717
rect 41834 296677 41840 296689
rect 43312 296677 43318 296689
rect 43370 296677 43376 296729
rect 674704 295419 674710 295471
rect 674762 295459 674768 295471
rect 675088 295459 675094 295471
rect 674762 295431 675094 295459
rect 674762 295419 674768 295431
rect 675088 295419 675094 295431
rect 675146 295419 675152 295471
rect 674608 294753 674614 294805
rect 674666 294793 674672 294805
rect 675088 294793 675094 294805
rect 674666 294765 675094 294793
rect 674666 294753 674672 294765
rect 675088 294753 675094 294765
rect 675146 294753 675152 294805
rect 53296 293865 53302 293917
rect 53354 293905 53360 293917
rect 59248 293905 59254 293917
rect 53354 293877 59254 293905
rect 53354 293865 53360 293877
rect 59248 293865 59254 293877
rect 59306 293865 59312 293917
rect 56176 293791 56182 293843
rect 56234 293831 56240 293843
rect 60304 293831 60310 293843
rect 56234 293803 60310 293831
rect 56234 293791 56240 293803
rect 60304 293791 60310 293803
rect 60362 293791 60368 293843
rect 39664 293717 39670 293769
rect 39722 293757 39728 293769
rect 58192 293757 58198 293769
rect 39722 293729 58198 293757
rect 39722 293717 39728 293729
rect 58192 293717 58198 293729
rect 58250 293717 58256 293769
rect 674416 292237 674422 292289
rect 674474 292277 674480 292289
rect 675472 292277 675478 292289
rect 674474 292249 675478 292277
rect 674474 292237 674480 292249
rect 675472 292237 675478 292249
rect 675530 292237 675536 292289
rect 674224 291571 674230 291623
rect 674282 291611 674288 291623
rect 675376 291611 675382 291623
rect 674282 291583 675382 291611
rect 674282 291571 674288 291583
rect 675376 291571 675382 291583
rect 675434 291571 675440 291623
rect 674896 291053 674902 291105
rect 674954 291093 674960 291105
rect 675376 291093 675382 291105
rect 674954 291065 675382 291093
rect 674954 291053 674960 291065
rect 675376 291053 675382 291065
rect 675434 291053 675440 291105
rect 48304 290979 48310 291031
rect 48362 291019 48368 291031
rect 59632 291019 59638 291031
rect 48362 290991 59638 291019
rect 48362 290979 48368 290991
rect 59632 290979 59638 290991
rect 59690 290979 59696 291031
rect 54640 290905 54646 290957
rect 54698 290945 54704 290957
rect 54698 290917 54782 290945
rect 54698 290905 54704 290917
rect 54754 290871 54782 290917
rect 58768 290871 58774 290883
rect 54754 290843 58774 290871
rect 58768 290831 58774 290843
rect 58826 290831 58832 290883
rect 41776 289351 41782 289403
rect 41834 289391 41840 289403
rect 43120 289391 43126 289403
rect 41834 289363 43126 289391
rect 41834 289351 41840 289363
rect 43120 289351 43126 289363
rect 43178 289351 43184 289403
rect 50704 288907 50710 288959
rect 50762 288947 50768 288959
rect 59536 288947 59542 288959
rect 50762 288919 59542 288947
rect 50762 288907 50768 288919
rect 59536 288907 59542 288919
rect 59594 288907 59600 288959
rect 41776 288167 41782 288219
rect 41834 288207 41840 288219
rect 42928 288207 42934 288219
rect 41834 288179 42934 288207
rect 41834 288167 41840 288179
rect 42928 288167 42934 288179
rect 42986 288167 42992 288219
rect 50320 288019 50326 288071
rect 50378 288059 50384 288071
rect 59152 288059 59158 288071
rect 50378 288031 59158 288059
rect 50378 288019 50384 288031
rect 59152 288019 59158 288031
rect 59210 288019 59216 288071
rect 41872 287723 41878 287775
rect 41930 287763 41936 287775
rect 45808 287763 45814 287775
rect 41930 287735 45814 287763
rect 41930 287723 41936 287735
rect 45808 287723 45814 287735
rect 45866 287723 45872 287775
rect 674320 287723 674326 287775
rect 674378 287763 674384 287775
rect 675376 287763 675382 287775
rect 674378 287735 675382 287763
rect 674378 287723 674384 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 674992 286761 674998 286813
rect 675050 286801 675056 286813
rect 675376 286801 675382 286813
rect 675050 286773 675382 286801
rect 675050 286761 675056 286773
rect 675376 286761 675382 286773
rect 675434 286761 675440 286813
rect 41584 285133 41590 285185
rect 41642 285173 41648 285185
rect 42928 285173 42934 285185
rect 41642 285145 42934 285173
rect 41642 285133 41648 285145
rect 42928 285133 42934 285145
rect 42986 285133 42992 285185
rect 53200 285133 53206 285185
rect 53258 285173 53264 285185
rect 59248 285173 59254 285185
rect 53258 285145 59254 285173
rect 53258 285133 53264 285145
rect 59248 285133 59254 285145
rect 59306 285133 59312 285185
rect 653776 284097 653782 284149
rect 653834 284137 653840 284149
rect 658000 284137 658006 284149
rect 653834 284109 658006 284137
rect 653834 284097 653840 284109
rect 658000 284097 658006 284109
rect 658058 284097 658064 284149
rect 41776 283801 41782 283853
rect 41834 283801 41840 283853
rect 41794 283557 41822 283801
rect 41776 283505 41782 283557
rect 41834 283505 41840 283557
rect 45328 282395 45334 282447
rect 45386 282435 45392 282447
rect 53008 282435 53014 282447
rect 45386 282407 53014 282435
rect 45386 282395 45392 282407
rect 53008 282395 53014 282407
rect 53066 282395 53072 282447
rect 56080 282395 56086 282447
rect 56138 282435 56144 282447
rect 57616 282435 57622 282447
rect 56138 282407 57622 282435
rect 56138 282395 56144 282407
rect 57616 282395 57622 282407
rect 57674 282395 57680 282447
rect 45520 282321 45526 282373
rect 45578 282361 45584 282373
rect 59632 282361 59638 282373
rect 45578 282333 59638 282361
rect 45578 282321 45584 282333
rect 59632 282321 59638 282333
rect 59690 282321 59696 282373
rect 48112 282247 48118 282299
rect 48170 282287 48176 282299
rect 58576 282287 58582 282299
rect 48170 282259 58582 282287
rect 48170 282247 48176 282259
rect 58576 282247 58582 282259
rect 58634 282247 58640 282299
rect 58768 282247 58774 282299
rect 58826 282287 58832 282299
rect 58826 282259 60542 282287
rect 58826 282247 58832 282259
rect 60514 282213 60542 282259
rect 63376 282213 63382 282225
rect 60514 282185 63382 282213
rect 63376 282173 63382 282185
rect 63434 282173 63440 282225
rect 42064 280101 42070 280153
rect 42122 280141 42128 280153
rect 42832 280141 42838 280153
rect 42122 280113 42838 280141
rect 42122 280101 42128 280113
rect 42832 280101 42838 280113
rect 42890 280101 42896 280153
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 42928 279919 42934 279931
rect 42218 279891 42934 279919
rect 42218 279879 42224 279891
rect 42928 279879 42934 279891
rect 42986 279879 42992 279931
rect 45328 279435 45334 279487
rect 45386 279475 45392 279487
rect 58384 279475 58390 279487
rect 45386 279447 58390 279475
rect 45386 279435 45392 279447
rect 58384 279435 58390 279447
rect 58442 279435 58448 279487
rect 654256 279435 654262 279487
rect 654314 279475 654320 279487
rect 663760 279475 663766 279487
rect 654314 279447 663766 279475
rect 654314 279435 654320 279447
rect 663760 279435 663766 279447
rect 663818 279435 663824 279487
rect 45616 279361 45622 279413
rect 45674 279401 45680 279413
rect 58576 279401 58582 279413
rect 45674 279373 58582 279401
rect 45674 279361 45680 279373
rect 58576 279361 58582 279373
rect 58634 279361 58640 279413
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 43024 278587 43030 278599
rect 42218 278559 43030 278587
rect 42218 278547 42224 278559
rect 43024 278547 43030 278559
rect 43082 278547 43088 278599
rect 42064 278473 42070 278525
rect 42122 278513 42128 278525
rect 42928 278513 42934 278525
rect 42122 278485 42934 278513
rect 42122 278473 42128 278485
rect 42928 278473 42934 278485
rect 42986 278473 42992 278525
rect 314896 278325 314902 278377
rect 314954 278365 314960 278377
rect 408304 278365 408310 278377
rect 314954 278337 408310 278365
rect 314954 278325 314960 278337
rect 408304 278325 408310 278337
rect 408362 278325 408368 278377
rect 381040 278251 381046 278303
rect 381098 278291 381104 278303
rect 571408 278291 571414 278303
rect 381098 278263 571414 278291
rect 381098 278251 381104 278263
rect 571408 278251 571414 278263
rect 571466 278251 571472 278303
rect 319504 278177 319510 278229
rect 319562 278217 319568 278229
rect 418960 278217 418966 278229
rect 319562 278189 418966 278217
rect 319562 278177 319568 278189
rect 418960 278177 418966 278189
rect 419018 278177 419024 278229
rect 320944 278103 320950 278155
rect 321002 278143 321008 278155
rect 422512 278143 422518 278155
rect 321002 278115 422518 278143
rect 321002 278103 321008 278115
rect 422512 278103 422518 278115
rect 422570 278103 422576 278155
rect 386512 278029 386518 278081
rect 386570 278069 386576 278081
rect 585616 278069 585622 278081
rect 386570 278041 585622 278069
rect 386570 278029 386576 278041
rect 585616 278029 585622 278041
rect 585674 278029 585680 278081
rect 53008 277955 53014 278007
rect 53066 277995 53072 278007
rect 138256 277995 138262 278007
rect 53066 277967 138262 277995
rect 53066 277955 53072 277967
rect 138256 277955 138262 277967
rect 138314 277955 138320 278007
rect 323824 277955 323830 278007
rect 323882 277995 323888 278007
rect 429616 277995 429622 278007
rect 323882 277967 429622 277995
rect 323882 277955 323888 277967
rect 429616 277955 429622 277967
rect 429674 277955 429680 278007
rect 63376 277881 63382 277933
rect 63434 277921 63440 277933
rect 382384 277921 382390 277933
rect 63434 277893 382390 277921
rect 63434 277881 63440 277893
rect 382384 277881 382390 277893
rect 382442 277881 382448 277933
rect 408880 277881 408886 277933
rect 408938 277921 408944 277933
rect 672496 277921 672502 277933
rect 408938 277893 672502 277921
rect 408938 277881 408944 277893
rect 672496 277881 672502 277893
rect 672554 277881 672560 277933
rect 326416 277807 326422 277859
rect 326474 277847 326480 277859
rect 437008 277847 437014 277859
rect 326474 277819 437014 277847
rect 326474 277807 326480 277819
rect 437008 277807 437014 277819
rect 437066 277807 437072 277859
rect 317872 277733 317878 277785
rect 317930 277773 317936 277785
rect 415696 277773 415702 277785
rect 317930 277745 415702 277773
rect 317930 277733 317936 277745
rect 415696 277733 415702 277745
rect 415754 277733 415760 277785
rect 329296 277659 329302 277711
rect 329354 277699 329360 277711
rect 444112 277699 444118 277711
rect 329354 277671 444118 277699
rect 329354 277659 329360 277671
rect 444112 277659 444118 277671
rect 444170 277659 444176 277711
rect 332368 277585 332374 277637
rect 332426 277625 332432 277637
rect 451216 277625 451222 277637
rect 332426 277597 451222 277625
rect 332426 277585 332432 277597
rect 451216 277585 451222 277597
rect 451274 277585 451280 277637
rect 334960 277511 334966 277563
rect 335018 277551 335024 277563
rect 458224 277551 458230 277563
rect 335018 277523 458230 277551
rect 335018 277511 335024 277523
rect 458224 277511 458230 277523
rect 458282 277511 458288 277563
rect 337840 277437 337846 277489
rect 337898 277477 337904 277489
rect 465328 277477 465334 277489
rect 337898 277449 465334 277477
rect 337898 277437 337904 277449
rect 465328 277437 465334 277449
rect 465386 277437 465392 277489
rect 341008 277363 341014 277415
rect 341066 277403 341072 277415
rect 472432 277403 472438 277415
rect 341066 277375 472438 277403
rect 341066 277363 341072 277375
rect 472432 277363 472438 277375
rect 472490 277363 472496 277415
rect 343888 277289 343894 277341
rect 343946 277329 343952 277341
rect 479536 277329 479542 277341
rect 343946 277301 479542 277329
rect 343946 277289 343952 277301
rect 479536 277289 479542 277301
rect 479594 277289 479600 277341
rect 42064 277215 42070 277267
rect 42122 277255 42128 277267
rect 43120 277255 43126 277267
rect 42122 277227 43126 277255
rect 42122 277215 42128 277227
rect 43120 277215 43126 277227
rect 43178 277215 43184 277267
rect 373840 277215 373846 277267
rect 373898 277255 373904 277267
rect 554032 277255 554038 277267
rect 373898 277227 554038 277255
rect 373898 277215 373904 277227
rect 554032 277215 554038 277227
rect 554090 277215 554096 277267
rect 375088 277141 375094 277193
rect 375146 277181 375152 277193
rect 557584 277181 557590 277193
rect 375146 277153 557590 277181
rect 375146 277141 375152 277153
rect 557584 277141 557590 277153
rect 557642 277141 557648 277193
rect 376816 277067 376822 277119
rect 376874 277107 376880 277119
rect 561136 277107 561142 277119
rect 376874 277079 561142 277107
rect 376874 277067 376880 277079
rect 561136 277067 561142 277079
rect 561194 277067 561200 277119
rect 377968 276993 377974 277045
rect 378026 277033 378032 277045
rect 564688 277033 564694 277045
rect 378026 277005 564694 277033
rect 378026 276993 378032 277005
rect 564688 276993 564694 277005
rect 564746 276993 564752 277045
rect 379408 276919 379414 276971
rect 379466 276959 379472 276971
rect 568240 276959 568246 276971
rect 379466 276931 568246 276959
rect 379466 276919 379472 276931
rect 568240 276919 568246 276931
rect 568298 276919 568304 276971
rect 316624 276845 316630 276897
rect 316682 276885 316688 276897
rect 412144 276885 412150 276897
rect 316682 276857 412150 276885
rect 316682 276845 316688 276857
rect 412144 276845 412150 276857
rect 412202 276845 412208 276897
rect 382288 276771 382294 276823
rect 382346 276811 382352 276823
rect 575248 276811 575254 276823
rect 382346 276783 575254 276811
rect 382346 276771 382352 276783
rect 575248 276771 575254 276783
rect 575306 276771 575312 276823
rect 383632 276697 383638 276749
rect 383690 276737 383696 276749
rect 578800 276737 578806 276749
rect 383690 276709 578806 276737
rect 383690 276697 383696 276709
rect 578800 276697 578806 276709
rect 578858 276697 578864 276749
rect 385360 276623 385366 276675
rect 385418 276663 385424 276675
rect 582352 276663 582358 276675
rect 385418 276635 582358 276663
rect 385418 276623 385424 276635
rect 582352 276623 582358 276635
rect 582410 276623 582416 276675
rect 675760 276623 675766 276675
rect 675818 276663 675824 276675
rect 679792 276663 679798 276675
rect 675818 276635 679798 276663
rect 675818 276623 675824 276635
rect 679792 276623 679798 276635
rect 679850 276623 679856 276675
rect 322096 276549 322102 276601
rect 322154 276589 322160 276601
rect 426352 276589 426358 276601
rect 322154 276561 426358 276589
rect 322154 276549 322160 276561
rect 426352 276549 426358 276561
rect 426410 276549 426416 276601
rect 387952 276475 387958 276527
rect 388010 276515 388016 276527
rect 589456 276515 589462 276527
rect 388010 276487 589462 276515
rect 388010 276475 388016 276487
rect 589456 276475 589462 276487
rect 589514 276475 589520 276527
rect 675280 276475 675286 276527
rect 675338 276515 675344 276527
rect 679696 276515 679702 276527
rect 675338 276487 679702 276515
rect 675338 276475 675344 276487
rect 679696 276475 679702 276487
rect 679754 276475 679760 276527
rect 42832 276401 42838 276453
rect 42890 276441 42896 276453
rect 53296 276441 53302 276453
rect 42890 276413 53302 276441
rect 42890 276401 42896 276413
rect 53296 276401 53302 276413
rect 53354 276401 53360 276453
rect 286096 276401 286102 276453
rect 286154 276441 286160 276453
rect 336496 276441 336502 276453
rect 286154 276413 336502 276441
rect 286154 276401 286160 276413
rect 336496 276401 336502 276413
rect 336554 276401 336560 276453
rect 356176 276401 356182 276453
rect 356234 276441 356240 276453
rect 510256 276441 510262 276453
rect 356234 276413 510262 276441
rect 356234 276401 356240 276413
rect 510256 276401 510262 276413
rect 510314 276401 510320 276453
rect 284464 276327 284470 276379
rect 284522 276367 284528 276379
rect 332944 276367 332950 276379
rect 284522 276339 332950 276367
rect 284522 276327 284528 276339
rect 332944 276327 332950 276339
rect 333002 276327 333008 276379
rect 359152 276327 359158 276379
rect 359210 276367 359216 276379
rect 517360 276367 517366 276379
rect 359210 276339 517366 276367
rect 359210 276327 359216 276339
rect 517360 276327 517366 276339
rect 517418 276327 517424 276379
rect 287344 276253 287350 276305
rect 287402 276293 287408 276305
rect 340048 276293 340054 276305
rect 287402 276265 340054 276293
rect 287402 276253 287408 276265
rect 340048 276253 340054 276265
rect 340106 276253 340112 276305
rect 361744 276253 361750 276305
rect 361802 276293 361808 276305
rect 524464 276293 524470 276305
rect 361802 276265 524470 276293
rect 361802 276253 361808 276265
rect 524464 276253 524470 276265
rect 524522 276253 524528 276305
rect 288688 276179 288694 276231
rect 288746 276219 288752 276231
rect 343600 276219 343606 276231
rect 288746 276191 343606 276219
rect 288746 276179 288752 276191
rect 343600 276179 343606 276191
rect 343658 276179 343664 276231
rect 364624 276179 364630 276231
rect 364682 276219 364688 276231
rect 531568 276219 531574 276231
rect 364682 276191 531574 276219
rect 364682 276179 364688 276191
rect 531568 276179 531574 276191
rect 531626 276179 531632 276231
rect 291856 276105 291862 276157
rect 291914 276145 291920 276157
rect 350704 276145 350710 276157
rect 291914 276117 350710 276145
rect 291914 276105 291920 276117
rect 350704 276105 350710 276117
rect 350762 276105 350768 276157
rect 367696 276105 367702 276157
rect 367754 276145 367760 276157
rect 538672 276145 538678 276157
rect 367754 276117 538678 276145
rect 367754 276105 367760 276117
rect 538672 276105 538678 276117
rect 538730 276105 538736 276157
rect 290320 276031 290326 276083
rect 290378 276071 290384 276083
rect 347152 276071 347158 276083
rect 290378 276043 347158 276071
rect 290378 276031 290384 276043
rect 347152 276031 347158 276043
rect 347210 276031 347216 276083
rect 371920 276031 371926 276083
rect 371978 276071 371984 276083
rect 549328 276071 549334 276083
rect 371978 276043 549334 276071
rect 371978 276031 371984 276043
rect 549328 276031 549334 276043
rect 549386 276031 549392 276083
rect 293008 275957 293014 276009
rect 293066 275997 293072 276009
rect 354256 275997 354262 276009
rect 293066 275969 354262 275997
rect 293066 275957 293072 275969
rect 354256 275957 354262 275969
rect 354314 275957 354320 276009
rect 371056 275957 371062 276009
rect 371114 275997 371120 276009
rect 546928 275997 546934 276009
rect 371114 275969 546934 275997
rect 371114 275957 371120 275969
rect 546928 275957 546934 275969
rect 546986 275957 546992 276009
rect 294640 275883 294646 275935
rect 294698 275923 294704 275935
rect 357808 275923 357814 275935
rect 294698 275895 357814 275923
rect 294698 275883 294704 275895
rect 357808 275883 357814 275895
rect 357866 275883 357872 275935
rect 370288 275883 370294 275935
rect 370346 275923 370352 275935
rect 545776 275923 545782 275935
rect 370346 275895 545782 275923
rect 370346 275883 370352 275895
rect 545776 275883 545782 275895
rect 545834 275883 545840 275935
rect 296464 275809 296470 275861
rect 296522 275849 296528 275861
rect 362512 275849 362518 275861
rect 296522 275821 362518 275849
rect 296522 275809 296528 275821
rect 362512 275809 362518 275821
rect 362570 275809 362576 275861
rect 373456 275809 373462 275861
rect 373514 275849 373520 275861
rect 552784 275849 552790 275861
rect 373514 275821 552790 275849
rect 373514 275809 373520 275821
rect 552784 275809 552790 275821
rect 552842 275809 552848 275861
rect 297328 275735 297334 275787
rect 297386 275775 297392 275787
rect 364912 275775 364918 275787
rect 297386 275747 364918 275775
rect 297386 275735 297392 275747
rect 364912 275735 364918 275747
rect 364970 275735 364976 275787
rect 374608 275735 374614 275787
rect 374666 275775 374672 275787
rect 556336 275775 556342 275787
rect 374666 275747 556342 275775
rect 374666 275735 374672 275747
rect 556336 275735 556342 275747
rect 556394 275735 556400 275787
rect 295888 275661 295894 275713
rect 295946 275701 295952 275713
rect 361360 275701 361366 275713
rect 295946 275673 361366 275701
rect 295946 275661 295952 275673
rect 361360 275661 361366 275673
rect 361418 275661 361424 275713
rect 377488 275661 377494 275713
rect 377546 275701 377552 275713
rect 563440 275701 563446 275713
rect 377546 275673 563446 275701
rect 377546 275661 377552 275673
rect 563440 275661 563446 275673
rect 563498 275661 563504 275713
rect 298960 275587 298966 275639
rect 299018 275627 299024 275639
rect 368464 275627 368470 275639
rect 299018 275599 368470 275627
rect 299018 275587 299024 275599
rect 368464 275587 368470 275599
rect 368522 275587 368528 275639
rect 376240 275587 376246 275639
rect 376298 275627 376304 275639
rect 559888 275627 559894 275639
rect 376298 275599 559894 275627
rect 376298 275587 376304 275599
rect 559888 275587 559894 275599
rect 559946 275587 559952 275639
rect 297808 275513 297814 275565
rect 297866 275553 297872 275565
rect 366064 275553 366070 275565
rect 297866 275525 366070 275553
rect 297866 275513 297872 275525
rect 366064 275513 366070 275525
rect 366122 275513 366128 275565
rect 380560 275513 380566 275565
rect 380618 275553 380624 275565
rect 570544 275553 570550 275565
rect 380618 275525 570550 275553
rect 380618 275513 380624 275525
rect 570544 275513 570550 275525
rect 570602 275513 570608 275565
rect 300208 275439 300214 275491
rect 300266 275479 300272 275491
rect 372016 275479 372022 275491
rect 300266 275451 372022 275479
rect 300266 275439 300272 275451
rect 372016 275439 372022 275451
rect 372074 275439 372080 275491
rect 381808 275439 381814 275491
rect 381866 275479 381872 275491
rect 574096 275479 574102 275491
rect 381866 275451 574102 275479
rect 381866 275439 381872 275451
rect 574096 275439 574102 275451
rect 574154 275439 574160 275491
rect 299152 275365 299158 275417
rect 299210 275405 299216 275417
rect 369616 275405 369622 275417
rect 299210 275377 369622 275405
rect 299210 275365 299216 275377
rect 369616 275365 369622 275377
rect 369674 275365 369680 275417
rect 388912 275365 388918 275417
rect 388970 275405 388976 275417
rect 591856 275405 591862 275417
rect 388970 275377 591862 275405
rect 388970 275365 388976 275377
rect 591856 275365 591862 275377
rect 591914 275365 591920 275417
rect 303280 275291 303286 275343
rect 303338 275331 303344 275343
rect 379120 275331 379126 275343
rect 303338 275303 379126 275331
rect 303338 275291 303344 275303
rect 379120 275291 379126 275303
rect 379178 275291 379184 275343
rect 389584 275291 389590 275343
rect 389642 275331 389648 275343
rect 593008 275331 593014 275343
rect 389642 275303 593014 275331
rect 389642 275291 389648 275303
rect 593008 275291 593014 275303
rect 593066 275291 593072 275343
rect 304432 275217 304438 275269
rect 304490 275257 304496 275269
rect 382576 275257 382582 275269
rect 304490 275229 382582 275257
rect 304490 275217 304496 275229
rect 382576 275217 382582 275229
rect 382634 275217 382640 275269
rect 391984 275217 391990 275269
rect 392042 275257 392048 275269
rect 598960 275257 598966 275269
rect 392042 275229 598966 275257
rect 392042 275217 392048 275229
rect 598960 275217 598966 275229
rect 599018 275217 599024 275269
rect 307312 275143 307318 275195
rect 307370 275183 307376 275195
rect 389680 275183 389686 275195
rect 307370 275155 389686 275183
rect 307370 275143 307376 275155
rect 389680 275143 389686 275155
rect 389738 275143 389744 275195
rect 396304 275143 396310 275195
rect 396362 275183 396368 275195
rect 609520 275183 609526 275195
rect 396362 275155 609526 275183
rect 396362 275143 396368 275155
rect 609520 275143 609526 275155
rect 609578 275143 609584 275195
rect 310384 275069 310390 275121
rect 310442 275109 310448 275121
rect 396784 275109 396790 275121
rect 310442 275081 396790 275109
rect 310442 275069 310448 275081
rect 396784 275069 396790 275081
rect 396842 275069 396848 275121
rect 401776 275069 401782 275121
rect 401834 275109 401840 275121
rect 623728 275109 623734 275121
rect 401834 275081 623734 275109
rect 401834 275069 401840 275081
rect 623728 275069 623734 275081
rect 623786 275069 623792 275121
rect 311632 274995 311638 275047
rect 311690 275035 311696 275047
rect 400336 275035 400342 275047
rect 311690 275007 400342 275035
rect 311690 274995 311696 275007
rect 400336 274995 400342 275007
rect 400394 274995 400400 275047
rect 404944 274995 404950 275047
rect 405002 275035 405008 275047
rect 630832 275035 630838 275047
rect 405002 275007 630838 275035
rect 405002 274995 405008 275007
rect 630832 274995 630838 275007
rect 630890 274995 630896 275047
rect 283024 274921 283030 274973
rect 283082 274961 283088 274973
rect 329392 274961 329398 274973
rect 283082 274933 329398 274961
rect 283082 274921 283088 274933
rect 329392 274921 329398 274933
rect 329450 274921 329456 274973
rect 344560 274921 344566 274973
rect 344618 274961 344624 274973
rect 481936 274961 481942 274973
rect 344618 274933 481942 274961
rect 344618 274921 344624 274933
rect 481936 274921 481942 274933
rect 481994 274921 482000 274973
rect 281776 274847 281782 274899
rect 281834 274887 281840 274899
rect 325840 274887 325846 274899
rect 281834 274859 325846 274887
rect 281834 274847 281840 274859
rect 325840 274847 325846 274859
rect 325898 274847 325904 274899
rect 339088 274847 339094 274899
rect 339146 274887 339152 274899
rect 467728 274887 467734 274899
rect 339146 274859 467734 274887
rect 339146 274847 339152 274859
rect 467728 274847 467734 274859
rect 467786 274847 467792 274899
rect 336016 274773 336022 274825
rect 336074 274813 336080 274825
rect 460624 274813 460630 274825
rect 336074 274785 460630 274813
rect 336074 274773 336080 274785
rect 460624 274773 460630 274785
rect 460682 274773 460688 274825
rect 333136 274699 333142 274751
rect 333194 274739 333200 274751
rect 453520 274739 453526 274751
rect 333194 274711 453526 274739
rect 333194 274699 333200 274711
rect 453520 274699 453526 274711
rect 453578 274699 453584 274751
rect 330448 274625 330454 274677
rect 330506 274665 330512 274677
rect 446416 274665 446422 274677
rect 330506 274637 446422 274665
rect 330506 274625 330512 274637
rect 446416 274625 446422 274637
rect 446474 274625 446480 274677
rect 328816 274551 328822 274603
rect 328874 274591 328880 274603
rect 442864 274591 442870 274603
rect 328874 274563 442870 274591
rect 328874 274551 328880 274563
rect 442864 274551 442870 274563
rect 442922 274551 442928 274603
rect 325936 274477 325942 274529
rect 325994 274517 326000 274529
rect 435856 274517 435862 274529
rect 325994 274489 435862 274517
rect 325994 274477 326000 274489
rect 435856 274477 435862 274489
rect 435914 274477 435920 274529
rect 323344 274403 323350 274455
rect 323402 274443 323408 274455
rect 428752 274443 428758 274455
rect 323402 274415 428758 274443
rect 323402 274403 323408 274415
rect 428752 274403 428758 274415
rect 428810 274403 428816 274455
rect 320176 274329 320182 274381
rect 320234 274369 320240 274381
rect 421648 274369 421654 274381
rect 320234 274341 421654 274369
rect 320234 274329 320240 274341
rect 421648 274329 421654 274341
rect 421706 274329 421712 274381
rect 315952 274255 315958 274307
rect 316010 274295 316016 274307
rect 410992 274295 410998 274307
rect 316010 274267 410998 274295
rect 316010 274255 316016 274267
rect 410992 274255 410998 274267
rect 411050 274255 411056 274307
rect 317296 274181 317302 274233
rect 317354 274221 317360 274233
rect 414544 274221 414550 274233
rect 317354 274193 414550 274221
rect 317354 274181 317360 274193
rect 414544 274181 414550 274193
rect 414602 274181 414608 274233
rect 314704 274107 314710 274159
rect 314762 274147 314768 274159
rect 407440 274147 407446 274159
rect 314762 274119 407446 274147
rect 314762 274107 314768 274119
rect 407440 274107 407446 274119
rect 407498 274107 407504 274159
rect 348496 274033 348502 274085
rect 348554 274073 348560 274085
rect 401488 274073 401494 274085
rect 348554 274045 401494 274073
rect 348554 274033 348560 274045
rect 401488 274033 401494 274045
rect 401546 274033 401552 274085
rect 341200 273959 341206 274011
rect 341258 273999 341264 274011
rect 387376 273999 387382 274011
rect 341258 273971 387382 273999
rect 341258 273959 341264 273971
rect 387376 273959 387382 273971
rect 387434 273959 387440 274011
rect 326800 273885 326806 273937
rect 326858 273925 326864 273937
rect 373168 273925 373174 273937
rect 326858 273897 373174 273925
rect 326858 273885 326864 273897
rect 373168 273885 373174 273897
rect 373226 273885 373232 273937
rect 334288 273811 334294 273863
rect 334346 273851 334352 273863
rect 380272 273851 380278 273863
rect 334346 273823 380278 273851
rect 334346 273811 334352 273823
rect 380272 273811 380278 273823
rect 380330 273811 380336 273863
rect 347056 273737 347062 273789
rect 347114 273777 347120 273789
rect 394480 273777 394486 273789
rect 347114 273749 394486 273777
rect 347114 273737 347120 273749
rect 394480 273737 394486 273749
rect 394538 273737 394544 273789
rect 331216 273663 331222 273715
rect 331274 273703 331280 273715
rect 376720 273703 376726 273715
rect 331274 273675 376726 273703
rect 331274 273663 331280 273675
rect 376720 273663 376726 273675
rect 376778 273663 376784 273715
rect 305218 273601 307070 273629
rect 42928 273515 42934 273567
rect 42986 273555 42992 273567
rect 56176 273555 56182 273567
rect 42986 273527 56182 273555
rect 42986 273515 42992 273527
rect 56176 273515 56182 273527
rect 56234 273515 56240 273567
rect 160432 273515 160438 273567
rect 160490 273555 160496 273567
rect 207472 273555 207478 273567
rect 160490 273527 207478 273555
rect 160490 273515 160496 273527
rect 207472 273515 207478 273527
rect 207530 273515 207536 273567
rect 230128 273515 230134 273567
rect 230186 273555 230192 273567
rect 242896 273555 242902 273567
rect 230186 273527 242902 273555
rect 230186 273515 230192 273527
rect 242896 273515 242902 273527
rect 242954 273515 242960 273567
rect 270256 273515 270262 273567
rect 270314 273555 270320 273567
rect 297520 273555 297526 273567
rect 270314 273527 297526 273555
rect 270314 273515 270320 273527
rect 297520 273515 297526 273527
rect 297578 273515 297584 273567
rect 299344 273515 299350 273567
rect 299402 273555 299408 273567
rect 305218 273555 305246 273601
rect 299402 273527 305246 273555
rect 299402 273515 299408 273527
rect 305296 273515 305302 273567
rect 305354 273555 305360 273567
rect 306928 273555 306934 273567
rect 305354 273527 306934 273555
rect 305354 273515 305360 273527
rect 306928 273515 306934 273527
rect 306986 273515 306992 273567
rect 307042 273555 307070 273601
rect 406576 273589 406582 273641
rect 406634 273629 406640 273641
rect 406634 273601 512702 273629
rect 406634 273589 406640 273601
rect 327088 273555 327094 273567
rect 307042 273527 327094 273555
rect 327088 273515 327094 273527
rect 327146 273515 327152 273567
rect 349456 273515 349462 273567
rect 349514 273555 349520 273567
rect 493744 273555 493750 273567
rect 349514 273527 493750 273555
rect 349514 273515 349520 273527
rect 493744 273515 493750 273527
rect 493802 273515 493808 273567
rect 512674 273555 512702 273601
rect 635536 273555 635542 273567
rect 512674 273527 635542 273555
rect 635536 273515 635542 273527
rect 635594 273515 635600 273567
rect 130864 273441 130870 273493
rect 130922 273481 130928 273493
rect 192976 273481 192982 273493
rect 130922 273453 192982 273481
rect 130922 273441 130928 273453
rect 192976 273441 192982 273453
rect 193034 273441 193040 273493
rect 195856 273441 195862 273493
rect 195914 273481 195920 273493
rect 221488 273481 221494 273493
rect 195914 273453 221494 273481
rect 195914 273441 195920 273453
rect 221488 273441 221494 273453
rect 221546 273441 221552 273493
rect 275344 273441 275350 273493
rect 275402 273481 275408 273493
rect 310480 273481 310486 273493
rect 275402 273453 310486 273481
rect 275402 273441 275408 273453
rect 310480 273441 310486 273453
rect 310538 273441 310544 273493
rect 310576 273441 310582 273493
rect 310634 273481 310640 273493
rect 344752 273481 344758 273493
rect 310634 273453 344758 273481
rect 310634 273441 310640 273453
rect 344752 273441 344758 273453
rect 344810 273441 344816 273493
rect 350032 273441 350038 273493
rect 350090 273481 350096 273493
rect 494896 273481 494902 273493
rect 350090 273453 494902 273481
rect 350090 273441 350096 273453
rect 494896 273441 494902 273453
rect 494954 273441 494960 273493
rect 526960 273441 526966 273493
rect 527018 273481 527024 273493
rect 624976 273481 624982 273493
rect 527018 273453 624982 273481
rect 527018 273441 527024 273453
rect 624976 273441 624982 273453
rect 625034 273441 625040 273493
rect 142672 273367 142678 273419
rect 142730 273407 142736 273419
rect 208144 273407 208150 273419
rect 142730 273379 208150 273407
rect 142730 273367 142736 273379
rect 208144 273367 208150 273379
rect 208202 273367 208208 273419
rect 219568 273367 219574 273419
rect 219626 273407 219632 273419
rect 238672 273407 238678 273419
rect 219626 273379 238678 273407
rect 219626 273367 219632 273379
rect 238672 273367 238678 273379
rect 238730 273367 238736 273419
rect 277072 273367 277078 273419
rect 277130 273407 277136 273419
rect 314032 273407 314038 273419
rect 277130 273379 314038 273407
rect 277130 273367 277136 273379
rect 314032 273367 314038 273379
rect 314090 273367 314096 273419
rect 352432 273367 352438 273419
rect 352490 273407 352496 273419
rect 500848 273407 500854 273419
rect 352490 273379 500854 273407
rect 352490 273367 352496 273379
rect 500848 273367 500854 273379
rect 500906 273367 500912 273419
rect 133264 273293 133270 273345
rect 133322 273333 133328 273345
rect 135280 273333 135286 273345
rect 133322 273305 135286 273333
rect 133322 273293 133328 273305
rect 135280 273293 135286 273305
rect 135338 273293 135344 273345
rect 135568 273293 135574 273345
rect 135626 273333 135632 273345
rect 209776 273333 209782 273345
rect 135626 273305 209782 273333
rect 135626 273293 135632 273305
rect 209776 273293 209782 273305
rect 209834 273293 209840 273345
rect 279664 273293 279670 273345
rect 279722 273333 279728 273345
rect 321136 273333 321142 273345
rect 279722 273305 321142 273333
rect 279722 273293 279728 273305
rect 321136 273293 321142 273305
rect 321194 273293 321200 273345
rect 352624 273293 352630 273345
rect 352682 273333 352688 273345
rect 502000 273333 502006 273345
rect 352682 273305 502006 273333
rect 352682 273293 352688 273305
rect 502000 273293 502006 273305
rect 502058 273293 502064 273345
rect 68272 273219 68278 273271
rect 68330 273259 68336 273271
rect 142576 273259 142582 273271
rect 68330 273231 142582 273259
rect 68330 273219 68336 273231
rect 142576 273219 142582 273231
rect 142634 273219 142640 273271
rect 153328 273219 153334 273271
rect 153386 273259 153392 273271
rect 207376 273259 207382 273271
rect 153386 273231 207382 273259
rect 153386 273219 153392 273231
rect 207376 273219 207382 273231
rect 207434 273219 207440 273271
rect 278224 273219 278230 273271
rect 278282 273259 278288 273271
rect 317584 273259 317590 273271
rect 278282 273231 317590 273259
rect 278282 273219 278288 273231
rect 317584 273219 317590 273231
rect 317642 273219 317648 273271
rect 355504 273219 355510 273271
rect 355562 273259 355568 273271
rect 509104 273259 509110 273271
rect 355562 273231 509110 273259
rect 355562 273219 355568 273231
rect 509104 273219 509110 273231
rect 509162 273219 509168 273271
rect 132016 273145 132022 273197
rect 132074 273185 132080 273197
rect 209872 273185 209878 273197
rect 132074 273157 209878 273185
rect 132074 273145 132080 273157
rect 209872 273145 209878 273157
rect 209930 273145 209936 273197
rect 218320 273145 218326 273197
rect 218378 273185 218384 273197
rect 238096 273185 238102 273197
rect 218378 273157 238102 273185
rect 218378 273145 218384 273157
rect 238096 273145 238102 273157
rect 238154 273145 238160 273197
rect 285616 273145 285622 273197
rect 285674 273185 285680 273197
rect 335344 273185 335350 273197
rect 285674 273157 335350 273185
rect 285674 273145 285680 273157
rect 335344 273145 335350 273157
rect 335402 273145 335408 273197
rect 355024 273145 355030 273197
rect 355082 273185 355088 273197
rect 507952 273185 507958 273197
rect 355082 273157 507958 273185
rect 355082 273145 355088 273157
rect 507952 273145 507958 273157
rect 508010 273145 508016 273197
rect 508240 273145 508246 273197
rect 508298 273185 508304 273197
rect 555184 273185 555190 273197
rect 508298 273157 555190 273185
rect 508298 273145 508304 273157
rect 555184 273145 555190 273157
rect 555242 273145 555248 273197
rect 127312 273071 127318 273123
rect 127370 273111 127376 273123
rect 209968 273111 209974 273123
rect 127370 273083 209974 273111
rect 127370 273071 127376 273083
rect 209968 273071 209974 273083
rect 210026 273071 210032 273123
rect 216016 273071 216022 273123
rect 216074 273111 216080 273123
rect 236944 273111 236950 273123
rect 216074 273083 236950 273111
rect 216074 273071 216080 273083
rect 236944 273071 236950 273083
rect 237002 273071 237008 273123
rect 286768 273071 286774 273123
rect 286826 273111 286832 273123
rect 286826 273083 306398 273111
rect 286826 273071 286832 273083
rect 128464 272997 128470 273049
rect 128522 273037 128528 273049
rect 210160 273037 210166 273049
rect 128522 273009 210166 273037
rect 128522 272997 128528 273009
rect 210160 272997 210166 273009
rect 210218 272997 210224 273049
rect 220720 272997 220726 273049
rect 220778 273037 220784 273049
rect 239152 273037 239158 273049
rect 220778 273009 239158 273037
rect 220778 272997 220784 273009
rect 239152 272997 239158 273009
rect 239210 272997 239216 273049
rect 289936 272997 289942 273049
rect 289994 273037 290000 273049
rect 306370 273037 306398 273083
rect 306640 273071 306646 273123
rect 306698 273111 306704 273123
rect 334192 273111 334198 273123
rect 306698 273083 334198 273111
rect 306698 273071 306704 273083
rect 334192 273071 334198 273083
rect 334250 273071 334256 273123
rect 358576 273071 358582 273123
rect 358634 273111 358640 273123
rect 358634 273083 375038 273111
rect 358634 273071 358640 273083
rect 338896 273037 338902 273049
rect 289994 273009 306302 273037
rect 306370 273009 338902 273037
rect 289994 272997 290000 273009
rect 123760 272923 123766 272975
rect 123818 272963 123824 272975
rect 209008 272963 209014 272975
rect 123818 272935 209014 272963
rect 123818 272923 123824 272935
rect 209008 272923 209014 272935
rect 209066 272923 209072 272975
rect 217168 272923 217174 272975
rect 217226 272963 217232 272975
rect 237616 272963 237622 272975
rect 217226 272935 237622 272963
rect 217226 272923 217232 272935
rect 237616 272923 237622 272935
rect 237674 272923 237680 272975
rect 274192 272923 274198 272975
rect 274250 272963 274256 272975
rect 305296 272963 305302 272975
rect 274250 272935 305302 272963
rect 274250 272923 274256 272935
rect 305296 272923 305302 272935
rect 305354 272923 305360 272975
rect 306274 272963 306302 273009
rect 338896 272997 338902 273009
rect 338954 272997 338960 273049
rect 360976 272997 360982 273049
rect 361034 273037 361040 273049
rect 375010 273037 375038 273083
rect 375184 273071 375190 273123
rect 375242 273111 375248 273123
rect 514960 273111 514966 273123
rect 375242 273083 514966 273111
rect 375242 273071 375248 273083
rect 514960 273071 514966 273083
rect 515018 273071 515024 273123
rect 516208 273037 516214 273049
rect 361034 273009 374942 273037
rect 375010 273009 516214 273037
rect 361034 272997 361040 273009
rect 306274 272935 306782 272963
rect 116656 272849 116662 272901
rect 116714 272889 116720 272901
rect 207088 272889 207094 272901
rect 116714 272861 207094 272889
rect 116714 272849 116720 272861
rect 207088 272849 207094 272861
rect 207146 272849 207152 272901
rect 213616 272849 213622 272901
rect 213674 272889 213680 272901
rect 236272 272889 236278 272901
rect 213674 272861 236278 272889
rect 213674 272849 213680 272861
rect 236272 272849 236278 272861
rect 236330 272849 236336 272901
rect 292240 272849 292246 272901
rect 292298 272889 292304 272901
rect 306754 272889 306782 272935
rect 306832 272923 306838 272975
rect 306890 272963 306896 272975
rect 358960 272963 358966 272975
rect 306890 272935 358966 272963
rect 306890 272923 306896 272935
rect 358960 272923 358966 272935
rect 359018 272923 359024 272975
rect 361264 272923 361270 272975
rect 361322 272963 361328 272975
rect 374914 272963 374942 273009
rect 516208 272997 516214 273009
rect 516266 272997 516272 273049
rect 522064 272963 522070 272975
rect 361322 272935 374846 272963
rect 374914 272935 522070 272963
rect 361322 272923 361328 272935
rect 346000 272889 346006 272901
rect 292298 272861 306686 272889
rect 306754 272861 346006 272889
rect 292298 272849 292304 272861
rect 120208 272775 120214 272827
rect 120266 272815 120272 272827
rect 207856 272815 207862 272827
rect 120266 272787 207862 272815
rect 120266 272775 120272 272787
rect 207856 272775 207862 272787
rect 207914 272775 207920 272827
rect 212464 272775 212470 272827
rect 212522 272815 212528 272827
rect 235696 272815 235702 272827
rect 212522 272787 235702 272815
rect 212522 272775 212528 272787
rect 235696 272775 235702 272787
rect 235754 272775 235760 272827
rect 292720 272775 292726 272827
rect 292778 272815 292784 272827
rect 306658 272815 306686 272861
rect 346000 272849 346006 272861
rect 346058 272849 346064 272901
rect 363568 272849 363574 272901
rect 363626 272889 363632 272901
rect 374818 272889 374846 272935
rect 522064 272923 522070 272935
rect 522122 272923 522128 272975
rect 523312 272889 523318 272901
rect 363626 272861 374750 272889
rect 374818 272861 523318 272889
rect 363626 272849 363632 272861
rect 351856 272815 351862 272827
rect 292778 272787 306590 272815
rect 306658 272787 351862 272815
rect 292778 272775 292784 272787
rect 113104 272701 113110 272753
rect 113162 272741 113168 272753
rect 206224 272741 206230 272753
rect 113162 272713 206230 272741
rect 113162 272701 113168 272713
rect 206224 272701 206230 272713
rect 206282 272701 206288 272753
rect 211216 272701 211222 272753
rect 211274 272741 211280 272753
rect 235024 272741 235030 272753
rect 211274 272713 235030 272741
rect 211274 272701 211280 272713
rect 235024 272701 235030 272713
rect 235082 272701 235088 272753
rect 295408 272701 295414 272753
rect 295466 272741 295472 272753
rect 295466 272713 296654 272741
rect 295466 272701 295472 272713
rect 110800 272627 110806 272679
rect 110858 272667 110864 272679
rect 205456 272667 205462 272679
rect 110858 272639 205462 272667
rect 110858 272627 110864 272639
rect 205456 272627 205462 272639
rect 205514 272627 205520 272679
rect 214768 272627 214774 272679
rect 214826 272667 214832 272679
rect 236464 272667 236470 272679
rect 214826 272639 236470 272667
rect 214826 272627 214832 272639
rect 236464 272627 236470 272639
rect 236522 272627 236528 272679
rect 296626 272667 296654 272713
rect 298288 272701 298294 272753
rect 298346 272741 298352 272753
rect 306562 272741 306590 272787
rect 351856 272775 351862 272787
rect 351914 272775 351920 272827
rect 364144 272775 364150 272827
rect 364202 272815 364208 272827
rect 374722 272815 374750 272861
rect 523312 272849 523318 272861
rect 523370 272849 523376 272901
rect 523984 272849 523990 272901
rect 524042 272889 524048 272901
rect 639088 272889 639094 272901
rect 524042 272861 639094 272889
rect 524042 272849 524048 272861
rect 639088 272849 639094 272861
rect 639146 272849 639152 272901
rect 529168 272815 529174 272827
rect 364202 272787 374654 272815
rect 374722 272787 529174 272815
rect 364202 272775 364208 272787
rect 353104 272741 353110 272753
rect 298346 272713 302174 272741
rect 306562 272713 353110 272741
rect 298346 272701 298352 272713
rect 302032 272667 302038 272679
rect 296626 272639 302038 272667
rect 302032 272627 302038 272639
rect 302090 272627 302096 272679
rect 106096 272553 106102 272605
rect 106154 272593 106160 272605
rect 204016 272593 204022 272605
rect 106154 272565 204022 272593
rect 106154 272553 106160 272565
rect 204016 272553 204022 272565
rect 204074 272553 204080 272605
rect 208912 272553 208918 272605
rect 208970 272593 208976 272605
rect 234352 272593 234358 272605
rect 208970 272565 234358 272593
rect 208970 272553 208976 272565
rect 234352 272553 234358 272565
rect 234410 272553 234416 272605
rect 270544 272553 270550 272605
rect 270602 272593 270608 272605
rect 298672 272593 298678 272605
rect 270602 272565 298678 272593
rect 270602 272553 270608 272565
rect 298672 272553 298678 272565
rect 298730 272553 298736 272605
rect 301360 272553 301366 272605
rect 301418 272593 301424 272605
rect 302146 272593 302174 272713
rect 353104 272701 353110 272713
rect 353162 272701 353168 272753
rect 366544 272701 366550 272753
rect 366602 272741 366608 272753
rect 374512 272741 374518 272753
rect 366602 272713 374518 272741
rect 366602 272701 366608 272713
rect 374512 272701 374518 272713
rect 374570 272701 374576 272753
rect 374626 272741 374654 272787
rect 529168 272775 529174 272787
rect 529226 272775 529232 272827
rect 530416 272741 530422 272753
rect 374626 272713 530422 272741
rect 530416 272701 530422 272713
rect 530474 272701 530480 272753
rect 532816 272701 532822 272753
rect 532874 272741 532880 272753
rect 611920 272741 611926 272753
rect 532874 272713 611926 272741
rect 532874 272701 532880 272713
rect 611920 272701 611926 272713
rect 611978 272701 611984 272753
rect 302320 272627 302326 272679
rect 302378 272667 302384 272679
rect 360208 272667 360214 272679
rect 302378 272639 360214 272667
rect 302378 272627 302384 272639
rect 360208 272627 360214 272639
rect 360266 272627 360272 272679
rect 367120 272627 367126 272679
rect 367178 272667 367184 272679
rect 537424 272667 537430 272679
rect 367178 272639 537430 272667
rect 367178 272627 367184 272639
rect 537424 272627 537430 272639
rect 537482 272627 537488 272679
rect 367216 272593 367222 272605
rect 301418 272565 302078 272593
rect 302146 272565 367222 272593
rect 301418 272553 301424 272565
rect 103696 272479 103702 272531
rect 103754 272519 103760 272531
rect 203536 272519 203542 272531
rect 103754 272491 203542 272519
rect 103754 272479 103760 272491
rect 203536 272479 203542 272491
rect 203594 272479 203600 272531
rect 210064 272479 210070 272531
rect 210122 272519 210128 272531
rect 234544 272519 234550 272531
rect 210122 272491 234550 272519
rect 210122 272479 210128 272491
rect 234544 272479 234550 272491
rect 234602 272479 234608 272531
rect 234928 272479 234934 272531
rect 234986 272519 234992 272531
rect 244816 272519 244822 272531
rect 234986 272491 244822 272519
rect 234986 272479 234992 272491
rect 244816 272479 244822 272491
rect 244874 272479 244880 272531
rect 272272 272479 272278 272531
rect 272330 272519 272336 272531
rect 301936 272519 301942 272531
rect 272330 272491 301942 272519
rect 272330 272479 272336 272491
rect 301936 272479 301942 272491
rect 301994 272479 302000 272531
rect 302050 272519 302078 272565
rect 367216 272553 367222 272565
rect 367274 272553 367280 272605
rect 372688 272553 372694 272605
rect 372746 272593 372752 272605
rect 372746 272565 374462 272593
rect 372746 272553 372752 272565
rect 374320 272519 374326 272531
rect 302050 272491 374326 272519
rect 374320 272479 374326 272491
rect 374378 272479 374384 272531
rect 374434 272519 374462 272565
rect 374512 272553 374518 272605
rect 374570 272593 374576 272605
rect 536272 272593 536278 272605
rect 374570 272565 536278 272593
rect 374570 272553 374576 272565
rect 536272 272553 536278 272565
rect 536330 272553 536336 272605
rect 551632 272519 551638 272531
rect 374434 272491 551638 272519
rect 551632 272479 551638 272491
rect 551690 272479 551696 272531
rect 98992 272405 98998 272457
rect 99050 272445 99056 272457
rect 199120 272445 199126 272457
rect 99050 272417 199126 272445
rect 99050 272405 99056 272417
rect 199120 272405 199126 272417
rect 199178 272405 199184 272457
rect 232528 272405 232534 272457
rect 232586 272445 232592 272457
rect 243664 272445 243670 272457
rect 232586 272417 243670 272445
rect 232586 272405 232592 272417
rect 243664 272405 243670 272417
rect 243722 272405 243728 272457
rect 272752 272405 272758 272457
rect 272810 272445 272816 272457
rect 303472 272445 303478 272457
rect 272810 272417 303478 272445
rect 272810 272405 272816 272417
rect 303472 272405 303478 272417
rect 303530 272405 303536 272457
rect 307120 272405 307126 272457
rect 307178 272445 307184 272457
rect 307178 272417 326846 272445
rect 307178 272405 307184 272417
rect 96592 272331 96598 272383
rect 96650 272371 96656 272383
rect 201616 272371 201622 272383
rect 96650 272343 201622 272371
rect 96650 272331 96656 272343
rect 201616 272331 201622 272343
rect 201674 272331 201680 272383
rect 207664 272331 207670 272383
rect 207722 272371 207728 272383
rect 233872 272371 233878 272383
rect 207722 272343 233878 272371
rect 207722 272331 207728 272343
rect 233872 272331 233878 272343
rect 233930 272331 233936 272383
rect 236080 272331 236086 272383
rect 236138 272371 236144 272383
rect 245296 272371 245302 272383
rect 236138 272343 245302 272371
rect 236138 272331 236144 272343
rect 245296 272331 245302 272343
rect 245354 272331 245360 272383
rect 273424 272331 273430 272383
rect 273482 272371 273488 272383
rect 305776 272371 305782 272383
rect 273482 272343 305782 272371
rect 273482 272331 273488 272343
rect 305776 272331 305782 272343
rect 305834 272331 305840 272383
rect 309904 272331 309910 272383
rect 309962 272371 309968 272383
rect 326818 272371 326846 272417
rect 326896 272405 326902 272457
rect 326954 272445 326960 272457
rect 381424 272445 381430 272457
rect 326954 272417 381430 272445
rect 326954 272405 326960 272417
rect 381424 272405 381430 272417
rect 381482 272405 381488 272457
rect 381520 272405 381526 272457
rect 381578 272445 381584 272457
rect 572944 272445 572950 272457
rect 381578 272417 572950 272445
rect 381578 272405 381584 272417
rect 572944 272405 572950 272417
rect 573002 272405 573008 272457
rect 388528 272371 388534 272383
rect 309962 272343 326750 272371
rect 326818 272343 388534 272371
rect 309962 272331 309968 272343
rect 84784 272257 84790 272309
rect 84842 272297 84848 272309
rect 86320 272297 86326 272309
rect 84842 272269 86326 272297
rect 84842 272257 84848 272269
rect 86320 272257 86326 272269
rect 86378 272257 86384 272309
rect 104848 272257 104854 272309
rect 104906 272297 104912 272309
rect 106480 272297 106486 272309
rect 104906 272269 106486 272297
rect 104906 272257 104912 272269
rect 106480 272257 106486 272269
rect 106538 272257 106544 272309
rect 198256 272257 198262 272309
rect 198314 272297 198320 272309
rect 224368 272297 224374 272309
rect 198314 272269 224374 272297
rect 198314 272257 198320 272269
rect 224368 272257 224374 272269
rect 224426 272257 224432 272309
rect 227824 272257 227830 272309
rect 227882 272297 227888 272309
rect 242128 272297 242134 272309
rect 227882 272269 242134 272297
rect 227882 272257 227888 272269
rect 242128 272257 242134 272269
rect 242186 272257 242192 272309
rect 275152 272257 275158 272309
rect 275210 272297 275216 272309
rect 309328 272297 309334 272309
rect 275210 272269 309334 272297
rect 275210 272257 275216 272269
rect 309328 272257 309334 272269
rect 309386 272257 309392 272309
rect 312784 272257 312790 272309
rect 312842 272297 312848 272309
rect 326722 272297 326750 272343
rect 388528 272331 388534 272343
rect 388586 272331 388592 272383
rect 407440 272331 407446 272383
rect 407498 272371 407504 272383
rect 587152 272371 587158 272383
rect 407498 272343 587158 272371
rect 407498 272331 407504 272343
rect 587152 272331 587158 272343
rect 587210 272331 587216 272383
rect 395632 272297 395638 272309
rect 312842 272269 316814 272297
rect 326722 272269 395638 272297
rect 312842 272257 312848 272269
rect 165136 272183 165142 272235
rect 165194 272223 165200 272235
rect 166960 272223 166966 272235
rect 165194 272195 166966 272223
rect 165194 272183 165200 272195
rect 166960 272183 166966 272195
rect 167018 272183 167024 272235
rect 192400 272223 192406 272235
rect 175666 272195 192406 272223
rect 65872 272109 65878 272161
rect 65930 272149 65936 272161
rect 175666 272149 175694 272195
rect 192400 272183 192406 272195
rect 192458 272183 192464 272235
rect 194704 272183 194710 272235
rect 194762 272223 194768 272235
rect 224464 272223 224470 272235
rect 194762 272195 224470 272223
rect 194762 272183 194768 272195
rect 224464 272183 224470 272195
rect 224522 272183 224528 272235
rect 276304 272183 276310 272235
rect 276362 272223 276368 272235
rect 312880 272223 312886 272235
rect 276362 272195 312886 272223
rect 276362 272183 276368 272195
rect 312880 272183 312886 272195
rect 312938 272183 312944 272235
rect 316432 272223 316438 272235
rect 312994 272195 316438 272223
rect 65930 272121 175694 272149
rect 65930 272109 65936 272121
rect 191152 272109 191158 272161
rect 191210 272149 191216 272161
rect 227152 272149 227158 272161
rect 191210 272121 227158 272149
rect 191210 272109 191216 272121
rect 227152 272109 227158 272121
rect 227210 272109 227216 272161
rect 228976 272109 228982 272161
rect 229034 272149 229040 272161
rect 242416 272149 242422 272161
rect 229034 272121 242422 272149
rect 229034 272109 229040 272121
rect 242416 272109 242422 272121
rect 242474 272109 242480 272161
rect 277744 272109 277750 272161
rect 277802 272149 277808 272161
rect 312994 272149 313022 272195
rect 316432 272183 316438 272195
rect 316490 272183 316496 272235
rect 316786 272223 316814 272269
rect 395632 272257 395638 272269
rect 395690 272257 395696 272309
rect 395920 272257 395926 272309
rect 395978 272297 395984 272309
rect 608368 272297 608374 272309
rect 395978 272269 608374 272297
rect 395978 272257 395984 272269
rect 608368 272257 608374 272269
rect 608426 272257 608432 272309
rect 402736 272223 402742 272235
rect 316786 272195 402742 272223
rect 402736 272183 402742 272195
rect 402794 272183 402800 272235
rect 402928 272183 402934 272235
rect 402986 272223 402992 272235
rect 622576 272223 622582 272235
rect 402986 272195 622582 272223
rect 402986 272183 402992 272195
rect 622576 272183 622582 272195
rect 622634 272183 622640 272235
rect 277802 272121 313022 272149
rect 277802 272109 277808 272121
rect 315472 272109 315478 272161
rect 315530 272149 315536 272161
rect 409840 272149 409846 272161
rect 315530 272121 409846 272149
rect 315530 272109 315536 272121
rect 409840 272109 409846 272121
rect 409898 272109 409904 272161
rect 413680 272109 413686 272161
rect 413738 272149 413744 272161
rect 643888 272149 643894 272161
rect 413738 272121 643894 272149
rect 413738 272109 413744 272121
rect 643888 272109 643894 272121
rect 643946 272109 643952 272161
rect 167536 272035 167542 272087
rect 167594 272075 167600 272087
rect 210640 272075 210646 272087
rect 167594 272047 210646 272075
rect 167594 272035 167600 272047
rect 210640 272035 210646 272047
rect 210698 272035 210704 272087
rect 271024 272035 271030 272087
rect 271082 272075 271088 272087
rect 299920 272075 299926 272087
rect 271082 272047 299926 272075
rect 271082 272035 271088 272047
rect 299920 272035 299926 272047
rect 299978 272035 299984 272087
rect 328240 272075 328246 272087
rect 300034 272047 328246 272075
rect 174640 271961 174646 272013
rect 174698 272001 174704 272013
rect 210544 272001 210550 272013
rect 174698 271973 210550 272001
rect 174698 271961 174704 271973
rect 210544 271961 210550 271973
rect 210602 271961 210608 272013
rect 231376 271961 231382 272013
rect 231434 272001 231440 272013
rect 243088 272001 243094 272013
rect 231434 271973 243094 272001
rect 231434 271961 231440 271973
rect 243088 271961 243094 271973
rect 243146 271961 243152 272013
rect 299440 271961 299446 272013
rect 299498 272001 299504 272013
rect 300034 272001 300062 272047
rect 328240 272035 328246 272047
rect 328298 272035 328304 272087
rect 346960 272035 346966 272087
rect 347018 272075 347024 272087
rect 487792 272075 487798 272087
rect 347018 272047 487798 272075
rect 347018 272035 347024 272047
rect 487792 272035 487798 272047
rect 487850 272035 487856 272087
rect 299498 271973 300062 272001
rect 299498 271961 299504 271973
rect 302320 271961 302326 272013
rect 302378 272001 302384 272013
rect 324688 272001 324694 272013
rect 302378 271973 324694 272001
rect 302378 271961 302384 271973
rect 324688 271961 324694 271973
rect 324746 271961 324752 272013
rect 346480 271961 346486 272013
rect 346538 272001 346544 272013
rect 486640 272001 486646 272013
rect 346538 271973 486646 272001
rect 346538 271961 346544 271973
rect 486640 271961 486646 271973
rect 486698 271961 486704 272013
rect 159280 271887 159286 271939
rect 159338 271927 159344 271939
rect 198640 271927 198646 271939
rect 159338 271899 198646 271927
rect 159338 271887 159344 271899
rect 198640 271887 198646 271899
rect 198698 271887 198704 271939
rect 201808 271887 201814 271939
rect 201866 271927 201872 271939
rect 223696 271927 223702 271939
rect 201866 271899 223702 271927
rect 201866 271887 201872 271899
rect 223696 271887 223702 271899
rect 223754 271887 223760 271939
rect 233680 271887 233686 271939
rect 233738 271927 233744 271939
rect 244048 271927 244054 271939
rect 233738 271899 244054 271927
rect 233738 271887 233744 271899
rect 244048 271887 244054 271899
rect 244106 271887 244112 271939
rect 303952 271887 303958 271939
rect 304010 271927 304016 271939
rect 326896 271927 326902 271939
rect 304010 271899 326902 271927
rect 304010 271887 304016 271899
rect 326896 271887 326902 271899
rect 326954 271887 326960 271939
rect 344080 271887 344086 271939
rect 344138 271927 344144 271939
rect 480688 271927 480694 271939
rect 344138 271899 480694 271927
rect 344138 271887 344144 271899
rect 480688 271887 480694 271899
rect 480746 271887 480752 271939
rect 147376 271813 147382 271865
rect 147434 271853 147440 271865
rect 149680 271853 149686 271865
rect 147434 271825 149686 271853
rect 147434 271813 147440 271825
rect 149680 271813 149686 271825
rect 149738 271813 149744 271865
rect 166288 271813 166294 271865
rect 166346 271853 166352 271865
rect 201520 271853 201526 271865
rect 166346 271825 201526 271853
rect 166346 271813 166352 271825
rect 201520 271813 201526 271825
rect 201578 271813 201584 271865
rect 205360 271813 205366 271865
rect 205418 271853 205424 271865
rect 232624 271853 232630 271865
rect 205418 271825 232630 271853
rect 205418 271813 205424 271825
rect 232624 271813 232630 271825
rect 232682 271813 232688 271865
rect 284944 271813 284950 271865
rect 285002 271853 285008 271865
rect 306640 271853 306646 271865
rect 285002 271825 306646 271853
rect 285002 271813 285008 271825
rect 306640 271813 306646 271825
rect 306698 271813 306704 271865
rect 351376 271813 351382 271865
rect 351434 271853 351440 271865
rect 355408 271853 355414 271865
rect 351434 271825 355414 271853
rect 351434 271813 351440 271825
rect 355408 271813 355414 271825
rect 355466 271813 355472 271865
rect 473680 271853 473686 271865
rect 355522 271825 473686 271853
rect 101296 271739 101302 271791
rect 101354 271779 101360 271791
rect 103600 271779 103606 271791
rect 101354 271751 103606 271779
rect 101354 271739 101360 271751
rect 103600 271739 103606 271751
rect 103658 271739 103664 271791
rect 173392 271739 173398 271791
rect 173450 271779 173456 271791
rect 206032 271779 206038 271791
rect 173450 271751 206038 271779
rect 173450 271739 173456 271751
rect 206032 271739 206038 271751
rect 206090 271739 206096 271791
rect 341488 271739 341494 271791
rect 341546 271779 341552 271791
rect 355522 271779 355550 271825
rect 473680 271813 473686 271825
rect 473738 271813 473744 271865
rect 341546 271751 355550 271779
rect 341546 271739 341552 271751
rect 355600 271739 355606 271791
rect 355658 271779 355664 271791
rect 466576 271779 466582 271791
rect 355658 271751 466582 271779
rect 355658 271739 355664 271751
rect 466576 271739 466582 271751
rect 466634 271739 466640 271791
rect 115504 271665 115510 271717
rect 115562 271705 115568 271717
rect 118000 271705 118006 271717
rect 115562 271677 118006 271705
rect 115562 271665 115568 271677
rect 118000 271665 118006 271677
rect 118058 271665 118064 271717
rect 192304 271665 192310 271717
rect 192362 271705 192368 271717
rect 224560 271705 224566 271717
rect 192362 271677 224566 271705
rect 192362 271665 192368 271677
rect 224560 271665 224566 271677
rect 224618 271665 224624 271717
rect 335440 271665 335446 271717
rect 335498 271705 335504 271717
rect 459472 271705 459478 271717
rect 335498 271677 459478 271705
rect 335498 271665 335504 271677
rect 459472 271665 459478 271677
rect 459530 271665 459536 271717
rect 75280 271591 75286 271643
rect 75338 271631 75344 271643
rect 77680 271631 77686 271643
rect 75338 271603 77686 271631
rect 75338 271591 75344 271603
rect 77680 271591 77686 271603
rect 77738 271591 77744 271643
rect 129712 271591 129718 271643
rect 129770 271631 129776 271643
rect 132400 271631 132406 271643
rect 129770 271603 132406 271631
rect 129770 271591 129776 271603
rect 132400 271591 132406 271603
rect 132458 271591 132464 271643
rect 150928 271591 150934 271643
rect 150986 271631 150992 271643
rect 152368 271631 152374 271643
rect 150986 271603 152374 271631
rect 150986 271591 150992 271603
rect 152368 271591 152374 271603
rect 152426 271591 152432 271643
rect 181744 271591 181750 271643
rect 181802 271631 181808 271643
rect 210448 271631 210454 271643
rect 181802 271603 210454 271631
rect 181802 271591 181808 271603
rect 210448 271591 210454 271603
rect 210506 271591 210512 271643
rect 332560 271591 332566 271643
rect 332618 271631 332624 271643
rect 452368 271631 452374 271643
rect 332618 271603 452374 271631
rect 332618 271591 332624 271603
rect 452368 271591 452374 271603
rect 452426 271591 452432 271643
rect 89488 271517 89494 271569
rect 89546 271557 89552 271569
rect 92080 271557 92086 271569
rect 89546 271529 92086 271557
rect 89546 271517 89552 271529
rect 92080 271517 92086 271529
rect 92138 271517 92144 271569
rect 180496 271517 180502 271569
rect 180554 271557 180560 271569
rect 205840 271557 205846 271569
rect 180554 271529 205846 271557
rect 180554 271517 180560 271529
rect 205840 271517 205846 271529
rect 205898 271517 205904 271569
rect 329968 271517 329974 271569
rect 330026 271557 330032 271569
rect 445264 271557 445270 271569
rect 330026 271529 445270 271557
rect 330026 271517 330032 271529
rect 445264 271517 445270 271529
rect 445322 271517 445328 271569
rect 185200 271443 185206 271495
rect 185258 271483 185264 271495
rect 210352 271483 210358 271495
rect 185258 271455 210358 271483
rect 185258 271443 185264 271455
rect 210352 271443 210358 271455
rect 210410 271443 210416 271495
rect 326896 271443 326902 271495
rect 326954 271483 326960 271495
rect 438160 271483 438166 271495
rect 326954 271455 438166 271483
rect 326954 271443 326960 271455
rect 438160 271443 438166 271455
rect 438218 271443 438224 271495
rect 193552 271369 193558 271421
rect 193610 271409 193616 271421
rect 221680 271409 221686 271421
rect 193610 271381 221686 271409
rect 193610 271369 193616 271381
rect 221680 271369 221686 271381
rect 221738 271369 221744 271421
rect 324016 271369 324022 271421
rect 324074 271409 324080 271421
rect 431056 271409 431062 271421
rect 324074 271381 431062 271409
rect 324074 271369 324080 271381
rect 431056 271369 431062 271381
rect 431114 271369 431120 271421
rect 161584 271295 161590 271347
rect 161642 271335 161648 271347
rect 163888 271335 163894 271347
rect 161642 271307 163894 271335
rect 161642 271295 161648 271307
rect 163888 271295 163894 271307
rect 163946 271295 163952 271347
rect 188752 271295 188758 271347
rect 188810 271335 188816 271347
rect 210256 271335 210262 271347
rect 188810 271307 210262 271335
rect 188810 271295 188816 271307
rect 210256 271295 210262 271307
rect 210314 271295 210320 271347
rect 321424 271295 321430 271347
rect 321482 271335 321488 271347
rect 423952 271335 423958 271347
rect 321482 271307 423958 271335
rect 321482 271295 321488 271307
rect 423952 271295 423958 271307
rect 424010 271295 424016 271347
rect 184048 271221 184054 271273
rect 184106 271261 184112 271273
rect 205744 271261 205750 271273
rect 184106 271233 205750 271261
rect 184106 271221 184112 271233
rect 205744 271221 205750 271233
rect 205802 271221 205808 271273
rect 237232 271221 237238 271273
rect 237290 271261 237296 271273
rect 245584 271261 245590 271273
rect 237290 271233 245590 271261
rect 237290 271221 237296 271233
rect 245584 271221 245590 271233
rect 245642 271221 245648 271273
rect 318352 271221 318358 271273
rect 318410 271261 318416 271273
rect 416944 271261 416950 271273
rect 318410 271233 416950 271261
rect 318410 271221 318416 271233
rect 416944 271221 416950 271233
rect 417002 271221 417008 271273
rect 76528 271147 76534 271199
rect 76586 271187 76592 271199
rect 76586 271159 175694 271187
rect 76586 271147 76592 271159
rect 175666 271113 175694 271159
rect 175792 271147 175798 271199
rect 175850 271187 175856 271199
rect 178288 271187 178294 271199
rect 175850 271159 178294 271187
rect 175850 271147 175856 271159
rect 178288 271147 178294 271159
rect 178346 271147 178352 271199
rect 195664 271187 195670 271199
rect 187522 271159 195670 271187
rect 187522 271113 187550 271159
rect 195664 271147 195670 271159
rect 195722 271147 195728 271199
rect 199408 271147 199414 271199
rect 199466 271187 199472 271199
rect 221584 271187 221590 271199
rect 199466 271159 221590 271187
rect 199466 271147 199472 271159
rect 221584 271147 221590 271159
rect 221642 271147 221648 271199
rect 238480 271147 238486 271199
rect 238538 271187 238544 271199
rect 246064 271187 246070 271199
rect 238538 271159 246070 271187
rect 238538 271147 238544 271159
rect 246064 271147 246070 271159
rect 246122 271147 246128 271199
rect 338608 271147 338614 271199
rect 338666 271187 338672 271199
rect 355600 271187 355606 271199
rect 338666 271159 355606 271187
rect 338666 271147 338672 271159
rect 355600 271147 355606 271159
rect 355658 271147 355664 271199
rect 357904 271147 357910 271199
rect 357962 271187 357968 271199
rect 375184 271187 375190 271199
rect 357962 271159 375190 271187
rect 357962 271147 357968 271159
rect 375184 271147 375190 271159
rect 375242 271147 375248 271199
rect 387280 271147 387286 271199
rect 387338 271187 387344 271199
rect 407440 271187 407446 271199
rect 387338 271159 407446 271187
rect 387338 271147 387344 271159
rect 407440 271147 407446 271159
rect 407498 271147 407504 271199
rect 175666 271085 187550 271113
rect 187600 271073 187606 271125
rect 187658 271113 187664 271125
rect 205936 271113 205942 271125
rect 187658 271085 205942 271113
rect 187658 271073 187664 271085
rect 205936 271073 205942 271085
rect 205994 271073 206000 271125
rect 240784 271073 240790 271125
rect 240842 271113 240848 271125
rect 247216 271113 247222 271125
rect 240842 271085 247222 271113
rect 240842 271073 240848 271085
rect 247216 271073 247222 271085
rect 247274 271073 247280 271125
rect 85936 270999 85942 271051
rect 85994 271039 86000 271051
rect 198544 271039 198550 271051
rect 85994 271011 198550 271039
rect 85994 270999 86000 271011
rect 198544 270999 198550 271011
rect 198602 270999 198608 271051
rect 221872 270999 221878 271051
rect 221930 271039 221936 271051
rect 239344 271039 239350 271051
rect 221930 271011 239350 271039
rect 221930 270999 221936 271011
rect 239344 270999 239350 271011
rect 239402 270999 239408 271051
rect 239536 270999 239542 271051
rect 239594 271039 239600 271051
rect 241264 271039 241270 271051
rect 239594 271011 241270 271039
rect 239594 270999 239600 271011
rect 241264 270999 241270 271011
rect 241322 270999 241328 271051
rect 241936 270999 241942 271051
rect 241994 271039 242000 271051
rect 247696 271039 247702 271051
rect 241994 271011 247702 271039
rect 241994 270999 242000 271011
rect 247696 270999 247702 271011
rect 247754 270999 247760 271051
rect 334096 270999 334102 271051
rect 334154 271039 334160 271051
rect 337744 271039 337750 271051
rect 334154 271011 337750 271039
rect 334154 270999 334160 271011
rect 337744 270999 337750 271011
rect 337802 270999 337808 271051
rect 223024 270925 223030 270977
rect 223082 270965 223088 270977
rect 240016 270965 240022 270977
rect 223082 270937 240022 270965
rect 223082 270925 223088 270937
rect 240016 270925 240022 270937
rect 240074 270925 240080 270977
rect 243184 270925 243190 270977
rect 243242 270965 243248 270977
rect 247984 270965 247990 270977
rect 243242 270937 247990 270965
rect 243242 270925 243248 270937
rect 247984 270925 247990 270937
rect 248042 270925 248048 270977
rect 224272 270851 224278 270903
rect 224330 270891 224336 270903
rect 240496 270891 240502 270903
rect 224330 270863 240502 270891
rect 224330 270851 224336 270863
rect 240496 270851 240502 270863
rect 240554 270851 240560 270903
rect 244336 270851 244342 270903
rect 244394 270891 244400 270903
rect 248656 270891 248662 270903
rect 244394 270863 248662 270891
rect 244394 270851 244400 270863
rect 248656 270851 248662 270863
rect 248714 270851 248720 270903
rect 338704 270851 338710 270903
rect 338762 270891 338768 270903
rect 341296 270891 341302 270903
rect 338762 270863 341302 270891
rect 338762 270851 338768 270863
rect 341296 270851 341302 270863
rect 341354 270851 341360 270903
rect 645232 270851 645238 270903
rect 645290 270891 645296 270903
rect 652336 270891 652342 270903
rect 645290 270863 652342 270891
rect 645290 270851 645296 270863
rect 652336 270851 652342 270863
rect 652394 270851 652400 270903
rect 225424 270777 225430 270829
rect 225482 270817 225488 270829
rect 241072 270817 241078 270829
rect 225482 270789 241078 270817
rect 225482 270777 225488 270789
rect 241072 270777 241078 270789
rect 241130 270777 241136 270829
rect 245488 270777 245494 270829
rect 245546 270817 245552 270829
rect 249136 270817 249142 270829
rect 245546 270789 249142 270817
rect 245546 270777 245552 270789
rect 249136 270777 249142 270789
rect 249194 270777 249200 270829
rect 342736 270777 342742 270829
rect 342794 270817 342800 270829
rect 348304 270817 348310 270829
rect 342794 270789 348310 270817
rect 342794 270777 342800 270789
rect 348304 270777 348310 270789
rect 348362 270777 348368 270829
rect 94192 270703 94198 270755
rect 94250 270743 94256 270755
rect 94960 270743 94966 270755
rect 94250 270715 94966 270743
rect 94250 270703 94256 270715
rect 94960 270703 94966 270715
rect 95018 270703 95024 270755
rect 108400 270703 108406 270755
rect 108458 270743 108464 270755
rect 109360 270743 109366 270755
rect 108458 270715 109366 270743
rect 108458 270703 108464 270715
rect 109360 270703 109366 270715
rect 109418 270703 109424 270755
rect 119056 270703 119062 270755
rect 119114 270743 119120 270755
rect 120880 270743 120886 270755
rect 119114 270715 120886 270743
rect 119114 270703 119120 270715
rect 120880 270703 120886 270715
rect 120938 270703 120944 270755
rect 122608 270703 122614 270755
rect 122666 270743 122672 270755
rect 123760 270743 123766 270755
rect 122666 270715 123766 270743
rect 122666 270703 122672 270715
rect 123760 270703 123766 270715
rect 123818 270703 123824 270755
rect 136816 270703 136822 270755
rect 136874 270743 136880 270755
rect 138160 270743 138166 270755
rect 136874 270715 138166 270743
rect 136874 270703 136880 270715
rect 138160 270703 138166 270715
rect 138218 270703 138224 270755
rect 138256 270703 138262 270755
rect 138314 270743 138320 270755
rect 151600 270743 151606 270755
rect 138314 270715 151606 270743
rect 138314 270703 138320 270715
rect 151600 270703 151606 270715
rect 151658 270703 151664 270755
rect 154480 270703 154486 270755
rect 154538 270743 154544 270755
rect 155440 270743 155446 270755
rect 154538 270715 155446 270743
rect 154538 270703 154544 270715
rect 155440 270703 155446 270715
rect 155498 270703 155504 270755
rect 168688 270703 168694 270755
rect 168746 270743 168752 270755
rect 169840 270743 169846 270755
rect 168746 270715 169846 270743
rect 168746 270703 168752 270715
rect 169840 270703 169846 270715
rect 169898 270703 169904 270755
rect 179344 270703 179350 270755
rect 179402 270743 179408 270755
rect 181360 270743 181366 270755
rect 179402 270715 181366 270743
rect 179402 270703 179408 270715
rect 181360 270703 181366 270715
rect 181418 270703 181424 270755
rect 182896 270703 182902 270755
rect 182954 270743 182960 270755
rect 184240 270743 184246 270755
rect 182954 270715 184246 270743
rect 182954 270703 182960 270715
rect 184240 270703 184246 270715
rect 184298 270703 184304 270755
rect 185488 270703 185494 270755
rect 185546 270743 185552 270755
rect 186448 270743 186454 270755
rect 185546 270715 186454 270743
rect 185546 270703 185552 270715
rect 186448 270703 186454 270715
rect 186506 270703 186512 270755
rect 226576 270703 226582 270755
rect 226634 270743 226640 270755
rect 239536 270743 239542 270755
rect 226634 270715 239542 270743
rect 226634 270703 226640 270715
rect 239536 270703 239542 270715
rect 239594 270703 239600 270755
rect 239632 270703 239638 270755
rect 239690 270743 239696 270755
rect 246448 270743 246454 270755
rect 239690 270715 246454 270743
rect 239690 270703 239696 270715
rect 246448 270703 246454 270715
rect 246506 270703 246512 270755
rect 246736 270703 246742 270755
rect 246794 270743 246800 270755
rect 249616 270743 249622 270755
rect 246794 270715 249622 270743
rect 246794 270703 246800 270715
rect 249616 270703 249622 270715
rect 249674 270703 249680 270755
rect 408976 270703 408982 270755
rect 409034 270743 409040 270755
rect 413392 270743 413398 270755
rect 409034 270715 413398 270743
rect 409034 270703 409040 270715
rect 413392 270703 413398 270715
rect 413450 270703 413456 270755
rect 145072 270629 145078 270681
rect 145130 270669 145136 270681
rect 214480 270669 214486 270681
rect 145130 270641 214486 270669
rect 145130 270629 145136 270641
rect 214480 270629 214486 270641
rect 214538 270629 214544 270681
rect 279280 270629 279286 270681
rect 279338 270669 279344 270681
rect 293296 270669 293302 270681
rect 279338 270641 293302 270669
rect 279338 270629 279344 270641
rect 293296 270629 293302 270641
rect 293354 270629 293360 270681
rect 293392 270629 293398 270681
rect 293450 270669 293456 270681
rect 318832 270669 318838 270681
rect 293450 270641 318838 270669
rect 293450 270629 293456 270641
rect 318832 270629 318838 270641
rect 318890 270629 318896 270681
rect 348112 270629 348118 270681
rect 348170 270669 348176 270681
rect 490192 270669 490198 270681
rect 348170 270641 490198 270669
rect 348170 270629 348176 270641
rect 490192 270629 490198 270641
rect 490250 270629 490256 270681
rect 141520 270555 141526 270607
rect 141578 270595 141584 270607
rect 213808 270595 213814 270607
rect 141578 270567 213814 270595
rect 141578 270555 141584 270567
rect 213808 270555 213814 270567
rect 213866 270555 213872 270607
rect 280144 270555 280150 270607
rect 280202 270595 280208 270607
rect 322384 270595 322390 270607
rect 280202 270567 322390 270595
rect 280202 270555 280208 270567
rect 322384 270555 322390 270567
rect 322442 270555 322448 270607
rect 348400 270555 348406 270607
rect 348458 270595 348464 270607
rect 491344 270595 491350 270607
rect 348458 270567 491350 270595
rect 348458 270555 348464 270567
rect 491344 270555 491350 270567
rect 491402 270555 491408 270607
rect 137968 270481 137974 270533
rect 138026 270521 138032 270533
rect 212656 270521 212662 270533
rect 138026 270493 212662 270521
rect 138026 270481 138032 270493
rect 212656 270481 212662 270493
rect 212714 270481 212720 270533
rect 264688 270481 264694 270533
rect 264746 270521 264752 270533
rect 283312 270521 283318 270533
rect 264746 270493 283318 270521
rect 264746 270481 264752 270493
rect 283312 270481 283318 270493
rect 283370 270481 283376 270533
rect 323536 270521 323542 270533
rect 283426 270493 323542 270521
rect 134416 270407 134422 270459
rect 134474 270447 134480 270459
rect 211888 270447 211894 270459
rect 134474 270419 211894 270447
rect 134474 270407 134480 270419
rect 211888 270407 211894 270419
rect 211946 270407 211952 270459
rect 253936 270407 253942 270459
rect 253994 270447 254000 270459
rect 257296 270447 257302 270459
rect 253994 270419 257302 270447
rect 253994 270407 254000 270419
rect 257296 270407 257302 270419
rect 257354 270407 257360 270459
rect 262000 270407 262006 270459
rect 262058 270447 262064 270459
rect 277456 270447 277462 270459
rect 262058 270419 277462 270447
rect 262058 270407 262064 270419
rect 277456 270407 277462 270419
rect 277514 270407 277520 270459
rect 280624 270407 280630 270459
rect 280682 270447 280688 270459
rect 283426 270447 283454 270493
rect 323536 270481 323542 270493
rect 323594 270481 323600 270533
rect 350704 270481 350710 270533
rect 350762 270521 350768 270533
rect 497296 270521 497302 270533
rect 350762 270493 497302 270521
rect 350762 270481 350768 270493
rect 497296 270481 497302 270493
rect 497354 270481 497360 270533
rect 280682 270419 283454 270447
rect 280682 270407 280688 270419
rect 283696 270407 283702 270459
rect 283754 270447 283760 270459
rect 283754 270419 293246 270447
rect 283754 270407 283760 270419
rect 125008 270333 125014 270385
rect 125066 270373 125072 270385
rect 209488 270373 209494 270385
rect 125066 270345 209494 270373
rect 125066 270333 125072 270345
rect 209488 270333 209494 270345
rect 209546 270333 209552 270385
rect 262480 270333 262486 270385
rect 262538 270373 262544 270385
rect 278608 270373 278614 270385
rect 262538 270345 278614 270373
rect 262538 270333 262544 270345
rect 278608 270333 278614 270345
rect 278666 270333 278672 270385
rect 284176 270333 284182 270385
rect 284234 270373 284240 270385
rect 293218 270373 293246 270419
rect 293296 270407 293302 270459
rect 293354 270447 293360 270459
rect 319984 270447 319990 270459
rect 293354 270419 319990 270447
rect 293354 270407 293360 270419
rect 319984 270407 319990 270419
rect 320042 270407 320048 270459
rect 351280 270407 351286 270459
rect 351338 270447 351344 270459
rect 498448 270447 498454 270459
rect 351338 270419 498454 270447
rect 351338 270407 351344 270419
rect 498448 270407 498454 270419
rect 498506 270407 498512 270459
rect 330640 270373 330646 270385
rect 284234 270345 293150 270373
rect 293218 270345 330646 270373
rect 284234 270333 284240 270345
rect 121456 270259 121462 270311
rect 121514 270299 121520 270311
rect 208336 270299 208342 270311
rect 121514 270271 208342 270299
rect 121514 270259 121520 270271
rect 208336 270259 208342 270271
rect 208394 270259 208400 270311
rect 210544 270259 210550 270311
rect 210602 270299 210608 270311
rect 222832 270299 222838 270311
rect 210602 270271 222838 270299
rect 210602 270259 210608 270271
rect 222832 270259 222838 270271
rect 222890 270259 222896 270311
rect 255280 270259 255286 270311
rect 255338 270299 255344 270311
rect 260848 270299 260854 270311
rect 255338 270271 260854 270299
rect 255338 270259 255344 270271
rect 260848 270259 260854 270271
rect 260906 270259 260912 270311
rect 262960 270259 262966 270311
rect 263018 270299 263024 270311
rect 279760 270299 279766 270311
rect 263018 270271 279766 270299
rect 263018 270259 263024 270271
rect 279760 270259 279766 270271
rect 279818 270259 279824 270311
rect 286288 270259 286294 270311
rect 286346 270299 286352 270311
rect 293122 270299 293150 270345
rect 330640 270333 330646 270345
rect 330698 270333 330704 270385
rect 354064 270333 354070 270385
rect 354122 270373 354128 270385
rect 505552 270373 505558 270385
rect 354122 270345 505558 270373
rect 354122 270333 354128 270345
rect 505552 270333 505558 270345
rect 505610 270333 505616 270385
rect 331792 270299 331798 270311
rect 286346 270271 293054 270299
rect 293122 270271 331798 270299
rect 286346 270259 286352 270271
rect 114352 270185 114358 270237
rect 114410 270225 114416 270237
rect 206416 270225 206422 270237
rect 114410 270197 206422 270225
rect 114410 270185 114416 270197
rect 206416 270185 206422 270197
rect 206474 270185 206480 270237
rect 264880 270185 264886 270237
rect 264938 270225 264944 270237
rect 284560 270225 284566 270237
rect 264938 270197 284566 270225
rect 264938 270185 264944 270197
rect 284560 270185 284566 270197
rect 284618 270185 284624 270237
rect 287920 270185 287926 270237
rect 287978 270225 287984 270237
rect 292912 270225 292918 270237
rect 287978 270197 292918 270225
rect 287978 270185 287984 270197
rect 292912 270185 292918 270197
rect 292970 270185 292976 270237
rect 293026 270225 293054 270271
rect 331792 270259 331798 270271
rect 331850 270259 331856 270311
rect 353680 270259 353686 270311
rect 353738 270299 353744 270311
rect 504400 270299 504406 270311
rect 353738 270271 504406 270299
rect 353738 270259 353744 270271
rect 504400 270259 504406 270271
rect 504458 270259 504464 270311
rect 334096 270225 334102 270237
rect 293026 270197 334102 270225
rect 334096 270185 334102 270197
rect 334154 270185 334160 270237
rect 356752 270185 356758 270237
rect 356810 270225 356816 270237
rect 511504 270225 511510 270237
rect 356810 270197 511510 270225
rect 356810 270185 356816 270197
rect 511504 270185 511510 270197
rect 511562 270185 511568 270237
rect 117904 270111 117910 270163
rect 117962 270151 117968 270163
rect 207568 270151 207574 270163
rect 117962 270123 207574 270151
rect 117962 270111 117968 270123
rect 207568 270111 207574 270123
rect 207626 270111 207632 270163
rect 210448 270111 210454 270163
rect 210506 270151 210512 270163
rect 224752 270151 224758 270163
rect 210506 270123 224758 270151
rect 210506 270111 210512 270123
rect 224752 270111 224758 270123
rect 224810 270111 224816 270163
rect 265360 270111 265366 270163
rect 265418 270151 265424 270163
rect 265418 270123 276446 270151
rect 265418 270111 265424 270123
rect 109552 270037 109558 270089
rect 109610 270077 109616 270089
rect 205264 270077 205270 270089
rect 109610 270049 205270 270077
rect 109610 270037 109616 270049
rect 205264 270037 205270 270049
rect 205322 270037 205328 270089
rect 210352 270037 210358 270089
rect 210410 270077 210416 270089
rect 225520 270077 225526 270089
rect 210410 270049 225526 270077
rect 210410 270037 210416 270049
rect 225520 270037 225526 270049
rect 225578 270037 225584 270089
rect 266512 270037 266518 270089
rect 266570 270077 266576 270089
rect 276418 270077 276446 270123
rect 288496 270111 288502 270163
rect 288554 270151 288560 270163
rect 342448 270151 342454 270163
rect 288554 270123 342454 270151
rect 288554 270111 288560 270123
rect 342448 270111 342454 270123
rect 342506 270111 342512 270163
rect 356944 270111 356950 270163
rect 357002 270151 357008 270163
rect 512656 270151 512662 270163
rect 357002 270123 512662 270151
rect 357002 270111 357008 270123
rect 512656 270111 512662 270123
rect 512714 270111 512720 270163
rect 285712 270077 285718 270089
rect 266570 270049 276350 270077
rect 276418 270049 285718 270077
rect 266570 270037 266576 270049
rect 107248 269963 107254 270015
rect 107306 270003 107312 270015
rect 204688 270003 204694 270015
rect 107306 269975 204694 270003
rect 107306 269963 107312 269975
rect 204688 269963 204694 269975
rect 204746 269963 204752 270015
rect 210256 269963 210262 270015
rect 210314 270003 210320 270015
rect 226672 270003 226678 270015
rect 210314 269975 226678 270003
rect 210314 269963 210320 269975
rect 226672 269963 226678 269975
rect 226730 269963 226736 270015
rect 276322 270003 276350 270049
rect 285712 270037 285718 270049
rect 285770 270037 285776 270089
rect 292816 270077 292822 270089
rect 288130 270049 292822 270077
rect 288016 270003 288022 270015
rect 276322 269975 288022 270003
rect 288016 269963 288022 269975
rect 288074 269963 288080 270015
rect 102544 269889 102550 269941
rect 102602 269929 102608 269941
rect 203344 269929 203350 269941
rect 102602 269901 203350 269929
rect 102602 269889 102608 269901
rect 203344 269889 203350 269901
rect 203402 269889 203408 269941
rect 205840 269889 205846 269941
rect 205898 269929 205904 269941
rect 224080 269929 224086 269941
rect 205898 269901 224086 269929
rect 205898 269889 205904 269901
rect 224080 269889 224086 269901
rect 224138 269889 224144 269941
rect 261808 269889 261814 269941
rect 261866 269929 261872 269941
rect 276208 269929 276214 269941
rect 261866 269901 276214 269929
rect 261866 269889 261872 269901
rect 276208 269889 276214 269901
rect 276266 269889 276272 269941
rect 276400 269889 276406 269941
rect 276458 269929 276464 269941
rect 288130 269929 288158 270049
rect 292816 270037 292822 270049
rect 292874 270037 292880 270089
rect 292912 270037 292918 270089
rect 292970 270077 292976 270089
rect 338704 270077 338710 270089
rect 292970 270049 338710 270077
rect 292970 270037 292976 270049
rect 338704 270037 338710 270049
rect 338762 270037 338768 270089
rect 359824 270037 359830 270089
rect 359882 270077 359888 270089
rect 519760 270077 519766 270089
rect 359882 270049 519766 270077
rect 359882 270037 359888 270049
rect 519760 270037 519766 270049
rect 519818 270037 519824 270089
rect 290608 269963 290614 270015
rect 290666 270003 290672 270015
rect 342736 270003 342742 270015
rect 290666 269975 342742 270003
rect 290666 269963 290672 269975
rect 342736 269963 342742 269975
rect 342794 269963 342800 270015
rect 359344 269963 359350 270015
rect 359402 270003 359408 270015
rect 518512 270003 518518 270015
rect 359402 269975 518518 270003
rect 359402 269963 359408 269975
rect 518512 269963 518518 269975
rect 518570 269963 518576 270015
rect 276458 269901 288158 269929
rect 276458 269889 276464 269901
rect 291088 269889 291094 269941
rect 291146 269929 291152 269941
rect 349552 269929 349558 269941
rect 291146 269901 349558 269929
rect 291146 269889 291152 269901
rect 349552 269889 349558 269901
rect 349610 269889 349616 269941
rect 362704 269889 362710 269941
rect 362762 269929 362768 269941
rect 526864 269929 526870 269941
rect 362762 269901 526870 269929
rect 362762 269889 362768 269901
rect 526864 269889 526870 269901
rect 526922 269889 526928 269941
rect 100144 269815 100150 269867
rect 100202 269855 100208 269867
rect 202864 269855 202870 269867
rect 100202 269827 202870 269855
rect 100202 269815 100208 269827
rect 202864 269815 202870 269827
rect 202922 269815 202928 269867
rect 206032 269815 206038 269867
rect 206090 269855 206096 269867
rect 222352 269855 222358 269867
rect 206090 269827 222358 269855
rect 206090 269815 206096 269827
rect 222352 269815 222358 269827
rect 222410 269815 222416 269867
rect 261232 269815 261238 269867
rect 261290 269855 261296 269867
rect 275056 269855 275062 269867
rect 261290 269827 275062 269855
rect 261290 269815 261296 269827
rect 275056 269815 275062 269827
rect 275114 269815 275120 269867
rect 275248 269815 275254 269867
rect 275306 269855 275312 269867
rect 289264 269855 289270 269867
rect 275306 269827 289270 269855
rect 275306 269815 275312 269827
rect 289264 269815 289270 269827
rect 289322 269815 289328 269867
rect 293968 269815 293974 269867
rect 294026 269855 294032 269867
rect 356656 269855 356662 269867
rect 294026 269827 356662 269855
rect 294026 269815 294032 269827
rect 356656 269815 356662 269827
rect 356714 269815 356720 269867
rect 362224 269815 362230 269867
rect 362282 269855 362288 269867
rect 525616 269855 525622 269867
rect 362282 269827 525622 269855
rect 362282 269815 362288 269827
rect 525616 269815 525622 269827
rect 525674 269815 525680 269867
rect 95440 269741 95446 269793
rect 95498 269781 95504 269793
rect 201136 269781 201142 269793
rect 95498 269753 201142 269781
rect 95498 269741 95504 269753
rect 201136 269741 201142 269753
rect 201194 269741 201200 269793
rect 201520 269741 201526 269793
rect 201578 269781 201584 269793
rect 220528 269781 220534 269793
rect 201578 269753 220534 269781
rect 201578 269741 201584 269753
rect 220528 269741 220534 269753
rect 220586 269741 220592 269793
rect 256240 269741 256246 269793
rect 256298 269781 256304 269793
rect 263248 269781 263254 269793
rect 256298 269753 263254 269781
rect 256298 269741 256304 269753
rect 263248 269741 263254 269753
rect 263306 269741 263312 269793
rect 267760 269741 267766 269793
rect 267818 269781 267824 269793
rect 291568 269781 291574 269793
rect 267818 269753 291574 269781
rect 267818 269741 267824 269753
rect 291568 269741 291574 269753
rect 291626 269741 291632 269793
rect 293488 269741 293494 269793
rect 293546 269781 293552 269793
rect 351376 269781 351382 269793
rect 293546 269753 351382 269781
rect 293546 269741 293552 269753
rect 351376 269741 351382 269753
rect 351434 269741 351440 269793
rect 365296 269741 365302 269793
rect 365354 269781 365360 269793
rect 532720 269781 532726 269793
rect 365354 269753 532726 269781
rect 365354 269741 365360 269753
rect 532720 269741 532726 269753
rect 532778 269741 532784 269793
rect 93040 269667 93046 269719
rect 93098 269707 93104 269719
rect 200944 269707 200950 269719
rect 93098 269679 200950 269707
rect 93098 269667 93104 269679
rect 200944 269667 200950 269679
rect 201002 269667 201008 269719
rect 205936 269667 205942 269719
rect 205994 269707 206000 269719
rect 226000 269707 226006 269719
rect 205994 269679 226006 269707
rect 205994 269667 206000 269679
rect 226000 269667 226006 269679
rect 226058 269667 226064 269719
rect 259888 269667 259894 269719
rect 259946 269707 259952 269719
rect 271504 269707 271510 269719
rect 259946 269679 271510 269707
rect 259946 269667 259952 269679
rect 271504 269667 271510 269679
rect 271562 269667 271568 269719
rect 296368 269707 296374 269719
rect 271618 269679 296374 269707
rect 90640 269593 90646 269645
rect 90698 269633 90704 269645
rect 199696 269633 199702 269645
rect 90698 269605 199702 269633
rect 90698 269593 90704 269605
rect 199696 269593 199702 269605
rect 199754 269593 199760 269645
rect 205744 269593 205750 269645
rect 205802 269633 205808 269645
rect 225232 269633 225238 269645
rect 205802 269605 225238 269633
rect 205802 269593 205808 269605
rect 225232 269593 225238 269605
rect 225290 269593 225296 269645
rect 249040 269593 249046 269645
rect 249098 269633 249104 269645
rect 250288 269633 250294 269645
rect 249098 269605 250294 269633
rect 249098 269593 249104 269605
rect 250288 269593 250294 269605
rect 250346 269593 250352 269645
rect 255760 269593 255766 269645
rect 255818 269633 255824 269645
rect 262096 269633 262102 269645
rect 255818 269605 262102 269633
rect 255818 269593 255824 269605
rect 262096 269593 262102 269605
rect 262154 269593 262160 269645
rect 269680 269593 269686 269645
rect 269738 269633 269744 269645
rect 271618 269633 271646 269679
rect 296368 269667 296374 269679
rect 296426 269667 296432 269719
rect 297040 269667 297046 269719
rect 297098 269707 297104 269719
rect 363664 269707 363670 269719
rect 297098 269679 363670 269707
rect 297098 269667 297104 269679
rect 363664 269667 363670 269679
rect 363722 269667 363728 269719
rect 365488 269667 365494 269719
rect 365546 269707 365552 269719
rect 533872 269707 533878 269719
rect 365546 269679 533878 269707
rect 365546 269667 365552 269679
rect 533872 269667 533878 269679
rect 533930 269667 533936 269719
rect 269738 269605 271646 269633
rect 269738 269593 269744 269605
rect 271696 269593 271702 269645
rect 271754 269633 271760 269645
rect 293776 269633 293782 269645
rect 271754 269605 293782 269633
rect 271754 269593 271760 269605
rect 293776 269593 293782 269605
rect 293834 269593 293840 269645
rect 299632 269593 299638 269645
rect 299690 269633 299696 269645
rect 370768 269633 370774 269645
rect 299690 269605 370774 269633
rect 299690 269593 299696 269605
rect 370768 269593 370774 269605
rect 370826 269593 370832 269645
rect 385072 269633 385078 269645
rect 379714 269605 385078 269633
rect 83632 269519 83638 269571
rect 83690 269559 83696 269571
rect 198064 269559 198070 269571
rect 83690 269531 198070 269559
rect 83690 269519 83696 269531
rect 198064 269519 198070 269531
rect 198122 269519 198128 269571
rect 206512 269519 206518 269571
rect 206570 269559 206576 269571
rect 233392 269559 233398 269571
rect 206570 269531 233398 269559
rect 206570 269519 206576 269531
rect 233392 269519 233398 269531
rect 233450 269519 233456 269571
rect 269200 269519 269206 269571
rect 269258 269559 269264 269571
rect 295120 269559 295126 269571
rect 269258 269531 295126 269559
rect 269258 269519 269264 269531
rect 295120 269519 295126 269531
rect 295178 269519 295184 269571
rect 302608 269519 302614 269571
rect 302666 269559 302672 269571
rect 377872 269559 377878 269571
rect 302666 269531 377878 269559
rect 302666 269519 302672 269531
rect 377872 269519 377878 269531
rect 377930 269519 377936 269571
rect 87184 269445 87190 269497
rect 87242 269485 87248 269497
rect 199024 269485 199030 269497
rect 87242 269457 199030 269485
rect 87242 269445 87248 269457
rect 199024 269445 199030 269457
rect 199082 269445 199088 269497
rect 202960 269445 202966 269497
rect 203018 269485 203024 269497
rect 231952 269485 231958 269497
rect 203018 269457 231958 269485
rect 203018 269445 203024 269457
rect 231952 269445 231958 269457
rect 232010 269445 232016 269497
rect 271504 269445 271510 269497
rect 271562 269485 271568 269497
rect 301072 269485 301078 269497
rect 271562 269457 301078 269485
rect 271562 269445 271568 269457
rect 301072 269445 301078 269457
rect 301130 269445 301136 269497
rect 305680 269445 305686 269497
rect 305738 269485 305744 269497
rect 379600 269485 379606 269497
rect 305738 269457 379606 269485
rect 305738 269445 305744 269457
rect 379600 269445 379606 269457
rect 379658 269445 379664 269497
rect 82384 269371 82390 269423
rect 82442 269411 82448 269423
rect 197392 269411 197398 269423
rect 82442 269383 197398 269411
rect 82442 269371 82448 269383
rect 197392 269371 197398 269383
rect 197450 269371 197456 269423
rect 204112 269371 204118 269423
rect 204170 269411 204176 269423
rect 232144 269411 232150 269423
rect 204170 269383 232150 269411
rect 204170 269371 204176 269383
rect 232144 269371 232150 269383
rect 232202 269371 232208 269423
rect 258640 269371 258646 269423
rect 258698 269411 258704 269423
rect 269104 269411 269110 269423
rect 258698 269383 269110 269411
rect 258698 269371 258704 269383
rect 269104 269371 269110 269383
rect 269162 269371 269168 269423
rect 272944 269371 272950 269423
rect 273002 269411 273008 269423
rect 304624 269411 304630 269423
rect 273002 269383 304630 269411
rect 273002 269371 273008 269383
rect 304624 269371 304630 269383
rect 304682 269371 304688 269423
rect 308272 269371 308278 269423
rect 308330 269411 308336 269423
rect 379714 269411 379742 269605
rect 385072 269593 385078 269605
rect 385130 269593 385136 269645
rect 387376 269593 387382 269645
rect 387434 269633 387440 269645
rect 399184 269633 399190 269645
rect 387434 269605 399190 269633
rect 387434 269593 387440 269605
rect 399184 269593 399190 269605
rect 399242 269593 399248 269645
rect 379888 269519 379894 269571
rect 379946 269559 379952 269571
rect 569392 269559 569398 269571
rect 379946 269531 569398 269559
rect 379946 269519 379952 269531
rect 569392 269519 569398 269531
rect 569450 269519 569456 269571
rect 384112 269445 384118 269497
rect 384170 269485 384176 269497
rect 580048 269485 580054 269497
rect 384170 269457 580054 269485
rect 384170 269445 384176 269457
rect 580048 269445 580054 269457
rect 580106 269445 580112 269497
rect 308330 269383 379742 269411
rect 308330 269371 308336 269383
rect 379792 269371 379798 269423
rect 379850 269411 379856 269423
rect 384976 269411 384982 269423
rect 379850 269383 384982 269411
rect 379850 269371 379856 269383
rect 384976 269371 384982 269383
rect 385034 269371 385040 269423
rect 385072 269371 385078 269423
rect 385130 269411 385136 269423
rect 392080 269411 392086 269423
rect 385130 269383 392086 269411
rect 385130 269371 385136 269383
rect 392080 269371 392086 269383
rect 392138 269371 392144 269423
rect 394384 269371 394390 269423
rect 394442 269411 394448 269423
rect 604816 269411 604822 269423
rect 394442 269383 604822 269411
rect 394442 269371 394448 269383
rect 604816 269371 604822 269383
rect 604874 269371 604880 269423
rect 81232 269297 81238 269349
rect 81290 269337 81296 269349
rect 196816 269337 196822 269349
rect 81290 269309 196822 269337
rect 81290 269297 81296 269309
rect 196816 269297 196822 269309
rect 196874 269297 196880 269349
rect 200656 269297 200662 269349
rect 200714 269337 200720 269349
rect 230992 269337 230998 269349
rect 200714 269309 230998 269337
rect 200714 269297 200720 269309
rect 230992 269297 230998 269309
rect 231050 269297 231056 269349
rect 268624 269297 268630 269349
rect 268682 269337 268688 269349
rect 271696 269337 271702 269349
rect 268682 269309 271702 269337
rect 268682 269297 268688 269309
rect 271696 269297 271702 269309
rect 271754 269297 271760 269349
rect 278896 269297 278902 269349
rect 278954 269337 278960 269349
rect 293392 269337 293398 269349
rect 278954 269309 293398 269337
rect 278954 269297 278960 269309
rect 293392 269297 293398 269309
rect 293450 269297 293456 269349
rect 311152 269297 311158 269349
rect 311210 269337 311216 269349
rect 387376 269337 387382 269349
rect 311210 269309 387382 269337
rect 311210 269297 311216 269309
rect 387376 269297 387382 269309
rect 387434 269297 387440 269349
rect 399952 269297 399958 269349
rect 400010 269337 400016 269349
rect 619024 269337 619030 269349
rect 400010 269309 619030 269337
rect 400010 269297 400016 269309
rect 619024 269297 619030 269309
rect 619082 269297 619088 269349
rect 74128 269223 74134 269275
rect 74186 269263 74192 269275
rect 194992 269263 194998 269275
rect 74186 269235 194998 269263
rect 74186 269223 74192 269235
rect 194992 269223 194998 269235
rect 195050 269223 195056 269275
rect 197104 269223 197110 269275
rect 197162 269263 197168 269275
rect 229552 269263 229558 269275
rect 197162 269235 229558 269263
rect 197162 269223 197168 269235
rect 229552 269223 229558 269235
rect 229610 269223 229616 269275
rect 260560 269223 260566 269275
rect 260618 269263 260624 269275
rect 273904 269263 273910 269275
rect 260618 269235 273910 269263
rect 260618 269223 260624 269235
rect 273904 269223 273910 269235
rect 273962 269223 273968 269275
rect 314224 269223 314230 269275
rect 314282 269263 314288 269275
rect 406288 269263 406294 269275
rect 314282 269235 406294 269263
rect 314282 269223 314288 269235
rect 406288 269223 406294 269235
rect 406346 269223 406352 269275
rect 146224 269149 146230 269201
rect 146282 269189 146288 269201
rect 214960 269189 214966 269201
rect 146282 269161 214966 269189
rect 146282 269149 146288 269161
rect 214960 269149 214966 269161
rect 215018 269149 215024 269201
rect 267088 269149 267094 269201
rect 267146 269189 267152 269201
rect 275248 269189 275254 269201
rect 267146 269161 275254 269189
rect 267146 269149 267152 269161
rect 275248 269149 275254 269161
rect 275306 269149 275312 269201
rect 277552 269149 277558 269201
rect 277610 269189 277616 269201
rect 315280 269189 315286 269201
rect 277610 269161 315286 269189
rect 277610 269149 277616 269161
rect 315280 269149 315286 269161
rect 315338 269149 315344 269201
rect 345424 269149 345430 269201
rect 345482 269189 345488 269201
rect 484240 269189 484246 269201
rect 345482 269161 484246 269189
rect 345482 269149 345488 269161
rect 484240 269149 484246 269161
rect 484298 269149 484304 269201
rect 148624 269075 148630 269127
rect 148682 269115 148688 269127
rect 215728 269115 215734 269127
rect 148682 269087 215734 269115
rect 148682 269075 148688 269087
rect 215728 269075 215734 269087
rect 215786 269075 215792 269127
rect 253360 269075 253366 269127
rect 253418 269115 253424 269127
rect 256144 269115 256150 269127
rect 253418 269087 256150 269115
rect 253418 269075 253424 269087
rect 256144 269075 256150 269087
rect 256202 269075 256208 269127
rect 257008 269075 257014 269127
rect 257066 269115 257072 269127
rect 264400 269115 264406 269127
rect 257066 269087 264406 269115
rect 257066 269075 257072 269087
rect 264400 269075 264406 269087
rect 264458 269075 264464 269127
rect 268432 269075 268438 269127
rect 268490 269115 268496 269127
rect 276400 269115 276406 269127
rect 268490 269087 276406 269115
rect 268490 269075 268496 269087
rect 276400 269075 276406 269087
rect 276458 269075 276464 269127
rect 281296 269075 281302 269127
rect 281354 269115 281360 269127
rect 302320 269115 302326 269127
rect 281354 269087 302326 269115
rect 281354 269075 281360 269087
rect 302320 269075 302326 269087
rect 302378 269075 302384 269127
rect 306352 269075 306358 269127
rect 306410 269115 306416 269127
rect 341200 269115 341206 269127
rect 306410 269087 341206 269115
rect 306410 269075 306416 269087
rect 341200 269075 341206 269087
rect 341258 269075 341264 269127
rect 345232 269075 345238 269127
rect 345290 269115 345296 269127
rect 483088 269115 483094 269127
rect 345290 269087 483094 269115
rect 345290 269075 345296 269087
rect 483088 269075 483094 269087
rect 483146 269075 483152 269127
rect 149776 269001 149782 269053
rect 149834 269041 149840 269053
rect 216208 269041 216214 269053
rect 149834 269013 216214 269041
rect 149834 269001 149840 269013
rect 216208 269001 216214 269013
rect 216266 269001 216272 269053
rect 266032 269001 266038 269053
rect 266090 269041 266096 269053
rect 286864 269041 286870 269053
rect 266090 269013 286870 269041
rect 266090 269001 266096 269013
rect 286864 269001 286870 269013
rect 286922 269001 286928 269053
rect 303760 269001 303766 269053
rect 303818 269041 303824 269053
rect 334288 269041 334294 269053
rect 303818 269013 334294 269041
rect 303818 269001 303824 269013
rect 334288 269001 334294 269013
rect 334346 269001 334352 269053
rect 342640 269001 342646 269053
rect 342698 269041 342704 269053
rect 477136 269041 477142 269053
rect 342698 269013 477142 269041
rect 342698 269001 342704 269013
rect 477136 269001 477142 269013
rect 477194 269001 477200 269053
rect 152176 268927 152182 268979
rect 152234 268967 152240 268979
rect 216688 268967 216694 268979
rect 152234 268939 216694 268967
rect 152234 268927 152240 268939
rect 216688 268927 216694 268939
rect 216746 268927 216752 268979
rect 260080 268927 260086 268979
rect 260138 268967 260144 268979
rect 272656 268967 272662 268979
rect 260138 268939 272662 268967
rect 260138 268927 260144 268939
rect 272656 268927 272662 268939
rect 272714 268927 272720 268979
rect 282064 268927 282070 268979
rect 282122 268967 282128 268979
rect 299344 268967 299350 268979
rect 282122 268939 299350 268967
rect 282122 268927 282128 268939
rect 299344 268927 299350 268939
rect 299402 268927 299408 268979
rect 302032 268927 302038 268979
rect 302090 268967 302096 268979
rect 331216 268967 331222 268979
rect 302090 268939 331222 268967
rect 302090 268927 302096 268939
rect 331216 268927 331222 268939
rect 331274 268927 331280 268979
rect 339760 268927 339766 268979
rect 339818 268967 339824 268979
rect 470128 268967 470134 268979
rect 339818 268939 470134 268967
rect 339818 268927 339824 268939
rect 470128 268927 470134 268939
rect 470186 268927 470192 268979
rect 155728 268853 155734 268905
rect 155786 268893 155792 268905
rect 217360 268893 217366 268905
rect 155786 268865 217366 268893
rect 155786 268853 155792 268865
rect 217360 268853 217366 268865
rect 217418 268853 217424 268905
rect 300688 268853 300694 268905
rect 300746 268893 300752 268905
rect 326800 268893 326806 268905
rect 300746 268865 326806 268893
rect 300746 268853 300752 268865
rect 326800 268853 326806 268865
rect 326858 268853 326864 268905
rect 336880 268853 336886 268905
rect 336938 268893 336944 268905
rect 463024 268893 463030 268905
rect 336938 268865 463030 268893
rect 336938 268853 336944 268865
rect 463024 268853 463030 268865
rect 463082 268853 463088 268905
rect 156880 268779 156886 268831
rect 156938 268819 156944 268831
rect 218128 268819 218134 268831
rect 156938 268791 218134 268819
rect 156938 268779 156944 268791
rect 218128 268779 218134 268791
rect 218186 268779 218192 268831
rect 258160 268779 258166 268831
rect 258218 268819 258224 268831
rect 267952 268819 267958 268831
rect 258218 268791 267958 268819
rect 258218 268779 258224 268791
rect 267952 268779 267958 268791
rect 268010 268779 268016 268831
rect 289168 268779 289174 268831
rect 289226 268819 289232 268831
rect 310576 268819 310582 268831
rect 289226 268791 310582 268819
rect 289226 268779 289232 268791
rect 310576 268779 310582 268791
rect 310634 268779 310640 268831
rect 334288 268779 334294 268831
rect 334346 268819 334352 268831
rect 455920 268819 455926 268831
rect 334346 268791 455926 268819
rect 334346 268779 334352 268791
rect 455920 268779 455926 268791
rect 455978 268779 455984 268831
rect 162832 268705 162838 268757
rect 162890 268745 162896 268757
rect 219280 268745 219286 268757
rect 162890 268717 219286 268745
rect 162890 268705 162896 268717
rect 219280 268705 219286 268717
rect 219338 268705 219344 268757
rect 257680 268705 257686 268757
rect 257738 268745 257744 268757
rect 266800 268745 266806 268757
rect 257738 268717 266806 268745
rect 257738 268705 257744 268717
rect 266800 268705 266806 268717
rect 266858 268705 266864 268757
rect 295216 268705 295222 268757
rect 295274 268745 295280 268757
rect 306832 268745 306838 268757
rect 295274 268717 306838 268745
rect 295274 268705 295280 268717
rect 306832 268705 306838 268717
rect 306890 268705 306896 268757
rect 331216 268705 331222 268757
rect 331274 268745 331280 268757
rect 448816 268745 448822 268757
rect 331274 268717 448822 268745
rect 331274 268705 331280 268717
rect 448816 268705 448822 268717
rect 448874 268705 448880 268757
rect 163984 268631 163990 268683
rect 164042 268671 164048 268683
rect 219952 268671 219958 268683
rect 164042 268643 219958 268671
rect 164042 268631 164048 268643
rect 219952 268631 219958 268643
rect 220010 268631 220016 268683
rect 254608 268631 254614 268683
rect 254666 268671 254672 268683
rect 258544 268671 258550 268683
rect 254666 268643 258550 268671
rect 254666 268631 254672 268643
rect 258544 268631 258550 268643
rect 258602 268631 258608 268683
rect 259408 268631 259414 268683
rect 259466 268671 259472 268683
rect 270352 268671 270358 268683
rect 259466 268643 270358 268671
rect 259466 268631 259472 268643
rect 270352 268631 270358 268643
rect 270410 268631 270416 268683
rect 275824 268631 275830 268683
rect 275882 268671 275888 268683
rect 311728 268671 311734 268683
rect 275882 268643 311734 268671
rect 275882 268631 275888 268643
rect 311728 268631 311734 268643
rect 311786 268631 311792 268683
rect 328336 268631 328342 268683
rect 328394 268671 328400 268683
rect 441712 268671 441718 268683
rect 328394 268643 441718 268671
rect 328394 268631 328400 268643
rect 441712 268631 441718 268643
rect 441770 268631 441776 268683
rect 42160 268557 42166 268609
rect 42218 268597 42224 268609
rect 48304 268597 48310 268609
rect 42218 268569 48310 268597
rect 42218 268557 42224 268569
rect 48304 268557 48310 268569
rect 48362 268557 48368 268609
rect 169744 268557 169750 268609
rect 169802 268597 169808 268609
rect 221200 268597 221206 268609
rect 169802 268569 221206 268597
rect 169802 268557 169808 268569
rect 221200 268557 221206 268569
rect 221258 268557 221264 268609
rect 274672 268557 274678 268609
rect 274730 268597 274736 268609
rect 308176 268597 308182 268609
rect 274730 268569 308182 268597
rect 274730 268557 274736 268569
rect 308176 268557 308182 268569
rect 308234 268557 308240 268609
rect 325744 268557 325750 268609
rect 325802 268597 325808 268609
rect 434608 268597 434614 268609
rect 325802 268569 434614 268597
rect 325802 268557 325808 268569
rect 434608 268557 434614 268569
rect 434666 268557 434672 268609
rect 171088 268483 171094 268535
rect 171146 268523 171152 268535
rect 221776 268523 221782 268535
rect 171146 268495 221782 268523
rect 171146 268483 171152 268495
rect 221776 268483 221782 268495
rect 221834 268483 221840 268535
rect 253168 268483 253174 268535
rect 253226 268523 253232 268535
rect 254992 268523 254998 268535
rect 253226 268495 254998 268523
rect 253226 268483 253232 268495
rect 254992 268483 254998 268495
rect 255050 268483 255056 268535
rect 267280 268483 267286 268535
rect 267338 268523 267344 268535
rect 290416 268523 290422 268535
rect 267338 268495 290422 268523
rect 267338 268483 267344 268495
rect 290416 268483 290422 268495
rect 290474 268483 290480 268535
rect 322576 268483 322582 268535
rect 322634 268523 322640 268535
rect 427504 268523 427510 268535
rect 322634 268495 427510 268523
rect 322634 268483 322640 268495
rect 427504 268483 427510 268495
rect 427562 268483 427568 268535
rect 176944 268409 176950 268461
rect 177002 268449 177008 268461
rect 223408 268449 223414 268461
rect 177002 268421 223414 268449
rect 177002 268409 177008 268421
rect 223408 268409 223414 268421
rect 223466 268409 223472 268461
rect 319696 268409 319702 268461
rect 319754 268449 319760 268461
rect 420496 268449 420502 268461
rect 319754 268421 420502 268449
rect 319754 268409 319760 268421
rect 420496 268409 420502 268421
rect 420554 268409 420560 268461
rect 178192 268335 178198 268387
rect 178250 268375 178256 268387
rect 223600 268375 223606 268387
rect 178250 268347 223606 268375
rect 178250 268335 178256 268347
rect 223600 268335 223606 268347
rect 223658 268335 223664 268387
rect 247888 268335 247894 268387
rect 247946 268375 247952 268387
rect 249808 268375 249814 268387
rect 247946 268347 249814 268375
rect 247946 268335 247952 268347
rect 249808 268335 249814 268347
rect 249866 268335 249872 268387
rect 255088 268335 255094 268387
rect 255146 268375 255152 268387
rect 259696 268375 259702 268387
rect 255146 268347 259702 268375
rect 255146 268335 255152 268347
rect 259696 268335 259702 268347
rect 259754 268335 259760 268387
rect 264112 268335 264118 268387
rect 264170 268375 264176 268387
rect 282160 268375 282166 268387
rect 264170 268347 282166 268375
rect 264170 268335 264176 268347
rect 282160 268335 282166 268347
rect 282218 268335 282224 268387
rect 317104 268335 317110 268387
rect 317162 268375 317168 268387
rect 408976 268375 408982 268387
rect 317162 268347 408982 268375
rect 317162 268335 317168 268347
rect 408976 268335 408982 268347
rect 409034 268335 409040 268387
rect 198640 268261 198646 268313
rect 198698 268301 198704 268313
rect 218608 268301 218614 268313
rect 198698 268273 218614 268301
rect 198698 268261 198704 268273
rect 218608 268261 218614 268273
rect 218666 268261 218672 268313
rect 221488 268261 221494 268313
rect 221546 268301 221552 268313
rect 229072 268301 229078 268313
rect 221546 268273 229078 268301
rect 221546 268261 221552 268273
rect 229072 268261 229078 268273
rect 229130 268261 229136 268313
rect 309232 268261 309238 268313
rect 309290 268301 309296 268313
rect 347056 268301 347062 268313
rect 309290 268273 347062 268301
rect 309290 268261 309296 268273
rect 347056 268261 347062 268273
rect 347114 268261 347120 268313
rect 192976 268187 192982 268239
rect 193034 268227 193040 268239
rect 210736 268227 210742 268239
rect 193034 268199 210742 268227
rect 193034 268187 193040 268199
rect 210736 268187 210742 268199
rect 210794 268187 210800 268239
rect 223696 268187 223702 268239
rect 223754 268227 223760 268239
rect 231472 268227 231478 268239
rect 223754 268199 231478 268227
rect 223754 268187 223760 268199
rect 231472 268187 231478 268199
rect 231530 268187 231536 268239
rect 257488 268187 257494 268239
rect 257546 268227 257552 268239
rect 265648 268227 265654 268239
rect 257546 268199 265654 268227
rect 257546 268187 257552 268199
rect 265648 268187 265654 268199
rect 265706 268187 265712 268239
rect 281008 268227 281014 268239
rect 276466 268199 281014 268227
rect 209776 268113 209782 268165
rect 209834 268153 209840 268165
rect 212368 268153 212374 268165
rect 209834 268125 212374 268153
rect 209834 268113 209840 268125
rect 212368 268113 212374 268125
rect 212426 268113 212432 268165
rect 212464 268113 212470 268165
rect 212522 268153 212528 268165
rect 218896 268153 218902 268165
rect 212522 268125 218902 268153
rect 212522 268113 212528 268125
rect 218896 268113 218902 268125
rect 218954 268113 218960 268165
rect 224368 268113 224374 268165
rect 224426 268153 224432 268165
rect 230032 268153 230038 268165
rect 224426 268125 230038 268153
rect 224426 268113 224432 268125
rect 230032 268113 230038 268125
rect 230090 268113 230096 268165
rect 263632 268113 263638 268165
rect 263690 268153 263696 268165
rect 276466 268153 276494 268199
rect 281008 268187 281014 268199
rect 281066 268187 281072 268239
rect 312304 268187 312310 268239
rect 312362 268227 312368 268239
rect 348496 268227 348502 268239
rect 312362 268199 348502 268227
rect 312362 268187 312368 268199
rect 348496 268187 348502 268199
rect 348554 268187 348560 268239
rect 408496 268187 408502 268239
rect 408554 268227 408560 268239
rect 640336 268227 640342 268239
rect 408554 268199 640342 268227
rect 408554 268187 408560 268199
rect 640336 268187 640342 268199
rect 640394 268187 640400 268239
rect 263690 268125 276494 268153
rect 263690 268113 263696 268125
rect 330736 268113 330742 268165
rect 330794 268153 330800 268165
rect 343792 268153 343798 268165
rect 330794 268125 343798 268153
rect 330794 268113 330800 268125
rect 343792 268113 343798 268125
rect 343850 268113 343856 268165
rect 371248 268113 371254 268165
rect 371306 268153 371312 268165
rect 548080 268153 548086 268165
rect 371306 268125 548086 268153
rect 371306 268113 371312 268125
rect 548080 268113 548086 268125
rect 548138 268113 548144 268165
rect 207376 268039 207382 268091
rect 207434 268079 207440 268091
rect 216880 268079 216886 268091
rect 207434 268051 216886 268079
rect 207434 268039 207440 268051
rect 216880 268039 216886 268051
rect 216938 268039 216944 268091
rect 224464 268039 224470 268091
rect 224522 268079 224528 268091
rect 228400 268079 228406 268091
rect 224522 268051 228406 268079
rect 224522 268039 224528 268051
rect 228400 268039 228406 268051
rect 228458 268039 228464 268091
rect 252688 268039 252694 268091
rect 252746 268079 252752 268091
rect 253744 268079 253750 268091
rect 252746 268051 253750 268079
rect 252746 268039 252752 268051
rect 253744 268039 253750 268051
rect 253802 268039 253808 268091
rect 333616 268039 333622 268091
rect 333674 268079 333680 268091
rect 351376 268079 351382 268091
rect 333674 268051 351382 268079
rect 333674 268039 333680 268051
rect 351376 268039 351382 268051
rect 351434 268039 351440 268091
rect 209872 267965 209878 268017
rect 209930 268005 209936 268017
rect 211408 268005 211414 268017
rect 209930 267977 211414 268005
rect 209930 267965 209936 267977
rect 211408 267965 211414 267977
rect 211466 267965 211472 268017
rect 221584 267965 221590 268017
rect 221642 268005 221648 268017
rect 230512 268005 230518 268017
rect 221642 267977 230518 268005
rect 221642 267965 221648 267977
rect 230512 267965 230518 267977
rect 230570 267965 230576 268017
rect 336688 267965 336694 268017
rect 336746 268005 336752 268017
rect 357616 268005 357622 268017
rect 336746 267977 357622 268005
rect 336746 267965 336752 267977
rect 357616 267965 357622 267977
rect 357674 267965 357680 268017
rect 210640 267891 210646 267943
rect 210698 267931 210704 267943
rect 221008 267931 221014 267943
rect 210698 267903 221014 267931
rect 210698 267891 210704 267903
rect 221008 267891 221014 267903
rect 221066 267891 221072 267943
rect 221680 267891 221686 267943
rect 221738 267931 221744 267943
rect 227824 267931 227830 267943
rect 221738 267903 227830 267931
rect 221738 267891 221744 267903
rect 227824 267891 227830 267903
rect 227882 267891 227888 267943
rect 339280 267891 339286 267943
rect 339338 267931 339344 267943
rect 362800 267931 362806 267943
rect 339338 267903 362806 267931
rect 339338 267891 339344 267903
rect 362800 267891 362806 267903
rect 362858 267891 362864 267943
rect 199120 267817 199126 267869
rect 199178 267857 199184 267869
rect 202288 267857 202294 267869
rect 199178 267829 202294 267857
rect 199178 267817 199184 267829
rect 202288 267817 202294 267829
rect 202346 267817 202352 267869
rect 207472 267817 207478 267869
rect 207530 267857 207536 267869
rect 212464 267857 212470 267869
rect 207530 267829 212470 267857
rect 207530 267817 207536 267829
rect 212464 267817 212470 267829
rect 212522 267817 212528 267869
rect 224560 267817 224566 267869
rect 224618 267857 224624 267869
rect 227632 267857 227638 267869
rect 224618 267829 227638 267857
rect 224618 267817 224624 267829
rect 227632 267817 227638 267829
rect 227690 267817 227696 267869
rect 282544 267817 282550 267869
rect 282602 267857 282608 267869
rect 299440 267857 299446 267869
rect 282602 267829 299446 267857
rect 282602 267817 282608 267829
rect 299440 267817 299446 267829
rect 299498 267817 299504 267869
rect 342160 267817 342166 267869
rect 342218 267857 342224 267869
rect 365680 267857 365686 267869
rect 342218 267829 365686 267857
rect 342218 267817 342224 267829
rect 365680 267817 365686 267829
rect 365738 267817 365744 267869
rect 401296 267817 401302 267869
rect 401354 267857 401360 267869
rect 402928 267857 402934 267869
rect 401354 267829 402934 267857
rect 401354 267817 401360 267829
rect 402928 267817 402934 267829
rect 402986 267817 402992 267869
rect 409936 267817 409942 267869
rect 409994 267857 410000 267869
rect 413680 267857 413686 267869
rect 409994 267829 413686 267857
rect 409994 267817 410000 267829
rect 413680 267817 413686 267829
rect 413738 267817 413744 267869
rect 388720 267743 388726 267795
rect 388778 267783 388784 267795
rect 645232 267783 645238 267795
rect 388778 267755 645238 267783
rect 388778 267743 388784 267755
rect 645232 267743 645238 267755
rect 645290 267743 645296 267795
rect 351952 267669 351958 267721
rect 352010 267709 352016 267721
rect 499600 267709 499606 267721
rect 352010 267681 499606 267709
rect 352010 267669 352016 267681
rect 499600 267669 499606 267681
rect 499658 267669 499664 267721
rect 354832 267595 354838 267647
rect 354890 267635 354896 267647
rect 506704 267635 506710 267647
rect 354890 267607 506710 267635
rect 354890 267595 354896 267607
rect 506704 267595 506710 267607
rect 506762 267595 506768 267647
rect 357424 267521 357430 267573
rect 357482 267561 357488 267573
rect 513808 267561 513814 267573
rect 357482 267533 513814 267561
rect 357482 267521 357488 267533
rect 513808 267521 513814 267533
rect 513866 267521 513872 267573
rect 360304 267447 360310 267499
rect 360362 267487 360368 267499
rect 520912 267487 520918 267499
rect 360362 267459 520918 267487
rect 360362 267447 360368 267459
rect 520912 267447 520918 267459
rect 520970 267447 520976 267499
rect 363376 267373 363382 267425
rect 363434 267413 363440 267425
rect 528016 267413 528022 267425
rect 363434 267385 528022 267413
rect 363434 267373 363440 267385
rect 528016 267373 528022 267385
rect 528074 267373 528080 267425
rect 365968 267299 365974 267351
rect 366026 267339 366032 267351
rect 535120 267339 535126 267351
rect 366026 267311 535126 267339
rect 366026 267299 366032 267311
rect 535120 267299 535126 267311
rect 535178 267299 535184 267351
rect 368944 267225 368950 267277
rect 369002 267265 369008 267277
rect 542224 267265 542230 267277
rect 369002 267237 542230 267265
rect 369002 267225 369008 267237
rect 542224 267225 542230 267237
rect 542282 267225 542288 267277
rect 372496 267151 372502 267203
rect 372554 267191 372560 267203
rect 550480 267191 550486 267203
rect 372554 267163 550486 267191
rect 372554 267151 372560 267163
rect 550480 267151 550486 267163
rect 550538 267151 550544 267203
rect 384880 267077 384886 267129
rect 384938 267117 384944 267129
rect 581200 267117 581206 267129
rect 384938 267089 581206 267117
rect 384938 267077 384944 267089
rect 581200 267077 581206 267089
rect 581258 267077 581264 267129
rect 386032 267003 386038 267055
rect 386090 267043 386096 267055
rect 584752 267043 584758 267055
rect 386090 267015 584758 267043
rect 386090 267003 386096 267015
rect 584752 267003 584758 267015
rect 584810 267003 584816 267055
rect 387760 266929 387766 266981
rect 387818 266969 387824 266981
rect 588304 266969 588310 266981
rect 387818 266941 588310 266969
rect 387818 266929 387824 266941
rect 588304 266929 588310 266941
rect 588362 266929 588368 266981
rect 301840 266855 301846 266907
rect 301898 266895 301904 266907
rect 375280 266895 375286 266907
rect 301898 266867 375286 266895
rect 301898 266855 301904 266867
rect 375280 266855 375286 266867
rect 375338 266855 375344 266907
rect 393232 266855 393238 266907
rect 393290 266895 393296 266907
rect 602512 266895 602518 266907
rect 393290 266867 602518 266895
rect 393290 266855 393296 266867
rect 602512 266855 602518 266867
rect 602570 266855 602576 266907
rect 305008 266781 305014 266833
rect 305066 266821 305072 266833
rect 383536 266821 383542 266833
rect 305066 266793 383542 266821
rect 305066 266781 305072 266793
rect 383536 266781 383542 266793
rect 383594 266781 383600 266833
rect 394672 266781 394678 266833
rect 394730 266821 394736 266833
rect 606064 266821 606070 266833
rect 394730 266793 606070 266821
rect 394730 266781 394736 266793
rect 606064 266781 606070 266793
rect 606122 266781 606128 266833
rect 306160 266707 306166 266759
rect 306218 266747 306224 266759
rect 386128 266747 386134 266759
rect 306218 266719 386134 266747
rect 306218 266707 306224 266719
rect 386128 266707 386134 266719
rect 386186 266707 386192 266759
rect 397552 266707 397558 266759
rect 397610 266747 397616 266759
rect 613072 266747 613078 266759
rect 397610 266719 613078 266747
rect 397610 266707 397616 266719
rect 613072 266707 613078 266719
rect 613130 266707 613136 266759
rect 308080 266633 308086 266685
rect 308138 266673 308144 266685
rect 390928 266673 390934 266685
rect 308138 266645 390934 266673
rect 308138 266633 308144 266645
rect 390928 266633 390934 266645
rect 390986 266633 390992 266685
rect 398224 266633 398230 266685
rect 398282 266673 398288 266685
rect 614320 266673 614326 266685
rect 398282 266645 614326 266673
rect 398282 266633 398288 266645
rect 614320 266633 614326 266645
rect 614378 266633 614384 266685
rect 308752 266559 308758 266611
rect 308810 266599 308816 266611
rect 392944 266599 392950 266611
rect 308810 266571 392950 266599
rect 308810 266559 308816 266571
rect 392944 266559 392950 266571
rect 393002 266559 393008 266611
rect 400624 266559 400630 266611
rect 400682 266599 400688 266611
rect 620176 266599 620182 266611
rect 400682 266571 620182 266599
rect 400682 266559 400688 266571
rect 620176 266559 620182 266571
rect 620234 266559 620240 266611
rect 310672 266485 310678 266537
rect 310730 266525 310736 266537
rect 398032 266525 398038 266537
rect 310730 266497 398038 266525
rect 310730 266485 310736 266497
rect 398032 266485 398038 266497
rect 398090 266485 398096 266537
rect 403216 266485 403222 266537
rect 403274 266525 403280 266537
rect 627280 266525 627286 266537
rect 403274 266497 627286 266525
rect 403274 266485 403280 266497
rect 627280 266485 627286 266497
rect 627338 266485 627344 266537
rect 313072 266411 313078 266463
rect 313130 266451 313136 266463
rect 403888 266451 403894 266463
rect 313130 266423 403894 266451
rect 313130 266411 313136 266423
rect 403888 266411 403894 266423
rect 403946 266411 403952 266463
rect 406096 266411 406102 266463
rect 406154 266451 406160 266463
rect 634384 266451 634390 266463
rect 406154 266423 634390 266451
rect 406154 266411 406160 266423
rect 634384 266411 634390 266423
rect 634442 266411 634448 266463
rect 313552 266337 313558 266389
rect 313610 266377 313616 266389
rect 405040 266377 405046 266389
rect 313610 266349 405046 266377
rect 313610 266337 313616 266349
rect 405040 266337 405046 266349
rect 405098 266337 405104 266389
rect 409168 266337 409174 266389
rect 409226 266377 409232 266389
rect 641488 266377 641494 266389
rect 409226 266349 641494 266377
rect 409226 266337 409232 266349
rect 641488 266337 641494 266349
rect 641546 266337 641552 266389
rect 348880 266263 348886 266315
rect 348938 266303 348944 266315
rect 492592 266303 492598 266315
rect 348938 266275 492598 266303
rect 348938 266263 348944 266275
rect 492592 266263 492598 266275
rect 492650 266263 492656 266315
rect 346000 266189 346006 266241
rect 346058 266229 346064 266241
rect 485488 266229 485494 266241
rect 346058 266201 485494 266229
rect 346058 266189 346064 266201
rect 485488 266189 485494 266201
rect 485546 266189 485552 266241
rect 343312 266115 343318 266167
rect 343370 266155 343376 266167
rect 478384 266155 478390 266167
rect 343370 266127 478390 266155
rect 343370 266115 343376 266127
rect 478384 266115 478390 266127
rect 478442 266115 478448 266167
rect 340240 266041 340246 266093
rect 340298 266081 340304 266093
rect 471280 266081 471286 266093
rect 340298 266053 471286 266081
rect 340298 266041 340304 266053
rect 471280 266041 471286 266053
rect 471338 266041 471344 266093
rect 337360 265967 337366 266019
rect 337418 266007 337424 266019
rect 464176 266007 464182 266019
rect 337418 265979 464182 266007
rect 337418 265967 337424 265979
rect 464176 265967 464182 265979
rect 464234 265967 464240 266019
rect 334768 265893 334774 265945
rect 334826 265933 334832 265945
rect 457072 265933 457078 265945
rect 334826 265905 457078 265933
rect 334826 265893 334832 265905
rect 457072 265893 457078 265905
rect 457130 265893 457136 265945
rect 331888 265819 331894 265871
rect 331946 265859 331952 265871
rect 449968 265859 449974 265871
rect 331946 265831 449974 265859
rect 331946 265819 331952 265831
rect 449968 265819 449974 265831
rect 450026 265819 450032 265871
rect 408016 265745 408022 265797
rect 408074 265785 408080 265797
rect 523984 265785 523990 265797
rect 408074 265757 523990 265785
rect 408074 265745 408080 265757
rect 523984 265745 523990 265757
rect 524042 265745 524048 265797
rect 327568 265671 327574 265723
rect 327626 265711 327632 265723
rect 439312 265711 439318 265723
rect 327626 265683 439318 265711
rect 327626 265671 327632 265683
rect 439312 265671 439318 265683
rect 439370 265671 439376 265723
rect 324496 265597 324502 265649
rect 324554 265637 324560 265649
rect 432304 265637 432310 265649
rect 324554 265609 432310 265637
rect 324554 265597 324560 265609
rect 432304 265597 432310 265609
rect 432362 265597 432368 265649
rect 321616 265523 321622 265575
rect 321674 265563 321680 265575
rect 425200 265563 425206 265575
rect 321674 265535 425206 265563
rect 321674 265523 321680 265535
rect 425200 265523 425206 265535
rect 425258 265523 425264 265575
rect 319024 265449 319030 265501
rect 319082 265489 319088 265501
rect 418096 265489 418102 265501
rect 319082 265461 418102 265489
rect 319082 265449 319088 265461
rect 418096 265449 418102 265461
rect 418154 265449 418160 265501
rect 656560 265375 656566 265427
rect 656618 265415 656624 265427
rect 676240 265415 676246 265427
rect 656618 265387 676246 265415
rect 656618 265375 656624 265387
rect 676240 265375 676246 265387
rect 676298 265375 676304 265427
rect 656464 265227 656470 265279
rect 656522 265267 656528 265279
rect 676144 265267 676150 265279
rect 656522 265239 676150 265267
rect 656522 265227 656528 265239
rect 676144 265227 676150 265239
rect 676202 265227 676208 265279
rect 656080 265079 656086 265131
rect 656138 265119 656144 265131
rect 676336 265119 676342 265131
rect 656138 265091 676342 265119
rect 656138 265079 656144 265091
rect 676336 265079 676342 265091
rect 676394 265079 676400 265131
rect 23152 265005 23158 265057
rect 23210 265045 23216 265057
rect 43504 265045 43510 265057
rect 23210 265017 43510 265045
rect 23210 265005 23216 265017
rect 43504 265005 43510 265017
rect 43562 265005 43568 265057
rect 671824 265005 671830 265057
rect 671882 265045 671888 265057
rect 673264 265045 673270 265057
rect 671882 265017 673270 265045
rect 671882 265005 671888 265017
rect 673264 265005 673270 265017
rect 673322 265045 673328 265057
rect 676240 265045 676246 265057
rect 673322 265017 676246 265045
rect 673322 265005 673328 265017
rect 676240 265005 676246 265017
rect 676298 265005 676304 265057
rect 43312 264931 43318 264983
rect 43370 264971 43376 264983
rect 44272 264971 44278 264983
rect 43370 264943 44278 264971
rect 43370 264931 43376 264943
rect 44272 264931 44278 264943
rect 44330 264971 44336 264983
rect 669808 264971 669814 264983
rect 44330 264943 669814 264971
rect 44330 264931 44336 264943
rect 669808 264931 669814 264943
rect 669866 264931 669872 264983
rect 43216 264857 43222 264909
rect 43274 264897 43280 264909
rect 44176 264897 44182 264909
rect 43274 264869 44182 264897
rect 43274 264857 43280 264869
rect 44176 264857 44182 264869
rect 44234 264897 44240 264909
rect 669616 264897 669622 264909
rect 44234 264869 669622 264897
rect 44234 264857 44240 264869
rect 669616 264857 669622 264869
rect 669674 264857 669680 264909
rect 365680 264783 365686 264835
rect 365738 264823 365744 264835
rect 475984 264823 475990 264835
rect 365738 264795 475990 264823
rect 365738 264783 365744 264795
rect 475984 264783 475990 264795
rect 476042 264783 476048 264835
rect 325360 264709 325366 264761
rect 325418 264749 325424 264761
rect 433456 264749 433462 264761
rect 325418 264721 433462 264749
rect 325418 264709 325424 264721
rect 433456 264709 433462 264721
rect 433514 264709 433520 264761
rect 362800 264635 362806 264687
rect 362858 264675 362864 264687
rect 468880 264675 468886 264687
rect 362858 264647 468886 264675
rect 362858 264635 362864 264647
rect 468880 264635 468886 264647
rect 468938 264635 468944 264687
rect 357616 264561 357622 264613
rect 357674 264601 357680 264613
rect 461776 264601 461782 264613
rect 357674 264573 461782 264601
rect 357674 264561 357680 264573
rect 461776 264561 461782 264573
rect 461834 264561 461840 264613
rect 328048 264487 328054 264539
rect 328106 264527 328112 264539
rect 440560 264527 440566 264539
rect 328106 264499 440566 264527
rect 328106 264487 328112 264499
rect 440560 264487 440566 264499
rect 440618 264487 440624 264539
rect 343792 264413 343798 264465
rect 343850 264453 343856 264465
rect 447664 264453 447670 264465
rect 343850 264425 447670 264453
rect 343850 264413 343856 264425
rect 447664 264413 447670 264425
rect 447722 264413 447728 264465
rect 351376 264339 351382 264391
rect 351434 264379 351440 264391
rect 454768 264379 454774 264391
rect 351434 264351 454774 264379
rect 351434 264339 351440 264351
rect 454768 264339 454774 264351
rect 454826 264339 454832 264391
rect 399376 264043 399382 264095
rect 399434 264083 399440 264095
rect 411664 264083 411670 264095
rect 399434 264055 411670 264083
rect 399434 264043 399440 264055
rect 411664 264043 411670 264055
rect 411722 264043 411728 264095
rect 390832 263969 390838 264021
rect 390890 264009 390896 264021
rect 596560 264009 596566 264021
rect 390890 263981 596566 264009
rect 390890 263969 390896 263981
rect 596560 263969 596566 263981
rect 596618 263969 596624 264021
rect 392272 263895 392278 263947
rect 392330 263935 392336 263947
rect 600112 263935 600118 263947
rect 392330 263907 600118 263935
rect 392330 263895 392336 263907
rect 600112 263895 600118 263907
rect 600170 263895 600176 263947
rect 395440 263821 395446 263873
rect 395498 263861 395504 263873
rect 607216 263861 607222 263873
rect 395498 263833 607222 263861
rect 395498 263821 395504 263833
rect 607216 263821 607222 263833
rect 607274 263821 607280 263873
rect 401104 263747 401110 263799
rect 401162 263787 401168 263799
rect 401162 263759 411614 263787
rect 401162 263747 401168 263759
rect 403984 263673 403990 263725
rect 404042 263713 404048 263725
rect 411586 263713 411614 263759
rect 411664 263747 411670 263799
rect 411722 263787 411728 263799
rect 617872 263787 617878 263799
rect 411722 263759 617878 263787
rect 411722 263747 411728 263759
rect 617872 263747 617878 263759
rect 617930 263747 617936 263799
rect 621424 263713 621430 263725
rect 404042 263685 411518 263713
rect 411586 263685 621430 263713
rect 404042 263673 404048 263685
rect 23536 263599 23542 263651
rect 23594 263639 23600 263651
rect 44176 263639 44182 263651
rect 23594 263611 44182 263639
rect 23594 263599 23600 263611
rect 44176 263599 44182 263611
rect 44234 263599 44240 263651
rect 405424 263599 405430 263651
rect 405482 263639 405488 263651
rect 411490 263639 411518 263685
rect 621424 263673 621430 263685
rect 621482 263673 621488 263725
rect 628432 263639 628438 263651
rect 405482 263611 411422 263639
rect 411490 263611 628438 263639
rect 405482 263599 405488 263611
rect 23056 263525 23062 263577
rect 23114 263565 23120 263577
rect 44272 263565 44278 263577
rect 23114 263537 44278 263565
rect 23114 263525 23120 263537
rect 44272 263525 44278 263537
rect 44330 263525 44336 263577
rect 409648 263525 409654 263577
rect 409706 263525 409712 263577
rect 411394 263565 411422 263611
rect 628432 263599 628438 263611
rect 628490 263599 628496 263651
rect 631984 263565 631990 263577
rect 411394 263537 631990 263565
rect 631984 263525 631990 263537
rect 632042 263525 632048 263577
rect 409666 263491 409694 263525
rect 642640 263491 642646 263503
rect 409666 263463 642646 263491
rect 642640 263451 642646 263463
rect 642698 263451 642704 263503
rect 23344 262119 23350 262171
rect 23402 262159 23408 262171
rect 43312 262159 43318 262171
rect 23402 262131 43318 262159
rect 23402 262119 23408 262131
rect 43312 262119 43318 262131
rect 43370 262119 43376 262171
rect 420400 262119 420406 262171
rect 420458 262159 420464 262171
rect 606160 262159 606166 262171
rect 420458 262131 606166 262159
rect 420458 262119 420464 262131
rect 606160 262119 606166 262131
rect 606218 262119 606224 262171
rect 675184 262119 675190 262171
rect 675242 262159 675248 262171
rect 676240 262159 676246 262171
rect 675242 262131 676246 262159
rect 675242 262119 675248 262131
rect 676240 262119 676246 262131
rect 676298 262119 676304 262171
rect 674800 259899 674806 259951
rect 674858 259939 674864 259951
rect 676240 259939 676246 259951
rect 674858 259911 676246 259939
rect 674858 259899 674864 259911
rect 676240 259899 676246 259911
rect 676298 259899 676304 259951
rect 673264 259529 673270 259581
rect 673322 259569 673328 259581
rect 673456 259569 673462 259581
rect 673322 259541 673462 259569
rect 673322 259529 673328 259541
rect 673456 259529 673462 259541
rect 673514 259529 673520 259581
rect 674704 259307 674710 259359
rect 674762 259347 674768 259359
rect 676048 259347 676054 259359
rect 674762 259319 676054 259347
rect 674762 259307 674768 259319
rect 676048 259307 676054 259319
rect 676106 259307 676112 259359
rect 420400 259233 420406 259285
rect 420458 259273 420464 259285
rect 606256 259273 606262 259285
rect 420458 259245 606262 259273
rect 420458 259233 420464 259245
rect 606256 259233 606262 259245
rect 606314 259233 606320 259285
rect 675280 259233 675286 259285
rect 675338 259273 675344 259285
rect 676240 259273 676246 259285
rect 675338 259245 676246 259273
rect 675338 259233 675344 259245
rect 676240 259233 676246 259245
rect 676298 259233 676304 259285
rect 151600 257753 151606 257805
rect 151658 257793 151664 257805
rect 169744 257793 169750 257805
rect 151658 257765 169750 257793
rect 151658 257753 151664 257765
rect 169744 257753 169750 257765
rect 169802 257753 169808 257805
rect 187216 257753 187222 257805
rect 187274 257793 187280 257805
rect 189712 257793 189718 257805
rect 187274 257765 189718 257793
rect 187274 257753 187280 257765
rect 189712 257753 189718 257765
rect 189770 257753 189776 257805
rect 41776 256421 41782 256473
rect 41834 256461 41840 256473
rect 56080 256461 56086 256473
rect 41834 256433 56086 256461
rect 41834 256421 41840 256433
rect 56080 256421 56086 256433
rect 56138 256421 56144 256473
rect 674608 256421 674614 256473
rect 674666 256461 674672 256473
rect 675952 256461 675958 256473
rect 674666 256433 675958 256461
rect 674666 256421 674672 256433
rect 675952 256421 675958 256433
rect 676010 256421 676016 256473
rect 41584 256347 41590 256399
rect 41642 256387 41648 256399
rect 58960 256387 58966 256399
rect 41642 256359 58966 256387
rect 41642 256347 41648 256359
rect 58960 256347 58966 256359
rect 59018 256347 59024 256399
rect 420400 256347 420406 256399
rect 420458 256387 420464 256399
rect 606352 256387 606358 256399
rect 420458 256359 606358 256387
rect 420458 256347 420464 256359
rect 606352 256347 606358 256359
rect 606410 256347 606416 256399
rect 674896 256347 674902 256399
rect 674954 256387 674960 256399
rect 676048 256387 676054 256399
rect 674954 256359 676054 256387
rect 674954 256347 674960 256359
rect 676048 256347 676054 256359
rect 676106 256347 676112 256399
rect 41776 255977 41782 256029
rect 41834 256017 41840 256029
rect 53200 256017 53206 256029
rect 41834 255989 53206 256017
rect 41834 255977 41840 255989
rect 53200 255977 53206 255989
rect 53258 255977 53264 256029
rect 41776 255533 41782 255585
rect 41834 255573 41840 255585
rect 43408 255573 43414 255585
rect 41834 255545 43414 255573
rect 41834 255533 41840 255545
rect 43408 255533 43414 255545
rect 43466 255533 43472 255585
rect 41776 255015 41782 255067
rect 41834 255055 41840 255067
rect 43408 255055 43414 255067
rect 41834 255027 43414 255055
rect 41834 255015 41840 255027
rect 43408 255015 43414 255027
rect 43466 255015 43472 255067
rect 47920 254941 47926 254993
rect 47978 254981 47984 254993
rect 186064 254981 186070 254993
rect 47978 254953 186070 254981
rect 47978 254941 47984 254953
rect 186064 254941 186070 254953
rect 186122 254941 186128 254993
rect 48016 254867 48022 254919
rect 48074 254907 48080 254919
rect 186256 254907 186262 254919
rect 48074 254879 186262 254907
rect 48074 254867 48080 254879
rect 186256 254867 186262 254879
rect 186314 254867 186320 254919
rect 420400 253461 420406 253513
rect 420458 253501 420464 253513
rect 603280 253501 603286 253513
rect 420458 253473 603286 253501
rect 420458 253461 420464 253473
rect 603280 253461 603286 253473
rect 603338 253461 603344 253513
rect 646672 253461 646678 253513
rect 646730 253501 646736 253513
rect 679792 253501 679798 253513
rect 646730 253473 679798 253501
rect 646730 253461 646736 253473
rect 679792 253461 679798 253473
rect 679850 253461 679856 253513
rect 141040 252499 141046 252551
rect 141098 252539 141104 252551
rect 171376 252539 171382 252551
rect 141098 252511 171382 252539
rect 141098 252499 141104 252511
rect 171376 252499 171382 252511
rect 171434 252499 171440 252551
rect 106480 252425 106486 252477
rect 106538 252465 106544 252477
rect 156880 252465 156886 252477
rect 106538 252437 156886 252465
rect 106538 252425 106544 252437
rect 156880 252425 156886 252437
rect 156938 252425 156944 252477
rect 97840 252351 97846 252403
rect 97898 252391 97904 252403
rect 154000 252391 154006 252403
rect 97898 252363 154006 252391
rect 97898 252351 97904 252363
rect 154000 252351 154006 252363
rect 154058 252351 154064 252403
rect 103600 252277 103606 252329
rect 103658 252317 103664 252329
rect 159760 252317 159766 252329
rect 103658 252289 159766 252317
rect 103658 252277 103664 252289
rect 159760 252277 159766 252289
rect 159818 252277 159824 252329
rect 109360 252203 109366 252255
rect 109418 252243 109424 252255
rect 177040 252243 177046 252255
rect 109418 252215 177046 252243
rect 109418 252203 109424 252215
rect 177040 252203 177046 252215
rect 177098 252203 177104 252255
rect 86320 252129 86326 252181
rect 86378 252169 86384 252181
rect 165520 252169 165526 252181
rect 86378 252141 165526 252169
rect 86378 252129 86384 252141
rect 165520 252129 165526 252141
rect 165578 252129 165584 252181
rect 94960 252055 94966 252107
rect 95018 252095 95024 252107
rect 174160 252095 174166 252107
rect 95018 252067 174166 252095
rect 95018 252055 95024 252067
rect 174160 252055 174166 252067
rect 174218 252055 174224 252107
rect 92080 251981 92086 252033
rect 92138 252021 92144 252033
rect 182800 252021 182806 252033
rect 92138 251993 182806 252021
rect 92138 251981 92144 251993
rect 182800 251981 182806 251993
rect 182858 251981 182864 252033
rect 670384 250649 670390 250701
rect 670442 250689 670448 250701
rect 675376 250689 675382 250701
rect 670442 250661 675382 250689
rect 670442 250649 670448 250661
rect 675376 250649 675382 250661
rect 675434 250649 675440 250701
rect 420400 250575 420406 250627
rect 420458 250615 420464 250627
rect 603376 250615 603382 250627
rect 420458 250587 603382 250615
rect 420458 250575 420464 250587
rect 603376 250575 603382 250587
rect 603434 250575 603440 250627
rect 120880 249835 120886 249887
rect 120938 249875 120944 249887
rect 145552 249875 145558 249887
rect 120938 249847 145558 249875
rect 120938 249835 120944 249847
rect 145552 249835 145558 249847
rect 145610 249835 145616 249887
rect 132400 249761 132406 249813
rect 132458 249801 132464 249813
rect 162736 249801 162742 249813
rect 132458 249773 162742 249801
rect 132458 249761 132464 249773
rect 162736 249761 162742 249773
rect 162794 249761 162800 249813
rect 135280 249687 135286 249739
rect 135338 249727 135344 249739
rect 168496 249727 168502 249739
rect 135338 249699 168502 249727
rect 135338 249687 135344 249699
rect 168496 249687 168502 249699
rect 168554 249687 168560 249739
rect 118000 249613 118006 249665
rect 118058 249653 118064 249665
rect 156976 249653 156982 249665
rect 118058 249625 156982 249653
rect 118058 249613 118064 249625
rect 156976 249613 156982 249625
rect 157034 249613 157040 249665
rect 138160 249539 138166 249591
rect 138218 249579 138224 249591
rect 180016 249579 180022 249591
rect 138218 249551 180022 249579
rect 138218 249539 138224 249551
rect 180016 249539 180022 249551
rect 180074 249539 180080 249591
rect 126640 249465 126646 249517
rect 126698 249505 126704 249517
rect 177232 249505 177238 249517
rect 126698 249477 177238 249505
rect 126698 249465 126704 249477
rect 177232 249465 177238 249477
rect 177290 249465 177296 249517
rect 123760 249391 123766 249443
rect 123818 249431 123824 249443
rect 174448 249431 174454 249443
rect 123818 249403 174454 249431
rect 123818 249391 123824 249403
rect 174448 249391 174454 249403
rect 174506 249391 174512 249443
rect 80560 249317 80566 249369
rect 80618 249357 80624 249369
rect 145456 249357 145462 249369
rect 80618 249329 145462 249357
rect 80618 249317 80624 249329
rect 145456 249317 145462 249329
rect 145514 249317 145520 249369
rect 77680 249243 77686 249295
rect 77738 249283 77744 249295
rect 145360 249283 145366 249295
rect 77738 249255 145366 249283
rect 77738 249243 77744 249255
rect 145360 249243 145366 249255
rect 145418 249243 145424 249295
rect 48208 249169 48214 249221
rect 48266 249209 48272 249221
rect 186736 249209 186742 249221
rect 48266 249181 186742 249209
rect 48266 249169 48272 249181
rect 186736 249169 186742 249181
rect 186794 249169 186800 249221
rect 47728 249095 47734 249147
rect 47786 249135 47792 249147
rect 186448 249135 186454 249147
rect 47786 249107 186454 249135
rect 47786 249095 47792 249107
rect 186448 249095 186454 249107
rect 186506 249095 186512 249147
rect 674800 247911 674806 247963
rect 674858 247951 674864 247963
rect 675376 247951 675382 247963
rect 674858 247923 675382 247951
rect 674858 247911 674864 247923
rect 675376 247911 675382 247923
rect 675434 247911 675440 247963
rect 420304 247763 420310 247815
rect 420362 247803 420368 247815
rect 603472 247803 603478 247815
rect 420362 247775 603478 247803
rect 420362 247763 420368 247775
rect 603472 247763 603478 247775
rect 603530 247763 603536 247815
rect 420400 247689 420406 247741
rect 420458 247729 420464 247741
rect 629200 247729 629206 247741
rect 420458 247701 629206 247729
rect 420458 247689 420464 247701
rect 629200 247689 629206 247701
rect 629258 247689 629264 247741
rect 655888 247615 655894 247667
rect 655946 247655 655952 247667
rect 670384 247655 670390 247667
rect 655946 247627 670390 247655
rect 655946 247615 655952 247627
rect 670384 247615 670390 247627
rect 670442 247615 670448 247667
rect 674800 247023 674806 247075
rect 674858 247063 674864 247075
rect 675472 247063 675478 247075
rect 674858 247035 675478 247063
rect 674858 247023 674864 247035
rect 675472 247023 675478 247035
rect 675530 247023 675536 247075
rect 112240 246653 112246 246705
rect 112298 246693 112304 246705
rect 185776 246693 185782 246705
rect 112298 246665 185782 246693
rect 112298 246653 112304 246665
rect 185776 246653 185782 246665
rect 185834 246653 185840 246705
rect 47536 246579 47542 246631
rect 47594 246619 47600 246631
rect 186352 246619 186358 246631
rect 47594 246591 186358 246619
rect 47594 246579 47600 246591
rect 186352 246579 186358 246591
rect 186410 246579 186416 246631
rect 47632 246505 47638 246557
rect 47690 246545 47696 246557
rect 186640 246545 186646 246557
rect 47690 246517 186646 246545
rect 47690 246505 47696 246517
rect 186640 246505 186646 246517
rect 186698 246505 186704 246557
rect 47440 246431 47446 246483
rect 47498 246471 47504 246483
rect 186544 246471 186550 246483
rect 47498 246443 186550 246471
rect 47498 246431 47504 246443
rect 186544 246431 186550 246443
rect 186602 246431 186608 246483
rect 45808 246357 45814 246409
rect 45866 246397 45872 246409
rect 186928 246397 186934 246409
rect 45866 246369 186934 246397
rect 45866 246357 45872 246369
rect 186928 246357 186934 246369
rect 186986 246357 186992 246409
rect 44848 246283 44854 246335
rect 44906 246323 44912 246335
rect 186160 246323 186166 246335
rect 44906 246295 186166 246323
rect 44906 246283 44912 246295
rect 186160 246283 186166 246295
rect 186218 246283 186224 246335
rect 44560 246209 44566 246261
rect 44618 246249 44624 246261
rect 185968 246249 185974 246261
rect 44618 246221 185974 246249
rect 44618 246209 44624 246221
rect 185968 246209 185974 246221
rect 186026 246209 186032 246261
rect 674896 245839 674902 245891
rect 674954 245879 674960 245891
rect 675376 245879 675382 245891
rect 674954 245851 675382 245879
rect 674954 245839 674960 245851
rect 675376 245839 675382 245851
rect 675434 245839 675440 245891
rect 41584 245469 41590 245521
rect 41642 245509 41648 245521
rect 43024 245509 43030 245521
rect 41642 245481 43030 245509
rect 41642 245469 41648 245481
rect 43024 245469 43030 245481
rect 43082 245469 43088 245521
rect 41680 245395 41686 245447
rect 41738 245435 41744 245447
rect 42832 245435 42838 245447
rect 41738 245407 42838 245435
rect 41738 245395 41744 245407
rect 42832 245395 42838 245407
rect 42890 245395 42896 245447
rect 41872 245025 41878 245077
rect 41930 245065 41936 245077
rect 42928 245065 42934 245077
rect 41930 245037 42934 245065
rect 41930 245025 41936 245037
rect 42928 245025 42934 245037
rect 42986 245025 42992 245077
rect 44656 244951 44662 245003
rect 44714 244991 44720 245003
rect 186832 244991 186838 245003
rect 44714 244963 186838 244991
rect 44714 244951 44720 244963
rect 186832 244951 186838 244963
rect 186890 244951 186896 245003
rect 41584 244877 41590 244929
rect 41642 244917 41648 244929
rect 142480 244917 142486 244929
rect 41642 244889 142486 244917
rect 41642 244877 41648 244889
rect 142480 244877 142486 244889
rect 142538 244877 142544 244929
rect 41680 244803 41686 244855
rect 41738 244843 41744 244855
rect 159952 244843 159958 244855
rect 41738 244815 159958 244843
rect 41738 244803 41744 244815
rect 159952 244803 159958 244815
rect 160010 244803 160016 244855
rect 420400 244803 420406 244855
rect 420458 244843 420464 244855
rect 629296 244843 629302 244855
rect 420458 244815 629302 244843
rect 420458 244803 420464 244815
rect 629296 244803 629302 244815
rect 629354 244803 629360 244855
rect 41488 244655 41494 244707
rect 41546 244695 41552 244707
rect 42736 244695 42742 244707
rect 41546 244667 42742 244695
rect 41546 244655 41552 244667
rect 42736 244655 42742 244667
rect 42794 244655 42800 244707
rect 169744 243027 169750 243079
rect 169802 243067 169808 243079
rect 180112 243067 180118 243079
rect 169802 243039 180118 243067
rect 169802 243027 169808 243039
rect 180112 243027 180118 243039
rect 180170 243027 180176 243079
rect 44752 242805 44758 242857
rect 44810 242845 44816 242857
rect 185680 242845 185686 242857
rect 44810 242817 185686 242845
rect 44810 242805 44816 242817
rect 185680 242805 185686 242817
rect 185738 242805 185744 242857
rect 44848 242731 44854 242783
rect 44906 242771 44912 242783
rect 185872 242771 185878 242783
rect 44906 242743 185878 242771
rect 44906 242731 44912 242743
rect 185872 242731 185878 242743
rect 185930 242731 185936 242783
rect 674608 242731 674614 242783
rect 674666 242771 674672 242783
rect 675376 242771 675382 242783
rect 674666 242743 675382 242771
rect 674666 242731 674672 242743
rect 675376 242731 675382 242743
rect 675434 242731 675440 242783
rect 44560 242657 44566 242709
rect 44618 242697 44624 242709
rect 187024 242697 187030 242709
rect 44618 242669 187030 242697
rect 44618 242657 44624 242669
rect 187024 242657 187030 242669
rect 187082 242657 187088 242709
rect 41584 242583 41590 242635
rect 41642 242623 41648 242635
rect 142672 242623 142678 242635
rect 41642 242595 142678 242623
rect 41642 242583 41648 242595
rect 142672 242583 142678 242595
rect 142730 242583 142736 242635
rect 420304 241917 420310 241969
rect 420362 241957 420368 241969
rect 600400 241957 600406 241969
rect 420362 241929 600406 241957
rect 420362 241917 420368 241929
rect 600400 241917 600406 241929
rect 600458 241917 600464 241969
rect 41776 240585 41782 240637
rect 41834 240585 41840 240637
rect 41794 240415 41822 240585
rect 41776 240363 41782 240415
rect 41834 240363 41840 240415
rect 368656 239919 368662 239971
rect 368714 239959 368720 239971
rect 412048 239959 412054 239971
rect 368714 239931 412054 239959
rect 368714 239919 368720 239931
rect 412048 239919 412054 239931
rect 412106 239919 412112 239971
rect 413008 239919 413014 239971
rect 413066 239959 413072 239971
rect 442192 239959 442198 239971
rect 413066 239931 442198 239959
rect 413066 239919 413072 239931
rect 442192 239919 442198 239931
rect 442250 239919 442256 239971
rect 409552 239845 409558 239897
rect 409610 239885 409616 239897
rect 412144 239885 412150 239897
rect 409610 239857 412150 239885
rect 409610 239845 409616 239857
rect 412144 239845 412150 239857
rect 412202 239845 412208 239897
rect 350704 239771 350710 239823
rect 350762 239811 350768 239823
rect 508624 239811 508630 239823
rect 350762 239783 508630 239811
rect 350762 239771 350768 239783
rect 508624 239771 508630 239783
rect 508682 239771 508688 239823
rect 360016 239697 360022 239749
rect 360074 239737 360080 239749
rect 434608 239737 434614 239749
rect 360074 239709 434614 239737
rect 360074 239697 360080 239709
rect 434608 239697 434614 239709
rect 434666 239697 434672 239749
rect 366544 239623 366550 239675
rect 366602 239663 366608 239675
rect 446704 239663 446710 239675
rect 366602 239635 446710 239663
rect 366602 239623 366608 239635
rect 446704 239623 446710 239635
rect 446762 239623 446768 239675
rect 396688 239549 396694 239601
rect 396746 239589 396752 239601
rect 412240 239589 412246 239601
rect 396746 239561 412246 239589
rect 396746 239549 396752 239561
rect 412240 239549 412246 239561
rect 412298 239549 412304 239601
rect 412912 239549 412918 239601
rect 412970 239589 412976 239601
rect 495760 239589 495766 239601
rect 412970 239561 495766 239589
rect 412970 239549 412976 239561
rect 495760 239549 495766 239561
rect 495818 239549 495824 239601
rect 383056 239475 383062 239527
rect 383114 239515 383120 239527
rect 470896 239515 470902 239527
rect 383114 239487 470902 239515
rect 383114 239475 383120 239487
rect 470896 239475 470902 239487
rect 470954 239475 470960 239527
rect 371632 239401 371638 239453
rect 371690 239441 371696 239453
rect 458800 239441 458806 239453
rect 371690 239413 458806 239441
rect 371690 239401 371696 239413
rect 458800 239401 458806 239413
rect 458858 239401 458864 239453
rect 406096 239327 406102 239379
rect 406154 239367 406160 239379
rect 412336 239367 412342 239379
rect 406154 239339 412342 239367
rect 406154 239327 406160 239339
rect 412336 239327 412342 239339
rect 412394 239327 412400 239379
rect 412816 239327 412822 239379
rect 412874 239367 412880 239379
rect 502576 239367 502582 239379
rect 412874 239339 502582 239367
rect 412874 239327 412880 239339
rect 502576 239327 502582 239339
rect 502634 239327 502640 239379
rect 378448 239253 378454 239305
rect 378506 239293 378512 239305
rect 488272 239293 488278 239305
rect 378506 239265 488278 239293
rect 378506 239253 378512 239265
rect 488272 239253 488278 239265
rect 488330 239253 488336 239305
rect 398416 239179 398422 239231
rect 398474 239219 398480 239231
rect 532816 239219 532822 239231
rect 398474 239191 532822 239219
rect 398474 239179 398480 239191
rect 532816 239179 532822 239191
rect 532874 239179 532880 239231
rect 411760 239105 411766 239157
rect 411818 239145 411824 239157
rect 412624 239145 412630 239157
rect 411818 239117 412630 239145
rect 411818 239105 411824 239117
rect 412624 239105 412630 239117
rect 412682 239105 412688 239157
rect 420304 239105 420310 239157
rect 420362 239145 420368 239157
rect 599056 239145 599062 239157
rect 420362 239117 599062 239145
rect 420362 239105 420368 239117
rect 599056 239105 599062 239117
rect 599114 239105 599120 239157
rect 380848 239031 380854 239083
rect 380906 239071 380912 239083
rect 412432 239071 412438 239083
rect 380906 239043 412438 239071
rect 380906 239031 380912 239043
rect 412432 239031 412438 239043
rect 412490 239031 412496 239083
rect 324400 238957 324406 239009
rect 324458 238997 324464 239009
rect 455152 238997 455158 239009
rect 324458 238969 455158 238997
rect 324458 238957 324464 238969
rect 455152 238957 455158 238969
rect 455210 238957 455216 239009
rect 323920 238883 323926 238935
rect 323978 238923 323984 238935
rect 455056 238923 455062 238935
rect 323978 238895 455062 238923
rect 323978 238883 323984 238895
rect 455056 238883 455062 238895
rect 455114 238883 455120 238935
rect 326704 238809 326710 238861
rect 326762 238849 326768 238861
rect 462544 238849 462550 238861
rect 326762 238821 462550 238849
rect 326762 238809 326768 238821
rect 462544 238809 462550 238821
rect 462602 238809 462608 238861
rect 328912 238735 328918 238787
rect 328970 238775 328976 238787
rect 464752 238775 464758 238787
rect 328970 238747 464758 238775
rect 328970 238735 328976 238747
rect 464752 238735 464758 238747
rect 464810 238735 464816 238787
rect 329872 238661 329878 238713
rect 329930 238701 329936 238713
rect 468592 238701 468598 238713
rect 329930 238673 468598 238701
rect 329930 238661 329936 238673
rect 468592 238661 468598 238673
rect 468650 238661 468656 238713
rect 332656 238587 332662 238639
rect 332714 238627 332720 238639
rect 474640 238627 474646 238639
rect 332714 238599 474646 238627
rect 332714 238587 332720 238599
rect 474640 238587 474646 238599
rect 474698 238587 474704 238639
rect 335728 238513 335734 238565
rect 335786 238553 335792 238565
rect 480688 238553 480694 238565
rect 335786 238525 480694 238553
rect 335786 238513 335792 238525
rect 480688 238513 480694 238525
rect 480746 238513 480752 238565
rect 336688 238439 336694 238491
rect 336746 238479 336752 238491
rect 479152 238479 479158 238491
rect 336746 238451 479158 238479
rect 336746 238439 336752 238451
rect 479152 238439 479158 238451
rect 479210 238439 479216 238491
rect 338992 238365 338998 238417
rect 339050 238405 339056 238417
rect 486736 238405 486742 238417
rect 339050 238377 486742 238405
rect 339050 238365 339056 238377
rect 486736 238365 486742 238377
rect 486794 238365 486800 238417
rect 341776 238291 341782 238343
rect 341834 238331 341840 238343
rect 492784 238331 492790 238343
rect 341834 238303 492790 238331
rect 341834 238291 341840 238303
rect 492784 238291 492790 238303
rect 492842 238291 492848 238343
rect 345328 238217 345334 238269
rect 345386 238257 345392 238269
rect 500272 238257 500278 238269
rect 345386 238229 500278 238257
rect 345386 238217 345392 238229
rect 500272 238217 500278 238229
rect 500330 238217 500336 238269
rect 346672 238143 346678 238195
rect 346730 238183 346736 238195
rect 503344 238183 503350 238195
rect 346730 238155 503350 238183
rect 346730 238143 346736 238155
rect 503344 238143 503350 238155
rect 503402 238143 503408 238195
rect 349936 238069 349942 238121
rect 349994 238109 350000 238121
rect 509392 238109 509398 238121
rect 349994 238081 509398 238109
rect 349994 238069 350000 238081
rect 509392 238069 509398 238081
rect 509450 238069 509456 238121
rect 353488 237995 353494 238047
rect 353546 238035 353552 238047
rect 514672 238035 514678 238047
rect 353546 238007 514678 238035
rect 353546 237995 353552 238007
rect 514672 237995 514678 238007
rect 514730 237995 514736 238047
rect 352720 237921 352726 237973
rect 352778 237961 352784 237973
rect 512752 237961 512758 237973
rect 352778 237933 512758 237961
rect 352778 237921 352784 237933
rect 512752 237921 512758 237933
rect 512810 237921 512816 237973
rect 355696 237847 355702 237899
rect 355754 237887 355760 237899
rect 521488 237887 521494 237899
rect 355754 237859 521494 237887
rect 355754 237847 355760 237859
rect 521488 237847 521494 237859
rect 521546 237847 521552 237899
rect 358576 237773 358582 237825
rect 358634 237813 358640 237825
rect 526000 237813 526006 237825
rect 358634 237785 526006 237813
rect 358634 237773 358640 237785
rect 526000 237773 526006 237785
rect 526058 237773 526064 237825
rect 363088 237699 363094 237751
rect 363146 237739 363152 237751
rect 535120 237739 535126 237751
rect 363146 237711 535126 237739
rect 363146 237699 363152 237711
rect 535120 237699 535126 237711
rect 535178 237699 535184 237751
rect 275344 237625 275350 237677
rect 275402 237665 275408 237677
rect 357712 237665 357718 237677
rect 275402 237637 357718 237665
rect 275402 237625 275408 237637
rect 357712 237625 357718 237637
rect 357770 237625 357776 237677
rect 361744 237625 361750 237677
rect 361802 237665 361808 237677
rect 533488 237665 533494 237677
rect 361802 237637 533494 237665
rect 361802 237625 361808 237637
rect 533488 237625 533494 237637
rect 533546 237625 533552 237677
rect 277072 237551 277078 237603
rect 277130 237591 277136 237603
rect 363664 237591 363670 237603
rect 277130 237563 363670 237591
rect 277130 237551 277136 237563
rect 363664 237551 363670 237563
rect 363722 237551 363728 237603
rect 364432 237551 364438 237603
rect 364490 237591 364496 237603
rect 535792 237591 535798 237603
rect 364490 237563 535798 237591
rect 364490 237551 364496 237563
rect 535792 237551 535798 237563
rect 535850 237551 535856 237603
rect 320848 237477 320854 237529
rect 320906 237517 320912 237529
rect 449296 237517 449302 237529
rect 320906 237489 449302 237517
rect 320906 237477 320912 237489
rect 449296 237477 449302 237489
rect 449354 237477 449360 237529
rect 317584 237403 317590 237455
rect 317642 237443 317648 237455
rect 444496 237443 444502 237455
rect 317642 237415 444502 237443
rect 317642 237403 317648 237415
rect 444496 237403 444502 237415
rect 444554 237403 444560 237455
rect 317104 237329 317110 237381
rect 317162 237369 317168 237381
rect 441424 237369 441430 237381
rect 317162 237341 441430 237369
rect 317162 237329 317168 237341
rect 441424 237329 441430 237341
rect 441482 237329 441488 237381
rect 314800 237255 314806 237307
rect 314858 237295 314864 237307
rect 438352 237295 438358 237307
rect 314858 237267 438358 237295
rect 314858 237255 314864 237267
rect 438352 237255 438358 237267
rect 438410 237255 438416 237307
rect 311536 237181 311542 237233
rect 311594 237221 311600 237233
rect 432400 237221 432406 237233
rect 311594 237193 432406 237221
rect 311594 237181 311600 237193
rect 432400 237181 432406 237193
rect 432458 237181 432464 237233
rect 308560 237107 308566 237159
rect 308618 237147 308624 237159
rect 411472 237147 411478 237159
rect 308618 237119 411478 237147
rect 308618 237107 308624 237119
rect 411472 237107 411478 237119
rect 411530 237107 411536 237159
rect 411664 237107 411670 237159
rect 411722 237147 411728 237159
rect 412720 237147 412726 237159
rect 411722 237119 412726 237147
rect 411722 237107 411728 237119
rect 412720 237107 412726 237119
rect 412778 237107 412784 237159
rect 310768 237033 310774 237085
rect 310826 237073 310832 237085
rect 411184 237073 411190 237085
rect 310826 237045 411190 237073
rect 310826 237033 310832 237045
rect 411184 237033 411190 237045
rect 411242 237033 411248 237085
rect 411568 237033 411574 237085
rect 411626 237073 411632 237085
rect 412816 237073 412822 237085
rect 411626 237045 412822 237073
rect 411626 237033 411632 237045
rect 412816 237033 412822 237045
rect 412874 237033 412880 237085
rect 305776 236959 305782 237011
rect 305834 236999 305840 237011
rect 420304 236999 420310 237011
rect 305834 236971 420310 236999
rect 305834 236959 305840 236971
rect 420304 236959 420310 236971
rect 420362 236959 420368 237011
rect 300208 236885 300214 236937
rect 300266 236925 300272 236937
rect 407152 236925 407158 236937
rect 300266 236897 407158 236925
rect 300266 236885 300272 236897
rect 407152 236885 407158 236897
rect 407210 236885 407216 236937
rect 408976 236885 408982 236937
rect 409034 236925 409040 236937
rect 413968 236925 413974 236937
rect 409034 236897 413974 236925
rect 409034 236885 409040 236897
rect 413968 236885 413974 236897
rect 414026 236885 414032 236937
rect 279856 236811 279862 236863
rect 279914 236851 279920 236863
rect 368848 236851 368854 236863
rect 279914 236823 368854 236851
rect 279914 236811 279920 236823
rect 368848 236811 368854 236823
rect 368906 236811 368912 236863
rect 382576 236811 382582 236863
rect 382634 236851 382640 236863
rect 388720 236851 388726 236863
rect 382634 236823 388726 236851
rect 382634 236811 382640 236823
rect 388720 236811 388726 236823
rect 388778 236811 388784 236863
rect 406000 236811 406006 236863
rect 406058 236851 406064 236863
rect 409168 236851 409174 236863
rect 406058 236823 409174 236851
rect 406058 236811 406064 236823
rect 409168 236811 409174 236823
rect 409226 236811 409232 236863
rect 411472 236811 411478 236863
rect 411530 236851 411536 236863
rect 426352 236851 426358 236863
rect 411530 236823 426358 236851
rect 411530 236811 411536 236823
rect 426352 236811 426358 236823
rect 426410 236811 426416 236863
rect 278416 236737 278422 236789
rect 278474 236777 278480 236789
rect 366736 236777 366742 236789
rect 278474 236749 366742 236777
rect 278474 236737 278480 236749
rect 366736 236737 366742 236749
rect 366794 236737 366800 236789
rect 388336 236737 388342 236789
rect 388394 236777 388400 236789
rect 389008 236777 389014 236789
rect 388394 236749 389014 236777
rect 388394 236737 388400 236749
rect 389008 236737 389014 236749
rect 389066 236737 389072 236789
rect 389392 236737 389398 236789
rect 389450 236777 389456 236789
rect 409360 236777 409366 236789
rect 389450 236749 409366 236777
rect 389450 236737 389456 236749
rect 409360 236737 409366 236749
rect 409418 236737 409424 236789
rect 411184 236737 411190 236789
rect 411242 236777 411248 236789
rect 428656 236777 428662 236789
rect 411242 236749 428662 236777
rect 411242 236737 411248 236749
rect 428656 236737 428662 236749
rect 428714 236737 428720 236789
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 42736 236703 42742 236715
rect 42218 236675 42742 236703
rect 42218 236663 42224 236675
rect 42736 236663 42742 236675
rect 42794 236663 42800 236715
rect 377776 236663 377782 236715
rect 377834 236703 377840 236715
rect 388624 236703 388630 236715
rect 377834 236675 388630 236703
rect 377834 236663 377840 236675
rect 388624 236663 388630 236675
rect 388682 236663 388688 236715
rect 408688 236663 408694 236715
rect 408746 236703 408752 236715
rect 413680 236703 413686 236715
rect 408746 236675 413686 236703
rect 408746 236663 408752 236675
rect 413680 236663 413686 236675
rect 413738 236663 413744 236715
rect 408784 236589 408790 236641
rect 408842 236629 408848 236641
rect 413392 236629 413398 236641
rect 408842 236601 413398 236629
rect 408842 236589 408848 236601
rect 413392 236589 413398 236601
rect 413450 236589 413456 236641
rect 42736 236515 42742 236567
rect 42794 236555 42800 236567
rect 43024 236555 43030 236567
rect 42794 236527 43030 236555
rect 42794 236515 42800 236527
rect 43024 236515 43030 236527
rect 43082 236515 43088 236567
rect 387952 236515 387958 236567
rect 388010 236555 388016 236567
rect 388624 236555 388630 236567
rect 388010 236527 388630 236555
rect 388010 236515 388016 236527
rect 388624 236515 388630 236527
rect 388682 236515 388688 236567
rect 405904 236515 405910 236567
rect 405962 236555 405968 236567
rect 412528 236555 412534 236567
rect 405962 236527 412534 236555
rect 405962 236515 405968 236527
rect 412528 236515 412534 236527
rect 412586 236515 412592 236567
rect 411472 236441 411478 236493
rect 411530 236481 411536 236493
rect 412912 236481 412918 236493
rect 411530 236453 412918 236481
rect 411530 236441 411536 236453
rect 412912 236441 412918 236453
rect 412970 236441 412976 236493
rect 414544 236367 414550 236419
rect 414602 236407 414608 236419
rect 430096 236407 430102 236419
rect 414602 236379 430102 236407
rect 414602 236367 414608 236379
rect 430096 236367 430102 236379
rect 430154 236367 430160 236419
rect 385936 236293 385942 236345
rect 385994 236333 386000 236345
rect 492016 236333 492022 236345
rect 385994 236305 492022 236333
rect 385994 236293 386000 236305
rect 492016 236293 492022 236305
rect 492074 236293 492080 236345
rect 397360 236219 397366 236271
rect 397418 236259 397424 236271
rect 505648 236259 505654 236271
rect 397418 236231 505654 236259
rect 397418 236219 397424 236231
rect 505648 236219 505654 236231
rect 505706 236219 505712 236271
rect 511600 236185 511606 236197
rect 398818 236157 511606 236185
rect 240208 236071 240214 236123
rect 240266 236111 240272 236123
rect 263728 236111 263734 236123
rect 240266 236083 263734 236111
rect 240266 236071 240272 236083
rect 263728 236071 263734 236083
rect 263786 236071 263792 236123
rect 273040 236071 273046 236123
rect 273098 236111 273104 236123
rect 305104 236111 305110 236123
rect 273098 236083 305110 236111
rect 273098 236071 273104 236083
rect 305104 236071 305110 236083
rect 305162 236071 305168 236123
rect 352144 236071 352150 236123
rect 352202 236111 352208 236123
rect 398818 236111 398846 236157
rect 511600 236145 511606 236157
rect 511658 236145 511664 236197
rect 352202 236083 398846 236111
rect 352202 236071 352208 236083
rect 410032 236071 410038 236123
rect 410090 236111 410096 236123
rect 528496 236111 528502 236123
rect 410090 236083 528502 236111
rect 410090 236071 410096 236083
rect 528496 236071 528502 236083
rect 528554 236071 528560 236123
rect 208432 235997 208438 236049
rect 208490 236037 208496 236049
rect 223216 236037 223222 236049
rect 208490 236009 223222 236037
rect 208490 235997 208496 236009
rect 223216 235997 223222 236009
rect 223274 235997 223280 236049
rect 247984 235997 247990 236049
rect 248042 236037 248048 236049
rect 273712 236037 273718 236049
rect 248042 236009 273718 236037
rect 248042 235997 248048 236009
rect 273712 235997 273718 236009
rect 273770 235997 273776 236049
rect 287056 235997 287062 236049
rect 287114 236037 287120 236049
rect 318256 236037 318262 236049
rect 287114 236009 318262 236037
rect 287114 235997 287120 236009
rect 318256 235997 318262 236009
rect 318314 235997 318320 236049
rect 362512 235997 362518 236049
rect 362570 236037 362576 236049
rect 392752 236037 392758 236049
rect 362570 236009 392758 236037
rect 362570 235997 362576 236009
rect 392752 235997 392758 236009
rect 392810 235997 392816 236049
rect 406000 236037 406006 236049
rect 392866 236009 406006 236037
rect 207472 235923 207478 235975
rect 207530 235963 207536 235975
rect 223984 235963 223990 235975
rect 207530 235935 223990 235963
rect 207530 235923 207536 235935
rect 223984 235923 223990 235935
rect 224042 235923 224048 235975
rect 243280 235923 243286 235975
rect 243338 235963 243344 235975
rect 270928 235963 270934 235975
rect 243338 235935 270934 235963
rect 243338 235923 243344 235935
rect 270928 235923 270934 235935
rect 270986 235923 270992 235975
rect 277552 235923 277558 235975
rect 277610 235963 277616 235975
rect 313936 235963 313942 235975
rect 277610 235935 313942 235963
rect 277610 235923 277616 235935
rect 313936 235923 313942 235935
rect 313994 235923 314000 235975
rect 319888 235923 319894 235975
rect 319946 235963 319952 235975
rect 366544 235963 366550 235975
rect 319946 235935 366550 235963
rect 319946 235923 319952 235935
rect 366544 235923 366550 235935
rect 366602 235923 366608 235975
rect 392866 235963 392894 236009
rect 406000 235997 406006 236009
rect 406058 235997 406064 236049
rect 406288 235997 406294 236049
rect 406346 236037 406352 236049
rect 414640 236037 414646 236049
rect 406346 236009 414646 236037
rect 406346 235997 406352 236009
rect 414640 235997 414646 236009
rect 414698 235997 414704 236049
rect 411664 235963 411670 235975
rect 371746 235935 392894 235963
rect 393058 235935 411670 235963
rect 209680 235849 209686 235901
rect 209738 235889 209744 235901
rect 226192 235889 226198 235901
rect 209738 235861 226198 235889
rect 209738 235849 209744 235861
rect 226192 235849 226198 235861
rect 226250 235849 226256 235901
rect 234256 235849 234262 235901
rect 234314 235889 234320 235901
rect 264688 235889 264694 235901
rect 234314 235861 264694 235889
rect 234314 235849 234320 235861
rect 264688 235849 264694 235861
rect 264746 235849 264752 235901
rect 276112 235849 276118 235901
rect 276170 235889 276176 235901
rect 310096 235889 310102 235901
rect 276170 235861 310102 235889
rect 276170 235849 276176 235861
rect 310096 235849 310102 235861
rect 310154 235849 310160 235901
rect 313840 235849 313846 235901
rect 313898 235889 313904 235901
rect 360016 235889 360022 235901
rect 313898 235861 360022 235889
rect 313898 235849 313904 235861
rect 360016 235849 360022 235861
rect 360074 235849 360080 235901
rect 371632 235889 371638 235901
rect 368626 235861 371638 235889
rect 208912 235775 208918 235827
rect 208970 235815 208976 235827
rect 226960 235815 226966 235827
rect 208970 235787 226966 235815
rect 208970 235775 208976 235787
rect 226960 235775 226966 235787
rect 227018 235775 227024 235827
rect 237520 235775 237526 235827
rect 237578 235815 237584 235827
rect 267952 235815 267958 235827
rect 237578 235787 267958 235815
rect 237578 235775 237584 235787
rect 267952 235775 267958 235787
rect 268010 235775 268016 235827
rect 279280 235775 279286 235827
rect 279338 235815 279344 235827
rect 318352 235815 318358 235827
rect 279338 235787 318358 235815
rect 279338 235775 279344 235787
rect 318352 235775 318358 235787
rect 318410 235775 318416 235827
rect 326128 235775 326134 235827
rect 326186 235815 326192 235827
rect 368626 235815 368654 235861
rect 371632 235849 371638 235861
rect 371690 235849 371696 235901
rect 326186 235787 368654 235815
rect 326186 235775 326192 235787
rect 211216 235701 211222 235753
rect 211274 235741 211280 235753
rect 229264 235741 229270 235753
rect 211274 235713 229270 235741
rect 211274 235701 211280 235713
rect 229264 235701 229270 235713
rect 229322 235701 229328 235753
rect 231184 235701 231190 235753
rect 231242 235741 231248 235753
rect 259024 235741 259030 235753
rect 231242 235713 259030 235741
rect 231242 235701 231248 235713
rect 259024 235701 259030 235713
rect 259082 235701 259088 235753
rect 262864 235701 262870 235753
rect 262922 235741 262928 235753
rect 305008 235741 305014 235753
rect 262922 235713 305014 235741
rect 262922 235701 262928 235713
rect 305008 235701 305014 235713
rect 305066 235701 305072 235753
rect 364048 235701 364054 235753
rect 364106 235741 364112 235753
rect 371746 235741 371774 235935
rect 371824 235849 371830 235901
rect 371882 235889 371888 235901
rect 392560 235889 392566 235901
rect 371882 235861 392566 235889
rect 371882 235849 371888 235861
rect 392560 235849 392566 235861
rect 392618 235849 392624 235901
rect 386704 235775 386710 235827
rect 386762 235815 386768 235827
rect 393058 235815 393086 235935
rect 411664 235923 411670 235935
rect 411722 235923 411728 235975
rect 401200 235849 401206 235901
rect 401258 235889 401264 235901
rect 411760 235889 411766 235901
rect 401258 235861 411766 235889
rect 401258 235849 401264 235861
rect 411760 235849 411766 235861
rect 411818 235849 411824 235901
rect 386762 235787 393086 235815
rect 386762 235775 386768 235787
rect 393136 235775 393142 235827
rect 393194 235815 393200 235827
rect 406096 235815 406102 235827
rect 393194 235787 406102 235815
rect 393194 235775 393200 235787
rect 406096 235775 406102 235787
rect 406154 235775 406160 235827
rect 410896 235775 410902 235827
rect 410954 235815 410960 235827
rect 413008 235815 413014 235827
rect 410954 235787 413014 235815
rect 410954 235775 410960 235787
rect 413008 235775 413014 235787
rect 413066 235775 413072 235827
rect 364106 235713 371774 235741
rect 364106 235701 364112 235713
rect 378832 235701 378838 235753
rect 378890 235741 378896 235753
rect 392848 235741 392854 235753
rect 378890 235713 392854 235741
rect 378890 235701 378896 235713
rect 392848 235701 392854 235713
rect 392906 235701 392912 235753
rect 392944 235701 392950 235753
rect 393002 235741 393008 235753
rect 398416 235741 398422 235753
rect 393002 235713 398422 235741
rect 393002 235701 393008 235713
rect 398416 235701 398422 235713
rect 398474 235701 398480 235753
rect 398608 235701 398614 235753
rect 398666 235741 398672 235753
rect 528400 235741 528406 235753
rect 398666 235713 528406 235741
rect 398666 235701 398672 235713
rect 528400 235701 528406 235713
rect 528458 235701 528464 235753
rect 210640 235627 210646 235679
rect 210698 235667 210704 235679
rect 230032 235667 230038 235679
rect 210698 235639 230038 235667
rect 210698 235627 210704 235639
rect 230032 235627 230038 235639
rect 230090 235627 230096 235679
rect 285136 235627 285142 235679
rect 285194 235667 285200 235679
rect 323344 235667 323350 235679
rect 285194 235639 323350 235667
rect 285194 235627 285200 235639
rect 323344 235627 323350 235639
rect 323402 235627 323408 235679
rect 326224 235627 326230 235679
rect 326282 235667 326288 235679
rect 460240 235667 460246 235679
rect 326282 235639 460246 235667
rect 326282 235627 326288 235639
rect 460240 235627 460246 235639
rect 460298 235627 460304 235679
rect 210064 235553 210070 235605
rect 210122 235593 210128 235605
rect 227824 235593 227830 235605
rect 210122 235565 227830 235593
rect 210122 235553 210128 235565
rect 227824 235553 227830 235565
rect 227882 235553 227888 235605
rect 236464 235553 236470 235605
rect 236522 235593 236528 235605
rect 282928 235593 282934 235605
rect 236522 235565 282934 235593
rect 236522 235553 236528 235565
rect 282928 235553 282934 235565
rect 282986 235553 282992 235605
rect 286672 235553 286678 235605
rect 286730 235593 286736 235605
rect 326800 235593 326806 235605
rect 286730 235565 326806 235593
rect 286730 235553 286736 235565
rect 326800 235553 326806 235565
rect 326858 235553 326864 235605
rect 332560 235553 332566 235605
rect 332618 235593 332624 235605
rect 472336 235593 472342 235605
rect 332618 235565 472342 235593
rect 332618 235553 332624 235565
rect 472336 235553 472342 235565
rect 472394 235553 472400 235605
rect 212944 235479 212950 235531
rect 213002 235519 213008 235531
rect 232336 235519 232342 235531
rect 213002 235491 232342 235519
rect 213002 235479 213008 235491
rect 232336 235479 232342 235491
rect 232394 235479 232400 235531
rect 238000 235479 238006 235531
rect 238058 235519 238064 235531
rect 285904 235519 285910 235531
rect 238058 235491 285910 235519
rect 238058 235479 238064 235491
rect 285904 235479 285910 235491
rect 285962 235479 285968 235531
rect 290320 235479 290326 235531
rect 290378 235519 290384 235531
rect 334288 235519 334294 235531
rect 290378 235491 334294 235519
rect 290378 235479 290384 235491
rect 334288 235479 334294 235491
rect 334346 235479 334352 235531
rect 348880 235479 348886 235531
rect 348938 235519 348944 235531
rect 397360 235519 397366 235531
rect 348938 235491 397366 235519
rect 348938 235479 348944 235491
rect 397360 235479 397366 235491
rect 397418 235479 397424 235531
rect 588976 235519 588982 235531
rect 402898 235491 588982 235519
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 42832 235445 42838 235457
rect 42218 235417 42838 235445
rect 42218 235405 42224 235417
rect 42832 235405 42838 235417
rect 42890 235405 42896 235457
rect 211984 235405 211990 235457
rect 212042 235445 212048 235457
rect 233008 235445 233014 235457
rect 212042 235417 233014 235445
rect 212042 235405 212048 235417
rect 233008 235405 233014 235417
rect 233066 235405 233072 235457
rect 242128 235405 242134 235457
rect 242186 235445 242192 235457
rect 293392 235445 293398 235457
rect 242186 235417 293398 235445
rect 242186 235405 242192 235417
rect 293392 235405 293398 235417
rect 293450 235405 293456 235457
rect 295216 235405 295222 235457
rect 295274 235445 295280 235457
rect 348688 235445 348694 235457
rect 295274 235417 348694 235445
rect 295274 235405 295280 235417
rect 348688 235405 348694 235417
rect 348746 235405 348752 235457
rect 392848 235405 392854 235457
rect 392906 235445 392912 235457
rect 396688 235445 396694 235457
rect 392906 235417 396694 235445
rect 392906 235405 392912 235417
rect 396688 235405 396694 235417
rect 396746 235405 396752 235457
rect 396784 235405 396790 235457
rect 396842 235445 396848 235457
rect 402898 235445 402926 235491
rect 588976 235479 588982 235491
rect 589034 235479 589040 235531
rect 396842 235417 402926 235445
rect 396842 235405 396848 235417
rect 403024 235405 403030 235457
rect 403082 235445 403088 235457
rect 588688 235445 588694 235457
rect 403082 235417 588694 235445
rect 403082 235405 403088 235417
rect 588688 235405 588694 235417
rect 588746 235405 588752 235457
rect 206992 235331 206998 235383
rect 207050 235371 207056 235383
rect 221776 235371 221782 235383
rect 207050 235343 221782 235371
rect 207050 235331 207056 235343
rect 221776 235331 221782 235343
rect 221834 235331 221840 235383
rect 223888 235331 223894 235383
rect 223946 235371 223952 235383
rect 244720 235371 244726 235383
rect 223946 235343 244726 235371
rect 223946 235331 223952 235343
rect 244720 235331 244726 235343
rect 244778 235331 244784 235383
rect 254224 235331 254230 235383
rect 254282 235371 254288 235383
rect 306736 235371 306742 235383
rect 254282 235343 306742 235371
rect 254282 235331 254288 235343
rect 306736 235331 306742 235343
rect 306794 235331 306800 235383
rect 339472 235331 339478 235383
rect 339530 235371 339536 235383
rect 395248 235371 395254 235383
rect 339530 235343 395254 235371
rect 339530 235331 339536 235343
rect 395248 235331 395254 235343
rect 395306 235331 395312 235383
rect 398512 235331 398518 235383
rect 398570 235371 398576 235383
rect 590416 235371 590422 235383
rect 398570 235343 590422 235371
rect 398570 235331 398576 235343
rect 590416 235331 590422 235343
rect 590474 235331 590480 235383
rect 214192 235257 214198 235309
rect 214250 235297 214256 235309
rect 235312 235297 235318 235309
rect 214250 235269 235318 235297
rect 214250 235257 214256 235269
rect 235312 235257 235318 235269
rect 235370 235257 235376 235309
rect 239344 235257 239350 235309
rect 239402 235297 239408 235309
rect 287344 235297 287350 235309
rect 239402 235269 287350 235297
rect 239402 235257 239408 235269
rect 287344 235257 287350 235269
rect 287402 235257 287408 235309
rect 288880 235257 288886 235309
rect 288938 235297 288944 235309
rect 345712 235297 345718 235309
rect 288938 235269 345718 235297
rect 288938 235257 288944 235269
rect 345712 235257 345718 235269
rect 345770 235257 345776 235309
rect 396304 235257 396310 235309
rect 396362 235297 396368 235309
rect 588880 235297 588886 235309
rect 396362 235269 588886 235297
rect 396362 235257 396368 235269
rect 588880 235257 588886 235269
rect 588938 235257 588944 235309
rect 220624 235183 220630 235235
rect 220682 235223 220688 235235
rect 241840 235223 241846 235235
rect 220682 235195 241846 235223
rect 220682 235183 220688 235195
rect 241840 235183 241846 235195
rect 241898 235183 241904 235235
rect 249712 235183 249718 235235
rect 249770 235223 249776 235235
rect 302320 235223 302326 235235
rect 249770 235195 302326 235223
rect 249770 235183 249776 235195
rect 302320 235183 302326 235195
rect 302378 235183 302384 235235
rect 305200 235183 305206 235235
rect 305258 235223 305264 235235
rect 365680 235223 365686 235235
rect 305258 235195 365686 235223
rect 305258 235183 305264 235195
rect 365680 235183 365686 235195
rect 365738 235183 365744 235235
rect 374512 235183 374518 235235
rect 374570 235223 374576 235235
rect 381616 235223 381622 235235
rect 374570 235195 381622 235223
rect 374570 235183 374576 235195
rect 381616 235183 381622 235195
rect 381674 235183 381680 235235
rect 394960 235183 394966 235235
rect 395018 235223 395024 235235
rect 403024 235223 403030 235235
rect 395018 235195 403030 235223
rect 395018 235183 395024 235195
rect 403024 235183 403030 235195
rect 403082 235183 403088 235235
rect 403120 235183 403126 235235
rect 403178 235223 403184 235235
rect 587920 235223 587926 235235
rect 403178 235195 587926 235223
rect 403178 235183 403184 235195
rect 587920 235183 587926 235195
rect 587978 235183 587984 235235
rect 206128 235109 206134 235161
rect 206186 235149 206192 235161
rect 215920 235149 215926 235161
rect 206186 235121 215926 235149
rect 206186 235109 206192 235121
rect 215920 235109 215926 235121
rect 215978 235109 215984 235161
rect 232912 235109 232918 235161
rect 232970 235149 232976 235161
rect 262000 235149 262006 235161
rect 232970 235121 262006 235149
rect 232970 235109 232976 235121
rect 262000 235109 262006 235121
rect 262058 235109 262064 235161
rect 266128 235109 266134 235161
rect 266186 235149 266192 235161
rect 324496 235149 324502 235161
rect 266186 235121 324502 235149
rect 266186 235109 266192 235121
rect 324496 235109 324502 235121
rect 324554 235109 324560 235161
rect 327664 235109 327670 235161
rect 327722 235149 327728 235161
rect 390352 235149 390358 235161
rect 327722 235121 390358 235149
rect 327722 235109 327728 235121
rect 390352 235109 390358 235121
rect 390410 235109 390416 235161
rect 392176 235109 392182 235161
rect 392234 235149 392240 235161
rect 592336 235149 592342 235161
rect 392234 235121 592342 235149
rect 392234 235109 392240 235121
rect 592336 235109 592342 235121
rect 592394 235109 592400 235161
rect 203248 235035 203254 235087
rect 203306 235075 203312 235087
rect 211504 235075 211510 235087
rect 203306 235047 211510 235075
rect 203306 235035 203312 235047
rect 211504 235035 211510 235047
rect 211562 235035 211568 235087
rect 213424 235035 213430 235087
rect 213482 235075 213488 235087
rect 233392 235075 233398 235087
rect 213482 235047 233398 235075
rect 213482 235035 213488 235047
rect 233392 235035 233398 235047
rect 233450 235035 233456 235087
rect 235696 235035 235702 235087
rect 235754 235075 235760 235087
rect 265264 235075 265270 235087
rect 235754 235047 265270 235075
rect 235754 235035 235760 235047
rect 265264 235035 265270 235047
rect 265322 235035 265328 235087
rect 268912 235035 268918 235087
rect 268970 235075 268976 235087
rect 331408 235075 331414 235087
rect 268970 235047 331414 235075
rect 268970 235035 268976 235047
rect 331408 235035 331414 235047
rect 331466 235035 331472 235087
rect 334960 235035 334966 235087
rect 335018 235075 335024 235087
rect 393520 235075 393526 235087
rect 335018 235047 393526 235075
rect 335018 235035 335024 235047
rect 393520 235035 393526 235047
rect 393578 235035 393584 235087
rect 394576 235035 394582 235087
rect 394634 235075 394640 235087
rect 597712 235075 597718 235087
rect 394634 235047 597718 235075
rect 394634 235035 394640 235047
rect 597712 235035 597718 235047
rect 597770 235035 597776 235087
rect 208816 234961 208822 235013
rect 208874 235001 208880 235013
rect 224752 235001 224758 235013
rect 208874 234973 224758 235001
rect 208874 234961 208880 234973
rect 224752 234961 224758 234973
rect 224810 234961 224816 235013
rect 225520 234961 225526 235013
rect 225578 235001 225584 235013
rect 260176 235001 260182 235013
rect 225578 234973 260182 235001
rect 225578 234961 225584 234973
rect 260176 234961 260182 234973
rect 260234 234961 260240 235013
rect 260272 234961 260278 235013
rect 260330 235001 260336 235013
rect 323248 235001 323254 235013
rect 260330 234973 323254 235001
rect 260330 234961 260336 234973
rect 323248 234961 323254 234973
rect 323306 234961 323312 235013
rect 333424 234961 333430 235013
rect 333482 235001 333488 235013
rect 333482 234973 378734 235001
rect 333482 234961 333488 234973
rect 211024 234887 211030 234939
rect 211082 234927 211088 234939
rect 231568 234927 231574 234939
rect 211082 234899 231574 234927
rect 211082 234887 211088 234899
rect 231568 234887 231574 234899
rect 231626 234887 231632 234939
rect 243856 234887 243862 234939
rect 243914 234927 243920 234939
rect 296464 234927 296470 234939
rect 243914 234899 296470 234927
rect 243914 234887 243920 234899
rect 296464 234887 296470 234899
rect 296522 234887 296528 234939
rect 296560 234887 296566 234939
rect 296618 234927 296624 234939
rect 361936 234927 361942 234939
rect 296618 234899 361942 234927
rect 296618 234887 296624 234899
rect 361936 234887 361942 234899
rect 361994 234887 362000 234939
rect 209296 234813 209302 234865
rect 209354 234853 209360 234865
rect 228496 234853 228502 234865
rect 209354 234825 228502 234853
rect 209354 234813 209360 234825
rect 228496 234813 228502 234825
rect 228554 234813 228560 234865
rect 229744 234813 229750 234865
rect 229802 234853 229808 234865
rect 253552 234853 253558 234865
rect 229802 234825 253558 234853
rect 229802 234813 229808 234825
rect 253552 234813 253558 234825
rect 253610 234813 253616 234865
rect 257488 234813 257494 234865
rect 257546 234853 257552 234865
rect 308176 234853 308182 234865
rect 257546 234825 308182 234853
rect 257546 234813 257552 234825
rect 308176 234813 308182 234825
rect 308234 234813 308240 234865
rect 321616 234813 321622 234865
rect 321674 234853 321680 234865
rect 378544 234853 378550 234865
rect 321674 234825 378550 234853
rect 321674 234813 321680 234825
rect 378544 234813 378550 234825
rect 378602 234813 378608 234865
rect 378706 234853 378734 234973
rect 389872 234961 389878 235013
rect 389930 235001 389936 235013
rect 403120 235001 403126 235013
rect 389930 234973 403126 235001
rect 389930 234961 389936 234973
rect 403120 234961 403126 234973
rect 403178 234961 403184 235013
rect 403600 234961 403606 235013
rect 403658 235001 403664 235013
rect 615856 235001 615862 235013
rect 403658 234973 615862 235001
rect 403658 234961 403664 234973
rect 615856 234961 615862 234973
rect 615914 234961 615920 235013
rect 381616 234887 381622 234939
rect 381674 234927 381680 234939
rect 398800 234927 398806 234939
rect 381674 234899 398806 234927
rect 381674 234887 381680 234899
rect 398800 234887 398806 234899
rect 398858 234887 398864 234939
rect 406672 234887 406678 234939
rect 406730 234927 406736 234939
rect 621808 234927 621814 234939
rect 406730 234899 621814 234927
rect 406730 234887 406736 234899
rect 621808 234887 621814 234899
rect 621866 234887 621872 234939
rect 395728 234853 395734 234865
rect 378706 234825 395734 234853
rect 395728 234813 395734 234825
rect 395786 234813 395792 234865
rect 398224 234813 398230 234865
rect 398282 234853 398288 234865
rect 405040 234853 405046 234865
rect 398282 234825 405046 234853
rect 398282 234813 398288 234825
rect 405040 234813 405046 234825
rect 405098 234813 405104 234865
rect 407920 234813 407926 234865
rect 407978 234853 407984 234865
rect 408784 234853 408790 234865
rect 407978 234825 408790 234853
rect 407978 234813 407984 234825
rect 408784 234813 408790 234825
rect 408842 234813 408848 234865
rect 409936 234813 409942 234865
rect 409994 234853 410000 234865
rect 627856 234853 627862 234865
rect 409994 234825 627862 234853
rect 409994 234813 410000 234825
rect 627856 234813 627862 234825
rect 627914 234813 627920 234865
rect 202864 234739 202870 234791
rect 202922 234779 202928 234791
rect 214768 234779 214774 234791
rect 202922 234751 214774 234779
rect 202922 234739 202928 234751
rect 214768 234739 214774 234751
rect 214826 234739 214832 234791
rect 225136 234739 225142 234791
rect 225194 234779 225200 234791
rect 247696 234779 247702 234791
rect 225194 234751 247702 234779
rect 225194 234739 225200 234751
rect 247696 234739 247702 234751
rect 247754 234739 247760 234791
rect 251152 234739 251158 234791
rect 251210 234779 251216 234791
rect 304144 234779 304150 234791
rect 251210 234751 304150 234779
rect 251210 234739 251216 234751
rect 304144 234739 304150 234751
rect 304202 234739 304208 234791
rect 315280 234739 315286 234791
rect 315338 234779 315344 234791
rect 396400 234779 396406 234791
rect 315338 234751 396406 234779
rect 315338 234739 315344 234751
rect 396400 234739 396406 234751
rect 396458 234739 396464 234791
rect 396496 234739 396502 234791
rect 396554 234779 396560 234791
rect 406864 234779 406870 234791
rect 396554 234751 406870 234779
rect 396554 234739 396560 234751
rect 406864 234739 406870 234751
rect 406922 234739 406928 234791
rect 412144 234739 412150 234791
rect 412202 234779 412208 234791
rect 632368 234779 632374 234791
rect 412202 234751 632374 234779
rect 412202 234739 412208 234751
rect 632368 234739 632374 234751
rect 632426 234739 632432 234791
rect 204784 234665 204790 234717
rect 204842 234705 204848 234717
rect 214864 234705 214870 234717
rect 204842 234677 214870 234705
rect 204842 234665 204848 234677
rect 214864 234665 214870 234677
rect 214922 234665 214928 234717
rect 222352 234665 222358 234717
rect 222410 234705 222416 234717
rect 243952 234705 243958 234717
rect 222410 234677 243958 234705
rect 222410 234665 222416 234677
rect 243952 234665 243958 234677
rect 244010 234665 244016 234717
rect 246640 234665 246646 234717
rect 246698 234705 246704 234717
rect 299344 234705 299350 234717
rect 246698 234677 299350 234705
rect 246698 234665 246704 234677
rect 299344 234665 299350 234677
rect 299402 234665 299408 234717
rect 301744 234665 301750 234717
rect 301802 234705 301808 234717
rect 398896 234705 398902 234717
rect 301802 234677 398902 234705
rect 301802 234665 301808 234677
rect 398896 234665 398902 234677
rect 398954 234665 398960 234717
rect 411280 234665 411286 234717
rect 411338 234705 411344 234717
rect 630928 234705 630934 234717
rect 411338 234677 630934 234705
rect 411338 234665 411344 234677
rect 630928 234665 630934 234677
rect 630986 234665 630992 234717
rect 42160 234591 42166 234643
rect 42218 234631 42224 234643
rect 42736 234631 42742 234643
rect 42218 234603 42742 234631
rect 42218 234591 42224 234603
rect 42736 234591 42742 234603
rect 42794 234591 42800 234643
rect 202000 234591 202006 234643
rect 202058 234631 202064 234643
rect 213424 234631 213430 234643
rect 202058 234603 213430 234631
rect 202058 234591 202064 234603
rect 213424 234591 213430 234603
rect 213482 234591 213488 234643
rect 251056 234591 251062 234643
rect 251114 234631 251120 234643
rect 273616 234631 273622 234643
rect 251114 234603 273622 234631
rect 251114 234591 251120 234603
rect 273616 234591 273622 234603
rect 273674 234591 273680 234643
rect 280624 234591 280630 234643
rect 280682 234631 280688 234643
rect 321040 234631 321046 234643
rect 280682 234603 321046 234631
rect 280682 234591 280688 234603
rect 321040 234591 321046 234603
rect 321098 234591 321104 234643
rect 323536 234591 323542 234643
rect 323594 234631 323600 234643
rect 434896 234631 434902 234643
rect 323594 234603 434902 234631
rect 323594 234591 323600 234603
rect 434896 234591 434902 234603
rect 434954 234591 434960 234643
rect 204208 234517 204214 234569
rect 204266 234557 204272 234569
rect 215536 234557 215542 234569
rect 204266 234529 215542 234557
rect 204266 234517 204272 234529
rect 215536 234517 215542 234529
rect 215594 234517 215600 234569
rect 237040 234517 237046 234569
rect 237098 234557 237104 234569
rect 258064 234557 258070 234569
rect 237098 234529 258070 234557
rect 237098 234517 237104 234529
rect 258064 234517 258070 234529
rect 258122 234517 258128 234569
rect 262480 234517 262486 234569
rect 262538 234557 262544 234569
rect 290896 234557 290902 234569
rect 262538 234529 290902 234557
rect 262538 234517 262544 234529
rect 290896 234517 290902 234529
rect 290954 234517 290960 234569
rect 295696 234517 295702 234569
rect 295754 234557 295760 234569
rect 341392 234557 341398 234569
rect 295754 234529 341398 234557
rect 295754 234517 295760 234529
rect 341392 234517 341398 234529
rect 341450 234517 341456 234569
rect 345904 234517 345910 234569
rect 345962 234557 345968 234569
rect 400336 234557 400342 234569
rect 345962 234529 400342 234557
rect 345962 234517 345968 234529
rect 400336 234517 400342 234529
rect 400394 234517 400400 234569
rect 410800 234517 410806 234569
rect 410858 234557 410864 234569
rect 522640 234557 522646 234569
rect 410858 234529 522646 234557
rect 410858 234517 410864 234529
rect 522640 234517 522646 234529
rect 522698 234517 522704 234569
rect 206512 234443 206518 234495
rect 206570 234483 206576 234495
rect 206570 234455 212126 234483
rect 206570 234443 206576 234455
rect 204400 234369 204406 234421
rect 204458 234409 204464 234421
rect 210160 234409 210166 234421
rect 204458 234381 210166 234409
rect 204458 234369 204464 234381
rect 210160 234369 210166 234381
rect 210218 234369 210224 234421
rect 201520 234295 201526 234347
rect 201578 234335 201584 234347
rect 211888 234335 211894 234347
rect 201578 234307 211894 234335
rect 201578 234295 201584 234307
rect 211888 234295 211894 234307
rect 211946 234295 211952 234347
rect 212098 234335 212126 234455
rect 250480 234443 250486 234495
rect 250538 234483 250544 234495
rect 269392 234483 269398 234495
rect 250538 234455 269398 234483
rect 250538 234443 250544 234455
rect 269392 234443 269398 234455
rect 269450 234443 269456 234495
rect 271600 234443 271606 234495
rect 271658 234483 271664 234495
rect 301264 234483 301270 234495
rect 271658 234455 301270 234483
rect 271658 234443 271664 234455
rect 301264 234443 301270 234455
rect 301322 234443 301328 234495
rect 306256 234443 306262 234495
rect 306314 234483 306320 234495
rect 358384 234483 358390 234495
rect 306314 234455 358390 234483
rect 306314 234443 306320 234455
rect 358384 234443 358390 234455
rect 358442 234443 358448 234495
rect 383632 234443 383638 234495
rect 383690 234483 383696 234495
rect 396496 234483 396502 234495
rect 383690 234455 396502 234483
rect 383690 234443 383696 234455
rect 396496 234443 396502 234455
rect 396554 234443 396560 234495
rect 396592 234443 396598 234495
rect 396650 234483 396656 234495
rect 408016 234483 408022 234495
rect 396650 234455 408022 234483
rect 396650 234443 396656 234455
rect 408016 234443 408022 234455
rect 408074 234443 408080 234495
rect 409264 234443 409270 234495
rect 409322 234483 409328 234495
rect 521200 234483 521206 234495
rect 409322 234455 521206 234483
rect 409322 234443 409328 234455
rect 521200 234443 521206 234455
rect 521258 234443 521264 234495
rect 215920 234369 215926 234421
rect 215978 234409 215984 234421
rect 221008 234409 221014 234421
rect 215978 234381 221014 234409
rect 215978 234369 215984 234381
rect 221008 234369 221014 234381
rect 221066 234369 221072 234421
rect 235600 234369 235606 234421
rect 235658 234409 235664 234421
rect 250576 234409 250582 234421
rect 235658 234381 250582 234409
rect 235658 234369 235664 234381
rect 250576 234369 250582 234381
rect 250634 234369 250640 234421
rect 255280 234369 255286 234421
rect 255338 234409 255344 234421
rect 277072 234409 277078 234421
rect 255338 234381 277078 234409
rect 255338 234369 255344 234381
rect 277072 234369 277078 234381
rect 277130 234369 277136 234421
rect 283984 234369 283990 234421
rect 284042 234409 284048 234421
rect 311344 234409 311350 234421
rect 284042 234381 311350 234409
rect 284042 234369 284048 234381
rect 311344 234369 311350 234381
rect 311402 234369 311408 234421
rect 314416 234369 314422 234421
rect 314474 234409 314480 234421
rect 423376 234409 423382 234421
rect 314474 234381 423382 234409
rect 314474 234369 314480 234381
rect 423376 234369 423382 234381
rect 423434 234369 423440 234421
rect 222448 234335 222454 234347
rect 212098 234307 222454 234335
rect 222448 234295 222454 234307
rect 222506 234295 222512 234347
rect 239824 234295 239830 234347
rect 239882 234335 239888 234347
rect 260464 234335 260470 234347
rect 239882 234307 260470 234335
rect 239882 234295 239888 234307
rect 260464 234295 260470 234307
rect 260522 234295 260528 234347
rect 261232 234295 261238 234347
rect 261290 234335 261296 234347
rect 288016 234335 288022 234347
rect 261290 234307 288022 234335
rect 261290 234295 261296 234307
rect 288016 234295 288022 234307
rect 288074 234295 288080 234347
rect 308464 234295 308470 234347
rect 308522 234335 308528 234347
rect 416368 234335 416374 234347
rect 308522 234307 416374 234335
rect 308522 234295 308528 234307
rect 416368 234295 416374 234307
rect 416426 234295 416432 234347
rect 207856 234221 207862 234273
rect 207914 234261 207920 234273
rect 207914 234233 214814 234261
rect 207914 234221 207920 234233
rect 200272 234147 200278 234199
rect 200330 234187 200336 234199
rect 210352 234187 210358 234199
rect 200330 234159 210358 234187
rect 200330 234147 200336 234159
rect 210352 234147 210358 234159
rect 210410 234147 210416 234199
rect 214786 234187 214814 234233
rect 214864 234221 214870 234273
rect 214922 234261 214928 234273
rect 219376 234261 219382 234273
rect 214922 234233 219382 234261
rect 214922 234221 214928 234233
rect 219376 234221 219382 234233
rect 219434 234221 219440 234273
rect 244336 234221 244342 234273
rect 244394 234261 244400 234273
rect 264880 234261 264886 234273
rect 244394 234233 264886 234261
rect 244394 234221 244400 234233
rect 264880 234221 264886 234233
rect 264938 234221 264944 234273
rect 268528 234221 268534 234273
rect 268586 234261 268592 234273
rect 293776 234261 293782 234273
rect 268586 234233 293782 234261
rect 268586 234221 268592 234233
rect 293776 234221 293782 234233
rect 293834 234221 293840 234273
rect 312688 234221 312694 234273
rect 312746 234261 312752 234273
rect 418288 234261 418294 234273
rect 312746 234233 418294 234261
rect 312746 234221 312752 234233
rect 418288 234221 418294 234233
rect 418346 234221 418352 234273
rect 225520 234187 225526 234199
rect 214786 234159 225526 234187
rect 225520 234147 225526 234159
rect 225578 234147 225584 234199
rect 256528 234147 256534 234199
rect 256586 234187 256592 234199
rect 279280 234187 279286 234199
rect 256586 234159 279286 234187
rect 256586 234147 256592 234159
rect 279280 234147 279286 234159
rect 279338 234147 279344 234199
rect 283888 234147 283894 234199
rect 283946 234187 283952 234199
rect 320752 234187 320758 234199
rect 283946 234159 320758 234187
rect 283946 234147 283952 234159
rect 320752 234147 320758 234159
rect 320810 234147 320816 234199
rect 330448 234147 330454 234199
rect 330506 234187 330512 234199
rect 374704 234187 374710 234199
rect 330506 234159 374710 234187
rect 330506 234147 330512 234159
rect 374704 234147 374710 234159
rect 374762 234147 374768 234199
rect 378544 234147 378550 234199
rect 378602 234187 378608 234199
rect 385936 234187 385942 234199
rect 378602 234159 385942 234187
rect 378602 234147 378608 234159
rect 385936 234147 385942 234159
rect 385994 234147 386000 234199
rect 395824 234147 395830 234199
rect 395882 234187 395888 234199
rect 403120 234187 403126 234199
rect 395882 234159 403126 234187
rect 395882 234147 395888 234159
rect 403120 234147 403126 234159
rect 403178 234147 403184 234199
rect 403216 234147 403222 234199
rect 403274 234187 403280 234199
rect 498544 234187 498550 234199
rect 403274 234159 498550 234187
rect 403274 234147 403280 234159
rect 498544 234147 498550 234159
rect 498602 234147 498608 234199
rect 200176 234073 200182 234125
rect 200234 234113 200240 234125
rect 208816 234113 208822 234125
rect 200234 234085 208822 234113
rect 200234 234073 200240 234085
rect 208816 234073 208822 234085
rect 208874 234073 208880 234125
rect 210160 234073 210166 234125
rect 210218 234113 210224 234125
rect 217936 234113 217942 234125
rect 210218 234085 217942 234113
rect 210218 234073 210224 234085
rect 217936 234073 217942 234085
rect 217994 234073 218000 234125
rect 247408 234073 247414 234125
rect 247466 234113 247472 234125
rect 266320 234113 266326 234125
rect 247466 234085 266326 234113
rect 247466 234073 247472 234085
rect 266320 234073 266326 234085
rect 266378 234073 266384 234125
rect 267088 234073 267094 234125
rect 267146 234113 267152 234125
rect 290992 234113 290998 234125
rect 267146 234085 290998 234113
rect 267146 234073 267152 234085
rect 290992 234073 290998 234085
rect 291050 234073 291056 234125
rect 294832 234073 294838 234125
rect 294890 234113 294896 234125
rect 339088 234113 339094 234125
rect 294890 234085 339094 234113
rect 294890 234073 294896 234085
rect 339088 234073 339094 234085
rect 339146 234073 339152 234125
rect 358000 234073 358006 234125
rect 358058 234113 358064 234125
rect 394864 234113 394870 234125
rect 358058 234085 394870 234113
rect 358058 234073 358064 234085
rect 394864 234073 394870 234085
rect 394922 234073 394928 234125
rect 401776 234073 401782 234125
rect 401834 234113 401840 234125
rect 486640 234113 486646 234125
rect 401834 234085 486646 234113
rect 401834 234073 401840 234085
rect 486640 234073 486646 234085
rect 486698 234073 486704 234125
rect 42064 233999 42070 234051
rect 42122 234039 42128 234051
rect 42928 234039 42934 234051
rect 42122 234011 42934 234039
rect 42122 233999 42128 234011
rect 42928 233999 42934 234011
rect 42986 233999 42992 234051
rect 198736 233999 198742 234051
rect 198794 234039 198800 234051
rect 207376 234039 207382 234051
rect 198794 234011 207382 234039
rect 198794 233999 198800 234011
rect 207376 233999 207382 234011
rect 207434 233999 207440 234051
rect 220240 234039 220246 234051
rect 211426 234011 220246 234039
rect 198352 233925 198358 233977
rect 198410 233965 198416 233977
rect 205936 233965 205942 233977
rect 198410 233937 205942 233965
rect 198410 233925 198416 233937
rect 205936 233925 205942 233937
rect 205994 233925 206000 233977
rect 206896 233925 206902 233977
rect 206954 233965 206960 233977
rect 211426 233965 211454 234011
rect 220240 233999 220246 234011
rect 220298 233999 220304 234051
rect 259792 233999 259798 234051
rect 259850 234039 259856 234051
rect 281872 234039 281878 234051
rect 259850 234011 281878 234039
rect 259850 233999 259856 234011
rect 281872 233999 281878 234011
rect 281930 233999 281936 234051
rect 299824 233999 299830 234051
rect 299882 234039 299888 234051
rect 344656 234039 344662 234051
rect 299882 234011 344662 234039
rect 299882 233999 299888 234011
rect 344656 233999 344662 234011
rect 344714 233999 344720 234051
rect 365872 233999 365878 234051
rect 365930 234039 365936 234051
rect 382768 234039 382774 234051
rect 365930 234011 382774 234039
rect 365930 233999 365936 234011
rect 382768 233999 382774 234011
rect 382826 233999 382832 234051
rect 399088 233999 399094 234051
rect 399146 234039 399152 234051
rect 400144 234039 400150 234051
rect 399146 234011 400150 234039
rect 399146 233999 399152 234011
rect 400144 233999 400150 234011
rect 400202 233999 400208 234051
rect 400240 233999 400246 234051
rect 400298 234039 400304 234051
rect 400298 234011 407966 234039
rect 400298 233999 400304 234011
rect 206954 233937 211454 233965
rect 206954 233925 206960 233937
rect 211504 233925 211510 233977
rect 211562 233965 211568 233977
rect 216496 233965 216502 233977
rect 211562 233937 216502 233965
rect 211562 233925 211568 233937
rect 216496 233925 216502 233937
rect 216554 233925 216560 233977
rect 296080 233925 296086 233977
rect 296138 233965 296144 233977
rect 339760 233965 339766 233977
rect 296138 233937 339766 233965
rect 296138 233925 296144 233937
rect 339760 233925 339766 233937
rect 339818 233925 339824 233977
rect 341200 233925 341206 233977
rect 341258 233965 341264 233977
rect 378448 233965 378454 233977
rect 341258 233937 378454 233965
rect 341258 233925 341264 233937
rect 378448 233925 378454 233937
rect 378506 233925 378512 233977
rect 382096 233925 382102 233977
rect 382154 233965 382160 233977
rect 400720 233965 400726 233977
rect 382154 233937 400726 233965
rect 382154 233925 382160 233937
rect 400720 233925 400726 233937
rect 400778 233925 400784 233977
rect 407938 233965 407966 234011
rect 408016 233999 408022 234051
rect 408074 234039 408080 234051
rect 475216 234039 475222 234051
rect 408074 234011 475222 234039
rect 408074 233999 408080 234011
rect 475216 233999 475222 234011
rect 475274 233999 475280 234051
rect 479248 233965 479254 233977
rect 407938 233937 479254 233965
rect 479248 233925 479254 233937
rect 479306 233925 479312 233977
rect 197488 233851 197494 233903
rect 197546 233891 197552 233903
rect 204304 233891 204310 233903
rect 197546 233863 204310 233891
rect 197546 233851 197552 233863
rect 204304 233851 204310 233863
rect 204362 233851 204368 233903
rect 214480 233891 214486 233903
rect 211522 233863 214486 233891
rect 196912 233777 196918 233829
rect 196970 233817 196976 233829
rect 202864 233817 202870 233829
rect 196970 233789 202870 233817
rect 196970 233777 196976 233789
rect 202864 233777 202870 233789
rect 202922 233777 202928 233829
rect 205168 233777 205174 233829
rect 205226 233817 205232 233829
rect 211522 233817 211550 233863
rect 214480 233851 214486 233863
rect 214538 233851 214544 233903
rect 253456 233851 253462 233903
rect 253514 233891 253520 233903
rect 270832 233891 270838 233903
rect 253514 233863 270838 233891
rect 253514 233851 253520 233863
rect 270832 233851 270838 233863
rect 270890 233851 270896 233903
rect 294448 233851 294454 233903
rect 294506 233891 294512 233903
rect 331216 233891 331222 233903
rect 294506 233863 331222 233891
rect 294506 233851 294512 233863
rect 331216 233851 331222 233863
rect 331274 233851 331280 233903
rect 339856 233851 339862 233903
rect 339914 233891 339920 233903
rect 351376 233891 351382 233903
rect 339914 233863 351382 233891
rect 339914 233851 339920 233863
rect 351376 233851 351382 233863
rect 351434 233851 351440 233903
rect 361264 233851 361270 233903
rect 361322 233891 361328 233903
rect 432016 233891 432022 233903
rect 361322 233863 392510 233891
rect 361322 233851 361328 233863
rect 205226 233789 211550 233817
rect 205226 233777 205232 233789
rect 211600 233777 211606 233829
rect 211658 233817 211664 233829
rect 230704 233817 230710 233829
rect 211658 233789 230710 233817
rect 211658 233777 211664 233789
rect 230704 233777 230710 233789
rect 230762 233777 230768 233829
rect 242896 233777 242902 233829
rect 242954 233817 242960 233829
rect 260848 233817 260854 233829
rect 242954 233789 260854 233817
rect 242954 233777 242960 233789
rect 260848 233777 260854 233789
rect 260906 233777 260912 233829
rect 267472 233777 267478 233829
rect 267530 233817 267536 233829
rect 285040 233817 285046 233829
rect 267530 233789 285046 233817
rect 267530 233777 267536 233789
rect 285040 233777 285046 233789
rect 285098 233777 285104 233829
rect 297232 233777 297238 233829
rect 297290 233817 297296 233829
rect 328336 233817 328342 233829
rect 297290 233789 328342 233817
rect 297290 233777 297296 233789
rect 328336 233777 328342 233789
rect 328394 233777 328400 233829
rect 332176 233777 332182 233829
rect 332234 233817 332240 233829
rect 383056 233817 383062 233829
rect 332234 233789 383062 233817
rect 332234 233777 332240 233789
rect 383056 233777 383062 233789
rect 383114 233777 383120 233829
rect 392482 233817 392510 233863
rect 400642 233863 432022 233891
rect 400642 233817 400670 233863
rect 432016 233851 432022 233863
rect 432074 233851 432080 233903
rect 392482 233789 400670 233817
rect 400720 233777 400726 233829
rect 400778 233817 400784 233829
rect 411760 233817 411766 233829
rect 400778 233789 411766 233817
rect 400778 233777 400784 233789
rect 411760 233777 411766 233789
rect 411818 233777 411824 233829
rect 197968 233703 197974 233755
rect 198026 233743 198032 233755
rect 203632 233743 203638 233755
rect 198026 233715 203638 233743
rect 198026 233703 198032 233715
rect 203632 233703 203638 233715
rect 203690 233703 203696 233755
rect 203920 233703 203926 233755
rect 203978 233743 203984 233755
rect 214192 233743 214198 233755
rect 203978 233715 214198 233743
rect 203978 233703 203984 233715
rect 214192 233703 214198 233715
rect 214250 233703 214256 233755
rect 218704 233743 218710 233755
rect 214402 233715 218710 233743
rect 195664 233629 195670 233681
rect 195722 233669 195728 233681
rect 201328 233669 201334 233681
rect 195722 233641 201334 233669
rect 195722 233629 195728 233641
rect 201328 233629 201334 233641
rect 201386 233629 201392 233681
rect 202480 233629 202486 233681
rect 202538 233669 202544 233681
rect 212560 233669 212566 233681
rect 202538 233641 212566 233669
rect 202538 233629 202544 233641
rect 212560 233629 212566 233641
rect 212618 233629 212624 233681
rect 192880 233555 192886 233607
rect 192938 233595 192944 233607
rect 195280 233595 195286 233607
rect 192938 233567 195286 233595
rect 192938 233555 192944 233567
rect 195280 233555 195286 233567
rect 195338 233555 195344 233607
rect 195568 233555 195574 233607
rect 195626 233595 195632 233607
rect 199792 233595 199798 233607
rect 195626 233567 199798 233595
rect 195626 233555 195632 233567
rect 199792 233555 199798 233567
rect 199850 233555 199856 233607
rect 201040 233555 201046 233607
rect 201098 233595 201104 233607
rect 209680 233595 209686 233607
rect 201098 233567 209686 233595
rect 201098 233555 201104 233567
rect 209680 233555 209686 233567
rect 209738 233555 209744 233607
rect 194224 233481 194230 233533
rect 194282 233521 194288 233533
rect 198352 233521 198358 233533
rect 194282 233493 198358 233521
rect 194282 233481 194288 233493
rect 198352 233481 198358 233493
rect 198410 233481 198416 233533
rect 199120 233481 199126 233533
rect 199178 233521 199184 233533
rect 205072 233521 205078 233533
rect 199178 233493 205078 233521
rect 199178 233481 199184 233493
rect 205072 233481 205078 233493
rect 205130 233481 205136 233533
rect 205552 233481 205558 233533
rect 205610 233521 205616 233533
rect 214402 233521 214430 233715
rect 218704 233703 218710 233715
rect 218762 233703 218768 233755
rect 258352 233703 258358 233755
rect 258410 233743 258416 233755
rect 278224 233743 278230 233755
rect 258410 233715 278230 233743
rect 258410 233703 258416 233715
rect 278224 233703 278230 233715
rect 278282 233703 278288 233755
rect 304816 233703 304822 233755
rect 304874 233743 304880 233755
rect 334096 233743 334102 233755
rect 304874 233715 334102 233743
rect 304874 233703 304880 233715
rect 334096 233703 334102 233715
rect 334154 233703 334160 233755
rect 338608 233703 338614 233755
rect 338666 233743 338672 233755
rect 464560 233743 464566 233755
rect 338666 233715 464566 233743
rect 338666 233703 338672 233715
rect 464560 233703 464566 233715
rect 464618 233703 464624 233755
rect 214480 233629 214486 233681
rect 214538 233669 214544 233681
rect 217168 233669 217174 233681
rect 214538 233641 217174 233669
rect 214538 233629 214544 233641
rect 217168 233629 217174 233641
rect 217226 233629 217232 233681
rect 287440 233629 287446 233681
rect 287498 233669 287504 233681
rect 311248 233669 311254 233681
rect 287498 233641 311254 233669
rect 287498 233629 287504 233641
rect 311248 233629 311254 233641
rect 311306 233629 311312 233681
rect 324784 233629 324790 233681
rect 324842 233669 324848 233681
rect 342640 233669 342646 233681
rect 324842 233641 342646 233669
rect 324842 233629 324848 233641
rect 342640 233629 342646 233641
rect 342698 233629 342704 233681
rect 343504 233629 343510 233681
rect 343562 233669 343568 233681
rect 411472 233669 411478 233681
rect 343562 233641 411478 233669
rect 343562 233629 343568 233641
rect 411472 233629 411478 233641
rect 411530 233629 411536 233681
rect 259888 233555 259894 233607
rect 259946 233595 259952 233607
rect 267760 233595 267766 233607
rect 259946 233567 267766 233595
rect 259946 233555 259952 233567
rect 267760 233555 267766 233567
rect 267818 233555 267824 233607
rect 288400 233555 288406 233607
rect 288458 233595 288464 233607
rect 313840 233595 313846 233607
rect 288458 233567 313846 233595
rect 288458 233555 288464 233567
rect 313840 233555 313846 233567
rect 313898 233555 313904 233607
rect 329296 233555 329302 233607
rect 329354 233595 329360 233607
rect 449296 233595 449302 233607
rect 329354 233567 449302 233595
rect 329354 233555 329360 233567
rect 449296 233555 449302 233567
rect 449354 233555 449360 233607
rect 205610 233493 214430 233521
rect 205610 233481 205616 233493
rect 240592 233481 240598 233533
rect 240650 233521 240656 233533
rect 290416 233521 290422 233533
rect 240650 233493 290422 233521
rect 240650 233481 240656 233493
rect 290416 233481 290422 233493
rect 290474 233481 290480 233533
rect 297136 233481 297142 233533
rect 297194 233521 297200 233533
rect 319600 233521 319606 233533
rect 297194 233493 319606 233521
rect 297194 233481 297200 233493
rect 319600 233481 319606 233493
rect 319658 233481 319664 233533
rect 335344 233481 335350 233533
rect 335402 233521 335408 233533
rect 463600 233521 463606 233533
rect 335402 233493 463606 233521
rect 335402 233481 335408 233493
rect 463600 233481 463606 233493
rect 463658 233481 463664 233533
rect 194608 233407 194614 233459
rect 194666 233447 194672 233459
rect 196048 233447 196054 233459
rect 194666 233419 196054 233447
rect 194666 233407 194672 233419
rect 196048 233407 196054 233419
rect 196106 233407 196112 233459
rect 196528 233407 196534 233459
rect 196586 233447 196592 233459
rect 200560 233447 200566 233459
rect 196586 233419 200566 233447
rect 196586 233407 196592 233419
rect 200560 233407 200566 233419
rect 200618 233407 200624 233459
rect 200656 233407 200662 233459
rect 200714 233447 200720 233459
rect 208144 233447 208150 233459
rect 200714 233419 208150 233447
rect 200714 233407 200720 233419
rect 208144 233407 208150 233419
rect 208202 233407 208208 233459
rect 233392 233407 233398 233459
rect 233450 233447 233456 233459
rect 235984 233447 235990 233459
rect 233450 233419 235990 233447
rect 233450 233407 233456 233419
rect 235984 233407 235990 233419
rect 236042 233407 236048 233459
rect 264400 233407 264406 233459
rect 264458 233447 264464 233459
rect 271888 233447 271894 233459
rect 264458 233419 271894 233447
rect 264458 233407 264464 233419
rect 271888 233407 271894 233419
rect 271946 233407 271952 233459
rect 292912 233407 292918 233459
rect 292970 233447 292976 233459
rect 311056 233447 311062 233459
rect 292970 233419 311062 233447
rect 292970 233407 292976 233419
rect 311056 233407 311062 233419
rect 311114 233407 311120 233459
rect 317200 233407 317206 233459
rect 317258 233447 317264 233459
rect 410896 233447 410902 233459
rect 317258 233419 410902 233447
rect 317258 233407 317264 233419
rect 410896 233407 410902 233419
rect 410954 233407 410960 233459
rect 192400 233333 192406 233385
rect 192458 233373 192464 233385
rect 193744 233373 193750 233385
rect 192458 233345 193750 233373
rect 192458 233333 192464 233345
rect 193744 233333 193750 233345
rect 193802 233333 193808 233385
rect 193840 233333 193846 233385
rect 193898 233373 193904 233385
rect 196816 233373 196822 233385
rect 193898 233345 196822 233373
rect 193898 233333 193904 233345
rect 196816 233333 196822 233345
rect 196874 233333 196880 233385
rect 197872 233333 197878 233385
rect 197930 233373 197936 233385
rect 202096 233373 202102 233385
rect 197930 233345 202102 233373
rect 197930 233333 197936 233345
rect 202096 233333 202102 233345
rect 202154 233333 202160 233385
rect 202384 233333 202390 233385
rect 202442 233373 202448 233385
rect 211120 233373 211126 233385
rect 202442 233345 211126 233373
rect 202442 233333 202448 233345
rect 211120 233333 211126 233345
rect 211178 233333 211184 233385
rect 228400 233333 228406 233385
rect 228458 233373 228464 233385
rect 236368 233373 236374 233385
rect 228458 233345 236374 233373
rect 228458 233333 228464 233345
rect 236368 233333 236374 233345
rect 236426 233333 236432 233385
rect 261616 233333 261622 233385
rect 261674 233373 261680 233385
rect 269008 233373 269014 233385
rect 261674 233345 269014 233373
rect 261674 233333 261680 233345
rect 269008 233333 269014 233345
rect 269066 233333 269072 233385
rect 270544 233333 270550 233385
rect 270602 233373 270608 233385
rect 274672 233373 274678 233385
rect 270602 233345 274678 233373
rect 270602 233333 270608 233345
rect 274672 233333 274678 233345
rect 274730 233333 274736 233385
rect 311152 233333 311158 233385
rect 311210 233373 311216 233385
rect 414544 233373 414550 233385
rect 311210 233345 414550 233373
rect 311210 233333 311216 233345
rect 414544 233333 414550 233345
rect 414602 233333 414608 233385
rect 193456 233259 193462 233311
rect 193514 233299 193520 233311
rect 194608 233299 194614 233311
rect 193514 233271 194614 233299
rect 193514 233259 193520 233271
rect 194608 233259 194614 233271
rect 194666 233259 194672 233311
rect 195184 233259 195190 233311
rect 195242 233299 195248 233311
rect 195856 233299 195862 233311
rect 195242 233271 195862 233299
rect 195242 233259 195248 233271
rect 195856 233259 195862 233271
rect 195914 233259 195920 233311
rect 196144 233259 196150 233311
rect 196202 233299 196208 233311
rect 199120 233299 199126 233311
rect 196202 233271 199126 233299
rect 196202 233259 196208 233271
rect 199120 233259 199126 233271
rect 199178 233259 199184 233311
rect 199696 233259 199702 233311
rect 199754 233299 199760 233311
rect 206608 233299 206614 233311
rect 199754 233271 206614 233299
rect 199754 233259 199760 233271
rect 206608 233259 206614 233271
rect 206666 233259 206672 233311
rect 226672 233259 226678 233311
rect 226730 233299 226736 233311
rect 238960 233299 238966 233311
rect 226730 233271 238966 233299
rect 226730 233259 226736 233271
rect 238960 233259 238966 233271
rect 239018 233259 239024 233311
rect 257968 233259 257974 233311
rect 258026 233299 258032 233311
rect 269104 233299 269110 233311
rect 258026 233271 269110 233299
rect 258026 233259 258032 233271
rect 269104 233259 269110 233271
rect 269162 233259 269168 233311
rect 270256 233259 270262 233311
rect 270314 233299 270320 233311
rect 273520 233299 273526 233311
rect 270314 233271 273526 233299
rect 270314 233259 270320 233271
rect 273520 233259 273526 233271
rect 273578 233259 273584 233311
rect 320272 233259 320278 233311
rect 320330 233299 320336 233311
rect 448240 233299 448246 233311
rect 320330 233271 448246 233299
rect 320330 233259 320336 233271
rect 448240 233259 448246 233271
rect 448298 233259 448304 233311
rect 262096 233185 262102 233237
rect 262154 233225 262160 233237
rect 334192 233225 334198 233237
rect 262154 233197 334198 233225
rect 262154 233185 262160 233197
rect 334192 233185 334198 233197
rect 334250 233185 334256 233237
rect 340816 233185 340822 233237
rect 340874 233225 340880 233237
rect 491248 233225 491254 233237
rect 340874 233197 491254 233225
rect 340874 233185 340880 233197
rect 491248 233185 491254 233197
rect 491306 233185 491312 233237
rect 495376 233185 495382 233237
rect 495434 233225 495440 233237
rect 622672 233225 622678 233237
rect 495434 233197 622678 233225
rect 495434 233185 495440 233197
rect 622672 233185 622678 233197
rect 622730 233185 622736 233237
rect 260656 233111 260662 233163
rect 260714 233151 260720 233163
rect 331312 233151 331318 233163
rect 260714 233123 331318 233151
rect 260714 233111 260720 233123
rect 331312 233111 331318 233123
rect 331370 233111 331376 233163
rect 347056 233111 347062 233163
rect 347114 233151 347120 233163
rect 501040 233151 501046 233163
rect 347114 233123 501046 233151
rect 347114 233111 347120 233123
rect 501040 233111 501046 233123
rect 501098 233111 501104 233163
rect 265744 233037 265750 233089
rect 265802 233077 265808 233089
rect 338032 233077 338038 233089
rect 265802 233049 338038 233077
rect 265802 233037 265808 233049
rect 338032 233037 338038 233049
rect 338090 233037 338096 233089
rect 350320 233037 350326 233089
rect 350378 233077 350384 233089
rect 507088 233077 507094 233089
rect 350378 233049 507094 233077
rect 350378 233037 350384 233049
rect 507088 233037 507094 233049
rect 507146 233037 507152 233089
rect 290800 232963 290806 233015
rect 290858 233003 290864 233015
rect 374608 233003 374614 233015
rect 290858 232975 374614 233003
rect 290858 232963 290864 232975
rect 374608 232963 374614 232975
rect 374666 232963 374672 233015
rect 398800 232963 398806 233015
rect 398858 233003 398864 233015
rect 557008 233003 557014 233015
rect 398858 232975 557014 233003
rect 398858 232963 398864 232975
rect 557008 232963 557014 232975
rect 557066 232963 557072 233015
rect 263920 232889 263926 232941
rect 263978 232929 263984 232941
rect 337264 232929 337270 232941
rect 263978 232901 337270 232929
rect 263978 232889 263984 232901
rect 337264 232889 337270 232901
rect 337322 232889 337328 232941
rect 353104 232889 353110 232941
rect 353162 232929 353168 232941
rect 513136 232929 513142 232941
rect 353162 232901 513142 232929
rect 353162 232889 353168 232901
rect 513136 232889 513142 232901
rect 513194 232889 513200 232941
rect 513232 232889 513238 232941
rect 513290 232929 513296 232941
rect 519184 232929 519190 232941
rect 513290 232901 519190 232929
rect 513290 232889 513296 232901
rect 519184 232889 519190 232901
rect 519242 232889 519248 232941
rect 237616 232815 237622 232867
rect 237674 232855 237680 232867
rect 284368 232855 284374 232867
rect 237674 232827 284374 232855
rect 237674 232815 237680 232827
rect 284368 232815 284374 232827
rect 284426 232815 284432 232867
rect 289936 232815 289942 232867
rect 289994 232855 290000 232867
rect 382864 232855 382870 232867
rect 289994 232827 382870 232855
rect 289994 232815 290000 232827
rect 382864 232815 382870 232827
rect 382922 232815 382928 232867
rect 411760 232815 411766 232867
rect 411818 232855 411824 232867
rect 572080 232855 572086 232867
rect 411818 232827 513182 232855
rect 411818 232815 411824 232827
rect 265168 232741 265174 232793
rect 265226 232781 265232 232793
rect 340240 232781 340246 232793
rect 265226 232753 340246 232781
rect 265226 232741 265232 232753
rect 340240 232741 340246 232753
rect 340298 232741 340304 232793
rect 346288 232781 346294 232793
rect 343714 232753 346294 232781
rect 216592 232667 216598 232719
rect 216650 232707 216656 232719
rect 242128 232707 242134 232719
rect 216650 232679 242134 232707
rect 216650 232667 216656 232679
rect 242128 232667 242134 232679
rect 242186 232667 242192 232719
rect 266608 232667 266614 232719
rect 266666 232707 266672 232719
rect 343216 232707 343222 232719
rect 266666 232679 343222 232707
rect 266666 232667 266672 232679
rect 343216 232667 343222 232679
rect 343274 232667 343280 232719
rect 219760 232593 219766 232645
rect 219818 232633 219824 232645
rect 248080 232633 248086 232645
rect 219818 232605 248086 232633
rect 219818 232593 219824 232605
rect 248080 232593 248086 232605
rect 248138 232593 248144 232645
rect 268432 232593 268438 232645
rect 268490 232633 268496 232645
rect 343714 232633 343742 232753
rect 346288 232741 346294 232753
rect 346346 232741 346352 232793
rect 356272 232741 356278 232793
rect 356330 232781 356336 232793
rect 513040 232781 513046 232793
rect 356330 232753 513046 232781
rect 356330 232741 356336 232753
rect 513040 232741 513046 232753
rect 513098 232741 513104 232793
rect 513154 232781 513182 232827
rect 518386 232827 572086 232855
rect 518386 232781 518414 232827
rect 572080 232815 572086 232827
rect 572138 232815 572144 232867
rect 513154 232753 518414 232781
rect 521200 232741 521206 232793
rect 521258 232781 521264 232793
rect 626416 232781 626422 232793
rect 521258 232753 626422 232781
rect 521258 232741 521264 232753
rect 626416 232741 626422 232753
rect 626474 232741 626480 232793
rect 268490 232605 343742 232633
rect 343810 232679 346910 232707
rect 268490 232593 268496 232605
rect 218032 232519 218038 232571
rect 218090 232559 218096 232571
rect 245104 232559 245110 232571
rect 218090 232531 245110 232559
rect 218090 232519 218096 232531
rect 245104 232519 245110 232531
rect 245162 232519 245168 232571
rect 274864 232519 274870 232571
rect 274922 232559 274928 232571
rect 343810 232559 343838 232679
rect 346882 232633 346910 232679
rect 346960 232667 346966 232719
rect 347018 232707 347024 232719
rect 361360 232707 361366 232719
rect 347018 232679 361366 232707
rect 347018 232667 347024 232679
rect 361360 232667 361366 232679
rect 361418 232667 361424 232719
rect 362128 232667 362134 232719
rect 362186 232707 362192 232719
rect 531280 232707 531286 232719
rect 362186 232679 531286 232707
rect 362186 232667 362192 232679
rect 531280 232667 531286 232679
rect 531338 232667 531344 232719
rect 356080 232633 356086 232645
rect 346882 232605 356086 232633
rect 356080 232593 356086 232605
rect 356138 232593 356144 232645
rect 365392 232593 365398 232645
rect 365450 232633 365456 232645
rect 537232 232633 537238 232645
rect 365450 232605 537238 232633
rect 365450 232593 365456 232605
rect 537232 232593 537238 232605
rect 537290 232593 537296 232645
rect 274922 232531 343838 232559
rect 274922 232519 274928 232531
rect 343888 232519 343894 232571
rect 343946 232559 343952 232571
rect 355312 232559 355318 232571
rect 343946 232531 355318 232559
rect 343946 232519 343952 232531
rect 355312 232519 355318 232531
rect 355370 232519 355376 232571
rect 365008 232519 365014 232571
rect 365066 232559 365072 232571
rect 539536 232559 539542 232571
rect 365066 232531 539542 232559
rect 365066 232519 365072 232531
rect 539536 232519 539542 232531
rect 539594 232519 539600 232571
rect 222544 232445 222550 232497
rect 222602 232485 222608 232497
rect 254224 232485 254230 232497
rect 222602 232457 254230 232485
rect 222602 232445 222608 232457
rect 254224 232445 254230 232457
rect 254282 232445 254288 232497
rect 269680 232445 269686 232497
rect 269738 232485 269744 232497
rect 349360 232485 349366 232497
rect 269738 232457 349366 232485
rect 269738 232445 269744 232457
rect 349360 232445 349366 232457
rect 349418 232445 349424 232497
rect 368176 232445 368182 232497
rect 368234 232485 368240 232497
rect 543376 232485 543382 232497
rect 368234 232457 543382 232485
rect 368234 232445 368240 232457
rect 543376 232445 543382 232457
rect 543434 232445 543440 232497
rect 221104 232371 221110 232423
rect 221162 232411 221168 232423
rect 251152 232411 251158 232423
rect 221162 232383 251158 232411
rect 221162 232371 221168 232383
rect 251152 232371 251158 232383
rect 251210 232371 251216 232423
rect 271216 232371 271222 232423
rect 271274 232411 271280 232423
rect 352336 232411 352342 232423
rect 271274 232383 352342 232411
rect 271274 232371 271280 232383
rect 352336 232371 352342 232383
rect 352394 232371 352400 232423
rect 366256 232371 366262 232423
rect 366314 232411 366320 232423
rect 542608 232411 542614 232423
rect 366314 232383 542614 232411
rect 366314 232371 366320 232383
rect 542608 232371 542614 232383
rect 542666 232371 542672 232423
rect 222928 232297 222934 232349
rect 222986 232337 222992 232349
rect 255664 232337 255670 232349
rect 222986 232309 255670 232337
rect 222986 232297 222992 232309
rect 255664 232297 255670 232309
rect 255722 232297 255728 232349
rect 272944 232297 272950 232349
rect 273002 232337 273008 232349
rect 343888 232337 343894 232349
rect 273002 232309 343894 232337
rect 273002 232297 273008 232309
rect 343888 232297 343894 232309
rect 343946 232297 343952 232349
rect 343984 232297 343990 232349
rect 344042 232337 344048 232349
rect 350512 232337 350518 232349
rect 344042 232309 350518 232337
rect 344042 232297 344048 232309
rect 350512 232297 350518 232309
rect 350570 232297 350576 232349
rect 371152 232297 371158 232349
rect 371210 232337 371216 232349
rect 549424 232337 549430 232349
rect 371210 232309 549430 232337
rect 371210 232297 371216 232309
rect 549424 232297 549430 232309
rect 549482 232297 549488 232349
rect 226288 232223 226294 232275
rect 226346 232263 226352 232275
rect 261712 232263 261718 232275
rect 226346 232235 261718 232263
rect 226346 232223 226352 232235
rect 261712 232223 261718 232235
rect 261770 232223 261776 232275
rect 274192 232223 274198 232275
rect 274250 232263 274256 232275
rect 358288 232263 358294 232275
rect 274250 232235 358294 232263
rect 274250 232223 274256 232235
rect 358288 232223 358294 232235
rect 358346 232223 358352 232275
rect 372688 232223 372694 232275
rect 372746 232263 372752 232275
rect 552400 232263 552406 232275
rect 372746 232235 552406 232263
rect 372746 232223 372752 232235
rect 552400 232223 552406 232235
rect 552458 232223 552464 232275
rect 224272 232149 224278 232201
rect 224330 232189 224336 232201
rect 257200 232189 257206 232201
rect 224330 232161 257206 232189
rect 224330 232149 224336 232161
rect 257200 232149 257206 232161
rect 257258 232149 257264 232201
rect 277456 232149 277462 232201
rect 277514 232189 277520 232201
rect 364432 232189 364438 232201
rect 277514 232161 364438 232189
rect 277514 232149 277520 232161
rect 364432 232149 364438 232161
rect 364490 232149 364496 232201
rect 368080 232149 368086 232201
rect 368138 232189 368144 232201
rect 545584 232189 545590 232201
rect 368138 232161 545590 232189
rect 368138 232149 368144 232161
rect 545584 232149 545590 232161
rect 545642 232149 545648 232201
rect 227056 232075 227062 232127
rect 227114 232115 227120 232127
rect 263248 232115 263254 232127
rect 227114 232087 263254 232115
rect 227114 232075 227120 232087
rect 263248 232075 263254 232087
rect 263306 232075 263312 232127
rect 275728 232075 275734 232127
rect 275786 232115 275792 232127
rect 346960 232115 346966 232127
rect 275786 232087 346966 232115
rect 275786 232075 275792 232087
rect 346960 232075 346966 232087
rect 347018 232075 347024 232127
rect 350512 232075 350518 232127
rect 350570 232115 350576 232127
rect 367120 232115 367126 232127
rect 350570 232087 367126 232115
rect 350570 232075 350576 232087
rect 367120 232075 367126 232087
rect 367178 232075 367184 232127
rect 369520 232075 369526 232127
rect 369578 232115 369584 232127
rect 548560 232115 548566 232127
rect 369578 232087 548566 232115
rect 369578 232075 369584 232087
rect 548560 232075 548566 232087
rect 548618 232075 548624 232127
rect 147664 232001 147670 232053
rect 147722 232041 147728 232053
rect 154096 232041 154102 232053
rect 147722 232013 154102 232041
rect 147722 232001 147728 232013
rect 154096 232001 154102 232013
rect 154154 232001 154160 232053
rect 233872 232001 233878 232053
rect 233930 232041 233936 232053
rect 274480 232041 274486 232053
rect 233930 232013 274486 232041
rect 233930 232001 233936 232013
rect 274480 232001 274486 232013
rect 274538 232001 274544 232053
rect 280240 232001 280246 232053
rect 280298 232041 280304 232053
rect 370384 232041 370390 232053
rect 280298 232013 370390 232041
rect 280298 232001 280304 232013
rect 370384 232001 370390 232013
rect 370442 232001 370448 232053
rect 375760 232001 375766 232053
rect 375818 232041 375824 232053
rect 558448 232041 558454 232053
rect 375818 232013 558454 232041
rect 375818 232001 375824 232013
rect 558448 232001 558454 232013
rect 558506 232001 558512 232053
rect 234832 231927 234838 231979
rect 234890 231967 234896 231979
rect 278320 231967 278326 231979
rect 234890 231939 278326 231967
rect 234890 231927 234896 231939
rect 278320 231927 278326 231939
rect 278378 231927 278384 231979
rect 278992 231927 278998 231979
rect 279050 231967 279056 231979
rect 367408 231967 367414 231979
rect 279050 231939 367414 231967
rect 279050 231927 279056 231939
rect 367408 231927 367414 231939
rect 367466 231927 367472 231979
rect 372304 231927 372310 231979
rect 372362 231967 372368 231979
rect 554704 231967 554710 231979
rect 372362 231939 554710 231967
rect 372362 231927 372368 231939
rect 554704 231927 554710 231939
rect 554762 231927 554768 231979
rect 233200 231853 233206 231905
rect 233258 231893 233264 231905
rect 275344 231893 275350 231905
rect 233258 231865 275350 231893
rect 233258 231853 233264 231865
rect 275344 231853 275350 231865
rect 275402 231853 275408 231905
rect 281968 231853 281974 231905
rect 282026 231893 282032 231905
rect 373456 231893 373462 231905
rect 282026 231865 373462 231893
rect 282026 231853 282032 231865
rect 373456 231853 373462 231865
rect 373514 231853 373520 231905
rect 374032 231853 374038 231905
rect 374090 231893 374096 231905
rect 557584 231893 557590 231905
rect 374090 231865 557590 231893
rect 374090 231853 374096 231865
rect 557584 231853 557590 231865
rect 557642 231853 557648 231905
rect 236080 231779 236086 231831
rect 236138 231819 236144 231831
rect 281296 231819 281302 231831
rect 236138 231791 281302 231819
rect 236138 231779 236144 231791
rect 281296 231779 281302 231791
rect 281354 231779 281360 231831
rect 295312 231779 295318 231831
rect 295370 231819 295376 231831
rect 400240 231819 400246 231831
rect 295370 231791 400246 231819
rect 295370 231779 295376 231791
rect 400240 231779 400246 231791
rect 400298 231779 400304 231831
rect 405040 231779 405046 231831
rect 405098 231819 405104 231831
rect 604528 231819 604534 231831
rect 405098 231791 604534 231819
rect 405098 231779 405104 231791
rect 604528 231779 604534 231791
rect 604586 231779 604592 231831
rect 259120 231705 259126 231757
rect 259178 231745 259184 231757
rect 328144 231745 328150 231757
rect 259178 231717 328150 231745
rect 259178 231705 259184 231717
rect 328144 231705 328150 231717
rect 328202 231705 328208 231757
rect 346960 231705 346966 231757
rect 347018 231745 347024 231757
rect 362128 231745 362134 231757
rect 347018 231717 362134 231745
rect 347018 231705 347024 231717
rect 362128 231705 362134 231717
rect 362186 231705 362192 231757
rect 367120 231705 367126 231757
rect 367178 231745 367184 231757
rect 495088 231745 495094 231757
rect 367178 231717 495094 231745
rect 367178 231705 367184 231717
rect 495088 231705 495094 231717
rect 495146 231705 495152 231757
rect 498544 231705 498550 231757
rect 498602 231745 498608 231757
rect 614992 231745 614998 231757
rect 498602 231717 614998 231745
rect 498602 231705 498608 231717
rect 614992 231705 614998 231717
rect 615050 231705 615056 231757
rect 258736 231631 258742 231683
rect 258794 231671 258800 231683
rect 326704 231671 326710 231683
rect 258794 231643 326710 231671
rect 258794 231631 258800 231643
rect 326704 231631 326710 231643
rect 326762 231631 326768 231683
rect 337552 231631 337558 231683
rect 337610 231671 337616 231683
rect 485200 231671 485206 231683
rect 337610 231643 485206 231671
rect 337610 231631 337616 231643
rect 485200 231631 485206 231643
rect 485258 231631 485264 231683
rect 255760 231557 255766 231609
rect 255818 231597 255824 231609
rect 320656 231597 320662 231609
rect 255818 231569 320662 231597
rect 255818 231557 255824 231569
rect 320656 231557 320662 231569
rect 320714 231557 320720 231609
rect 327088 231557 327094 231609
rect 327146 231597 327152 231609
rect 464080 231597 464086 231609
rect 327146 231569 464086 231597
rect 327146 231557 327152 231569
rect 464080 231557 464086 231569
rect 464138 231557 464144 231609
rect 248368 231483 248374 231535
rect 248426 231523 248432 231535
rect 305488 231523 305494 231535
rect 248426 231495 305494 231523
rect 248426 231483 248432 231495
rect 305488 231483 305494 231495
rect 305546 231483 305552 231535
rect 312208 231483 312214 231535
rect 312266 231523 312272 231535
rect 433840 231523 433846 231535
rect 312266 231495 433846 231523
rect 312266 231483 312272 231495
rect 433840 231483 433846 231495
rect 433898 231483 433904 231535
rect 292528 231409 292534 231461
rect 292586 231449 292592 231461
rect 379984 231449 379990 231461
rect 292586 231421 379990 231449
rect 292586 231409 292592 231421
rect 379984 231409 379990 231421
rect 380042 231409 380048 231461
rect 400432 231409 400438 231461
rect 400490 231449 400496 231461
rect 520720 231449 520726 231461
rect 400490 231421 520726 231449
rect 400490 231409 400496 231421
rect 520720 231409 520726 231421
rect 520778 231409 520784 231461
rect 293104 231335 293110 231387
rect 293162 231375 293168 231387
rect 371632 231375 371638 231387
rect 293162 231347 371638 231375
rect 293162 231335 293168 231347
rect 371632 231335 371638 231347
rect 371690 231335 371696 231387
rect 400336 231335 400342 231387
rect 400394 231375 400400 231387
rect 499600 231375 499606 231387
rect 400394 231347 499606 231375
rect 400394 231335 400400 231347
rect 499600 231335 499606 231347
rect 499658 231335 499664 231387
rect 281200 231261 281206 231313
rect 281258 231301 281264 231313
rect 289264 231301 289270 231313
rect 281258 231273 289270 231301
rect 281258 231261 281264 231273
rect 289264 231261 289270 231273
rect 289322 231261 289328 231313
rect 293488 231261 293494 231313
rect 293546 231301 293552 231313
rect 364240 231301 364246 231313
rect 293546 231273 364246 231301
rect 293546 231261 293552 231273
rect 364240 231261 364246 231273
rect 364298 231261 364304 231313
rect 395248 231261 395254 231313
rect 395306 231301 395312 231313
rect 485968 231301 485974 231313
rect 395306 231273 485974 231301
rect 395306 231261 395312 231273
rect 485968 231261 485974 231273
rect 486026 231261 486032 231313
rect 257584 231187 257590 231239
rect 257642 231227 257648 231239
rect 325168 231227 325174 231239
rect 257642 231199 325174 231227
rect 257642 231187 257648 231199
rect 325168 231187 325174 231199
rect 325226 231187 325232 231239
rect 334096 231187 334102 231239
rect 334154 231227 334160 231239
rect 416464 231227 416470 231239
rect 334154 231199 416470 231227
rect 334154 231187 334160 231199
rect 416464 231187 416470 231199
rect 416522 231187 416528 231239
rect 256144 231113 256150 231165
rect 256202 231153 256208 231165
rect 322096 231153 322102 231165
rect 256202 231125 322102 231153
rect 256202 231113 256208 231125
rect 322096 231113 322102 231125
rect 322154 231113 322160 231165
rect 331216 231113 331222 231165
rect 331274 231153 331280 231165
rect 395344 231153 395350 231165
rect 331274 231125 395350 231153
rect 331274 231113 331280 231125
rect 395344 231113 395350 231125
rect 395402 231113 395408 231165
rect 395728 231113 395734 231165
rect 395786 231153 395792 231165
rect 473872 231153 473878 231165
rect 395786 231125 473878 231153
rect 395786 231113 395792 231125
rect 473872 231113 473878 231125
rect 473930 231113 473936 231165
rect 149392 231039 149398 231091
rect 149450 231079 149456 231091
rect 159856 231079 159862 231091
rect 149450 231051 159862 231079
rect 149450 231039 149456 231051
rect 159856 231039 159862 231051
rect 159914 231039 159920 231091
rect 252976 231039 252982 231091
rect 253034 231079 253040 231091
rect 314512 231079 314518 231091
rect 253034 231051 314518 231079
rect 253034 231039 253040 231051
rect 314512 231039 314518 231051
rect 314570 231039 314576 231091
rect 328336 231039 328342 231091
rect 328394 231079 328400 231091
rect 368752 231079 368758 231091
rect 328394 231051 368758 231079
rect 328394 231039 328400 231051
rect 368752 231039 368758 231051
rect 368810 231039 368816 231091
rect 245200 230965 245206 231017
rect 245258 231005 245264 231017
rect 299440 231005 299446 231017
rect 245258 230977 299446 231005
rect 245258 230965 245264 230977
rect 299440 230965 299446 230977
rect 299498 230965 299504 231017
rect 308176 230965 308182 231017
rect 308234 231005 308240 231017
rect 323632 231005 323638 231017
rect 308234 230977 323638 231005
rect 308234 230965 308240 230977
rect 323632 230965 323638 230977
rect 323690 230965 323696 231017
rect 344656 230965 344662 231017
rect 344714 231005 344720 231017
rect 409648 231005 409654 231017
rect 344714 230977 409654 231005
rect 344714 230965 344720 230977
rect 409648 230965 409654 230977
rect 409706 230965 409712 231017
rect 416368 230965 416374 231017
rect 416426 231005 416432 231017
rect 424048 231005 424054 231017
rect 416426 230977 424054 231005
rect 416426 230965 416432 230977
rect 424048 230965 424054 230977
rect 424106 230965 424112 231017
rect 326800 230891 326806 230943
rect 326858 230931 326864 230943
rect 380272 230931 380278 230943
rect 326858 230903 380278 230931
rect 326858 230891 326864 230903
rect 380272 230891 380278 230903
rect 380330 230891 380336 230943
rect 385936 230891 385942 230943
rect 385994 230931 386000 230943
rect 449680 230931 449686 230943
rect 385994 230903 449686 230931
rect 385994 230891 386000 230903
rect 449680 230891 449686 230903
rect 449738 230891 449744 230943
rect 290704 230817 290710 230869
rect 290762 230857 290768 230869
rect 297424 230857 297430 230869
rect 290762 230829 297430 230857
rect 290762 230817 290768 230829
rect 297424 230817 297430 230829
rect 297482 230817 297488 230869
rect 313936 230817 313942 230869
rect 313994 230857 314000 230869
rect 346960 230857 346966 230869
rect 313994 230829 346966 230857
rect 313994 230817 314000 230829
rect 346960 230817 346966 230829
rect 347018 230817 347024 230869
rect 358384 230817 358390 230869
rect 358442 230857 358448 230869
rect 419536 230857 419542 230869
rect 358442 230829 419542 230857
rect 358442 230817 358448 230829
rect 419536 230817 419542 230829
rect 419594 230817 419600 230869
rect 323344 230743 323350 230795
rect 323402 230783 323408 230795
rect 377104 230783 377110 230795
rect 323402 230755 377110 230783
rect 323402 230743 323408 230755
rect 377104 230743 377110 230755
rect 377162 230743 377168 230795
rect 320752 230669 320758 230721
rect 320810 230709 320816 230721
rect 368560 230709 368566 230721
rect 320810 230681 368566 230709
rect 320810 230669 320816 230681
rect 368560 230669 368566 230681
rect 368618 230669 368624 230721
rect 368752 230669 368758 230721
rect 368810 230709 368816 230721
rect 401392 230709 401398 230721
rect 368810 230681 401398 230709
rect 368810 230669 368816 230681
rect 401392 230669 401398 230681
rect 401450 230669 401456 230721
rect 302320 230595 302326 230647
rect 302378 230635 302384 230647
rect 308560 230635 308566 230647
rect 302378 230607 308566 230635
rect 302378 230595 302384 230607
rect 308560 230595 308566 230607
rect 308618 230595 308624 230647
rect 323248 230595 323254 230647
rect 323306 230635 323312 230647
rect 329584 230635 329590 230647
rect 323306 230607 329590 230635
rect 323306 230595 323312 230607
rect 329584 230595 329590 230607
rect 329642 230595 329648 230647
rect 354256 230595 354262 230647
rect 354314 230635 354320 230647
rect 404464 230635 404470 230647
rect 354314 230607 368510 230635
rect 354314 230595 354320 230607
rect 306736 230521 306742 230573
rect 306794 230561 306800 230573
rect 317584 230561 317590 230573
rect 306794 230533 317590 230561
rect 306794 230521 306800 230533
rect 317584 230521 317590 230533
rect 317642 230521 317648 230573
rect 321040 230521 321046 230573
rect 321098 230561 321104 230573
rect 368176 230561 368182 230573
rect 321098 230533 368182 230561
rect 321098 230521 321104 230533
rect 368176 230521 368182 230533
rect 368234 230521 368240 230573
rect 368482 230561 368510 230607
rect 383026 230607 404470 230635
rect 383026 230561 383054 230607
rect 404464 230595 404470 230607
rect 404522 230595 404528 230647
rect 368482 230533 383054 230561
rect 299344 230447 299350 230499
rect 299402 230487 299408 230499
rect 302512 230487 302518 230499
rect 299402 230459 302518 230487
rect 299402 230447 299408 230459
rect 302512 230447 302518 230459
rect 302570 230447 302576 230499
rect 304144 230447 304150 230499
rect 304202 230487 304208 230499
rect 311632 230487 311638 230499
rect 304202 230459 311638 230487
rect 304202 230447 304208 230459
rect 311632 230447 311638 230459
rect 311690 230447 311696 230499
rect 318352 230447 318358 230499
rect 318410 230487 318416 230499
rect 365104 230487 365110 230499
rect 318410 230459 365110 230487
rect 318410 230447 318416 230459
rect 365104 230447 365110 230459
rect 365162 230447 365168 230499
rect 398896 230447 398902 230499
rect 398954 230487 398960 230499
rect 410512 230487 410518 230499
rect 398954 230459 410518 230487
rect 398954 230447 398960 230459
rect 410512 230447 410518 230459
rect 410570 230447 410576 230499
rect 423376 230447 423382 230499
rect 423434 230487 423440 230499
rect 436144 230487 436150 230499
rect 423434 230459 436150 230487
rect 423434 230447 423440 230459
rect 436144 230447 436150 230459
rect 436202 230447 436208 230499
rect 248944 230373 248950 230425
rect 249002 230413 249008 230425
rect 304816 230413 304822 230425
rect 249002 230385 304822 230413
rect 249002 230373 249008 230385
rect 304816 230373 304822 230385
rect 304874 230373 304880 230425
rect 321232 230373 321238 230425
rect 321290 230413 321296 230425
rect 451984 230413 451990 230425
rect 321290 230385 451990 230413
rect 321290 230373 321296 230385
rect 451984 230373 451990 230385
rect 452042 230373 452048 230425
rect 228880 230299 228886 230351
rect 228938 230339 228944 230351
rect 267856 230339 267862 230351
rect 228938 230311 267862 230339
rect 228938 230299 228944 230311
rect 267856 230299 267862 230311
rect 267914 230299 267920 230351
rect 269104 230299 269110 230351
rect 269162 230339 269168 230351
rect 322960 230339 322966 230351
rect 269162 230311 322966 230339
rect 269162 230299 269168 230311
rect 322960 230299 322966 230311
rect 323018 230299 323024 230351
rect 325744 230299 325750 230351
rect 325802 230339 325808 230351
rect 461008 230339 461014 230351
rect 325802 230311 461014 230339
rect 325802 230299 325808 230311
rect 461008 230299 461014 230311
rect 461066 230299 461072 230351
rect 463600 230299 463606 230351
rect 463658 230339 463664 230351
rect 478384 230339 478390 230351
rect 463658 230311 478390 230339
rect 463658 230299 463664 230311
rect 478384 230299 478390 230311
rect 478442 230299 478448 230351
rect 247024 230225 247030 230277
rect 247082 230265 247088 230277
rect 303952 230265 303958 230277
rect 247082 230237 303958 230265
rect 247082 230225 247088 230237
rect 303952 230225 303958 230237
rect 304010 230225 304016 230277
rect 305104 230225 305110 230277
rect 305162 230265 305168 230277
rect 326800 230265 326806 230277
rect 305162 230237 326806 230265
rect 305162 230225 305168 230237
rect 326800 230225 326806 230237
rect 326858 230225 326864 230277
rect 458032 230265 458038 230277
rect 328450 230237 458038 230265
rect 248752 230151 248758 230203
rect 248810 230191 248816 230203
rect 307024 230191 307030 230203
rect 248810 230163 307030 230191
rect 248810 230151 248816 230163
rect 307024 230151 307030 230163
rect 307082 230151 307088 230203
rect 324016 230151 324022 230203
rect 324074 230191 324080 230203
rect 328450 230191 328478 230237
rect 458032 230225 458038 230237
rect 458090 230225 458096 230277
rect 464560 230225 464566 230277
rect 464618 230265 464624 230277
rect 484432 230265 484438 230277
rect 464618 230237 484438 230265
rect 464618 230225 464624 230237
rect 484432 230225 484438 230237
rect 484490 230225 484496 230277
rect 324074 230163 328478 230191
rect 324074 230151 324080 230163
rect 328528 230151 328534 230203
rect 328586 230191 328592 230203
rect 467056 230191 467062 230203
rect 328586 230163 467062 230191
rect 328586 230151 328592 230163
rect 467056 230151 467062 230163
rect 467114 230151 467120 230203
rect 475216 230151 475222 230203
rect 475274 230191 475280 230203
rect 601456 230191 601462 230203
rect 475274 230163 601462 230191
rect 475274 230151 475280 230163
rect 601456 230151 601462 230163
rect 601514 230151 601520 230203
rect 251920 230077 251926 230129
rect 251978 230117 251984 230129
rect 310768 230117 310774 230129
rect 251978 230089 310774 230117
rect 251978 230077 251984 230089
rect 310768 230077 310774 230089
rect 310826 230077 310832 230129
rect 331600 230077 331606 230129
rect 331658 230117 331664 230129
rect 473104 230117 473110 230129
rect 331658 230089 473110 230117
rect 331658 230077 331664 230089
rect 473104 230077 473110 230089
rect 473162 230077 473168 230129
rect 479248 230077 479254 230129
rect 479306 230117 479312 230129
rect 609040 230117 609046 230129
rect 479306 230089 609046 230117
rect 479306 230077 479312 230089
rect 609040 230077 609046 230089
rect 609098 230077 609104 230129
rect 251536 230003 251542 230055
rect 251594 230043 251600 230055
rect 313072 230043 313078 230055
rect 251594 230015 313078 230043
rect 251594 230003 251600 230015
rect 313072 230003 313078 230015
rect 313130 230003 313136 230055
rect 336304 230003 336310 230055
rect 336362 230043 336368 230055
rect 482128 230043 482134 230055
rect 336362 230015 482134 230043
rect 336362 230003 336368 230015
rect 482128 230003 482134 230015
rect 482186 230003 482192 230055
rect 486640 230003 486646 230055
rect 486698 230043 486704 230055
rect 612112 230043 612118 230055
rect 486698 230015 612118 230043
rect 486698 230003 486704 230015
rect 612112 230003 612118 230015
rect 612170 230003 612176 230055
rect 227440 229929 227446 229981
rect 227498 229969 227504 229981
rect 264784 229969 264790 229981
rect 227498 229941 264790 229969
rect 227498 229929 227504 229941
rect 264784 229929 264790 229941
rect 264842 229929 264848 229981
rect 290896 229929 290902 229981
rect 290954 229969 290960 229981
rect 331888 229969 331894 229981
rect 290954 229941 331894 229969
rect 290954 229929 290960 229941
rect 331888 229929 331894 229941
rect 331946 229929 331952 229981
rect 348496 229929 348502 229981
rect 348554 229969 348560 229981
rect 504016 229969 504022 229981
rect 348554 229941 504022 229969
rect 348554 229929 348560 229941
rect 504016 229929 504022 229941
rect 504074 229929 504080 229981
rect 253072 229855 253078 229907
rect 253130 229895 253136 229907
rect 316144 229895 316150 229907
rect 253130 229867 316150 229895
rect 253130 229855 253136 229867
rect 316144 229855 316150 229867
rect 316202 229855 316208 229907
rect 351760 229855 351766 229907
rect 351818 229895 351824 229907
rect 510160 229895 510166 229907
rect 351818 229867 510166 229895
rect 351818 229855 351824 229867
rect 510160 229855 510166 229867
rect 510218 229855 510224 229907
rect 512176 229855 512182 229907
rect 512234 229895 512240 229907
rect 625552 229895 625558 229907
rect 512234 229867 625558 229895
rect 512234 229855 512240 229867
rect 625552 229855 625558 229867
rect 625610 229855 625616 229907
rect 146896 229781 146902 229833
rect 146954 229821 146960 229833
rect 151216 229821 151222 229833
rect 146954 229793 151222 229821
rect 146954 229781 146960 229793
rect 151216 229781 151222 229793
rect 151274 229781 151280 229833
rect 239728 229781 239734 229833
rect 239786 229821 239792 229833
rect 288880 229821 288886 229833
rect 239786 229793 288886 229821
rect 239786 229781 239792 229793
rect 288880 229781 288886 229793
rect 288938 229781 288944 229833
rect 291184 229781 291190 229833
rect 291242 229821 291248 229833
rect 382960 229821 382966 229833
rect 291242 229793 382966 229821
rect 291242 229781 291248 229793
rect 382960 229781 382966 229793
rect 383018 229781 383024 229833
rect 389104 229781 389110 229833
rect 389162 229821 389168 229833
rect 396976 229821 396982 229833
rect 389162 229793 396982 229821
rect 389162 229781 389168 229793
rect 396976 229781 396982 229793
rect 397034 229781 397040 229833
rect 406960 229781 406966 229833
rect 407018 229821 407024 229833
rect 565936 229821 565942 229833
rect 407018 229793 565942 229821
rect 407018 229781 407024 229793
rect 565936 229781 565942 229793
rect 565994 229781 566000 229833
rect 220144 229707 220150 229759
rect 220202 229747 220208 229759
rect 249712 229747 249718 229759
rect 220202 229719 249718 229747
rect 220202 229707 220208 229719
rect 249712 229707 249718 229719
rect 249770 229707 249776 229759
rect 255184 229707 255190 229759
rect 255242 229747 255248 229759
rect 316816 229747 316822 229759
rect 255242 229719 316822 229747
rect 255242 229707 255248 229719
rect 316816 229707 316822 229719
rect 316874 229707 316880 229759
rect 354832 229707 354838 229759
rect 354890 229747 354896 229759
rect 516112 229747 516118 229759
rect 354890 229719 516118 229747
rect 354890 229707 354896 229719
rect 516112 229707 516118 229719
rect 516170 229707 516176 229759
rect 528400 229707 528406 229759
rect 528458 229747 528464 229759
rect 605968 229747 605974 229759
rect 528458 229719 605974 229747
rect 528458 229707 528464 229719
rect 605968 229707 605974 229719
rect 606026 229707 606032 229759
rect 221584 229633 221590 229685
rect 221642 229673 221648 229685
rect 252592 229673 252598 229685
rect 221642 229645 252598 229673
rect 221642 229633 221648 229645
rect 252592 229633 252598 229645
rect 252650 229633 252656 229685
rect 254800 229633 254806 229685
rect 254858 229673 254864 229685
rect 319120 229673 319126 229685
rect 254858 229645 319126 229673
rect 254858 229633 254864 229645
rect 319120 229633 319126 229645
rect 319178 229633 319184 229685
rect 360880 229633 360886 229685
rect 360938 229673 360944 229685
rect 360938 229645 368654 229673
rect 360938 229633 360944 229645
rect 241072 229559 241078 229611
rect 241130 229599 241136 229611
rect 291952 229599 291958 229611
rect 241130 229571 291958 229599
rect 241130 229559 241136 229571
rect 291952 229559 291958 229571
rect 292010 229559 292016 229611
rect 298096 229559 298102 229611
rect 298154 229599 298160 229611
rect 362800 229599 362806 229611
rect 298154 229571 362806 229599
rect 298154 229559 298160 229571
rect 362800 229559 362806 229571
rect 362858 229559 362864 229611
rect 368626 229599 368654 229645
rect 369904 229633 369910 229685
rect 369962 229673 369968 229685
rect 378544 229673 378550 229685
rect 369962 229645 378550 229673
rect 369962 229633 369968 229645
rect 378544 229633 378550 229645
rect 378602 229633 378608 229685
rect 378640 229633 378646 229685
rect 378698 229673 378704 229685
rect 522160 229673 522166 229685
rect 378698 229645 522166 229673
rect 378698 229633 378704 229645
rect 522160 229633 522166 229645
rect 522218 229633 522224 229685
rect 522640 229633 522646 229685
rect 522698 229673 522704 229685
rect 630160 229673 630166 229685
rect 522698 229645 630166 229673
rect 522698 229633 522704 229645
rect 630160 229633 630166 229645
rect 630218 229633 630224 229685
rect 528304 229599 528310 229611
rect 368626 229571 528310 229599
rect 528304 229559 528310 229571
rect 528362 229559 528368 229611
rect 528496 229559 528502 229611
rect 528554 229599 528560 229611
rect 628624 229599 628630 229611
rect 528554 229571 628630 229599
rect 528554 229559 528560 229571
rect 628624 229559 628630 229571
rect 628682 229559 628688 229611
rect 215248 229485 215254 229537
rect 215306 229525 215312 229537
rect 239056 229525 239062 229537
rect 215306 229497 239062 229525
rect 215306 229485 215312 229497
rect 239056 229485 239062 229497
rect 239114 229485 239120 229537
rect 244240 229485 244246 229537
rect 244298 229525 244304 229537
rect 298000 229525 298006 229537
rect 244298 229497 298006 229525
rect 244298 229485 244304 229497
rect 298000 229485 298006 229497
rect 298058 229485 298064 229537
rect 298384 229485 298390 229537
rect 298442 229525 298448 229537
rect 406768 229525 406774 229537
rect 298442 229497 406774 229525
rect 298442 229485 298448 229497
rect 406768 229485 406774 229497
rect 406826 229485 406832 229537
rect 406864 229485 406870 229537
rect 406922 229525 406928 229537
rect 575056 229525 575062 229537
rect 406922 229497 575062 229525
rect 406922 229485 406928 229497
rect 575056 229485 575062 229497
rect 575114 229485 575120 229537
rect 264304 229411 264310 229463
rect 264362 229451 264368 229463
rect 334960 229451 334966 229463
rect 264362 229423 334966 229451
rect 264362 229411 264368 229423
rect 334960 229411 334966 229423
rect 335018 229411 335024 229463
rect 366640 229411 366646 229463
rect 366698 229451 366704 229463
rect 540304 229451 540310 229463
rect 366698 229423 540310 229451
rect 366698 229411 366704 229423
rect 540304 229411 540310 229423
rect 540362 229411 540368 229463
rect 231856 229337 231862 229389
rect 231914 229377 231920 229389
rect 272272 229377 272278 229389
rect 231914 229349 272278 229377
rect 231914 229337 231920 229349
rect 272272 229337 272278 229349
rect 272330 229337 272336 229389
rect 273520 229337 273526 229389
rect 273578 229377 273584 229389
rect 347056 229377 347062 229389
rect 273578 229349 347062 229377
rect 273578 229337 273584 229349
rect 347056 229337 347062 229349
rect 347114 229337 347120 229389
rect 357616 229337 357622 229389
rect 357674 229377 357680 229389
rect 378640 229377 378646 229389
rect 357674 229349 378646 229377
rect 357674 229337 357680 229349
rect 378640 229337 378646 229349
rect 378698 229337 378704 229389
rect 378736 229337 378742 229389
rect 378794 229377 378800 229389
rect 546352 229377 546358 229389
rect 378794 229349 546358 229377
rect 378794 229337 378800 229349
rect 546352 229337 546358 229349
rect 546410 229337 546416 229389
rect 230800 229263 230806 229315
rect 230858 229303 230864 229315
rect 270736 229303 270742 229315
rect 230858 229275 270742 229303
rect 230858 229263 230864 229275
rect 270736 229263 270742 229275
rect 270794 229263 270800 229315
rect 283504 229263 283510 229315
rect 283562 229303 283568 229315
rect 367504 229303 367510 229315
rect 283562 229275 367510 229303
rect 283562 229263 283568 229275
rect 367504 229263 367510 229275
rect 367562 229263 367568 229315
rect 374128 229263 374134 229315
rect 374186 229303 374192 229315
rect 555376 229303 555382 229315
rect 374186 229275 555382 229303
rect 374186 229263 374192 229275
rect 555376 229263 555382 229275
rect 555434 229263 555440 229315
rect 233488 229189 233494 229241
rect 233546 229229 233552 229241
rect 276784 229229 276790 229241
rect 233546 229201 276790 229229
rect 233546 229189 233552 229201
rect 276784 229189 276790 229201
rect 276842 229189 276848 229241
rect 282160 229189 282166 229241
rect 282218 229229 282224 229241
rect 371248 229229 371254 229241
rect 282218 229201 371254 229229
rect 282218 229189 282224 229201
rect 371248 229189 371254 229201
rect 371306 229189 371312 229241
rect 377200 229189 377206 229241
rect 377258 229229 377264 229241
rect 561424 229229 561430 229241
rect 377258 229201 561430 229229
rect 377258 229189 377264 229201
rect 561424 229189 561430 229201
rect 561482 229189 561488 229241
rect 231952 229115 231958 229167
rect 232010 229155 232016 229167
rect 273808 229155 273814 229167
rect 232010 229127 273814 229155
rect 232010 229115 232016 229127
rect 273808 229115 273814 229127
rect 273866 229115 273872 229167
rect 284752 229115 284758 229167
rect 284810 229155 284816 229167
rect 371536 229155 371542 229167
rect 284810 229127 371542 229155
rect 284810 229115 284816 229127
rect 371536 229115 371542 229127
rect 371594 229115 371600 229167
rect 376816 229115 376822 229167
rect 376874 229155 376880 229167
rect 563632 229155 563638 229167
rect 376874 229127 563638 229155
rect 376874 229115 376880 229127
rect 563632 229115 563638 229127
rect 563690 229115 563696 229167
rect 235216 229041 235222 229093
rect 235274 229081 235280 229093
rect 279856 229081 279862 229093
rect 235274 229053 279862 229081
rect 235274 229041 235280 229053
rect 279856 229041 279862 229053
rect 279914 229041 279920 229093
rect 286288 229041 286294 229093
rect 286346 229081 286352 229093
rect 374512 229081 374518 229093
rect 286346 229053 374518 229081
rect 286346 229041 286352 229053
rect 374512 229041 374518 229053
rect 374570 229041 374576 229093
rect 380464 229041 380470 229093
rect 380522 229081 380528 229093
rect 567472 229081 567478 229093
rect 380522 229053 567478 229081
rect 380522 229041 380528 229053
rect 567472 229041 567478 229053
rect 567530 229041 567536 229093
rect 238384 228967 238390 229019
rect 238442 229007 238448 229019
rect 283600 229007 283606 229019
rect 238442 228979 283606 229007
rect 238442 228967 238448 228979
rect 283600 228967 283606 228979
rect 283658 228967 283664 229019
rect 287920 228967 287926 229019
rect 287978 229007 287984 229019
rect 374416 229007 374422 229019
rect 287978 228979 374422 229007
rect 287978 228967 287984 228979
rect 374416 228967 374422 228979
rect 374474 228967 374480 229019
rect 379888 228967 379894 229019
rect 379946 229007 379952 229019
rect 569776 229007 569782 229019
rect 379946 228979 569782 229007
rect 379946 228967 379952 228979
rect 569776 228967 569782 228979
rect 569834 228967 569840 229019
rect 245776 228893 245782 228945
rect 245834 228933 245840 228945
rect 300976 228933 300982 228945
rect 245834 228905 300982 228933
rect 245834 228893 245840 228905
rect 300976 228893 300982 228905
rect 301034 228893 301040 228945
rect 317968 228893 317974 228945
rect 318026 228933 318032 228945
rect 445936 228933 445942 228945
rect 318026 228905 445942 228933
rect 318026 228893 318032 228905
rect 445936 228893 445942 228905
rect 445994 228893 446000 228945
rect 449296 228893 449302 228945
rect 449354 228933 449360 228945
rect 466384 228933 466390 228945
rect 449354 228905 466390 228933
rect 449354 228893 449360 228905
rect 466384 228893 466390 228905
rect 466442 228893 466448 228945
rect 246160 228819 246166 228871
rect 246218 228859 246224 228871
rect 298672 228859 298678 228871
rect 246218 228831 298678 228859
rect 246218 228819 246224 228831
rect 298672 228819 298678 228831
rect 298730 228819 298736 228871
rect 314896 228819 314902 228871
rect 314954 228859 314960 228871
rect 439984 228859 439990 228871
rect 314954 228831 439990 228859
rect 314954 228819 314960 228831
rect 439984 228819 439990 228831
rect 440042 228819 440048 228871
rect 242512 228745 242518 228797
rect 242570 228785 242576 228797
rect 294928 228785 294934 228797
rect 242570 228757 294934 228785
rect 242570 228745 242576 228757
rect 294928 228745 294934 228757
rect 294986 228745 294992 228797
rect 308944 228745 308950 228797
rect 309002 228785 309008 228797
rect 427792 228785 427798 228797
rect 309002 228757 427798 228785
rect 309002 228745 309008 228757
rect 427792 228745 427798 228757
rect 427850 228745 427856 228797
rect 428272 228745 428278 228797
rect 428330 228785 428336 228797
rect 547888 228785 547894 228797
rect 428330 228757 547894 228785
rect 428330 228745 428336 228757
rect 547888 228745 547894 228757
rect 547946 228745 547952 228797
rect 241648 228671 241654 228723
rect 241706 228711 241712 228723
rect 289744 228711 289750 228723
rect 241706 228683 289750 228711
rect 241706 228671 241712 228683
rect 289744 228671 289750 228683
rect 289802 228671 289808 228723
rect 306160 228671 306166 228723
rect 306218 228711 306224 228723
rect 306218 228683 309278 228711
rect 306218 228671 306224 228683
rect 230320 228597 230326 228649
rect 230378 228637 230384 228649
rect 269296 228637 269302 228649
rect 230378 228609 269302 228637
rect 230378 228597 230384 228609
rect 269296 228597 269302 228609
rect 269354 228597 269360 228649
rect 269392 228597 269398 228649
rect 269450 228637 269456 228649
rect 307696 228637 307702 228649
rect 269450 228609 307702 228637
rect 269450 228597 269456 228609
rect 307696 228597 307702 228609
rect 307754 228597 307760 228649
rect 309250 228637 309278 228683
rect 309328 228671 309334 228723
rect 309386 228711 309392 228723
rect 425584 228711 425590 228723
rect 309386 228683 425590 228711
rect 309386 228671 309392 228683
rect 425584 228671 425590 228683
rect 425642 228671 425648 228723
rect 432016 228671 432022 228723
rect 432074 228711 432080 228723
rect 529744 228711 529750 228723
rect 432074 228683 529750 228711
rect 432074 228671 432080 228683
rect 529744 228671 529750 228683
rect 529802 228671 529808 228723
rect 421840 228637 421846 228649
rect 309250 228609 421846 228637
rect 421840 228597 421846 228609
rect 421898 228597 421904 228649
rect 434896 228597 434902 228649
rect 434954 228637 434960 228649
rect 454288 228637 454294 228649
rect 434954 228609 454294 228637
rect 434954 228597 434960 228609
rect 454288 228597 454294 228609
rect 454346 228597 454352 228649
rect 190192 228523 190198 228575
rect 190250 228563 190256 228575
rect 192304 228563 192310 228575
rect 190250 228535 192310 228563
rect 190250 228523 190256 228535
rect 192304 228523 192310 228535
rect 192362 228523 192368 228575
rect 228784 228523 228790 228575
rect 228842 228563 228848 228575
rect 266224 228563 266230 228575
rect 228842 228535 266230 228563
rect 228842 228523 228848 228535
rect 266224 228523 266230 228535
rect 266282 228523 266288 228575
rect 266320 228523 266326 228575
rect 266378 228563 266384 228575
rect 301744 228563 301750 228575
rect 266378 228535 301750 228563
rect 266378 228523 266384 228535
rect 301744 228523 301750 228535
rect 301802 228523 301808 228575
rect 304432 228523 304438 228575
rect 304490 228563 304496 228575
rect 418768 228563 418774 228575
rect 304490 228535 418774 228563
rect 304490 228523 304496 228535
rect 418768 228523 418774 228535
rect 418826 228523 418832 228575
rect 455056 228523 455062 228575
rect 455114 228563 455120 228575
rect 456496 228563 456502 228575
rect 455114 228535 456502 228563
rect 455114 228523 455120 228535
rect 456496 228523 456502 228535
rect 456554 228523 456560 228575
rect 535792 228523 535798 228575
rect 535850 228563 535856 228575
rect 538000 228563 538006 228575
rect 535850 228535 538006 228563
rect 535850 228523 535856 228535
rect 538000 228523 538006 228535
rect 538058 228523 538064 228575
rect 544336 228523 544342 228575
rect 544394 228563 544400 228575
rect 547120 228563 547126 228575
rect 544394 228535 547126 228563
rect 544394 228523 544400 228535
rect 547120 228523 547126 228535
rect 547178 228523 547184 228575
rect 556144 228523 556150 228575
rect 556202 228563 556208 228575
rect 557680 228563 557686 228575
rect 556202 228535 557686 228563
rect 556202 228523 556208 228535
rect 557680 228523 557686 228535
rect 557738 228523 557744 228575
rect 567376 228523 567382 228575
rect 567434 228563 567440 228575
rect 569008 228563 569014 228575
rect 567434 228535 569014 228563
rect 567434 228523 567440 228535
rect 569008 228523 569014 228535
rect 569066 228523 569072 228575
rect 224368 228449 224374 228501
rect 224426 228489 224432 228501
rect 258736 228489 258742 228501
rect 224426 228461 258742 228489
rect 224426 228449 224432 228461
rect 258736 228449 258742 228461
rect 258794 228449 258800 228501
rect 260464 228449 260470 228501
rect 260522 228489 260528 228501
rect 286672 228489 286678 228501
rect 260522 228461 286678 228489
rect 260522 228449 260528 228461
rect 286672 228449 286678 228461
rect 286730 228449 286736 228501
rect 289360 228449 289366 228501
rect 289418 228489 289424 228501
rect 380080 228489 380086 228501
rect 289418 228461 380086 228489
rect 289418 228449 289424 228461
rect 380080 228449 380086 228461
rect 380138 228449 380144 228501
rect 403312 228449 403318 228501
rect 403370 228489 403376 228501
rect 517648 228489 517654 228501
rect 403370 228461 517654 228489
rect 403370 228449 403376 228461
rect 517648 228449 517654 228461
rect 517706 228449 517712 228501
rect 264880 228375 264886 228427
rect 264938 228415 264944 228427
rect 295696 228415 295702 228427
rect 264938 228387 295702 228415
rect 264938 228375 264944 228387
rect 295696 228375 295702 228387
rect 295754 228375 295760 228427
rect 303472 228375 303478 228427
rect 303530 228415 303536 228427
rect 413488 228415 413494 228427
rect 303530 228387 413494 228415
rect 303530 228375 303536 228387
rect 413488 228375 413494 228387
rect 413546 228375 413552 228427
rect 535792 228375 535798 228427
rect 535850 228415 535856 228427
rect 537904 228415 537910 228427
rect 535850 228387 537910 228415
rect 535850 228375 535856 228387
rect 537904 228375 537910 228387
rect 537962 228375 537968 228427
rect 260848 228301 260854 228353
rect 260906 228341 260912 228353
rect 292624 228341 292630 228353
rect 260906 228313 292630 228341
rect 260906 228301 260912 228313
rect 292624 228301 292630 228313
rect 292682 228301 292688 228353
rect 293872 228301 293878 228353
rect 293930 228341 293936 228353
rect 381712 228341 381718 228353
rect 293930 228313 381718 228341
rect 293930 228301 293936 228313
rect 381712 228301 381718 228313
rect 381770 228301 381776 228353
rect 393520 228301 393526 228353
rect 393578 228341 393584 228353
rect 476944 228341 476950 228353
rect 393578 228313 476950 228341
rect 393578 228301 393584 228313
rect 476944 228301 476950 228313
rect 477002 228301 477008 228353
rect 250576 228227 250582 228279
rect 250634 228267 250640 228279
rect 276496 228267 276502 228279
rect 250634 228239 276502 228267
rect 250634 228227 250640 228239
rect 276496 228227 276502 228239
rect 276554 228227 276560 228279
rect 288016 228227 288022 228279
rect 288074 228267 288080 228279
rect 328912 228267 328918 228279
rect 288074 228239 328918 228267
rect 288074 228227 288080 228239
rect 328912 228227 328918 228239
rect 328970 228227 328976 228279
rect 357712 228227 357718 228279
rect 357770 228267 357776 228279
rect 359920 228267 359926 228279
rect 357770 228239 359926 228267
rect 357770 228227 357776 228239
rect 359920 228227 359926 228239
rect 359978 228227 359984 228279
rect 270832 228153 270838 228205
rect 270890 228193 270896 228205
rect 313840 228193 313846 228205
rect 270890 228165 313846 228193
rect 270890 228153 270896 228165
rect 313840 228153 313846 228165
rect 313898 228153 313904 228205
rect 392368 228193 392374 228205
rect 313954 228165 392374 228193
rect 258064 228079 258070 228131
rect 258122 228119 258128 228131
rect 280624 228119 280630 228131
rect 258122 228091 280630 228119
rect 258122 228079 258128 228091
rect 280624 228079 280630 228091
rect 280682 228079 280688 228131
rect 311056 228079 311062 228131
rect 311114 228119 311120 228131
rect 313954 228119 313982 228165
rect 392368 228153 392374 228165
rect 392426 228153 392432 228205
rect 396400 228153 396406 228205
rect 396458 228193 396464 228205
rect 437680 228193 437686 228205
rect 396458 228165 437686 228193
rect 396458 228153 396464 228165
rect 437680 228153 437686 228165
rect 437738 228153 437744 228205
rect 311114 228091 313982 228119
rect 311114 228079 311120 228091
rect 314032 228079 314038 228131
rect 314090 228119 314096 228131
rect 383248 228119 383254 228131
rect 314090 228091 383254 228119
rect 314090 228079 314096 228091
rect 383248 228079 383254 228091
rect 383306 228079 383312 228131
rect 390352 228079 390358 228131
rect 390410 228119 390416 228131
rect 461872 228119 461878 228131
rect 390410 228091 461878 228119
rect 390410 228079 390416 228091
rect 461872 228079 461878 228091
rect 461930 228079 461936 228131
rect 290992 228005 290998 228057
rect 291050 228045 291056 228057
rect 341008 228045 341014 228057
rect 291050 228017 341014 228045
rect 291050 228005 291056 228017
rect 341008 228005 341014 228017
rect 341066 228005 341072 228057
rect 344176 228005 344182 228057
rect 344234 228045 344240 228057
rect 412720 228045 412726 228057
rect 344234 228017 412726 228045
rect 344234 228005 344240 228017
rect 412720 228005 412726 228017
rect 412778 228005 412784 228057
rect 281872 227931 281878 227983
rect 281930 227971 281936 227983
rect 325840 227971 325846 227983
rect 281930 227943 325846 227971
rect 281930 227931 281936 227943
rect 325840 227931 325846 227943
rect 325898 227931 325904 227983
rect 341392 227931 341398 227983
rect 341450 227971 341456 227983
rect 398320 227971 398326 227983
rect 341450 227943 398326 227971
rect 341450 227931 341456 227943
rect 398320 227931 398326 227943
rect 398378 227931 398384 227983
rect 250192 227857 250198 227909
rect 250250 227897 250256 227909
rect 310000 227897 310006 227909
rect 250250 227869 310006 227897
rect 250250 227857 250256 227869
rect 310000 227857 310006 227869
rect 310058 227857 310064 227909
rect 310096 227857 310102 227909
rect 310154 227897 310160 227909
rect 359152 227897 359158 227909
rect 310154 227869 359158 227897
rect 310154 227857 310160 227869
rect 359152 227857 359158 227869
rect 359210 227857 359216 227909
rect 293776 227783 293782 227835
rect 293834 227823 293840 227835
rect 343984 227823 343990 227835
rect 293834 227795 343990 227823
rect 293834 227783 293840 227795
rect 343984 227783 343990 227795
rect 344042 227783 344048 227835
rect 301264 227709 301270 227761
rect 301322 227749 301328 227761
rect 350032 227749 350038 227761
rect 301322 227721 350038 227749
rect 301322 227709 301328 227721
rect 350032 227709 350038 227721
rect 350090 227709 350096 227761
rect 319600 227635 319606 227687
rect 319658 227675 319664 227687
rect 319658 227647 320030 227675
rect 319658 227635 319664 227647
rect 149392 227561 149398 227613
rect 149450 227601 149456 227613
rect 182896 227601 182902 227613
rect 149450 227573 182902 227601
rect 149450 227561 149456 227573
rect 182896 227561 182902 227573
rect 182954 227561 182960 227613
rect 279280 227561 279286 227613
rect 279338 227601 279344 227613
rect 319888 227601 319894 227613
rect 279338 227573 319894 227601
rect 279338 227561 279344 227573
rect 319888 227561 319894 227573
rect 319946 227561 319952 227613
rect 320002 227601 320030 227647
rect 326800 227635 326806 227687
rect 326858 227675 326864 227687
rect 353104 227675 353110 227687
rect 326858 227647 353110 227675
rect 326858 227635 326864 227647
rect 353104 227635 353110 227647
rect 353162 227635 353168 227687
rect 403696 227601 403702 227613
rect 320002 227573 403702 227601
rect 403696 227561 403702 227573
rect 403754 227561 403760 227613
rect 418288 227561 418294 227613
rect 418346 227601 418352 227613
rect 433168 227601 433174 227613
rect 418346 227573 433174 227601
rect 418346 227561 418352 227573
rect 433168 227561 433174 227573
rect 433226 227561 433232 227613
rect 187120 227487 187126 227539
rect 187178 227527 187184 227539
rect 190768 227527 190774 227539
rect 187178 227499 190774 227527
rect 187178 227487 187184 227499
rect 190768 227487 190774 227499
rect 190826 227487 190832 227539
rect 213808 227487 213814 227539
rect 213866 227527 213872 227539
rect 237520 227527 237526 227539
rect 213866 227499 237526 227527
rect 213866 227487 213872 227499
rect 237520 227487 237526 227499
rect 237578 227487 237584 227539
rect 249328 227487 249334 227539
rect 249386 227527 249392 227539
rect 306256 227527 306262 227539
rect 249386 227499 306262 227527
rect 249386 227487 249392 227499
rect 306256 227487 306262 227499
rect 306314 227487 306320 227539
rect 311344 227487 311350 227539
rect 311402 227527 311408 227539
rect 375760 227527 375766 227539
rect 311402 227499 375766 227527
rect 311402 227487 311408 227499
rect 375760 227487 375766 227499
rect 375818 227487 375824 227539
rect 390064 227487 390070 227539
rect 390122 227527 390128 227539
rect 588592 227527 588598 227539
rect 390122 227499 588598 227527
rect 390122 227487 390128 227499
rect 588592 227487 588598 227499
rect 588650 227487 588656 227539
rect 596176 227487 596182 227539
rect 596234 227527 596240 227539
rect 616624 227527 616630 227539
rect 596234 227499 616630 227527
rect 596234 227487 596240 227499
rect 616624 227487 616630 227499
rect 616682 227487 616688 227539
rect 629296 227487 629302 227539
rect 629354 227527 629360 227539
rect 634000 227527 634006 227539
rect 629354 227499 634006 227527
rect 629354 227487 629360 227499
rect 634000 227487 634006 227499
rect 634058 227487 634064 227539
rect 216112 227413 216118 227465
rect 216170 227453 216176 227465
rect 239824 227453 239830 227465
rect 216170 227425 239830 227453
rect 216170 227413 216176 227425
rect 239824 227413 239830 227425
rect 239882 227413 239888 227465
rect 253840 227413 253846 227465
rect 253898 227453 253904 227465
rect 315376 227453 315382 227465
rect 253898 227425 315382 227453
rect 253898 227413 253904 227425
rect 315376 227413 315382 227425
rect 315434 227413 315440 227465
rect 318256 227413 318262 227465
rect 318314 227453 318320 227465
rect 381808 227453 381814 227465
rect 318314 227425 381814 227453
rect 318314 227413 318320 227425
rect 381808 227413 381814 227425
rect 381866 227413 381872 227465
rect 390832 227413 390838 227465
rect 390890 227453 390896 227465
rect 590128 227453 590134 227465
rect 390890 227425 590134 227453
rect 390890 227413 390896 227425
rect 590128 227413 590134 227425
rect 590186 227413 590192 227465
rect 593008 227413 593014 227465
rect 593066 227453 593072 227465
rect 611248 227453 611254 227465
rect 593066 227425 611254 227453
rect 593066 227413 593072 227425
rect 611248 227413 611254 227425
rect 611306 227413 611312 227465
rect 215728 227339 215734 227391
rect 215786 227379 215792 227391
rect 238384 227379 238390 227391
rect 215786 227351 238390 227379
rect 215786 227339 215792 227351
rect 238384 227339 238390 227351
rect 238442 227339 238448 227391
rect 284656 227339 284662 227391
rect 284714 227379 284720 227391
rect 306640 227379 306646 227391
rect 284714 227351 306646 227379
rect 284714 227339 284720 227351
rect 306640 227339 306646 227351
rect 306698 227339 306704 227391
rect 311248 227339 311254 227391
rect 311306 227379 311312 227391
rect 384016 227379 384022 227391
rect 311306 227351 384022 227379
rect 311306 227339 311312 227351
rect 384016 227339 384022 227351
rect 384074 227339 384080 227391
rect 388240 227339 388246 227391
rect 388298 227379 388304 227391
rect 585616 227379 585622 227391
rect 388298 227351 585622 227379
rect 388298 227339 388304 227351
rect 585616 227339 585622 227351
rect 585674 227339 585680 227391
rect 595888 227339 595894 227391
rect 595946 227379 595952 227391
rect 614320 227379 614326 227391
rect 595946 227351 614326 227379
rect 595946 227339 595952 227351
rect 614320 227339 614326 227351
rect 614378 227339 614384 227391
rect 274672 227265 274678 227317
rect 274730 227305 274736 227317
rect 348592 227305 348598 227317
rect 274730 227277 348598 227305
rect 274730 227265 274736 227277
rect 348592 227265 348598 227277
rect 348650 227265 348656 227317
rect 392272 227265 392278 227317
rect 392330 227305 392336 227317
rect 593104 227305 593110 227317
rect 392330 227277 593110 227305
rect 392330 227265 392336 227277
rect 593104 227265 593110 227277
rect 593162 227265 593168 227317
rect 597424 227265 597430 227317
rect 597482 227305 597488 227317
rect 619600 227305 619606 227317
rect 597482 227277 619606 227305
rect 597482 227265 597488 227277
rect 619600 227265 619606 227277
rect 619658 227265 619664 227317
rect 220336 227191 220342 227243
rect 220394 227231 220400 227243
rect 247408 227231 247414 227243
rect 220394 227203 247414 227231
rect 220394 227191 220400 227203
rect 247408 227191 247414 227203
rect 247466 227191 247472 227243
rect 247696 227191 247702 227243
rect 247754 227231 247760 227243
rect 257968 227231 257974 227243
rect 247754 227203 257974 227231
rect 247754 227191 247760 227203
rect 257968 227191 257974 227203
rect 258026 227191 258032 227243
rect 271984 227191 271990 227243
rect 272042 227231 272048 227243
rect 351568 227231 351574 227243
rect 272042 227203 351574 227231
rect 272042 227191 272048 227203
rect 351568 227191 351574 227203
rect 351626 227191 351632 227243
rect 603472 227191 603478 227243
rect 603530 227231 603536 227243
rect 636208 227231 636214 227243
rect 603530 227203 636214 227231
rect 603530 227191 603536 227203
rect 636208 227191 636214 227203
rect 636266 227191 636272 227243
rect 219472 227117 219478 227169
rect 219530 227157 219536 227169
rect 245872 227157 245878 227169
rect 219530 227129 245878 227157
rect 219530 227117 219536 227129
rect 245872 227117 245878 227129
rect 245930 227117 245936 227169
rect 263728 227117 263734 227169
rect 263786 227157 263792 227169
rect 288112 227157 288118 227169
rect 263786 227129 288118 227157
rect 263786 227117 263792 227129
rect 288112 227117 288118 227129
rect 288170 227117 288176 227169
rect 289264 227117 289270 227169
rect 289322 227157 289328 227169
rect 369616 227157 369622 227169
rect 289322 227129 369622 227157
rect 289322 227117 289328 227129
rect 369616 227117 369622 227129
rect 369674 227117 369680 227169
rect 388144 227117 388150 227169
rect 388202 227157 388208 227169
rect 584848 227157 584854 227169
rect 388202 227129 584854 227157
rect 388202 227117 388208 227129
rect 584848 227117 584854 227129
rect 584906 227117 584912 227169
rect 606352 227117 606358 227169
rect 606410 227157 606416 227169
rect 638512 227157 638518 227169
rect 606410 227129 638518 227157
rect 606410 227117 606416 227129
rect 638512 227117 638518 227129
rect 638570 227117 638576 227169
rect 238768 227043 238774 227095
rect 238826 227083 238832 227095
rect 254896 227083 254902 227095
rect 238826 227055 254902 227083
rect 238826 227043 238832 227055
rect 254896 227043 254902 227055
rect 254954 227043 254960 227095
rect 259024 227043 259030 227095
rect 259082 227083 259088 227095
rect 269968 227083 269974 227095
rect 259082 227055 269974 227083
rect 259082 227043 259088 227055
rect 269968 227043 269974 227055
rect 270026 227043 270032 227095
rect 275248 227043 275254 227095
rect 275306 227083 275312 227095
rect 357616 227083 357622 227095
rect 275306 227055 357622 227083
rect 275306 227043 275312 227055
rect 357616 227043 357622 227055
rect 357674 227043 357680 227095
rect 392656 227043 392662 227095
rect 392714 227083 392720 227095
rect 593968 227083 593974 227095
rect 392714 227055 593974 227083
rect 392714 227043 392720 227055
rect 593968 227043 593974 227055
rect 594026 227043 594032 227095
rect 599056 227043 599062 227095
rect 599114 227083 599120 227095
rect 633136 227083 633142 227095
rect 599114 227055 633142 227083
rect 599114 227043 599120 227055
rect 633136 227043 633142 227055
rect 633194 227043 633200 227095
rect 212368 226969 212374 227021
rect 212426 227009 212432 227021
rect 234544 227009 234550 227021
rect 212426 226981 234550 227009
rect 212426 226969 212432 226981
rect 234544 226969 234550 226981
rect 234602 226969 234608 227021
rect 236368 226969 236374 227021
rect 236426 227009 236432 227021
rect 264016 227009 264022 227021
rect 236426 226981 264022 227009
rect 236426 226969 236432 226981
rect 264016 226969 264022 226981
rect 264074 226969 264080 227021
rect 276688 226969 276694 227021
rect 276746 227009 276752 227021
rect 360592 227009 360598 227021
rect 276746 226981 360598 227009
rect 276746 226969 276752 226981
rect 360592 226969 360598 226981
rect 360650 226969 360656 227021
rect 391216 226969 391222 227021
rect 391274 227009 391280 227021
rect 590896 227009 590902 227021
rect 391274 226981 590902 227009
rect 391274 226969 391280 226981
rect 590896 226969 590902 226981
rect 590954 226969 590960 227021
rect 603664 227009 603670 227021
rect 599026 226981 603670 227009
rect 221680 226895 221686 226947
rect 221738 226935 221744 226947
rect 250384 226935 250390 226947
rect 221738 226907 250390 226935
rect 221738 226895 221744 226907
rect 250384 226895 250390 226907
rect 250442 226895 250448 226947
rect 253552 226895 253558 226947
rect 253610 226935 253616 226947
rect 266992 226935 266998 226947
rect 253610 226907 266998 226935
rect 253610 226895 253616 226907
rect 266992 226895 266998 226907
rect 267050 226895 267056 226947
rect 273424 226895 273430 226947
rect 273482 226935 273488 226947
rect 354544 226935 354550 226947
rect 273482 226907 354550 226935
rect 273482 226895 273488 226907
rect 354544 226895 354550 226907
rect 354602 226895 354608 226947
rect 359824 226895 359830 226947
rect 359882 226935 359888 226947
rect 393136 226935 393142 226947
rect 359882 226907 393142 226935
rect 359882 226895 359888 226907
rect 393136 226895 393142 226907
rect 393194 226895 393200 226947
rect 395536 226895 395542 226947
rect 395594 226935 395600 226947
rect 395594 226907 397454 226935
rect 395594 226895 395600 226907
rect 224848 226821 224854 226873
rect 224906 226861 224912 226873
rect 256432 226861 256438 226873
rect 224906 226833 256438 226861
rect 224906 226821 224912 226833
rect 256432 226821 256438 226833
rect 256490 226821 256496 226873
rect 277936 226821 277942 226873
rect 277994 226861 278000 226873
rect 363760 226861 363766 226873
rect 277994 226833 363766 226861
rect 277994 226821 278000 226833
rect 363760 226821 363766 226833
rect 363818 226821 363824 226873
rect 364240 226821 364246 226873
rect 364298 226861 364304 226873
rect 396112 226861 396118 226873
rect 364298 226833 396118 226861
rect 364298 226821 364304 226833
rect 396112 226821 396118 226833
rect 396170 226821 396176 226873
rect 397426 226861 397454 226907
rect 397648 226895 397654 226947
rect 397706 226935 397712 226947
rect 599026 226935 599054 226981
rect 603664 226969 603670 226981
rect 603722 226969 603728 227021
rect 606256 226969 606262 227021
rect 606314 227009 606320 227021
rect 639184 227009 639190 227021
rect 606314 226981 639190 227009
rect 606314 226969 606320 226981
rect 639184 226969 639190 226981
rect 639242 226969 639248 227021
rect 397706 226907 599054 226935
rect 397706 226895 397712 226907
rect 603376 226895 603382 226947
rect 603434 226935 603440 226947
rect 636880 226935 636886 226947
rect 603434 226907 636886 226935
rect 603434 226895 603440 226907
rect 636880 226895 636886 226907
rect 636938 226895 636944 226947
rect 599152 226861 599158 226873
rect 397426 226833 599158 226861
rect 599152 226821 599158 226833
rect 599210 226821 599216 226873
rect 600400 226821 600406 226873
rect 600458 226861 600464 226873
rect 634672 226861 634678 226873
rect 600458 226833 634678 226861
rect 600458 226821 600464 226833
rect 634672 226821 634678 226833
rect 634730 226821 634736 226873
rect 223312 226747 223318 226799
rect 223370 226787 223376 226799
rect 253456 226787 253462 226799
rect 223370 226759 253462 226787
rect 223370 226747 223376 226759
rect 253456 226747 253462 226759
rect 253514 226747 253520 226799
rect 279760 226747 279766 226799
rect 279818 226787 279824 226799
rect 366736 226787 366742 226799
rect 279818 226759 366742 226787
rect 279818 226747 279824 226759
rect 366736 226747 366742 226759
rect 366794 226747 366800 226799
rect 374608 226747 374614 226799
rect 374666 226787 374672 226799
rect 391504 226787 391510 226799
rect 374666 226759 391510 226787
rect 374666 226747 374672 226759
rect 391504 226747 391510 226759
rect 391562 226747 391568 226799
rect 397168 226747 397174 226799
rect 397226 226787 397232 226799
rect 602992 226787 602998 226799
rect 397226 226759 602998 226787
rect 397226 226747 397232 226759
rect 602992 226747 602998 226759
rect 603050 226747 603056 226799
rect 603280 226747 603286 226799
rect 603338 226787 603344 226799
rect 637744 226787 637750 226799
rect 603338 226759 637750 226787
rect 603338 226747 603344 226759
rect 637744 226747 637750 226759
rect 637802 226747 637808 226799
rect 226576 226673 226582 226725
rect 226634 226713 226640 226725
rect 259408 226713 259414 226725
rect 226634 226685 259414 226713
rect 226634 226673 226640 226685
rect 259408 226673 259414 226685
rect 259466 226673 259472 226725
rect 271888 226673 271894 226725
rect 271946 226713 271952 226725
rect 336400 226713 336406 226725
rect 271946 226685 336406 226713
rect 271946 226673 271952 226685
rect 336400 226673 336406 226685
rect 336458 226673 336464 226725
rect 371632 226673 371638 226725
rect 371690 226713 371696 226725
rect 393808 226713 393814 226725
rect 371690 226685 393814 226713
rect 371690 226673 371696 226685
rect 393808 226673 393814 226685
rect 393866 226673 393872 226725
rect 400816 226673 400822 226725
rect 400874 226713 400880 226725
rect 609808 226713 609814 226725
rect 400874 226685 609814 226713
rect 400874 226673 400880 226685
rect 609808 226673 609814 226685
rect 609866 226673 609872 226725
rect 227920 226599 227926 226651
rect 227978 226639 227984 226651
rect 262480 226639 262486 226651
rect 227978 226611 262486 226639
rect 227978 226599 227984 226611
rect 262480 226599 262486 226611
rect 262538 226599 262544 226651
rect 264688 226599 264694 226651
rect 264746 226639 264752 226651
rect 276112 226639 276118 226651
rect 264746 226611 276118 226639
rect 264746 226599 264752 226611
rect 276112 226599 276118 226611
rect 276170 226599 276176 226651
rect 285712 226599 285718 226651
rect 285770 226639 285776 226651
rect 378736 226639 378742 226651
rect 285770 226611 378742 226639
rect 285770 226599 285776 226611
rect 378736 226599 378742 226611
rect 378794 226599 378800 226651
rect 381712 226599 381718 226651
rect 381770 226639 381776 226651
rect 397648 226639 397654 226651
rect 381770 226611 397654 226639
rect 381770 226599 381776 226611
rect 397648 226599 397654 226611
rect 397706 226599 397712 226651
rect 588880 226599 588886 226651
rect 588938 226639 588944 226651
rect 600784 226639 600790 226651
rect 588938 226611 600790 226639
rect 588938 226599 588944 226611
rect 600784 226599 600790 226611
rect 600842 226599 600848 226651
rect 606160 226599 606166 226651
rect 606218 226639 606224 226651
rect 639952 226639 639958 226651
rect 606218 226611 639958 226639
rect 606218 226599 606224 226611
rect 639952 226599 639958 226611
rect 640010 226599 640016 226651
rect 231088 226525 231094 226577
rect 231146 226565 231152 226577
rect 268528 226565 268534 226577
rect 231146 226537 268534 226565
rect 231146 226525 231152 226537
rect 268528 226525 268534 226537
rect 268586 226525 268592 226577
rect 270928 226525 270934 226577
rect 270986 226565 270992 226577
rect 294256 226565 294262 226577
rect 270986 226537 294262 226565
rect 270986 226525 270992 226537
rect 294256 226525 294262 226537
rect 294314 226525 294320 226577
rect 297424 226525 297430 226577
rect 297482 226565 297488 226577
rect 390064 226565 390070 226577
rect 297482 226537 390070 226565
rect 297482 226525 297488 226537
rect 390064 226525 390070 226537
rect 390122 226525 390128 226577
rect 402160 226525 402166 226577
rect 402218 226565 402224 226577
rect 612784 226565 612790 226577
rect 402218 226537 612790 226565
rect 402218 226525 402224 226537
rect 612784 226525 612790 226537
rect 612842 226525 612848 226577
rect 229552 226451 229558 226503
rect 229610 226491 229616 226503
rect 265552 226491 265558 226503
rect 229610 226463 265558 226491
rect 229610 226451 229616 226463
rect 265552 226451 265558 226463
rect 265610 226451 265616 226503
rect 288496 226451 288502 226503
rect 288554 226491 288560 226503
rect 384784 226491 384790 226503
rect 288554 226463 384790 226491
rect 288554 226451 288560 226463
rect 384784 226451 384790 226463
rect 384842 226451 384848 226503
rect 385744 226451 385750 226503
rect 385802 226491 385808 226503
rect 392080 226491 392086 226503
rect 385802 226463 392086 226491
rect 385802 226451 385808 226463
rect 392080 226451 392086 226463
rect 392138 226451 392144 226503
rect 404368 226451 404374 226503
rect 404426 226491 404432 226503
rect 617296 226491 617302 226503
rect 404426 226463 617302 226491
rect 404426 226451 404432 226463
rect 617296 226451 617302 226463
rect 617354 226451 617360 226503
rect 232528 226377 232534 226429
rect 232586 226417 232592 226429
rect 271600 226417 271606 226429
rect 232586 226389 271606 226417
rect 232586 226377 232592 226389
rect 271600 226377 271606 226389
rect 271658 226377 271664 226429
rect 291568 226377 291574 226429
rect 291626 226417 291632 226429
rect 291626 226389 296654 226417
rect 291626 226377 291632 226389
rect 214576 226303 214582 226355
rect 214634 226343 214640 226355
rect 236848 226343 236854 226355
rect 214634 226315 236854 226343
rect 214634 226303 214640 226315
rect 236848 226303 236854 226315
rect 236906 226303 236912 226355
rect 241744 226303 241750 226355
rect 241802 226343 241808 226355
rect 241802 226315 254846 226343
rect 241802 226303 241808 226315
rect 217840 226229 217846 226281
rect 217898 226269 217904 226281
rect 242896 226269 242902 226281
rect 217898 226241 242902 226269
rect 217898 226229 217904 226241
rect 242896 226229 242902 226241
rect 242954 226229 242960 226281
rect 215632 226155 215638 226207
rect 215690 226195 215696 226207
rect 240592 226195 240598 226207
rect 215690 226167 240598 226195
rect 215690 226155 215696 226167
rect 240592 226155 240598 226167
rect 240650 226155 240656 226207
rect 246544 226155 246550 226207
rect 246602 226195 246608 226207
rect 254818 226195 254846 226315
rect 254896 226303 254902 226355
rect 254954 226343 254960 226355
rect 285136 226343 285142 226355
rect 254954 226315 285142 226343
rect 254954 226303 254960 226315
rect 285136 226303 285142 226315
rect 285194 226303 285200 226355
rect 296626 226343 296654 226389
rect 306640 226377 306646 226429
rect 306698 226417 306704 226429
rect 378064 226417 378070 226429
rect 306698 226389 378070 226417
rect 306698 226377 306704 226389
rect 378064 226377 378070 226389
rect 378122 226377 378128 226429
rect 379984 226377 379990 226429
rect 380042 226417 380048 226429
rect 394576 226417 394582 226429
rect 380042 226389 394582 226417
rect 380042 226377 380048 226389
rect 394576 226377 394582 226389
rect 394634 226377 394640 226429
rect 402640 226377 402646 226429
rect 402698 226417 402704 226429
rect 613552 226417 613558 226429
rect 402698 226389 613558 226417
rect 402698 226377 402704 226389
rect 613552 226377 613558 226389
rect 613610 226377 613616 226429
rect 629200 226377 629206 226429
rect 629258 226417 629264 226429
rect 635440 226417 635446 226429
rect 629258 226389 635446 226417
rect 629258 226377 629264 226389
rect 635440 226377 635446 226389
rect 635498 226377 635504 226429
rect 390832 226343 390838 226355
rect 296626 226315 390838 226343
rect 390832 226303 390838 226315
rect 390890 226303 390896 226355
rect 404944 226303 404950 226355
rect 405002 226343 405008 226355
rect 618064 226343 618070 226355
rect 405002 226315 618070 226343
rect 405002 226303 405008 226315
rect 618064 226303 618070 226315
rect 618122 226303 618128 226355
rect 254992 226229 254998 226281
rect 255050 226269 255056 226281
rect 297232 226269 297238 226281
rect 255050 226241 297238 226269
rect 255050 226229 255056 226241
rect 297232 226229 297238 226241
rect 297290 226229 297296 226281
rect 297616 226229 297622 226281
rect 297674 226269 297680 226281
rect 402832 226269 402838 226281
rect 297674 226241 402838 226269
rect 297674 226229 297680 226241
rect 402832 226229 402838 226241
rect 402890 226229 402896 226281
rect 407728 226229 407734 226281
rect 407786 226269 407792 226281
rect 624112 226269 624118 226281
rect 407786 226241 624118 226269
rect 407786 226229 407792 226241
rect 624112 226229 624118 226241
rect 624170 226229 624176 226281
rect 291184 226195 291190 226207
rect 246602 226167 254750 226195
rect 254818 226167 291190 226195
rect 246602 226155 246608 226167
rect 151120 226081 151126 226133
rect 151178 226121 151184 226133
rect 187120 226121 187126 226133
rect 151178 226093 187126 226121
rect 151178 226081 151184 226093
rect 187120 226081 187126 226093
rect 187178 226081 187184 226133
rect 218320 226081 218326 226133
rect 218378 226121 218384 226133
rect 246640 226121 246646 226133
rect 218378 226093 246646 226121
rect 218378 226081 218384 226093
rect 246640 226081 246646 226093
rect 246698 226081 246704 226133
rect 254722 226121 254750 226167
rect 291184 226155 291190 226167
rect 291242 226155 291248 226207
rect 300688 226155 300694 226207
rect 300746 226195 300752 226207
rect 408976 226195 408982 226207
rect 300746 226167 408982 226195
rect 300746 226155 300752 226167
rect 408976 226155 408982 226167
rect 409034 226155 409040 226207
rect 300208 226121 300214 226133
rect 254722 226093 300214 226121
rect 300208 226081 300214 226093
rect 300266 226081 300272 226133
rect 301360 226081 301366 226133
rect 301418 226121 301424 226133
rect 411280 226121 411286 226133
rect 301418 226093 411286 226121
rect 301418 226081 301424 226093
rect 411280 226081 411286 226093
rect 411338 226081 411344 226133
rect 411376 226081 411382 226133
rect 411434 226121 411440 226133
rect 631696 226121 631702 226133
rect 411434 226093 631702 226121
rect 411434 226081 411440 226093
rect 631696 226081 631702 226093
rect 631754 226081 631760 226133
rect 213040 226007 213046 226059
rect 213098 226047 213104 226059
rect 233776 226047 233782 226059
rect 213098 226019 233782 226047
rect 213098 226007 213104 226019
rect 233776 226007 233782 226019
rect 233834 226007 233840 226059
rect 238960 226007 238966 226059
rect 239018 226047 239024 226059
rect 239018 226019 241406 226047
rect 239018 226007 239024 226019
rect 217456 225933 217462 225985
rect 217514 225973 217520 225985
rect 241264 225973 241270 225985
rect 217514 225945 241270 225973
rect 217514 225933 217520 225945
rect 241264 225933 241270 225945
rect 241322 225933 241328 225985
rect 241378 225973 241406 226019
rect 244816 226007 244822 226059
rect 244874 226047 244880 226059
rect 254992 226047 254998 226059
rect 244874 226019 254998 226047
rect 244874 226007 244880 226019
rect 254992 226007 254998 226019
rect 255050 226007 255056 226059
rect 257104 226007 257110 226059
rect 257162 226047 257168 226059
rect 257162 226019 267854 226047
rect 257162 226007 257168 226019
rect 261040 225973 261046 225985
rect 241378 225945 261046 225973
rect 261040 225933 261046 225945
rect 261098 225933 261104 225985
rect 267826 225973 267854 226019
rect 324496 226007 324502 226059
rect 324554 226047 324560 226059
rect 339472 226047 339478 226059
rect 324554 226019 339478 226047
rect 324554 226007 324560 226019
rect 339472 226007 339478 226019
rect 339530 226007 339536 226059
rect 341506 226019 387230 226047
rect 321328 225973 321334 225985
rect 267826 225945 321334 225973
rect 321328 225933 321334 225945
rect 321386 225933 321392 225985
rect 334288 225933 334294 225985
rect 334346 225973 334352 225985
rect 341506 225973 341534 226019
rect 334346 225945 341534 225973
rect 334346 225933 334352 225945
rect 345712 225933 345718 225985
rect 345770 225973 345776 225985
rect 386992 225973 386998 225985
rect 345770 225945 386998 225973
rect 345770 225933 345776 225945
rect 386992 225933 386998 225945
rect 387050 225933 387056 225985
rect 387202 225973 387230 226019
rect 387280 226007 387286 226059
rect 387338 226047 387344 226059
rect 582640 226047 582646 226059
rect 387338 226019 582646 226047
rect 387338 226007 387344 226019
rect 582640 226007 582646 226019
rect 582698 226007 582704 226059
rect 591472 226007 591478 226059
rect 591530 226047 591536 226059
rect 608272 226047 608278 226059
rect 591530 226019 608278 226047
rect 591530 226007 591536 226019
rect 608272 226007 608278 226019
rect 608330 226007 608336 226059
rect 387760 225973 387766 225985
rect 387202 225945 387766 225973
rect 387760 225933 387766 225945
rect 387818 225933 387824 225985
rect 388048 225933 388054 225985
rect 388106 225973 388112 225985
rect 584080 225973 584086 225985
rect 388106 225945 584086 225973
rect 388106 225933 388112 225945
rect 584080 225933 584086 225945
rect 584138 225933 584144 225985
rect 590416 225933 590422 225985
rect 590474 225973 590480 225985
rect 590474 225945 599054 225973
rect 590474 225933 590480 225945
rect 218800 225859 218806 225911
rect 218858 225899 218864 225911
rect 244336 225899 244342 225911
rect 218858 225871 244342 225899
rect 218858 225859 218864 225871
rect 244336 225859 244342 225871
rect 244394 225859 244400 225911
rect 244720 225859 244726 225911
rect 244778 225899 244784 225911
rect 254896 225899 254902 225911
rect 244778 225871 254902 225899
rect 244778 225859 244784 225871
rect 254896 225859 254902 225871
rect 254954 225859 254960 225911
rect 269008 225859 269014 225911
rect 269066 225899 269072 225911
rect 330448 225899 330454 225911
rect 269066 225871 330454 225899
rect 269066 225859 269072 225871
rect 330448 225859 330454 225871
rect 330506 225859 330512 225911
rect 331408 225859 331414 225911
rect 331466 225899 331472 225911
rect 345520 225899 345526 225911
rect 331466 225871 345526 225899
rect 331466 225859 331472 225871
rect 345520 225859 345526 225871
rect 345578 225859 345584 225911
rect 365680 225859 365686 225911
rect 365738 225899 365744 225911
rect 382672 225899 382678 225911
rect 365738 225871 382678 225899
rect 365738 225859 365744 225871
rect 382672 225859 382678 225871
rect 382730 225859 382736 225911
rect 382960 225859 382966 225911
rect 383018 225899 383024 225911
rect 388720 225899 388726 225911
rect 383018 225871 388726 225899
rect 383018 225859 383024 225871
rect 388720 225859 388726 225871
rect 388778 225859 388784 225911
rect 389488 225859 389494 225911
rect 389546 225899 389552 225911
rect 587152 225899 587158 225911
rect 389546 225871 587158 225899
rect 389546 225859 389552 225871
rect 587152 225859 587158 225871
rect 587210 225859 587216 225911
rect 588688 225859 588694 225911
rect 588746 225899 588752 225911
rect 598480 225899 598486 225911
rect 588746 225871 598486 225899
rect 588746 225859 588752 225871
rect 598480 225859 598486 225871
rect 598538 225859 598544 225911
rect 599026 225899 599054 225945
rect 605296 225899 605302 225911
rect 599026 225871 605302 225899
rect 605296 225859 605302 225871
rect 605354 225859 605360 225911
rect 217072 225785 217078 225837
rect 217130 225825 217136 225837
rect 243568 225825 243574 225837
rect 217130 225797 243574 225825
rect 217130 225785 217136 225797
rect 243568 225785 243574 225797
rect 243626 225785 243632 225837
rect 267760 225785 267766 225837
rect 267818 225825 267824 225837
rect 327376 225825 327382 225837
rect 267818 225797 327382 225825
rect 267818 225785 267824 225797
rect 327376 225785 327382 225797
rect 327434 225785 327440 225837
rect 368560 225785 368566 225837
rect 368618 225825 368624 225837
rect 374224 225825 374230 225837
rect 368618 225797 374230 225825
rect 368618 225785 368624 225797
rect 374224 225785 374230 225797
rect 374282 225785 374288 225837
rect 374416 225785 374422 225837
rect 374474 225825 374480 225837
rect 385552 225825 385558 225837
rect 374474 225797 385558 225825
rect 374474 225785 374480 225797
rect 385552 225785 385558 225797
rect 385610 225785 385616 225837
rect 386608 225785 386614 225837
rect 386666 225825 386672 225837
rect 386666 225797 392030 225825
rect 386666 225785 386672 225797
rect 285040 225711 285046 225763
rect 285098 225751 285104 225763
rect 342544 225751 342550 225763
rect 285098 225723 342550 225751
rect 285098 225711 285104 225723
rect 342544 225711 342550 225723
rect 342602 225711 342608 225763
rect 371344 225711 371350 225763
rect 371402 225751 371408 225763
rect 376432 225751 376438 225763
rect 371402 225723 376438 225751
rect 371402 225711 371408 225723
rect 376432 225711 376438 225723
rect 376490 225711 376496 225763
rect 380080 225711 380086 225763
rect 380138 225751 380144 225763
rect 388624 225751 388630 225763
rect 380138 225723 388630 225751
rect 380138 225711 380144 225723
rect 388624 225711 388630 225723
rect 388682 225711 388688 225763
rect 388720 225711 388726 225763
rect 388778 225751 388784 225763
rect 389296 225751 389302 225763
rect 388778 225723 389302 225751
rect 388778 225711 388784 225723
rect 389296 225711 389302 225723
rect 389354 225711 389360 225763
rect 392002 225751 392030 225797
rect 392080 225785 392086 225837
rect 392138 225825 392144 225837
rect 579568 225825 579574 225837
rect 392138 225797 579574 225825
rect 392138 225785 392144 225797
rect 579568 225785 579574 225797
rect 579626 225785 579632 225837
rect 581104 225751 581110 225763
rect 392002 225723 581110 225751
rect 581104 225711 581110 225723
rect 581162 225711 581168 225763
rect 588976 225711 588982 225763
rect 589034 225751 589040 225763
rect 602224 225751 602230 225763
rect 589034 225723 602230 225751
rect 589034 225711 589040 225723
rect 602224 225711 602230 225723
rect 602282 225711 602288 225763
rect 278224 225637 278230 225689
rect 278282 225677 278288 225689
rect 324400 225677 324406 225689
rect 278282 225649 324406 225677
rect 278282 225637 278288 225649
rect 324400 225637 324406 225649
rect 324458 225637 324464 225689
rect 339088 225637 339094 225689
rect 339146 225677 339152 225689
rect 396880 225677 396886 225689
rect 339146 225649 396886 225677
rect 339146 225637 339152 225649
rect 396880 225637 396886 225649
rect 396938 225637 396944 225689
rect 396976 225637 396982 225689
rect 397034 225677 397040 225689
rect 586384 225677 586390 225689
rect 397034 225649 586390 225677
rect 397034 225637 397040 225649
rect 586384 225637 586390 225649
rect 586442 225637 586448 225689
rect 273616 225563 273622 225615
rect 273674 225603 273680 225615
rect 309328 225603 309334 225615
rect 273674 225575 309334 225603
rect 273674 225563 273680 225575
rect 309328 225563 309334 225575
rect 309386 225563 309392 225615
rect 315760 225563 315766 225615
rect 315818 225603 315824 225615
rect 439120 225603 439126 225615
rect 315818 225575 439126 225603
rect 315818 225563 315824 225575
rect 439120 225563 439126 225575
rect 439178 225563 439184 225615
rect 265264 225489 265270 225541
rect 265322 225529 265328 225541
rect 279088 225529 279094 225541
rect 265322 225501 279094 225529
rect 265322 225489 265328 225501
rect 279088 225489 279094 225501
rect 279146 225489 279152 225541
rect 303184 225529 303190 225541
rect 287986 225501 303190 225529
rect 243952 225415 243958 225467
rect 244010 225455 244016 225467
rect 251920 225455 251926 225467
rect 244010 225427 251926 225455
rect 244010 225415 244016 225427
rect 251920 225415 251926 225427
rect 251978 225415 251984 225467
rect 262000 225415 262006 225467
rect 262058 225455 262064 225467
rect 273040 225455 273046 225467
rect 262058 225427 273046 225455
rect 262058 225415 262064 225427
rect 273040 225415 273046 225427
rect 273098 225415 273104 225467
rect 273712 225415 273718 225467
rect 273770 225455 273776 225467
rect 287986 225455 288014 225501
rect 303184 225489 303190 225501
rect 303242 225489 303248 225541
rect 309904 225489 309910 225541
rect 309962 225529 309968 225541
rect 427024 225529 427030 225541
rect 309962 225501 427030 225529
rect 309962 225489 309968 225501
rect 427024 225489 427030 225501
rect 427082 225489 427088 225541
rect 273770 225427 288014 225455
rect 273770 225415 273776 225427
rect 306736 225415 306742 225467
rect 306794 225455 306800 225467
rect 420976 225455 420982 225467
rect 306794 225427 420982 225455
rect 306794 225415 306800 225427
rect 420976 225415 420982 225427
rect 421034 225415 421040 225467
rect 241840 225341 241846 225393
rect 241898 225381 241904 225393
rect 248848 225381 248854 225393
rect 241898 225353 248854 225381
rect 241898 225341 241904 225353
rect 248848 225341 248854 225353
rect 248906 225341 248912 225393
rect 303856 225341 303862 225393
rect 303914 225381 303920 225393
rect 415024 225381 415030 225393
rect 303914 225353 415030 225381
rect 303914 225341 303920 225353
rect 415024 225341 415030 225353
rect 415082 225341 415088 225393
rect 302128 225267 302134 225319
rect 302186 225307 302192 225319
rect 411952 225307 411958 225319
rect 302186 225279 411958 225307
rect 302186 225267 302192 225279
rect 411952 225267 411958 225279
rect 412010 225267 412016 225319
rect 277072 225193 277078 225245
rect 277130 225233 277136 225245
rect 318352 225233 318358 225245
rect 277130 225205 318358 225233
rect 277130 225193 277136 225205
rect 318352 225193 318358 225205
rect 318410 225193 318416 225245
rect 339760 225193 339766 225245
rect 339818 225233 339824 225245
rect 399952 225233 399958 225245
rect 339818 225205 399958 225233
rect 339818 225193 339824 225205
rect 399952 225193 399958 225205
rect 400010 225193 400016 225245
rect 400144 225193 400150 225245
rect 400202 225233 400208 225245
rect 606736 225233 606742 225245
rect 400202 225205 606742 225233
rect 400202 225193 400208 225205
rect 606736 225193 606742 225205
rect 606794 225193 606800 225245
rect 305008 225119 305014 225171
rect 305066 225159 305072 225171
rect 333520 225159 333526 225171
rect 305066 225131 333526 225159
rect 305066 225119 305072 225131
rect 333520 225119 333526 225131
rect 333578 225119 333584 225171
rect 349744 225119 349750 225171
rect 349802 225159 349808 225171
rect 405904 225159 405910 225171
rect 349802 225131 405910 225159
rect 349802 225119 349808 225131
rect 405904 225119 405910 225131
rect 405962 225119 405968 225171
rect 410416 225119 410422 225171
rect 410474 225159 410480 225171
rect 629392 225159 629398 225171
rect 410474 225131 629398 225159
rect 410474 225119 410480 225131
rect 629392 225119 629398 225131
rect 629450 225119 629456 225171
rect 252688 225045 252694 225097
rect 252746 225085 252752 225097
rect 312304 225085 312310 225097
rect 252746 225057 312310 225085
rect 252746 225045 252752 225057
rect 312304 225045 312310 225057
rect 312362 225045 312368 225097
rect 367504 225045 367510 225097
rect 367562 225085 367568 225097
rect 371344 225085 371350 225097
rect 367562 225057 371350 225085
rect 367562 225045 367568 225057
rect 371344 225045 371350 225057
rect 371402 225045 371408 225097
rect 371440 225045 371446 225097
rect 371498 225085 371504 225097
rect 372688 225085 372694 225097
rect 371498 225057 372694 225085
rect 371498 225045 371504 225057
rect 372688 225045 372694 225057
rect 372746 225045 372752 225097
rect 374512 225045 374518 225097
rect 374570 225085 374576 225097
rect 382576 225085 382582 225097
rect 374570 225057 382582 225085
rect 374570 225045 374576 225057
rect 382576 225045 382582 225057
rect 382634 225045 382640 225097
rect 382672 225045 382678 225097
rect 382730 225085 382736 225097
rect 418000 225085 418006 225097
rect 382730 225057 418006 225085
rect 382730 225045 382736 225057
rect 418000 225045 418006 225057
rect 418058 225045 418064 225097
rect 354352 224971 354358 225023
rect 354410 225011 354416 225023
rect 408208 225011 408214 225023
rect 354410 224983 408214 225011
rect 354410 224971 354416 224983
rect 408208 224971 408214 224983
rect 408266 224971 408272 225023
rect 348688 224897 348694 224949
rect 348746 224937 348752 224949
rect 399088 224937 399094 224949
rect 348746 224909 399094 224937
rect 348746 224897 348752 224909
rect 399088 224897 399094 224909
rect 399146 224897 399152 224949
rect 149296 224823 149302 224875
rect 149354 224863 149360 224875
rect 165616 224863 165622 224875
rect 149354 224835 165622 224863
rect 149354 224823 149360 224835
rect 165616 224823 165622 224835
rect 165674 224823 165680 224875
rect 362800 224823 362806 224875
rect 362858 224863 362864 224875
rect 405136 224863 405142 224875
rect 362858 224835 405142 224863
rect 362858 224823 362864 224835
rect 405136 224823 405142 224835
rect 405194 224823 405200 224875
rect 149392 224749 149398 224801
rect 149450 224789 149456 224801
rect 171280 224789 171286 224801
rect 149450 224761 171286 224789
rect 149450 224749 149456 224761
rect 171280 224749 171286 224761
rect 171338 224749 171344 224801
rect 361936 224749 361942 224801
rect 361994 224789 362000 224801
rect 402160 224789 402166 224801
rect 361994 224761 402166 224789
rect 361994 224749 362000 224761
rect 402160 224749 402166 224761
rect 402218 224749 402224 224801
rect 149488 224675 149494 224727
rect 149546 224715 149552 224727
rect 174256 224715 174262 224727
rect 149546 224687 174262 224715
rect 149546 224675 149552 224687
rect 174256 224675 174262 224687
rect 174314 224675 174320 224727
rect 267952 224675 267958 224727
rect 268010 224715 268016 224727
rect 282064 224715 282070 224727
rect 268010 224687 282070 224715
rect 268010 224675 268016 224687
rect 282064 224675 282070 224687
rect 282122 224675 282128 224727
rect 282544 224675 282550 224727
rect 282602 224715 282608 224727
rect 371440 224715 371446 224727
rect 282602 224687 371446 224715
rect 282602 224675 282608 224687
rect 371440 224675 371446 224687
rect 371498 224675 371504 224727
rect 371536 224675 371542 224727
rect 371594 224715 371600 224727
rect 379504 224715 379510 224727
rect 371594 224687 379510 224715
rect 371594 224675 371600 224687
rect 379504 224675 379510 224687
rect 379562 224675 379568 224727
rect 382864 224675 382870 224727
rect 382922 224715 382928 224727
rect 386320 224715 386326 224727
rect 382922 224687 386326 224715
rect 382922 224675 382928 224687
rect 386320 224675 386326 224687
rect 386378 224675 386384 224727
rect 390448 224675 390454 224727
rect 390506 224715 390512 224727
rect 589360 224715 589366 224727
rect 390506 224687 589366 224715
rect 390506 224675 390512 224687
rect 589360 224675 589366 224687
rect 589418 224675 589424 224727
rect 323152 224601 323158 224653
rect 323210 224641 323216 224653
rect 452752 224641 452758 224653
rect 323210 224613 452758 224641
rect 323210 224601 323216 224613
rect 452752 224601 452758 224613
rect 452810 224601 452816 224653
rect 319408 224527 319414 224579
rect 319466 224567 319472 224579
rect 447472 224567 447478 224579
rect 319466 224539 447478 224567
rect 319466 224527 319472 224539
rect 447472 224527 447478 224539
rect 447530 224527 447536 224579
rect 322288 224453 322294 224505
rect 322346 224493 322352 224505
rect 453424 224493 453430 224505
rect 322346 224465 453430 224493
rect 322346 224453 322352 224465
rect 453424 224453 453430 224465
rect 453482 224453 453488 224505
rect 325072 224379 325078 224431
rect 325130 224419 325136 224431
rect 459568 224419 459574 224431
rect 325130 224391 459574 224419
rect 325130 224379 325136 224391
rect 459568 224379 459574 224391
rect 459626 224379 459632 224431
rect 328240 224305 328246 224357
rect 328298 224345 328304 224357
rect 465616 224345 465622 224357
rect 328298 224317 465622 224345
rect 328298 224305 328304 224317
rect 465616 224305 465622 224317
rect 465674 224305 465680 224357
rect 331504 224231 331510 224283
rect 331562 224271 331568 224283
rect 471568 224271 471574 224283
rect 331562 224243 471574 224271
rect 331562 224231 331568 224243
rect 471568 224231 471574 224243
rect 471626 224231 471632 224283
rect 276496 224157 276502 224209
rect 276554 224197 276560 224209
rect 277552 224197 277558 224209
rect 276554 224169 277558 224197
rect 276554 224157 276560 224169
rect 277552 224157 277558 224169
rect 277610 224157 277616 224209
rect 338128 224157 338134 224209
rect 338186 224197 338192 224209
rect 482896 224197 482902 224209
rect 338186 224169 482902 224197
rect 338186 224157 338192 224169
rect 482896 224157 482902 224169
rect 482954 224157 482960 224209
rect 334480 224083 334486 224135
rect 334538 224123 334544 224135
rect 477616 224123 477622 224135
rect 334538 224095 477622 224123
rect 334538 224083 334544 224095
rect 477616 224083 477622 224095
rect 477674 224083 477680 224135
rect 337168 224009 337174 224061
rect 337226 224049 337232 224061
rect 483760 224049 483766 224061
rect 337226 224021 483766 224049
rect 337226 224009 337232 224021
rect 483760 224009 483766 224021
rect 483818 224009 483824 224061
rect 340432 223935 340438 223987
rect 340490 223975 340496 223987
rect 489712 223975 489718 223987
rect 340490 223947 489718 223975
rect 340490 223935 340496 223947
rect 489712 223935 489718 223947
rect 489770 223935 489776 223987
rect 343600 223861 343606 223913
rect 343658 223901 343664 223913
rect 497296 223901 497302 223913
rect 343658 223873 497302 223901
rect 343658 223861 343664 223873
rect 497296 223861 497302 223873
rect 497354 223861 497360 223913
rect 263536 223787 263542 223839
rect 263594 223827 263600 223839
rect 335728 223827 335734 223839
rect 263594 223799 335734 223827
rect 263594 223787 263600 223799
rect 335728 223787 335734 223799
rect 335786 223787 335792 223839
rect 346576 223787 346582 223839
rect 346634 223827 346640 223839
rect 501808 223827 501814 223839
rect 346634 223799 501814 223827
rect 346634 223787 346640 223799
rect 501808 223787 501814 223799
rect 501866 223787 501872 223839
rect 261904 223713 261910 223765
rect 261962 223753 261968 223765
rect 332656 223753 332662 223765
rect 261962 223725 332662 223753
rect 261962 223713 261968 223725
rect 332656 223713 332662 223725
rect 332714 223713 332720 223765
rect 348016 223713 348022 223765
rect 348074 223753 348080 223765
rect 504784 223753 504790 223765
rect 348074 223725 504790 223753
rect 348074 223713 348080 223725
rect 504784 223713 504790 223725
rect 504842 223713 504848 223765
rect 266512 223639 266518 223691
rect 266570 223679 266576 223691
rect 341776 223679 341782 223691
rect 266570 223651 341782 223679
rect 266570 223639 266576 223651
rect 341776 223639 341782 223651
rect 341834 223639 341840 223691
rect 349552 223639 349558 223691
rect 349610 223679 349616 223691
rect 507856 223679 507862 223691
rect 349610 223651 507862 223679
rect 349610 223639 349616 223651
rect 507856 223639 507862 223651
rect 507914 223639 507920 223691
rect 268048 223565 268054 223617
rect 268106 223605 268112 223617
rect 344848 223605 344854 223617
rect 268106 223577 344854 223605
rect 268106 223565 268112 223577
rect 344848 223565 344854 223577
rect 344906 223565 344912 223617
rect 350800 223565 350806 223617
rect 350858 223605 350864 223617
rect 510832 223605 510838 223617
rect 350858 223577 510838 223605
rect 350858 223565 350864 223577
rect 510832 223565 510838 223577
rect 510890 223565 510896 223617
rect 264592 223491 264598 223543
rect 264650 223531 264656 223543
rect 338704 223531 338710 223543
rect 264650 223503 338710 223531
rect 264650 223491 264656 223503
rect 338704 223491 338710 223503
rect 338762 223491 338768 223543
rect 348112 223491 348118 223543
rect 348170 223531 348176 223543
rect 506320 223531 506326 223543
rect 348170 223503 506326 223531
rect 348170 223491 348176 223503
rect 506320 223491 506326 223503
rect 506378 223491 506384 223543
rect 269488 223417 269494 223469
rect 269546 223457 269552 223469
rect 347728 223457 347734 223469
rect 269546 223429 347734 223457
rect 269546 223417 269552 223429
rect 347728 223417 347734 223429
rect 347786 223417 347792 223469
rect 351184 223417 351190 223469
rect 351242 223457 351248 223469
rect 512368 223457 512374 223469
rect 351242 223429 512374 223457
rect 351242 223417 351248 223429
rect 512368 223417 512374 223429
rect 512426 223417 512432 223469
rect 271120 223343 271126 223395
rect 271178 223383 271184 223395
rect 350800 223383 350806 223395
rect 271178 223355 350806 223383
rect 271178 223343 271184 223355
rect 350800 223343 350806 223355
rect 350858 223343 350864 223395
rect 352528 223343 352534 223395
rect 352586 223383 352592 223395
rect 513904 223383 513910 223395
rect 352586 223355 513910 223383
rect 352586 223343 352592 223355
rect 513904 223343 513910 223355
rect 513962 223343 513968 223395
rect 354064 223269 354070 223321
rect 354122 223309 354128 223321
rect 516976 223309 516982 223321
rect 354122 223281 516982 223309
rect 354122 223269 354128 223281
rect 516976 223269 516982 223281
rect 517034 223269 517040 223321
rect 272560 223195 272566 223247
rect 272618 223235 272624 223247
rect 353872 223235 353878 223247
rect 272618 223207 353878 223235
rect 272618 223195 272624 223207
rect 353872 223195 353878 223207
rect 353930 223195 353936 223247
rect 355600 223195 355606 223247
rect 355658 223235 355664 223247
rect 519856 223235 519862 223247
rect 355658 223207 519862 223235
rect 355658 223195 355664 223207
rect 519856 223195 519862 223207
rect 519914 223195 519920 223247
rect 286192 223121 286198 223173
rect 286250 223161 286256 223173
rect 381040 223161 381046 223173
rect 286250 223133 381046 223161
rect 286250 223121 286256 223133
rect 381040 223121 381046 223133
rect 381098 223121 381104 223173
rect 394864 223121 394870 223173
rect 394922 223161 394928 223173
rect 523792 223161 523798 223173
rect 394922 223133 523798 223161
rect 394922 223121 394928 223133
rect 523792 223121 523798 223133
rect 523850 223121 523856 223173
rect 316336 223047 316342 223099
rect 316394 223087 316400 223099
rect 441424 223087 441430 223099
rect 316394 223059 441430 223087
rect 316394 223047 316400 223059
rect 441424 223047 441430 223059
rect 441482 223047 441488 223099
rect 318544 222973 318550 223025
rect 318602 223013 318608 223025
rect 443728 223013 443734 223025
rect 318602 222985 443734 223013
rect 318602 222973 318608 222985
rect 443728 222973 443734 222985
rect 443786 222973 443792 223025
rect 313360 222899 313366 222951
rect 313418 222939 313424 222951
rect 435376 222939 435382 222951
rect 313418 222911 435382 222939
rect 313418 222899 313424 222911
rect 435376 222899 435382 222911
rect 435434 222899 435440 222951
rect 310288 222825 310294 222877
rect 310346 222865 310352 222877
rect 429328 222865 429334 222877
rect 310346 222837 429334 222865
rect 310346 222825 310352 222837
rect 429328 222825 429334 222837
rect 429386 222825 429392 222877
rect 307984 222751 307990 222803
rect 308042 222791 308048 222803
rect 422512 222791 422518 222803
rect 308042 222763 422518 222791
rect 308042 222751 308048 222763
rect 422512 222751 422518 222763
rect 422570 222751 422576 222803
rect 312592 222677 312598 222729
rect 312650 222717 312656 222729
rect 431536 222717 431542 222729
rect 312650 222689 431542 222717
rect 312650 222677 312656 222689
rect 431536 222677 431542 222689
rect 431594 222677 431600 222729
rect 307216 222603 307222 222655
rect 307274 222643 307280 222655
rect 423280 222643 423286 222655
rect 307274 222615 423286 222643
rect 307274 222603 307280 222615
rect 423280 222603 423286 222615
rect 423338 222603 423344 222655
rect 304240 222529 304246 222581
rect 304298 222569 304304 222581
rect 417232 222569 417238 222581
rect 304298 222541 417238 222569
rect 304298 222529 304304 222541
rect 417232 222529 417238 222541
rect 417290 222529 417296 222581
rect 302800 222455 302806 222507
rect 302858 222495 302864 222507
rect 414256 222495 414262 222507
rect 302858 222467 414262 222495
rect 302858 222455 302864 222467
rect 414256 222455 414262 222467
rect 414314 222455 414320 222507
rect 283120 222381 283126 222433
rect 283178 222421 283184 222433
rect 374992 222421 374998 222433
rect 283178 222393 374998 222421
rect 283178 222381 283184 222393
rect 374992 222381 374998 222393
rect 375050 222381 375056 222433
rect 391792 222381 391798 222433
rect 391850 222421 391856 222433
rect 496528 222421 496534 222433
rect 391850 222393 496534 222421
rect 391850 222381 391856 222393
rect 496528 222381 496534 222393
rect 496586 222381 496592 222433
rect 281584 222307 281590 222359
rect 281642 222347 281648 222359
rect 371920 222347 371926 222359
rect 281642 222319 371926 222347
rect 281642 222307 281648 222319
rect 371920 222307 371926 222319
rect 371978 222307 371984 222359
rect 374704 222307 374710 222359
rect 374762 222347 374768 222359
rect 467824 222347 467830 222359
rect 374762 222319 467830 222347
rect 374762 222307 374768 222319
rect 467824 222307 467830 222319
rect 467882 222307 467888 222359
rect 274096 222233 274102 222285
rect 274154 222273 274160 222285
rect 356848 222273 356854 222285
rect 274154 222245 356854 222273
rect 274154 222233 274160 222245
rect 356848 222233 356854 222245
rect 356906 222233 356912 222285
rect 656176 222011 656182 222063
rect 656234 222051 656240 222063
rect 676240 222051 676246 222063
rect 656234 222023 676246 222051
rect 656234 222011 656240 222023
rect 676240 222011 676246 222023
rect 676298 222011 676304 222063
rect 149488 221863 149494 221915
rect 149546 221903 149552 221915
rect 162640 221903 162646 221915
rect 149546 221875 162646 221903
rect 149546 221863 149552 221875
rect 162640 221863 162646 221875
rect 162698 221863 162704 221915
rect 655984 221863 655990 221915
rect 656042 221903 656048 221915
rect 676240 221903 676246 221915
rect 656042 221875 676246 221903
rect 656042 221863 656048 221875
rect 676240 221863 676246 221875
rect 676298 221863 676304 221915
rect 149392 221789 149398 221841
rect 149450 221829 149456 221841
rect 168400 221829 168406 221841
rect 149450 221801 168406 221829
rect 149450 221789 149456 221801
rect 168400 221789 168406 221801
rect 168458 221789 168464 221841
rect 42064 221715 42070 221767
rect 42122 221755 42128 221767
rect 50320 221755 50326 221767
rect 42122 221727 50326 221755
rect 42122 221715 42128 221727
rect 50320 221715 50326 221727
rect 50378 221715 50384 221767
rect 159952 221715 159958 221767
rect 160010 221755 160016 221767
rect 184336 221755 184342 221767
rect 160010 221727 184342 221755
rect 160010 221715 160016 221727
rect 184336 221715 184342 221727
rect 184394 221715 184400 221767
rect 195760 221715 195766 221767
rect 195818 221715 195824 221767
rect 197536 221715 197542 221767
rect 197594 221715 197600 221767
rect 512752 221715 512758 221767
rect 512810 221755 512816 221767
rect 515392 221755 515398 221767
rect 512810 221727 515398 221755
rect 512810 221715 512816 221727
rect 515392 221715 515398 221727
rect 515450 221715 515456 221767
rect 195778 221681 195806 221715
rect 197554 221681 197582 221715
rect 195778 221653 197582 221681
rect 673456 219865 673462 219917
rect 673514 219905 673520 219917
rect 676240 219905 676246 219917
rect 673514 219877 676246 219905
rect 673514 219865 673520 219877
rect 676240 219865 676246 219877
rect 676298 219865 676304 219917
rect 147664 219051 147670 219103
rect 147722 219091 147728 219103
rect 174352 219091 174358 219103
rect 147722 219063 174358 219091
rect 147722 219051 147728 219063
rect 174352 219051 174358 219063
rect 174410 219051 174416 219103
rect 655792 219051 655798 219103
rect 655850 219091 655856 219103
rect 676048 219091 676054 219103
rect 655850 219063 676054 219091
rect 655850 219051 655856 219063
rect 676048 219051 676054 219063
rect 676106 219051 676112 219103
rect 149392 218977 149398 219029
rect 149450 219017 149456 219029
rect 177136 219017 177142 219029
rect 149450 218989 177142 219017
rect 149450 218977 149456 218989
rect 177136 218977 177142 218989
rect 177194 218977 177200 219029
rect 149488 218903 149494 218955
rect 149546 218943 149552 218955
rect 179920 218943 179926 218955
rect 149546 218915 179926 218943
rect 149546 218903 149552 218915
rect 179920 218903 179926 218915
rect 179978 218903 179984 218955
rect 143056 218829 143062 218881
rect 143114 218869 143120 218881
rect 184336 218869 184342 218881
rect 143114 218841 184342 218869
rect 143114 218829 143120 218841
rect 184336 218829 184342 218841
rect 184394 218829 184400 218881
rect 673360 218755 673366 218807
rect 673418 218795 673424 218807
rect 676048 218795 676054 218807
rect 673418 218767 676054 218795
rect 673418 218755 673424 218767
rect 676048 218755 676054 218767
rect 676106 218755 676112 218807
rect 147280 217719 147286 217771
rect 147338 217759 147344 217771
rect 151792 217759 151798 217771
rect 147338 217731 151798 217759
rect 147338 217719 147344 217731
rect 151792 217719 151798 217731
rect 151850 217719 151856 217771
rect 149392 216387 149398 216439
rect 149450 216427 149456 216439
rect 159952 216427 159958 216439
rect 149450 216399 159958 216427
rect 149450 216387 149456 216399
rect 159952 216387 159958 216399
rect 160010 216387 160016 216439
rect 41776 213649 41782 213701
rect 41834 213689 41840 213701
rect 45328 213689 45334 213701
rect 41834 213661 45334 213689
rect 41834 213649 41840 213661
rect 45328 213649 45334 213661
rect 45386 213649 45392 213701
rect 147568 213279 147574 213331
rect 147626 213319 147632 213331
rect 151696 213319 151702 213331
rect 147626 213291 151702 213319
rect 147626 213279 147632 213291
rect 151696 213279 151702 213291
rect 151754 213279 151760 213331
rect 674800 213205 674806 213257
rect 674858 213245 674864 213257
rect 676048 213245 676054 213257
rect 674858 213217 676054 213245
rect 674858 213205 674864 213217
rect 676048 213205 676054 213217
rect 676106 213205 676112 213257
rect 41776 213131 41782 213183
rect 41834 213171 41840 213183
rect 45616 213171 45622 213183
rect 41834 213143 45622 213171
rect 41834 213131 41840 213143
rect 45616 213131 45622 213143
rect 45674 213131 45680 213183
rect 147376 213131 147382 213183
rect 147434 213171 147440 213183
rect 151504 213171 151510 213183
rect 147434 213143 151510 213171
rect 147434 213131 147440 213143
rect 151504 213131 151510 213143
rect 151562 213131 151568 213183
rect 675088 213131 675094 213183
rect 675146 213171 675152 213183
rect 676240 213171 676246 213183
rect 675146 213143 676246 213171
rect 675146 213131 675152 213143
rect 676240 213131 676246 213143
rect 676298 213131 676304 213183
rect 146896 212835 146902 212887
rect 146954 212875 146960 212887
rect 152080 212875 152086 212887
rect 146954 212847 152086 212875
rect 146954 212835 146960 212847
rect 152080 212835 152086 212847
rect 152138 212835 152144 212887
rect 180112 212835 180118 212887
rect 180170 212875 180176 212887
rect 187024 212875 187030 212887
rect 180170 212847 187030 212875
rect 180170 212835 180176 212847
rect 187024 212835 187030 212847
rect 187082 212835 187088 212887
rect 41584 212761 41590 212813
rect 41642 212801 41648 212813
rect 45520 212801 45526 212813
rect 41642 212773 45526 212801
rect 41642 212761 41648 212773
rect 45520 212761 45526 212773
rect 45578 212761 45584 212813
rect 41776 212169 41782 212221
rect 41834 212209 41840 212221
rect 43408 212209 43414 212221
rect 41834 212181 43414 212209
rect 41834 212169 41840 212181
rect 43408 212169 43414 212181
rect 43466 212169 43472 212221
rect 674608 211873 674614 211925
rect 674666 211913 674672 211925
rect 676048 211913 676054 211925
rect 674666 211885 676054 211913
rect 674666 211873 674672 211885
rect 676048 211873 676054 211885
rect 676106 211873 676112 211925
rect 41776 211651 41782 211703
rect 41834 211691 41840 211703
rect 44848 211691 44854 211703
rect 41834 211663 44854 211691
rect 41834 211651 41840 211663
rect 44848 211651 44854 211663
rect 44906 211651 44912 211703
rect 41584 211281 41590 211333
rect 41642 211321 41648 211333
rect 50608 211321 50614 211333
rect 41642 211293 50614 211321
rect 41642 211281 41648 211293
rect 50608 211281 50614 211293
rect 50666 211281 50672 211333
rect 41776 210689 41782 210741
rect 41834 210729 41840 210741
rect 43312 210729 43318 210741
rect 41834 210701 43318 210729
rect 41834 210689 41840 210701
rect 43312 210689 43318 210701
rect 43370 210689 43376 210741
rect 147376 210467 147382 210519
rect 147434 210507 147440 210519
rect 151600 210507 151606 210519
rect 147434 210479 151606 210507
rect 147434 210467 147440 210479
rect 151600 210467 151606 210479
rect 151658 210467 151664 210519
rect 674704 210393 674710 210445
rect 674762 210433 674768 210445
rect 675952 210433 675958 210445
rect 674762 210405 675958 210433
rect 674762 210393 674768 210405
rect 675952 210393 675958 210405
rect 676010 210393 676016 210445
rect 147376 210319 147382 210371
rect 147434 210359 147440 210371
rect 151408 210359 151414 210371
rect 147434 210331 151414 210359
rect 147434 210319 147440 210331
rect 151408 210319 151414 210331
rect 151466 210319 151472 210371
rect 674896 210319 674902 210371
rect 674954 210359 674960 210371
rect 676048 210359 676054 210371
rect 674954 210331 676054 210359
rect 674954 210319 674960 210331
rect 676048 210319 676054 210331
rect 676106 210319 676112 210371
rect 674992 210245 674998 210297
rect 675050 210285 675056 210297
rect 676240 210285 676246 210297
rect 675050 210257 676246 210285
rect 675050 210245 675056 210257
rect 676240 210245 676246 210257
rect 676298 210245 676304 210297
rect 41776 210097 41782 210149
rect 41834 210137 41840 210149
rect 50416 210137 50422 210149
rect 41834 210109 50422 210137
rect 41834 210097 41840 210109
rect 50416 210097 50422 210109
rect 50474 210097 50480 210149
rect 41584 209801 41590 209853
rect 41642 209841 41648 209853
rect 43504 209841 43510 209853
rect 41642 209813 43510 209841
rect 41642 209801 41648 209813
rect 43504 209801 43510 209813
rect 43562 209801 43568 209853
rect 146896 208321 146902 208373
rect 146954 208361 146960 208373
rect 151984 208361 151990 208373
rect 146954 208333 151990 208361
rect 146954 208321 146960 208333
rect 151984 208321 151990 208333
rect 152042 208321 152048 208373
rect 146992 207359 146998 207411
rect 147050 207399 147056 207411
rect 151312 207399 151318 207411
rect 147050 207371 151318 207399
rect 147050 207359 147056 207371
rect 151312 207359 151318 207371
rect 151370 207359 151376 207411
rect 646768 207359 646774 207411
rect 646826 207399 646832 207411
rect 679984 207399 679990 207411
rect 646826 207371 679990 207399
rect 646826 207359 646832 207371
rect 679984 207359 679990 207371
rect 680042 207359 680048 207411
rect 147088 206249 147094 206301
rect 147146 206289 147152 206301
rect 151888 206289 151894 206301
rect 147146 206261 151894 206289
rect 147146 206249 147152 206261
rect 151888 206249 151894 206261
rect 151946 206249 151952 206301
rect 675760 206101 675766 206153
rect 675818 206101 675824 206153
rect 675088 205657 675094 205709
rect 675146 205697 675152 205709
rect 675472 205697 675478 205709
rect 675146 205669 675478 205697
rect 675146 205657 675152 205669
rect 675472 205657 675478 205669
rect 675530 205657 675536 205709
rect 675778 205635 675806 206101
rect 675760 205583 675766 205635
rect 675818 205583 675824 205635
rect 149392 204547 149398 204599
rect 149450 204587 149456 204599
rect 157072 204587 157078 204599
rect 149450 204559 157078 204587
rect 149450 204547 149456 204559
rect 157072 204547 157078 204559
rect 157130 204547 157136 204599
rect 147664 204029 147670 204081
rect 147722 204069 147728 204081
rect 154192 204069 154198 204081
rect 147722 204041 154198 204069
rect 147722 204029 147728 204041
rect 154192 204029 154198 204041
rect 154250 204029 154256 204081
rect 41776 203289 41782 203341
rect 41834 203329 41840 203341
rect 43024 203329 43030 203341
rect 41834 203301 43030 203329
rect 41834 203289 41840 203301
rect 43024 203289 43030 203301
rect 43082 203289 43088 203341
rect 41776 202771 41782 202823
rect 41834 202811 41840 202823
rect 42928 202811 42934 202823
rect 41834 202783 42934 202811
rect 41834 202771 41840 202783
rect 42928 202771 42934 202783
rect 42986 202771 42992 202823
rect 41968 202105 41974 202157
rect 42026 202145 42032 202157
rect 44656 202145 44662 202157
rect 42026 202117 44662 202145
rect 42026 202105 42032 202117
rect 44656 202105 44662 202117
rect 44714 202105 44720 202157
rect 675184 201883 675190 201935
rect 675242 201923 675248 201935
rect 675472 201923 675478 201935
rect 675242 201895 675478 201923
rect 675242 201883 675248 201895
rect 675472 201883 675478 201895
rect 675530 201883 675536 201935
rect 41968 201661 41974 201713
rect 42026 201701 42032 201713
rect 44752 201701 44758 201713
rect 42026 201673 44758 201701
rect 42026 201661 42032 201673
rect 44752 201661 44758 201673
rect 44810 201661 44816 201713
rect 149488 201661 149494 201713
rect 149546 201701 149552 201713
rect 180112 201701 180118 201713
rect 149546 201673 180118 201701
rect 149546 201661 149552 201673
rect 180112 201661 180118 201673
rect 180170 201661 180176 201713
rect 41776 201587 41782 201639
rect 41834 201627 41840 201639
rect 42736 201627 42742 201639
rect 41834 201599 42742 201627
rect 41834 201587 41840 201599
rect 42736 201587 42742 201599
rect 42794 201587 42800 201639
rect 149392 201587 149398 201639
rect 149450 201627 149456 201639
rect 182992 201627 182998 201639
rect 149450 201599 182998 201627
rect 149450 201587 149456 201599
rect 182992 201587 182998 201599
rect 183050 201587 183056 201639
rect 143056 201513 143062 201565
rect 143114 201553 143120 201565
rect 184336 201553 184342 201565
rect 143114 201525 184342 201553
rect 143114 201513 143120 201525
rect 184336 201513 184342 201525
rect 184394 201513 184400 201565
rect 655600 201513 655606 201565
rect 655658 201553 655664 201565
rect 675088 201553 675094 201565
rect 655658 201525 675094 201553
rect 655658 201513 655664 201525
rect 675088 201513 675094 201525
rect 675146 201513 675152 201565
rect 674800 201291 674806 201343
rect 674858 201331 674864 201343
rect 675376 201331 675382 201343
rect 674858 201303 675382 201331
rect 674858 201291 674864 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 41776 201217 41782 201269
rect 41834 201257 41840 201269
rect 44560 201257 44566 201269
rect 41834 201229 44566 201257
rect 41834 201217 41840 201229
rect 44560 201217 44566 201229
rect 44618 201217 44624 201269
rect 674992 200847 674998 200899
rect 675050 200887 675056 200899
rect 675376 200887 675382 200899
rect 675050 200859 675382 200887
rect 675050 200847 675056 200859
rect 675376 200847 675382 200859
rect 675434 200847 675440 200899
rect 41584 198849 41590 198901
rect 41642 198889 41648 198901
rect 42832 198889 42838 198901
rect 41642 198861 42838 198889
rect 41642 198849 41648 198861
rect 42832 198849 42838 198861
rect 42890 198849 42896 198901
rect 147472 198775 147478 198827
rect 147530 198815 147536 198827
rect 152176 198815 152182 198827
rect 147530 198787 152182 198815
rect 147530 198775 147536 198787
rect 152176 198775 152182 198787
rect 152234 198775 152240 198827
rect 149392 198701 149398 198753
rect 149450 198741 149456 198753
rect 165712 198741 165718 198753
rect 149450 198713 165718 198741
rect 149450 198701 149456 198713
rect 165712 198701 165718 198713
rect 165770 198701 165776 198753
rect 181360 198627 181366 198679
rect 181418 198667 181424 198679
rect 184432 198667 184438 198679
rect 181418 198639 184438 198667
rect 181418 198627 181424 198639
rect 184432 198627 184438 198639
rect 184490 198627 184496 198679
rect 178288 198553 178294 198605
rect 178346 198593 178352 198605
rect 184336 198593 184342 198605
rect 178346 198565 184342 198593
rect 178346 198553 178352 198565
rect 184336 198553 184342 198565
rect 184394 198553 184400 198605
rect 674896 197739 674902 197791
rect 674954 197779 674960 197791
rect 675376 197779 675382 197791
rect 674954 197751 675382 197779
rect 674954 197739 674960 197751
rect 675376 197739 675382 197751
rect 675434 197739 675440 197791
rect 41872 197369 41878 197421
rect 41930 197369 41936 197421
rect 41890 197199 41918 197369
rect 41872 197147 41878 197199
rect 41930 197147 41936 197199
rect 674608 196999 674614 197051
rect 674666 197039 674672 197051
rect 675472 197039 675478 197051
rect 674666 197011 675478 197039
rect 674666 196999 674672 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 674704 196555 674710 196607
rect 674762 196595 674768 196607
rect 675376 196595 675382 196607
rect 674762 196567 675382 196595
rect 674762 196555 674768 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 147280 195963 147286 196015
rect 147338 196003 147344 196015
rect 168592 196003 168598 196015
rect 147338 195975 168598 196003
rect 147338 195963 147344 195975
rect 168592 195963 168598 195975
rect 168650 195963 168656 196015
rect 149392 195889 149398 195941
rect 149450 195929 149456 195941
rect 171472 195929 171478 195941
rect 149450 195901 171478 195929
rect 149450 195889 149456 195901
rect 171472 195889 171478 195901
rect 171530 195889 171536 195941
rect 149296 195815 149302 195867
rect 149354 195855 149360 195867
rect 177328 195855 177334 195867
rect 149354 195827 177334 195855
rect 149354 195815 149360 195827
rect 177328 195815 177334 195827
rect 177386 195815 177392 195867
rect 166960 195741 166966 195793
rect 167018 195781 167024 195793
rect 184528 195781 184534 195793
rect 167018 195753 184534 195781
rect 167018 195741 167024 195753
rect 184528 195741 184534 195753
rect 184586 195741 184592 195793
rect 169840 195667 169846 195719
rect 169898 195707 169904 195719
rect 184432 195707 184438 195719
rect 169898 195679 184438 195707
rect 169898 195667 169904 195679
rect 184432 195667 184438 195679
rect 184490 195667 184496 195719
rect 172720 195593 172726 195645
rect 172778 195633 172784 195645
rect 184336 195633 184342 195645
rect 172778 195605 184342 195633
rect 172778 195593 172784 195605
rect 184336 195593 184342 195605
rect 184394 195593 184400 195645
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 42832 193487 42838 193499
rect 42122 193459 42838 193487
rect 42122 193447 42128 193459
rect 42832 193447 42838 193459
rect 42890 193447 42896 193499
rect 149392 193151 149398 193203
rect 149450 193191 149456 193203
rect 160048 193191 160054 193203
rect 149450 193163 160054 193191
rect 149450 193151 149456 193163
rect 160048 193151 160054 193163
rect 160106 193151 160112 193203
rect 149488 193003 149494 193055
rect 149546 193043 149552 193055
rect 162832 193043 162838 193055
rect 149546 193015 162838 193043
rect 149546 193003 149552 193015
rect 162832 193003 162838 193015
rect 162890 193003 162896 193055
rect 152368 192929 152374 192981
rect 152426 192969 152432 192981
rect 184624 192969 184630 192981
rect 152426 192941 184630 192969
rect 152426 192929 152432 192941
rect 184624 192929 184630 192941
rect 184682 192929 184688 192981
rect 155440 192855 155446 192907
rect 155498 192895 155504 192907
rect 184528 192895 184534 192907
rect 155498 192867 184534 192895
rect 155498 192855 155504 192867
rect 184528 192855 184534 192867
rect 184586 192855 184592 192907
rect 158128 192781 158134 192833
rect 158186 192821 158192 192833
rect 184336 192821 184342 192833
rect 158186 192793 184342 192821
rect 158186 192781 158192 192793
rect 184336 192781 184342 192793
rect 184394 192781 184400 192833
rect 163888 192707 163894 192759
rect 163946 192747 163952 192759
rect 184432 192747 184438 192759
rect 163946 192719 184438 192747
rect 163946 192707 163952 192719
rect 184432 192707 184438 192719
rect 184490 192707 184496 192759
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 42736 192229 42742 192241
rect 42218 192201 42742 192229
rect 42218 192189 42224 192201
rect 42736 192189 42742 192201
rect 42794 192189 42800 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 43024 191489 43030 191501
rect 42122 191461 43030 191489
rect 42122 191449 42128 191461
rect 43024 191449 43030 191461
rect 43082 191449 43088 191501
rect 149392 191079 149398 191131
rect 149450 191119 149456 191131
rect 157168 191119 157174 191131
rect 149450 191091 157174 191119
rect 149450 191079 149456 191091
rect 157168 191079 157174 191091
rect 157226 191079 157232 191131
rect 42160 191005 42166 191057
rect 42218 191045 42224 191057
rect 42928 191045 42934 191057
rect 42218 191017 42934 191045
rect 42218 191005 42224 191017
rect 42928 191005 42934 191017
rect 42986 191005 42992 191057
rect 147280 190117 147286 190169
rect 147338 190157 147344 190169
rect 154288 190157 154294 190169
rect 147338 190129 154294 190157
rect 147338 190117 147344 190129
rect 154288 190117 154294 190129
rect 154346 190117 154352 190169
rect 143920 190043 143926 190095
rect 143978 190083 143984 190095
rect 184528 190083 184534 190095
rect 143978 190055 184534 190083
rect 143978 190043 143984 190055
rect 184528 190043 184534 190055
rect 184586 190043 184592 190095
rect 149680 189969 149686 190021
rect 149738 190009 149744 190021
rect 184336 190009 184342 190021
rect 149738 189981 184342 190009
rect 149738 189969 149744 189981
rect 184336 189969 184342 189981
rect 184394 189969 184400 190021
rect 171376 189895 171382 189947
rect 171434 189935 171440 189947
rect 184432 189935 184438 189947
rect 171434 189907 184438 189935
rect 171434 189895 171440 189907
rect 184432 189895 184438 189907
rect 184490 189895 184496 189947
rect 180016 189821 180022 189873
rect 180074 189861 180080 189873
rect 184336 189861 184342 189873
rect 180074 189833 184342 189861
rect 180074 189821 180080 189833
rect 184336 189821 184342 189833
rect 184394 189821 184400 189873
rect 162736 187157 162742 187209
rect 162794 187197 162800 187209
rect 184432 187197 184438 187209
rect 162794 187169 184438 187197
rect 162794 187157 162800 187169
rect 184432 187157 184438 187169
rect 184490 187157 184496 187209
rect 168496 187083 168502 187135
rect 168554 187123 168560 187135
rect 184336 187123 184342 187135
rect 168554 187095 184342 187123
rect 168554 187083 168560 187095
rect 184336 187083 184342 187095
rect 184394 187083 184400 187135
rect 174448 187009 174454 187061
rect 174506 187049 174512 187061
rect 184528 187049 184534 187061
rect 174506 187021 184534 187049
rect 174506 187009 174512 187021
rect 184528 187009 184534 187021
rect 184586 187009 184592 187061
rect 177232 186935 177238 186987
rect 177290 186975 177296 186987
rect 184624 186975 184630 186987
rect 177290 186947 184630 186975
rect 177290 186935 177296 186947
rect 184624 186935 184630 186947
rect 184682 186935 184688 186987
rect 149392 185751 149398 185803
rect 149450 185791 149456 185803
rect 186064 185791 186070 185803
rect 149450 185763 186070 185791
rect 149450 185751 149456 185763
rect 186064 185751 186070 185763
rect 186122 185751 186128 185803
rect 145552 184271 145558 184323
rect 145610 184311 145616 184323
rect 184336 184311 184342 184323
rect 145610 184283 184342 184311
rect 145610 184271 145616 184283
rect 184336 184271 184342 184283
rect 184394 184271 184400 184323
rect 156976 184197 156982 184249
rect 157034 184237 157040 184249
rect 184432 184237 184438 184249
rect 157034 184209 184438 184237
rect 157034 184197 157040 184209
rect 184432 184197 184438 184209
rect 184490 184197 184496 184249
rect 177040 184123 177046 184175
rect 177098 184163 177104 184175
rect 184528 184163 184534 184175
rect 177098 184135 184534 184163
rect 177098 184123 177104 184135
rect 184528 184123 184534 184135
rect 184586 184123 184592 184175
rect 645136 183087 645142 183139
rect 645194 183127 645200 183139
rect 649360 183127 649366 183139
rect 645194 183099 649366 183127
rect 645194 183087 645200 183099
rect 649360 183087 649366 183099
rect 649418 183087 649424 183139
rect 149296 182939 149302 182991
rect 149354 182979 149360 182991
rect 185968 182979 185974 182991
rect 149354 182951 185974 182979
rect 149354 182939 149360 182951
rect 185968 182939 185974 182951
rect 186026 182939 186032 182991
rect 149584 182865 149590 182917
rect 149642 182905 149648 182917
rect 186160 182905 186166 182917
rect 149642 182877 186166 182905
rect 149642 182865 149648 182877
rect 186160 182865 186166 182877
rect 186218 182865 186224 182917
rect 42160 182199 42166 182251
rect 42218 182239 42224 182251
rect 48112 182239 48118 182251
rect 42218 182211 48118 182239
rect 42218 182199 42224 182211
rect 48112 182199 48118 182211
rect 48170 182199 48176 182251
rect 149392 181533 149398 181585
rect 149450 181573 149456 181585
rect 165808 181573 165814 181585
rect 149450 181545 165814 181573
rect 149450 181533 149456 181545
rect 165808 181533 165814 181545
rect 165866 181533 165872 181585
rect 149488 181459 149494 181511
rect 149546 181499 149552 181511
rect 174448 181499 174454 181511
rect 149546 181471 174454 181499
rect 149546 181459 149552 181471
rect 174448 181459 174454 181471
rect 174506 181459 174512 181511
rect 154000 181385 154006 181437
rect 154058 181425 154064 181437
rect 184624 181425 184630 181437
rect 154058 181397 184630 181425
rect 154058 181385 154064 181397
rect 184624 181385 184630 181397
rect 184682 181385 184688 181437
rect 156880 181311 156886 181363
rect 156938 181351 156944 181363
rect 184336 181351 184342 181363
rect 156938 181323 184342 181351
rect 156938 181311 156944 181323
rect 184336 181311 184342 181323
rect 184394 181311 184400 181363
rect 159760 181237 159766 181289
rect 159818 181277 159824 181289
rect 184432 181277 184438 181289
rect 159818 181249 184438 181277
rect 159818 181237 159824 181249
rect 184432 181237 184438 181249
rect 184490 181237 184496 181289
rect 174160 181163 174166 181215
rect 174218 181203 174224 181215
rect 184528 181203 184534 181215
rect 174218 181175 184534 181203
rect 174218 181163 174224 181175
rect 184528 181163 184534 181175
rect 184586 181163 184592 181215
rect 149200 179979 149206 180031
rect 149258 180019 149264 180031
rect 185488 180019 185494 180031
rect 149258 179991 185494 180019
rect 149258 179979 149264 179991
rect 185488 179979 185494 179991
rect 185546 179979 185552 180031
rect 645136 179387 645142 179439
rect 645194 179427 645200 179439
rect 649456 179427 649462 179439
rect 645194 179399 649462 179427
rect 645194 179387 645200 179399
rect 649456 179387 649462 179399
rect 649514 179387 649520 179439
rect 149488 178721 149494 178773
rect 149546 178761 149552 178773
rect 162736 178761 162742 178773
rect 149546 178733 162742 178761
rect 149546 178721 149552 178733
rect 162736 178721 162742 178733
rect 162794 178721 162800 178773
rect 149392 178647 149398 178699
rect 149450 178687 149456 178699
rect 171376 178687 171382 178699
rect 149450 178659 171382 178687
rect 149450 178647 149456 178659
rect 171376 178647 171382 178659
rect 171434 178647 171440 178699
rect 149296 178573 149302 178625
rect 149354 178613 149360 178625
rect 183088 178613 183094 178625
rect 149354 178585 183094 178613
rect 149354 178573 149360 178585
rect 183088 178573 183094 178585
rect 183146 178573 183152 178625
rect 145456 178499 145462 178551
rect 145514 178539 145520 178551
rect 184432 178539 184438 178551
rect 145514 178511 184438 178539
rect 145514 178499 145520 178511
rect 184432 178499 184438 178511
rect 184490 178499 184496 178551
rect 165520 178425 165526 178477
rect 165578 178465 165584 178477
rect 184336 178465 184342 178477
rect 165578 178437 184342 178465
rect 165578 178425 165584 178437
rect 184336 178425 184342 178437
rect 184394 178425 184400 178477
rect 182800 178351 182806 178403
rect 182858 178391 182864 178403
rect 186736 178391 186742 178403
rect 182858 178363 186742 178391
rect 182858 178351 182864 178363
rect 186736 178351 186742 178363
rect 186794 178351 186800 178403
rect 655696 176131 655702 176183
rect 655754 176171 655760 176183
rect 676144 176171 676150 176183
rect 655754 176143 676150 176171
rect 655754 176131 655760 176143
rect 676144 176131 676150 176143
rect 676202 176131 676208 176183
rect 655504 175983 655510 176035
rect 655562 176023 655568 176035
rect 676240 176023 676246 176035
rect 655562 175995 676246 176023
rect 655562 175983 655568 175995
rect 676240 175983 676246 175995
rect 676298 175983 676304 176035
rect 655408 175835 655414 175887
rect 655466 175875 655472 175887
rect 676336 175875 676342 175887
rect 655466 175847 676342 175875
rect 655466 175835 655472 175847
rect 676336 175835 676342 175847
rect 676394 175835 676400 175887
rect 149392 175761 149398 175813
rect 149450 175801 149456 175813
rect 156880 175801 156886 175813
rect 149450 175773 156886 175801
rect 149450 175761 149456 175773
rect 156880 175761 156886 175773
rect 156938 175761 156944 175813
rect 149488 175687 149494 175739
rect 149546 175727 149552 175739
rect 168496 175727 168502 175739
rect 149546 175699 168502 175727
rect 149546 175687 149552 175699
rect 168496 175687 168502 175699
rect 168554 175687 168560 175739
rect 143056 175613 143062 175665
rect 143114 175653 143120 175665
rect 184432 175653 184438 175665
rect 143114 175625 184438 175653
rect 143114 175613 143120 175625
rect 184432 175613 184438 175625
rect 184490 175613 184496 175665
rect 145360 175539 145366 175591
rect 145418 175579 145424 175591
rect 184336 175579 184342 175591
rect 145418 175551 184342 175579
rect 145418 175539 145424 175551
rect 184336 175539 184342 175551
rect 184394 175539 184400 175591
rect 147664 175021 147670 175073
rect 147722 175061 147728 175073
rect 154000 175061 154006 175073
rect 147722 175033 154006 175061
rect 147722 175021 147728 175033
rect 154000 175021 154006 175033
rect 154058 175021 154064 175073
rect 645136 174873 645142 174925
rect 645194 174913 645200 174925
rect 649552 174913 649558 174925
rect 645194 174885 649558 174913
rect 645194 174873 645200 174885
rect 649552 174873 649558 174885
rect 649610 174873 649616 174925
rect 149200 174207 149206 174259
rect 149258 174247 149264 174259
rect 186256 174247 186262 174259
rect 149258 174219 186262 174247
rect 149258 174207 149264 174219
rect 186256 174207 186262 174219
rect 186314 174207 186320 174259
rect 148912 174059 148918 174111
rect 148970 174099 148976 174111
rect 149392 174099 149398 174111
rect 148970 174071 149398 174099
rect 148970 174059 148976 174071
rect 149392 174059 149398 174071
rect 149450 174059 149456 174111
rect 148528 172727 148534 172779
rect 148586 172767 148592 172779
rect 184528 172767 184534 172779
rect 148586 172739 184534 172767
rect 148586 172727 148592 172739
rect 184528 172727 184534 172739
rect 184586 172727 184592 172779
rect 148720 172653 148726 172705
rect 148778 172693 148784 172705
rect 184624 172693 184630 172705
rect 148778 172665 184630 172693
rect 148778 172653 148784 172665
rect 184624 172653 184630 172665
rect 184682 172653 184688 172705
rect 148336 172579 148342 172631
rect 148394 172619 148400 172631
rect 184336 172619 184342 172631
rect 148394 172591 184342 172619
rect 148394 172579 148400 172591
rect 184336 172579 184342 172591
rect 184394 172579 184400 172631
rect 149008 172505 149014 172557
rect 149066 172545 149072 172557
rect 184432 172545 184438 172557
rect 149066 172517 184438 172545
rect 149066 172505 149072 172517
rect 184432 172505 184438 172517
rect 184490 172505 184496 172557
rect 645136 171025 645142 171077
rect 645194 171065 645200 171077
rect 649648 171065 649654 171077
rect 645194 171037 649654 171065
rect 645194 171025 645200 171037
rect 649648 171025 649654 171037
rect 649706 171025 649712 171077
rect 674800 170285 674806 170337
rect 674858 170325 674864 170337
rect 676048 170325 676054 170337
rect 674858 170297 676054 170325
rect 674858 170285 674864 170297
rect 676048 170285 676054 170297
rect 676106 170285 676112 170337
rect 675280 169915 675286 169967
rect 675338 169955 675344 169967
rect 676048 169955 676054 169967
rect 675338 169927 676054 169955
rect 675338 169915 675344 169927
rect 676048 169915 676054 169927
rect 676106 169915 676112 169967
rect 148624 169841 148630 169893
rect 148682 169881 148688 169893
rect 184624 169881 184630 169893
rect 148682 169853 184630 169881
rect 148682 169841 148688 169853
rect 184624 169841 184630 169853
rect 184682 169841 184688 169893
rect 148816 169767 148822 169819
rect 148874 169807 148880 169819
rect 184432 169807 184438 169819
rect 148874 169779 184438 169807
rect 148874 169767 148880 169779
rect 184432 169767 184438 169779
rect 184490 169767 184496 169819
rect 148240 169693 148246 169745
rect 148298 169733 148304 169745
rect 184336 169733 184342 169745
rect 148298 169705 184342 169733
rect 148298 169693 148304 169705
rect 184336 169693 184342 169705
rect 184394 169693 184400 169745
rect 149296 169619 149302 169671
rect 149354 169659 149360 169671
rect 184528 169659 184534 169671
rect 149354 169631 184534 169659
rect 149354 169619 149360 169631
rect 184528 169619 184534 169631
rect 184586 169619 184592 169671
rect 645136 168213 645142 168265
rect 645194 168253 645200 168265
rect 649840 168253 649846 168265
rect 645194 168225 649846 168253
rect 645194 168213 645200 168225
rect 649840 168213 649846 168225
rect 649898 168213 649904 168265
rect 674896 167695 674902 167747
rect 674954 167735 674960 167747
rect 676048 167735 676054 167747
rect 674954 167707 676054 167735
rect 674954 167695 674960 167707
rect 676048 167695 676054 167707
rect 676106 167695 676112 167747
rect 675184 167103 675190 167155
rect 675242 167143 675248 167155
rect 676240 167143 676246 167155
rect 675242 167115 676246 167143
rect 675242 167103 675248 167115
rect 676240 167103 676246 167115
rect 676298 167103 676304 167155
rect 674992 167029 674998 167081
rect 675050 167069 675056 167081
rect 676048 167069 676054 167081
rect 675050 167041 676054 167069
rect 675050 167029 675056 167041
rect 676048 167029 676054 167041
rect 676106 167029 676112 167081
rect 148432 166955 148438 167007
rect 148490 166995 148496 167007
rect 184336 166995 184342 167007
rect 148490 166967 184342 166995
rect 148490 166955 148496 166967
rect 184336 166955 184342 166967
rect 184394 166955 184400 167007
rect 149392 166881 149398 166933
rect 149450 166921 149456 166933
rect 184432 166921 184438 166933
rect 149450 166893 184438 166921
rect 149450 166881 149456 166893
rect 184432 166881 184438 166893
rect 184490 166881 184496 166933
rect 154096 166807 154102 166859
rect 154154 166847 154160 166859
rect 184528 166847 184534 166859
rect 154154 166819 184534 166847
rect 154154 166807 154160 166819
rect 184528 166807 184534 166819
rect 184586 166807 184592 166859
rect 148720 166659 148726 166711
rect 148778 166699 148784 166711
rect 149104 166699 149110 166711
rect 148778 166671 149110 166699
rect 148778 166659 148784 166671
rect 149104 166659 149110 166671
rect 149162 166659 149168 166711
rect 674704 166215 674710 166267
rect 674762 166255 674768 166267
rect 676048 166255 676054 166267
rect 674762 166227 676054 166255
rect 674762 166215 674768 166227
rect 676048 166215 676054 166227
rect 676106 166215 676112 166267
rect 646864 164365 646870 164417
rect 646922 164405 646928 164417
rect 676048 164405 676054 164417
rect 646922 164377 676054 164405
rect 646922 164365 646928 164377
rect 676048 164365 676054 164377
rect 676106 164365 676112 164417
rect 647056 164291 647062 164343
rect 647114 164331 647120 164343
rect 676240 164331 676246 164343
rect 647114 164303 676246 164331
rect 647114 164291 647120 164303
rect 676240 164291 676246 164303
rect 676298 164291 676304 164343
rect 646960 164217 646966 164269
rect 647018 164257 647024 164269
rect 676144 164257 676150 164269
rect 647018 164229 676150 164257
rect 647018 164217 647024 164229
rect 676144 164217 676150 164229
rect 676202 164217 676208 164269
rect 182896 164069 182902 164121
rect 182954 164109 182960 164121
rect 185296 164109 185302 164121
rect 182954 164081 185302 164109
rect 182954 164069 182960 164081
rect 185296 164069 185302 164081
rect 185354 164069 185360 164121
rect 159856 163995 159862 164047
rect 159914 164035 159920 164047
rect 184336 164035 184342 164047
rect 159914 164007 184342 164035
rect 159914 163995 159920 164007
rect 184336 163995 184342 164007
rect 184394 163995 184400 164047
rect 165616 163921 165622 163973
rect 165674 163961 165680 163973
rect 184432 163961 184438 163973
rect 165674 163933 184438 163961
rect 165674 163921 165680 163933
rect 184432 163921 184438 163933
rect 184490 163921 184496 163973
rect 151216 163847 151222 163899
rect 151274 163887 151280 163899
rect 184336 163887 184342 163899
rect 151274 163859 184342 163887
rect 151274 163847 151280 163859
rect 184336 163847 184342 163859
rect 184394 163847 184400 163899
rect 645136 163329 645142 163381
rect 645194 163369 645200 163381
rect 649936 163369 649942 163381
rect 645194 163341 649942 163369
rect 645194 163329 645200 163341
rect 649936 163329 649942 163341
rect 649994 163329 650000 163381
rect 162640 161183 162646 161235
rect 162698 161223 162704 161235
rect 184528 161223 184534 161235
rect 162698 161195 184534 161223
rect 162698 161183 162704 161195
rect 184528 161183 184534 161195
rect 184586 161183 184592 161235
rect 168400 161109 168406 161161
rect 168458 161149 168464 161161
rect 184624 161149 184630 161161
rect 168458 161121 184630 161149
rect 168458 161109 168464 161121
rect 184624 161109 184630 161121
rect 184682 161109 184688 161161
rect 675664 161109 675670 161161
rect 675722 161109 675728 161161
rect 171280 161035 171286 161087
rect 171338 161075 171344 161087
rect 184336 161075 184342 161087
rect 171338 161047 184342 161075
rect 171338 161035 171344 161047
rect 184336 161035 184342 161047
rect 184394 161035 184400 161087
rect 174256 160961 174262 161013
rect 174314 161001 174320 161013
rect 184432 161001 184438 161013
rect 174314 160973 184438 161001
rect 174314 160961 174320 160973
rect 184432 160961 184438 160973
rect 184490 160961 184496 161013
rect 675682 160643 675710 161109
rect 675664 160591 675670 160643
rect 675722 160591 675728 160643
rect 670384 160443 670390 160495
rect 670442 160483 670448 160495
rect 675376 160483 675382 160495
rect 670442 160455 675382 160483
rect 670442 160443 670448 160455
rect 675376 160443 675382 160455
rect 675434 160443 675440 160495
rect 645136 159703 645142 159755
rect 645194 159743 645200 159755
rect 650032 159743 650038 159755
rect 645194 159715 650038 159743
rect 645194 159703 645200 159715
rect 650032 159703 650038 159715
rect 650090 159703 650096 159755
rect 146896 159111 146902 159163
rect 146954 159151 146960 159163
rect 151216 159151 151222 159163
rect 146954 159123 151222 159151
rect 146954 159111 146960 159123
rect 151216 159111 151222 159123
rect 151274 159111 151280 159163
rect 151792 158371 151798 158423
rect 151850 158411 151856 158423
rect 184432 158411 184438 158423
rect 151850 158383 184438 158411
rect 151850 158371 151856 158383
rect 184432 158371 184438 158383
rect 184490 158371 184496 158423
rect 174352 158297 174358 158349
rect 174410 158337 174416 158349
rect 184336 158337 184342 158349
rect 174410 158309 184342 158337
rect 174410 158297 174416 158309
rect 184336 158297 184342 158309
rect 184394 158297 184400 158349
rect 179920 158223 179926 158275
rect 179978 158263 179984 158275
rect 184528 158263 184534 158275
rect 179978 158235 184534 158263
rect 179978 158223 179984 158235
rect 184528 158223 184534 158235
rect 184586 158223 184592 158275
rect 177136 158149 177142 158201
rect 177194 158189 177200 158201
rect 184624 158189 184630 158201
rect 177194 158161 184630 158189
rect 177194 158149 177200 158161
rect 184624 158149 184630 158161
rect 184682 158149 184688 158201
rect 674800 157705 674806 157757
rect 674858 157745 674864 157757
rect 675376 157745 675382 157757
rect 674858 157717 675382 157745
rect 674858 157705 674864 157717
rect 675376 157705 675382 157717
rect 675434 157705 675440 157757
rect 674896 157039 674902 157091
rect 674954 157079 674960 157091
rect 675472 157079 675478 157091
rect 674954 157051 675478 157079
rect 674954 157039 674960 157051
rect 675472 157039 675478 157051
rect 675530 157039 675536 157091
rect 675184 156521 675190 156573
rect 675242 156561 675248 156573
rect 675376 156561 675382 156573
rect 675242 156533 675382 156561
rect 675242 156521 675248 156533
rect 675376 156521 675382 156533
rect 675434 156521 675440 156573
rect 645136 156003 645142 156055
rect 645194 156043 645200 156055
rect 650128 156043 650134 156055
rect 645194 156015 650134 156043
rect 645194 156003 645200 156015
rect 650128 156003 650134 156015
rect 650186 156003 650192 156055
rect 674992 155855 674998 155907
rect 675050 155895 675056 155907
rect 675376 155895 675382 155907
rect 675050 155867 675382 155895
rect 675050 155855 675056 155867
rect 675376 155855 675382 155867
rect 675434 155855 675440 155907
rect 149296 155707 149302 155759
rect 149354 155747 149360 155759
rect 174544 155747 174550 155759
rect 149354 155719 174550 155747
rect 149354 155707 149360 155719
rect 174544 155707 174550 155719
rect 174602 155707 174608 155759
rect 148816 155633 148822 155685
rect 148874 155673 148880 155685
rect 180016 155673 180022 155685
rect 148874 155645 180022 155673
rect 148874 155633 148880 155645
rect 180016 155633 180022 155645
rect 180074 155633 180080 155685
rect 148912 155559 148918 155611
rect 148970 155599 148976 155611
rect 149296 155599 149302 155611
rect 148970 155571 149302 155599
rect 148970 155559 148976 155571
rect 149296 155559 149302 155571
rect 149354 155559 149360 155611
rect 149680 155559 149686 155611
rect 149738 155599 149744 155611
rect 182800 155599 182806 155611
rect 149738 155571 182806 155599
rect 149738 155559 149744 155571
rect 182800 155559 182806 155571
rect 182858 155559 182864 155611
rect 151696 155485 151702 155537
rect 151754 155525 151760 155537
rect 184528 155525 184534 155537
rect 151754 155497 184534 155525
rect 151754 155485 151760 155497
rect 184528 155485 184534 155497
rect 184586 155485 184592 155537
rect 658000 155485 658006 155537
rect 658058 155525 658064 155537
rect 670384 155525 670390 155537
rect 658058 155497 670390 155525
rect 658058 155485 658064 155497
rect 670384 155485 670390 155497
rect 670442 155485 670448 155537
rect 151504 155411 151510 155463
rect 151562 155451 151568 155463
rect 184432 155451 184438 155463
rect 151562 155423 184438 155451
rect 151562 155411 151568 155423
rect 184432 155411 184438 155423
rect 184490 155411 184496 155463
rect 152080 155337 152086 155389
rect 152138 155377 152144 155389
rect 184624 155377 184630 155389
rect 152138 155349 184630 155377
rect 152138 155337 152144 155349
rect 184624 155337 184630 155349
rect 184682 155337 184688 155389
rect 159952 155263 159958 155315
rect 160010 155303 160016 155315
rect 184336 155303 184342 155315
rect 160010 155275 184342 155303
rect 160010 155263 160016 155275
rect 184336 155263 184342 155275
rect 184394 155263 184400 155315
rect 149200 152747 149206 152799
rect 149258 152787 149264 152799
rect 177040 152787 177046 152799
rect 149258 152759 177046 152787
rect 149258 152747 149264 152759
rect 177040 152747 177046 152759
rect 177098 152747 177104 152799
rect 149680 152673 149686 152725
rect 149738 152713 149744 152725
rect 177136 152713 177142 152725
rect 149738 152685 177142 152713
rect 149738 152673 149744 152685
rect 177136 152673 177142 152685
rect 177194 152673 177200 152725
rect 151408 152599 151414 152651
rect 151466 152639 151472 152651
rect 184528 152639 184534 152651
rect 151466 152611 184534 152639
rect 151466 152599 151472 152611
rect 184528 152599 184534 152611
rect 184586 152599 184592 152651
rect 151600 152525 151606 152577
rect 151658 152565 151664 152577
rect 184336 152565 184342 152577
rect 151658 152537 184342 152565
rect 151658 152525 151664 152537
rect 184336 152525 184342 152537
rect 184394 152525 184400 152577
rect 645136 152525 645142 152577
rect 645194 152565 645200 152577
rect 650224 152565 650230 152577
rect 645194 152537 650230 152565
rect 645194 152525 645200 152537
rect 650224 152525 650230 152537
rect 650282 152525 650288 152577
rect 151984 152451 151990 152503
rect 152042 152491 152048 152503
rect 184432 152491 184438 152503
rect 152042 152463 184438 152491
rect 152042 152451 152048 152463
rect 184432 152451 184438 152463
rect 184490 152451 184496 152503
rect 149200 151785 149206 151837
rect 149258 151825 149264 151837
rect 159952 151825 159958 151837
rect 149258 151797 159958 151825
rect 149258 151785 149264 151797
rect 159952 151785 159958 151797
rect 160010 151785 160016 151837
rect 674704 151415 674710 151467
rect 674762 151455 674768 151467
rect 675376 151455 675382 151467
rect 674762 151427 675382 151455
rect 674762 151415 674768 151427
rect 675376 151415 675382 151427
rect 675434 151415 675440 151467
rect 149200 149861 149206 149913
rect 149258 149901 149264 149913
rect 174160 149901 174166 149913
rect 149258 149873 174166 149901
rect 149258 149861 149264 149873
rect 174160 149861 174166 149873
rect 174218 149861 174224 149913
rect 149680 149787 149686 149839
rect 149738 149827 149744 149839
rect 179920 149827 179926 149839
rect 149738 149799 179926 149827
rect 149738 149787 149744 149799
rect 179920 149787 179926 149799
rect 179978 149787 179984 149839
rect 151312 149713 151318 149765
rect 151370 149753 151376 149765
rect 184336 149753 184342 149765
rect 151370 149725 184342 149753
rect 151370 149713 151376 149725
rect 184336 149713 184342 149725
rect 184394 149713 184400 149765
rect 151888 149639 151894 149691
rect 151946 149679 151952 149691
rect 184432 149679 184438 149691
rect 151946 149651 184438 149679
rect 151946 149639 151952 149651
rect 184432 149639 184438 149651
rect 184490 149639 184496 149691
rect 154192 149565 154198 149617
rect 154250 149605 154256 149617
rect 184528 149605 184534 149617
rect 154250 149577 184534 149605
rect 154250 149565 154256 149577
rect 184528 149565 184534 149577
rect 184586 149565 184592 149617
rect 157072 149491 157078 149543
rect 157130 149531 157136 149543
rect 184336 149531 184342 149543
rect 157130 149503 184342 149531
rect 157130 149491 157136 149503
rect 184336 149491 184342 149503
rect 184394 149491 184400 149543
rect 645136 148159 645142 148211
rect 645194 148199 645200 148211
rect 650320 148199 650326 148211
rect 645194 148171 650326 148199
rect 645194 148159 645200 148171
rect 650320 148159 650326 148171
rect 650378 148159 650384 148211
rect 149200 146975 149206 147027
rect 149258 147015 149264 147027
rect 168400 147015 168406 147027
rect 149258 146987 168406 147015
rect 149258 146975 149264 146987
rect 168400 146975 168406 146987
rect 168458 146975 168464 147027
rect 149680 146901 149686 146953
rect 149738 146941 149744 146953
rect 171568 146941 171574 146953
rect 149738 146913 171574 146941
rect 149738 146901 149744 146913
rect 171568 146901 171574 146913
rect 171626 146901 171632 146953
rect 182992 146827 182998 146879
rect 183050 146867 183056 146879
rect 186736 146867 186742 146879
rect 183050 146839 186742 146867
rect 183050 146827 183056 146839
rect 186736 146827 186742 146839
rect 186794 146827 186800 146879
rect 165712 146753 165718 146805
rect 165770 146793 165776 146805
rect 184336 146793 184342 146805
rect 165770 146765 184342 146793
rect 165770 146753 165776 146765
rect 184336 146753 184342 146765
rect 184394 146753 184400 146805
rect 180112 146679 180118 146731
rect 180170 146719 180176 146731
rect 185392 146719 185398 146731
rect 180170 146691 185398 146719
rect 180170 146679 180176 146691
rect 185392 146679 185398 146691
rect 185450 146679 185456 146731
rect 152176 146605 152182 146657
rect 152234 146645 152240 146657
rect 184432 146645 184438 146657
rect 152234 146617 184438 146645
rect 152234 146605 152240 146617
rect 184432 146605 184438 146617
rect 184490 146605 184496 146657
rect 148624 145495 148630 145547
rect 148682 145495 148688 145547
rect 147856 145421 147862 145473
rect 147914 145461 147920 145473
rect 148336 145461 148342 145473
rect 147914 145433 148342 145461
rect 147914 145421 147920 145433
rect 148336 145421 148342 145433
rect 148394 145421 148400 145473
rect 148336 145273 148342 145325
rect 148394 145313 148400 145325
rect 148642 145313 148670 145495
rect 148394 145285 148670 145313
rect 148394 145273 148400 145285
rect 149200 144089 149206 144141
rect 149258 144129 149264 144141
rect 162928 144129 162934 144141
rect 149258 144101 162934 144129
rect 149258 144089 149264 144101
rect 162928 144089 162934 144101
rect 162986 144089 162992 144141
rect 149680 144015 149686 144067
rect 149738 144055 149744 144067
rect 165616 144055 165622 144067
rect 149738 144027 165622 144055
rect 149738 144015 149744 144027
rect 165616 144015 165622 144027
rect 165674 144015 165680 144067
rect 162832 143941 162838 143993
rect 162890 143981 162896 143993
rect 184528 143981 184534 143993
rect 162890 143953 184534 143981
rect 162890 143941 162896 143953
rect 184528 143941 184534 143953
rect 184586 143941 184592 143993
rect 168592 143867 168598 143919
rect 168650 143907 168656 143919
rect 184432 143907 184438 143919
rect 168650 143879 184438 143907
rect 168650 143867 168656 143879
rect 184432 143867 184438 143879
rect 184490 143867 184496 143919
rect 171472 143793 171478 143845
rect 171530 143833 171536 143845
rect 184336 143833 184342 143845
rect 171530 143805 184342 143833
rect 171530 143793 171536 143805
rect 184336 143793 184342 143805
rect 184394 143793 184400 143845
rect 177328 143719 177334 143771
rect 177386 143759 177392 143771
rect 184624 143759 184630 143771
rect 177386 143731 184630 143759
rect 177386 143719 177392 143731
rect 184624 143719 184630 143731
rect 184682 143719 184688 143771
rect 149680 142313 149686 142365
rect 149738 142353 149744 142365
rect 159856 142353 159862 142365
rect 149738 142325 159862 142353
rect 149738 142313 149744 142325
rect 159856 142313 159862 142325
rect 159914 142313 159920 142365
rect 149200 142239 149206 142291
rect 149258 142279 149264 142291
rect 156976 142279 156982 142291
rect 149258 142251 156982 142279
rect 149258 142239 149264 142251
rect 156976 142239 156982 142251
rect 157034 142239 157040 142291
rect 148816 141203 148822 141255
rect 148874 141243 148880 141255
rect 154096 141243 154102 141255
rect 148874 141215 154102 141243
rect 148874 141203 148880 141215
rect 154096 141203 154102 141215
rect 154154 141203 154160 141255
rect 154288 141055 154294 141107
rect 154346 141095 154352 141107
rect 184528 141095 184534 141107
rect 154346 141067 184534 141095
rect 154346 141055 154352 141067
rect 184528 141055 184534 141067
rect 184586 141055 184592 141107
rect 157168 140981 157174 141033
rect 157226 141021 157232 141033
rect 184432 141021 184438 141033
rect 157226 140993 184438 141021
rect 157226 140981 157232 140993
rect 184432 140981 184438 140993
rect 184490 140981 184496 141033
rect 160048 140907 160054 140959
rect 160106 140947 160112 140959
rect 184336 140947 184342 140959
rect 160106 140919 184342 140947
rect 160106 140907 160112 140919
rect 184336 140907 184342 140919
rect 184394 140907 184400 140959
rect 147088 140167 147094 140219
rect 147146 140207 147152 140219
rect 151120 140207 151126 140219
rect 147146 140179 151126 140207
rect 147146 140167 147152 140179
rect 151120 140167 151126 140179
rect 151178 140167 151184 140219
rect 149200 138243 149206 138295
rect 149258 138283 149264 138295
rect 165520 138283 165526 138295
rect 149258 138255 165526 138283
rect 149258 138243 149264 138255
rect 165520 138243 165526 138255
rect 165578 138243 165584 138295
rect 149200 135431 149206 135483
rect 149258 135471 149264 135483
rect 159760 135471 159766 135483
rect 149258 135443 159766 135471
rect 149258 135431 149264 135443
rect 159760 135431 159766 135443
rect 159818 135431 159824 135483
rect 149680 135357 149686 135409
rect 149738 135397 149744 135409
rect 162640 135397 162646 135409
rect 149738 135369 162646 135397
rect 149738 135357 149744 135369
rect 162640 135357 162646 135369
rect 162698 135357 162704 135409
rect 162736 135283 162742 135335
rect 162794 135323 162800 135335
rect 184528 135323 184534 135335
rect 162794 135295 184534 135323
rect 162794 135283 162800 135295
rect 184528 135283 184534 135295
rect 184586 135283 184592 135335
rect 165808 135209 165814 135261
rect 165866 135249 165872 135261
rect 184432 135249 184438 135261
rect 165866 135221 184438 135249
rect 165866 135209 165872 135221
rect 184432 135209 184438 135221
rect 184490 135209 184496 135261
rect 149488 135135 149494 135187
rect 149546 135175 149552 135187
rect 149680 135175 149686 135187
rect 149546 135147 149686 135175
rect 149546 135135 149552 135147
rect 149680 135135 149686 135147
rect 149738 135135 149744 135187
rect 174448 135135 174454 135187
rect 174506 135175 174512 135187
rect 184336 135175 184342 135187
rect 174506 135147 184342 135175
rect 174506 135135 174512 135147
rect 184336 135135 184342 135147
rect 184394 135135 184400 135187
rect 174544 133951 174550 134003
rect 174602 133991 174608 134003
rect 185680 133991 185686 134003
rect 174602 133963 185686 133991
rect 174602 133951 174608 133963
rect 185680 133951 185686 133963
rect 185738 133951 185744 134003
rect 159952 133877 159958 133929
rect 160010 133917 160016 133929
rect 185584 133917 185590 133929
rect 160010 133889 185590 133917
rect 160010 133877 160016 133889
rect 185584 133877 185590 133889
rect 185642 133877 185648 133929
rect 149392 132545 149398 132597
rect 149450 132585 149456 132597
rect 171280 132585 171286 132597
rect 149450 132557 171286 132585
rect 149450 132545 149456 132557
rect 171280 132545 171286 132557
rect 171338 132545 171344 132597
rect 149488 132471 149494 132523
rect 149546 132511 149552 132523
rect 174256 132511 174262 132523
rect 149546 132483 174262 132511
rect 149546 132471 149552 132483
rect 174256 132471 174262 132483
rect 174314 132471 174320 132523
rect 183088 132397 183094 132449
rect 183146 132437 183152 132449
rect 184624 132437 184630 132449
rect 183146 132409 184630 132437
rect 183146 132397 183152 132409
rect 184624 132397 184630 132409
rect 184682 132397 184688 132449
rect 168496 132323 168502 132375
rect 168554 132363 168560 132375
rect 184528 132363 184534 132375
rect 168554 132335 184534 132363
rect 168554 132323 168560 132335
rect 184528 132323 184534 132335
rect 184586 132323 184592 132375
rect 171376 132249 171382 132301
rect 171434 132289 171440 132301
rect 184336 132289 184342 132301
rect 171434 132261 184342 132289
rect 171434 132249 171440 132261
rect 184336 132249 184342 132261
rect 184394 132249 184400 132301
rect 156880 132175 156886 132227
rect 156938 132215 156944 132227
rect 184432 132215 184438 132227
rect 156938 132187 184438 132215
rect 156938 132175 156944 132187
rect 184432 132175 184438 132187
rect 184490 132175 184496 132227
rect 147184 130251 147190 130303
rect 147242 130291 147248 130303
rect 151120 130291 151126 130303
rect 147242 130263 151126 130291
rect 147242 130251 147248 130263
rect 151120 130251 151126 130263
rect 151178 130251 151184 130303
rect 655312 130103 655318 130155
rect 655370 130143 655376 130155
rect 676144 130143 676150 130155
rect 655370 130115 676150 130143
rect 655370 130103 655376 130115
rect 676144 130103 676150 130115
rect 676202 130103 676208 130155
rect 655216 129955 655222 130007
rect 655274 129995 655280 130007
rect 676240 129995 676246 130007
rect 655274 129967 676246 129995
rect 655274 129955 655280 129967
rect 676240 129955 676246 129967
rect 676298 129955 676304 130007
rect 655120 129807 655126 129859
rect 655178 129847 655184 129859
rect 676336 129847 676342 129859
rect 655178 129819 676342 129847
rect 655178 129807 655184 129819
rect 676336 129807 676342 129819
rect 676394 129807 676400 129859
rect 645712 129585 645718 129637
rect 645770 129625 645776 129637
rect 676240 129625 676246 129637
rect 645770 129597 676246 129625
rect 645770 129585 645776 129597
rect 676240 129585 676246 129597
rect 676298 129585 676304 129637
rect 149296 129511 149302 129563
rect 149354 129551 149360 129563
rect 184624 129551 184630 129563
rect 149354 129523 184630 129551
rect 149354 129511 149360 129523
rect 184624 129511 184630 129523
rect 184682 129511 184688 129563
rect 149200 129437 149206 129489
rect 149258 129477 149264 129489
rect 184432 129477 184438 129489
rect 149258 129449 184438 129477
rect 149258 129437 149264 129449
rect 184432 129437 184438 129449
rect 184490 129437 184496 129489
rect 148240 129363 148246 129415
rect 148298 129403 148304 129415
rect 148432 129403 148438 129415
rect 148298 129375 148438 129403
rect 148298 129363 148304 129375
rect 148432 129363 148438 129375
rect 148490 129363 148496 129415
rect 149584 129363 149590 129415
rect 149642 129403 149648 129415
rect 184528 129403 184534 129415
rect 149642 129375 184534 129403
rect 149642 129363 149648 129375
rect 184528 129363 184534 129375
rect 184586 129363 184592 129415
rect 154000 129289 154006 129341
rect 154058 129329 154064 129341
rect 184336 129329 184342 129341
rect 154058 129301 184342 129329
rect 154058 129289 154064 129301
rect 184336 129289 184342 129301
rect 184394 129289 184400 129341
rect 646480 126847 646486 126899
rect 646538 126887 646544 126899
rect 676240 126887 676246 126899
rect 646538 126859 676246 126887
rect 646538 126847 646544 126859
rect 676240 126847 676246 126859
rect 676298 126847 676304 126899
rect 646576 126773 646582 126825
rect 646634 126813 646640 126825
rect 676144 126813 676150 126825
rect 646634 126785 676150 126813
rect 646634 126773 646640 126785
rect 676144 126773 676150 126785
rect 676202 126773 676208 126825
rect 674128 126699 674134 126751
rect 674186 126739 674192 126751
rect 676048 126739 676054 126751
rect 674186 126711 676054 126739
rect 674186 126699 674192 126711
rect 676048 126699 676054 126711
rect 676106 126699 676112 126751
rect 149008 126625 149014 126677
rect 149066 126665 149072 126677
rect 184432 126665 184438 126677
rect 149066 126637 184438 126665
rect 149066 126625 149072 126637
rect 184432 126625 184438 126637
rect 184490 126625 184496 126677
rect 148720 126551 148726 126603
rect 148778 126591 148784 126603
rect 184528 126591 184534 126603
rect 148778 126563 184534 126591
rect 148778 126551 148784 126563
rect 184528 126551 184534 126563
rect 184586 126551 184592 126603
rect 149680 126477 149686 126529
rect 149738 126517 149744 126529
rect 184336 126517 184342 126529
rect 149738 126489 184342 126517
rect 149738 126477 149744 126489
rect 184336 126477 184342 126489
rect 184394 126477 184400 126529
rect 674224 124627 674230 124679
rect 674282 124667 674288 124679
rect 676048 124667 676054 124679
rect 674282 124639 676054 124667
rect 674282 124627 674288 124639
rect 676048 124627 676054 124639
rect 676106 124627 676112 124679
rect 674032 124035 674038 124087
rect 674090 124075 674096 124087
rect 675952 124075 675958 124087
rect 674090 124047 675958 124075
rect 674090 124035 674096 124047
rect 675952 124035 675958 124047
rect 676010 124035 676016 124087
rect 674608 123961 674614 124013
rect 674666 124001 674672 124013
rect 676048 124001 676054 124013
rect 674666 123973 676054 124001
rect 674666 123961 674672 123973
rect 676048 123961 676054 123973
rect 676106 123961 676112 124013
rect 675184 123887 675190 123939
rect 675242 123927 675248 123939
rect 676240 123927 676246 123939
rect 675242 123899 676246 123927
rect 675242 123887 675248 123899
rect 676240 123887 676246 123899
rect 676298 123887 676304 123939
rect 148624 123813 148630 123865
rect 148682 123853 148688 123865
rect 184336 123853 184342 123865
rect 148682 123825 184342 123853
rect 148682 123813 148688 123825
rect 184336 123813 184342 123825
rect 184394 123813 184400 123865
rect 148432 123739 148438 123791
rect 148490 123779 148496 123791
rect 184432 123779 184438 123791
rect 148490 123751 184438 123779
rect 148490 123739 148496 123751
rect 184432 123739 184438 123751
rect 184490 123739 184496 123791
rect 147856 123665 147862 123717
rect 147914 123705 147920 123717
rect 184336 123705 184342 123717
rect 147914 123677 184342 123705
rect 147914 123665 147920 123677
rect 184336 123665 184342 123677
rect 184394 123665 184400 123717
rect 148336 123591 148342 123643
rect 148394 123631 148400 123643
rect 184528 123631 184534 123643
rect 148394 123603 184534 123631
rect 148394 123591 148400 123603
rect 184528 123591 184534 123603
rect 184586 123591 184592 123643
rect 179920 123517 179926 123569
rect 179978 123557 179984 123569
rect 186160 123557 186166 123569
rect 179978 123529 186166 123557
rect 179978 123517 179984 123529
rect 186160 123517 186166 123529
rect 186218 123517 186224 123569
rect 674416 122111 674422 122163
rect 674474 122151 674480 122163
rect 676048 122151 676054 122163
rect 674474 122123 676054 122151
rect 674474 122111 674480 122123
rect 676048 122111 676054 122123
rect 676106 122111 676112 122163
rect 674704 121149 674710 121201
rect 674762 121189 674768 121201
rect 676048 121189 676054 121201
rect 674762 121161 676054 121189
rect 674762 121149 674768 121161
rect 676048 121149 676054 121161
rect 676106 121149 676112 121201
rect 674320 121075 674326 121127
rect 674378 121115 674384 121127
rect 676240 121115 676246 121127
rect 674378 121087 676246 121115
rect 674378 121075 674384 121087
rect 676240 121075 676246 121087
rect 676298 121075 676304 121127
rect 674800 121001 674806 121053
rect 674858 121041 674864 121053
rect 676048 121041 676054 121053
rect 674858 121013 676054 121041
rect 674858 121001 674864 121013
rect 676048 121001 676054 121013
rect 676106 121001 676112 121053
rect 147952 120927 147958 120979
rect 148010 120967 148016 120979
rect 184432 120967 184438 120979
rect 148010 120939 184438 120967
rect 148010 120927 148016 120939
rect 184432 120927 184438 120939
rect 184490 120927 184496 120979
rect 148240 120853 148246 120905
rect 148298 120893 148304 120905
rect 184528 120893 184534 120905
rect 148298 120865 184534 120893
rect 148298 120853 148304 120865
rect 184528 120853 184534 120865
rect 184586 120853 184592 120905
rect 171568 120779 171574 120831
rect 171626 120819 171632 120831
rect 184624 120819 184630 120831
rect 171626 120791 184630 120819
rect 171626 120779 171632 120791
rect 184624 120779 184630 120791
rect 184682 120779 184688 120831
rect 174160 120705 174166 120757
rect 174218 120745 174224 120757
rect 184336 120745 184342 120757
rect 174218 120717 184342 120745
rect 174218 120705 174224 120717
rect 184336 120705 184342 120717
rect 184394 120705 184400 120757
rect 647824 118337 647830 118389
rect 647882 118377 647888 118389
rect 676240 118377 676246 118389
rect 647882 118349 676246 118377
rect 647882 118337 647888 118349
rect 676240 118337 676246 118349
rect 676298 118337 676304 118389
rect 149392 118263 149398 118315
rect 149450 118303 149456 118315
rect 168496 118303 168502 118315
rect 149450 118275 168502 118303
rect 149450 118263 149456 118275
rect 168496 118263 168502 118275
rect 168554 118263 168560 118315
rect 149488 118189 149494 118241
rect 149546 118229 149552 118241
rect 174352 118229 174358 118241
rect 149546 118201 174358 118229
rect 149546 118189 149552 118201
rect 174352 118189 174358 118201
rect 174410 118189 174416 118241
rect 647920 118189 647926 118241
rect 647978 118229 647984 118241
rect 676144 118229 676150 118241
rect 647978 118201 676150 118229
rect 647978 118189 647984 118201
rect 676144 118189 676150 118201
rect 676202 118189 676208 118241
rect 149392 118115 149398 118167
rect 149450 118155 149456 118167
rect 182896 118155 182902 118167
rect 149450 118127 182902 118155
rect 149450 118115 149456 118127
rect 182896 118115 182902 118127
rect 182954 118115 182960 118167
rect 645232 118115 645238 118167
rect 645290 118155 645296 118167
rect 676048 118155 676054 118167
rect 645290 118127 676054 118155
rect 645290 118115 645296 118127
rect 676048 118115 676054 118127
rect 676106 118115 676112 118167
rect 159856 118041 159862 118093
rect 159914 118081 159920 118093
rect 184624 118081 184630 118093
rect 159914 118053 184630 118081
rect 159914 118041 159920 118053
rect 184624 118041 184630 118053
rect 184682 118041 184688 118093
rect 162928 117967 162934 118019
rect 162986 118007 162992 118019
rect 184528 118007 184534 118019
rect 162986 117979 184534 118007
rect 162986 117967 162992 117979
rect 184528 117967 184534 117979
rect 184586 117967 184592 118019
rect 165616 117893 165622 117945
rect 165674 117933 165680 117945
rect 184432 117933 184438 117945
rect 165674 117905 184438 117933
rect 165674 117893 165680 117905
rect 184432 117893 184438 117905
rect 184490 117893 184496 117945
rect 168400 117819 168406 117871
rect 168458 117859 168464 117871
rect 184336 117859 184342 117871
rect 168458 117831 184342 117859
rect 168458 117819 168464 117831
rect 184336 117819 184342 117831
rect 184394 117819 184400 117871
rect 675088 115377 675094 115429
rect 675146 115417 675152 115429
rect 675280 115417 675286 115429
rect 675146 115389 675286 115417
rect 675146 115377 675152 115389
rect 675280 115377 675286 115389
rect 675338 115377 675344 115429
rect 149392 115303 149398 115355
rect 149450 115343 149456 115355
rect 165712 115343 165718 115355
rect 149450 115315 165718 115343
rect 149450 115303 149456 115315
rect 165712 115303 165718 115315
rect 165770 115303 165776 115355
rect 149488 115229 149494 115281
rect 149546 115269 149552 115281
rect 179920 115269 179926 115281
rect 149546 115241 179926 115269
rect 149546 115229 149552 115241
rect 179920 115229 179926 115241
rect 179978 115229 179984 115281
rect 647920 115229 647926 115281
rect 647978 115269 647984 115281
rect 665296 115269 665302 115281
rect 647978 115241 665302 115269
rect 647978 115229 647984 115241
rect 665296 115229 665302 115241
rect 665354 115229 665360 115281
rect 151216 115155 151222 115207
rect 151274 115195 151280 115207
rect 184528 115195 184534 115207
rect 151274 115167 184534 115195
rect 151274 115155 151280 115167
rect 184528 115155 184534 115167
rect 184586 115155 184592 115207
rect 663760 115155 663766 115207
rect 663818 115195 663824 115207
rect 665200 115195 665206 115207
rect 663818 115167 665206 115195
rect 663818 115155 663824 115167
rect 665200 115155 665206 115167
rect 665258 115155 665264 115207
rect 154096 115081 154102 115133
rect 154154 115121 154160 115133
rect 184432 115121 184438 115133
rect 154154 115093 184438 115121
rect 154154 115081 154160 115093
rect 184432 115081 184438 115093
rect 184490 115081 184496 115133
rect 156976 115007 156982 115059
rect 157034 115047 157040 115059
rect 184336 115047 184342 115059
rect 157034 115019 184342 115047
rect 157034 115007 157040 115019
rect 184336 115007 184342 115019
rect 184394 115007 184400 115059
rect 674608 114785 674614 114837
rect 674666 114825 674672 114837
rect 675184 114825 675190 114837
rect 674666 114797 675190 114825
rect 674666 114785 674672 114797
rect 675184 114785 675190 114797
rect 675242 114785 675248 114837
rect 674128 114119 674134 114171
rect 674186 114159 674192 114171
rect 675376 114159 675382 114171
rect 674186 114131 675382 114159
rect 674186 114119 674192 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 148720 113675 148726 113727
rect 148778 113715 148784 113727
rect 149008 113715 149014 113727
rect 148778 113687 149014 113715
rect 148778 113675 148784 113687
rect 149008 113675 149014 113687
rect 149066 113675 149072 113727
rect 149008 113527 149014 113579
rect 149066 113567 149072 113579
rect 149200 113567 149206 113579
rect 149066 113539 149206 113567
rect 149066 113527 149072 113539
rect 149200 113527 149206 113539
rect 149258 113527 149264 113579
rect 149392 112861 149398 112913
rect 149450 112901 149456 112913
rect 159856 112901 159862 112913
rect 149450 112873 159862 112901
rect 149450 112861 149456 112873
rect 159856 112861 159862 112873
rect 159914 112861 159920 112913
rect 674224 112491 674230 112543
rect 674282 112531 674288 112543
rect 675376 112531 675382 112543
rect 674282 112503 675382 112531
rect 674282 112491 674288 112503
rect 675376 112491 675382 112503
rect 675434 112491 675440 112543
rect 149488 112343 149494 112395
rect 149546 112383 149552 112395
rect 162736 112383 162742 112395
rect 149546 112355 162742 112383
rect 149546 112343 149552 112355
rect 162736 112343 162742 112355
rect 162794 112343 162800 112395
rect 182800 112269 182806 112321
rect 182858 112309 182864 112321
rect 184336 112309 184342 112321
rect 182858 112281 184342 112309
rect 182858 112269 182864 112281
rect 184336 112269 184342 112281
rect 184394 112269 184400 112321
rect 665200 112269 665206 112321
rect 665258 112309 665264 112321
rect 675088 112309 675094 112321
rect 665258 112281 675094 112309
rect 665258 112269 665264 112281
rect 675088 112269 675094 112281
rect 675146 112269 675152 112321
rect 180016 112195 180022 112247
rect 180074 112235 180080 112247
rect 184432 112235 184438 112247
rect 180074 112207 184438 112235
rect 180074 112195 180080 112207
rect 184432 112195 184438 112207
rect 184490 112195 184496 112247
rect 177136 112121 177142 112173
rect 177194 112161 177200 112173
rect 184528 112161 184534 112173
rect 177194 112133 184534 112161
rect 177194 112121 177200 112133
rect 184528 112121 184534 112133
rect 184586 112121 184592 112173
rect 674032 111677 674038 111729
rect 674090 111717 674096 111729
rect 675376 111717 675382 111729
rect 674090 111689 675382 111717
rect 674090 111677 674096 111689
rect 675376 111677 675382 111689
rect 675434 111677 675440 111729
rect 674416 111307 674422 111359
rect 674474 111347 674480 111359
rect 675376 111347 675382 111359
rect 674474 111319 675382 111347
rect 674474 111307 674480 111319
rect 675376 111307 675382 111319
rect 675434 111307 675440 111359
rect 674704 110641 674710 110693
rect 674762 110681 674768 110693
rect 675376 110681 675382 110693
rect 674762 110653 675382 110681
rect 674762 110641 674768 110653
rect 675376 110641 675382 110653
rect 675434 110641 675440 110693
rect 149392 109531 149398 109583
rect 149450 109571 149456 109583
rect 156880 109571 156886 109583
rect 149450 109543 156886 109571
rect 149450 109531 149456 109543
rect 156880 109531 156886 109543
rect 156938 109531 156944 109583
rect 165520 109383 165526 109435
rect 165578 109423 165584 109435
rect 184336 109423 184342 109435
rect 165578 109395 184342 109423
rect 165578 109383 165584 109395
rect 184336 109383 184342 109395
rect 184394 109383 184400 109435
rect 177040 109309 177046 109361
rect 177098 109349 177104 109361
rect 184432 109349 184438 109361
rect 177098 109321 184438 109349
rect 177098 109309 177104 109321
rect 184432 109309 184438 109321
rect 184490 109309 184496 109361
rect 147664 108347 147670 108399
rect 147722 108387 147728 108399
rect 154000 108387 154006 108399
rect 147722 108359 154006 108387
rect 147722 108347 147728 108359
rect 154000 108347 154006 108359
rect 154058 108347 154064 108399
rect 674320 107311 674326 107363
rect 674378 107351 674384 107363
rect 675376 107351 675382 107363
rect 674378 107323 675382 107351
rect 674378 107311 674384 107323
rect 675376 107311 675382 107323
rect 675434 107311 675440 107363
rect 146992 106571 146998 106623
rect 147050 106611 147056 106623
rect 151216 106611 151222 106623
rect 147050 106583 151222 106611
rect 147050 106571 147056 106583
rect 151216 106571 151222 106583
rect 151274 106571 151280 106623
rect 159760 106497 159766 106549
rect 159818 106537 159824 106549
rect 184528 106537 184534 106549
rect 159818 106509 184534 106537
rect 159818 106497 159824 106509
rect 184528 106497 184534 106509
rect 184586 106497 184592 106549
rect 162640 106423 162646 106475
rect 162698 106463 162704 106475
rect 184336 106463 184342 106475
rect 162698 106435 184342 106463
rect 162698 106423 162704 106435
rect 184336 106423 184342 106435
rect 184394 106423 184400 106475
rect 171280 106349 171286 106401
rect 171338 106389 171344 106401
rect 184624 106389 184630 106401
rect 171338 106361 184630 106389
rect 171338 106349 171344 106361
rect 184624 106349 184630 106361
rect 184682 106349 184688 106401
rect 674800 106349 674806 106401
rect 674858 106389 674864 106401
rect 675376 106389 675382 106401
rect 674858 106361 675382 106389
rect 674858 106349 674864 106361
rect 675376 106349 675382 106361
rect 675434 106349 675440 106401
rect 174256 106275 174262 106327
rect 174314 106315 174320 106327
rect 184432 106315 184438 106327
rect 174314 106287 184438 106315
rect 174314 106275 174320 106287
rect 184432 106275 184438 106287
rect 184490 106275 184496 106327
rect 151120 105091 151126 105143
rect 151178 105131 151184 105143
rect 184720 105131 184726 105143
rect 151178 105103 184726 105131
rect 151178 105091 151184 105103
rect 184720 105091 184726 105103
rect 184778 105091 184784 105143
rect 647920 103759 647926 103811
rect 647978 103799 647984 103811
rect 661168 103799 661174 103811
rect 647978 103771 661174 103799
rect 647978 103759 647984 103771
rect 661168 103759 661174 103771
rect 661226 103759 661232 103811
rect 645712 103685 645718 103737
rect 645770 103725 645776 103737
rect 657520 103725 657526 103737
rect 645770 103697 657526 103725
rect 645770 103685 645776 103697
rect 657520 103685 657526 103697
rect 657578 103685 657584 103737
rect 148912 103611 148918 103663
rect 148970 103651 148976 103663
rect 184432 103651 184438 103663
rect 148970 103623 184438 103651
rect 148970 103611 148976 103623
rect 184432 103611 184438 103623
rect 184490 103611 184496 103663
rect 148816 103537 148822 103589
rect 148874 103577 148880 103589
rect 184336 103577 184342 103589
rect 148874 103549 184342 103577
rect 148874 103537 148880 103549
rect 184336 103537 184342 103549
rect 184394 103537 184400 103589
rect 149296 103463 149302 103515
rect 149354 103503 149360 103515
rect 184528 103503 184534 103515
rect 149354 103475 184534 103503
rect 149354 103463 149360 103475
rect 184528 103463 184534 103475
rect 184586 103463 184592 103515
rect 645136 102057 645142 102109
rect 645194 102097 645200 102109
rect 652432 102097 652438 102109
rect 645194 102069 652438 102097
rect 645194 102057 645200 102069
rect 652432 102057 652438 102069
rect 652490 102057 652496 102109
rect 149392 100799 149398 100851
rect 149450 100839 149456 100851
rect 168400 100839 168406 100851
rect 149450 100811 168406 100839
rect 149450 100799 149456 100811
rect 168400 100799 168406 100811
rect 168458 100799 168464 100851
rect 148144 100725 148150 100777
rect 148202 100765 148208 100777
rect 184528 100765 184534 100777
rect 148202 100737 184534 100765
rect 148202 100725 148208 100737
rect 184528 100725 184534 100737
rect 184586 100725 184592 100777
rect 149200 100651 149206 100703
rect 149258 100691 149264 100703
rect 184624 100691 184630 100703
rect 149258 100663 184630 100691
rect 149258 100651 149264 100663
rect 184624 100651 184630 100663
rect 184682 100651 184688 100703
rect 149104 100577 149110 100629
rect 149162 100617 149168 100629
rect 184336 100617 184342 100629
rect 149162 100589 184342 100617
rect 149162 100577 149168 100589
rect 184336 100577 184342 100589
rect 184394 100577 184400 100629
rect 149680 100503 149686 100555
rect 149738 100543 149744 100555
rect 184432 100543 184438 100555
rect 149738 100515 184438 100543
rect 149738 100503 149744 100515
rect 184432 100503 184438 100515
rect 184490 100503 184496 100555
rect 149392 97987 149398 98039
rect 149450 98027 149456 98039
rect 184240 98027 184246 98039
rect 149450 97999 184246 98027
rect 149450 97987 149456 97999
rect 184240 97987 184246 97999
rect 184298 97987 184304 98039
rect 149488 97913 149494 97965
rect 149546 97953 149552 97965
rect 186160 97953 186166 97965
rect 149546 97925 186166 97953
rect 149546 97913 149552 97925
rect 186160 97913 186166 97925
rect 186218 97913 186224 97965
rect 647920 97913 647926 97965
rect 647978 97953 647984 97965
rect 662512 97953 662518 97965
rect 647978 97925 662518 97953
rect 647978 97913 647984 97925
rect 662512 97913 662518 97925
rect 662570 97913 662576 97965
rect 148720 97839 148726 97891
rect 148778 97879 148784 97891
rect 184336 97879 184342 97891
rect 148778 97851 184342 97879
rect 148778 97839 148784 97851
rect 184336 97839 184342 97851
rect 184394 97839 184400 97891
rect 149008 97765 149014 97817
rect 149066 97805 149072 97817
rect 184432 97805 184438 97817
rect 149066 97777 184438 97805
rect 149066 97765 149072 97777
rect 184432 97765 184438 97777
rect 184490 97765 184496 97817
rect 168496 97691 168502 97743
rect 168554 97731 168560 97743
rect 184528 97731 184534 97743
rect 168554 97703 184534 97731
rect 168554 97691 168560 97703
rect 184528 97691 184534 97703
rect 184586 97691 184592 97743
rect 645424 95915 645430 95967
rect 645482 95955 645488 95967
rect 653680 95955 653686 95967
rect 645482 95927 653686 95955
rect 645482 95915 645488 95927
rect 653680 95915 653686 95927
rect 653738 95915 653744 95967
rect 149488 95101 149494 95153
rect 149546 95141 149552 95153
rect 165520 95141 165526 95153
rect 149546 95113 165526 95141
rect 149546 95101 149552 95113
rect 165520 95101 165526 95113
rect 165578 95101 165584 95153
rect 149392 95027 149398 95079
rect 149450 95067 149456 95079
rect 180016 95067 180022 95079
rect 149450 95039 180022 95067
rect 149450 95027 149456 95039
rect 180016 95027 180022 95039
rect 180074 95027 180080 95079
rect 174352 94879 174358 94931
rect 174410 94919 174416 94931
rect 184336 94919 184342 94931
rect 174410 94891 184342 94919
rect 174410 94879 174416 94891
rect 184336 94879 184342 94891
rect 184394 94879 184400 94931
rect 165712 94731 165718 94783
rect 165770 94771 165776 94783
rect 184336 94771 184342 94783
rect 165770 94743 184342 94771
rect 165770 94731 165776 94743
rect 184336 94731 184342 94743
rect 184394 94731 184400 94783
rect 182896 94657 182902 94709
rect 182954 94697 182960 94709
rect 186256 94697 186262 94709
rect 182954 94669 186262 94697
rect 182954 94657 182960 94669
rect 186256 94657 186262 94669
rect 186314 94657 186320 94709
rect 179920 94583 179926 94635
rect 179978 94623 179984 94635
rect 184624 94623 184630 94635
rect 179978 94595 184630 94623
rect 179978 94583 179984 94595
rect 184624 94583 184630 94595
rect 184682 94583 184688 94635
rect 646768 92659 646774 92711
rect 646826 92699 646832 92711
rect 663088 92699 663094 92711
rect 646826 92671 663094 92699
rect 646826 92659 646832 92671
rect 663088 92659 663094 92671
rect 663146 92659 663152 92711
rect 149392 92363 149398 92415
rect 149450 92403 149456 92415
rect 159568 92403 159574 92415
rect 149450 92375 159574 92403
rect 149450 92363 149456 92375
rect 159568 92363 159574 92375
rect 159626 92363 159632 92415
rect 645520 92363 645526 92415
rect 645578 92403 645584 92415
rect 661744 92403 661750 92415
rect 645578 92375 661750 92403
rect 645578 92363 645584 92375
rect 661744 92363 661750 92375
rect 661802 92363 661808 92415
rect 646480 92289 646486 92341
rect 646538 92329 646544 92341
rect 660688 92329 660694 92341
rect 646538 92301 660694 92329
rect 646538 92289 646544 92301
rect 660688 92289 660694 92301
rect 660746 92289 660752 92341
rect 646864 92215 646870 92267
rect 646922 92255 646928 92267
rect 659824 92255 659830 92267
rect 646922 92227 659830 92255
rect 646922 92215 646928 92227
rect 659824 92215 659830 92227
rect 659882 92215 659888 92267
rect 149488 92141 149494 92193
rect 149546 92181 149552 92193
rect 162352 92181 162358 92193
rect 149546 92153 162358 92181
rect 149546 92141 149552 92153
rect 162352 92141 162358 92153
rect 162410 92141 162416 92193
rect 647152 92141 647158 92193
rect 647210 92181 647216 92193
rect 658864 92181 658870 92193
rect 647210 92153 658870 92181
rect 647210 92141 647216 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 148432 92067 148438 92119
rect 148490 92107 148496 92119
rect 184624 92107 184630 92119
rect 148490 92079 184630 92107
rect 148490 92067 148496 92079
rect 184624 92067 184630 92079
rect 184682 92067 184688 92119
rect 148240 91993 148246 92045
rect 148298 92033 148304 92045
rect 184528 92033 184534 92045
rect 148298 92005 184534 92033
rect 148298 91993 148304 92005
rect 184528 91993 184534 92005
rect 184586 91993 184592 92045
rect 159856 91919 159862 91971
rect 159914 91959 159920 91971
rect 184432 91959 184438 91971
rect 159914 91931 184438 91959
rect 159914 91919 159920 91931
rect 184432 91919 184438 91931
rect 184490 91919 184496 91971
rect 162736 91845 162742 91897
rect 162794 91885 162800 91897
rect 184336 91885 184342 91897
rect 162794 91857 184342 91885
rect 162794 91845 162800 91857
rect 184336 91845 184342 91857
rect 184394 91845 184400 91897
rect 148528 89181 148534 89233
rect 148586 89221 148592 89233
rect 184624 89221 184630 89233
rect 148586 89193 184630 89221
rect 148586 89181 148592 89193
rect 184624 89181 184630 89193
rect 184682 89181 184688 89233
rect 151216 89107 151222 89159
rect 151274 89147 151280 89159
rect 184528 89147 184534 89159
rect 151274 89119 184534 89147
rect 151274 89107 151280 89119
rect 184528 89107 184534 89119
rect 184586 89107 184592 89159
rect 154000 89033 154006 89085
rect 154058 89073 154064 89085
rect 184432 89073 184438 89085
rect 154058 89045 184438 89073
rect 154058 89033 154064 89045
rect 184432 89033 184438 89045
rect 184490 89033 184496 89085
rect 156880 88959 156886 89011
rect 156938 88999 156944 89011
rect 184336 88999 184342 89011
rect 156938 88971 184342 88999
rect 156938 88959 156944 88971
rect 184336 88959 184342 88971
rect 184394 88959 184400 89011
rect 645904 87479 645910 87531
rect 645962 87519 645968 87531
rect 650896 87519 650902 87531
rect 645962 87491 650902 87519
rect 645962 87479 645968 87491
rect 650896 87479 650902 87491
rect 650954 87479 650960 87531
rect 647920 87257 647926 87309
rect 647978 87297 647984 87309
rect 658000 87297 658006 87309
rect 647978 87269 658006 87297
rect 647978 87257 647984 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 149488 87035 149494 87087
rect 149546 87075 149552 87087
rect 156400 87075 156406 87087
rect 149546 87047 156406 87075
rect 149546 87035 149552 87047
rect 156400 87035 156406 87047
rect 156458 87035 156464 87087
rect 647056 87035 647062 87087
rect 647114 87075 647120 87087
rect 663280 87075 663286 87087
rect 647114 87047 663286 87075
rect 647114 87035 647120 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 148720 86443 148726 86495
rect 148778 86483 148784 86495
rect 154096 86483 154102 86495
rect 148778 86455 154102 86483
rect 148778 86443 148784 86455
rect 154096 86443 154102 86455
rect 154154 86443 154160 86495
rect 148336 86369 148342 86421
rect 148394 86409 148400 86421
rect 184432 86409 184438 86421
rect 148394 86381 184438 86409
rect 148394 86369 148400 86381
rect 184432 86369 184438 86381
rect 184490 86369 184496 86421
rect 148624 86295 148630 86347
rect 148682 86335 148688 86347
rect 184528 86335 184534 86347
rect 148682 86307 184534 86335
rect 148682 86295 148688 86307
rect 184528 86295 184534 86307
rect 184586 86295 184592 86347
rect 149584 86221 149590 86273
rect 149642 86261 149648 86273
rect 184336 86261 184342 86273
rect 149642 86233 184342 86261
rect 149642 86221 149648 86233
rect 184336 86221 184342 86233
rect 184394 86221 184400 86273
rect 645904 84149 645910 84201
rect 645962 84189 645968 84201
rect 657040 84189 657046 84201
rect 645962 84161 657046 84189
rect 645962 84149 645968 84161
rect 657040 84149 657046 84161
rect 657098 84149 657104 84201
rect 147088 83557 147094 83609
rect 147146 83597 147152 83609
rect 151120 83597 151126 83609
rect 147146 83569 151126 83597
rect 147146 83557 147152 83569
rect 151120 83557 151126 83569
rect 151178 83557 151184 83609
rect 646768 83557 646774 83609
rect 646826 83597 646832 83609
rect 651760 83597 651766 83609
rect 646826 83569 651766 83597
rect 646826 83557 646832 83569
rect 651760 83557 651766 83569
rect 651818 83557 651824 83609
rect 165520 83483 165526 83535
rect 165578 83523 165584 83535
rect 184432 83523 184438 83535
rect 165578 83495 184438 83523
rect 165578 83483 165584 83495
rect 184432 83483 184438 83495
rect 184490 83483 184496 83535
rect 168400 83409 168406 83461
rect 168458 83449 168464 83461
rect 184336 83449 184342 83461
rect 168458 83421 184342 83449
rect 168458 83409 168464 83421
rect 184336 83409 184342 83421
rect 184394 83409 184400 83461
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 647824 81781 647830 81833
rect 647882 81821 647888 81833
rect 663376 81821 663382 81833
rect 647882 81793 663382 81821
rect 647882 81781 647888 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 657040 81633 657046 81685
rect 657098 81673 657104 81685
rect 658576 81673 658582 81685
rect 657098 81645 658582 81673
rect 657098 81633 657104 81645
rect 658576 81633 658582 81645
rect 658634 81633 658640 81685
rect 647728 81559 647734 81611
rect 647786 81599 647792 81611
rect 662416 81599 662422 81611
rect 647786 81571 662422 81599
rect 647786 81559 647792 81571
rect 662416 81559 662422 81571
rect 662474 81559 662480 81611
rect 660880 80967 660886 81019
rect 660938 81007 660944 81019
rect 668368 81007 668374 81019
rect 660938 80979 668374 81007
rect 660938 80967 660944 80979
rect 668368 80967 668374 80979
rect 668426 80967 668432 81019
rect 647920 80745 647926 80797
rect 647978 80785 647984 80797
rect 662512 80785 662518 80797
rect 647978 80757 662518 80785
rect 647978 80745 647984 80757
rect 662512 80745 662518 80757
rect 662570 80745 662576 80797
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 149680 80597 149686 80649
rect 149738 80637 149744 80649
rect 184432 80637 184438 80649
rect 149738 80609 184438 80637
rect 149738 80597 149744 80609
rect 184432 80597 184438 80609
rect 184490 80597 184496 80649
rect 159568 80523 159574 80575
rect 159626 80563 159632 80575
rect 184528 80563 184534 80575
rect 159626 80535 184534 80563
rect 159626 80523 159632 80535
rect 184528 80523 184534 80535
rect 184586 80523 184592 80575
rect 162352 80449 162358 80501
rect 162410 80489 162416 80501
rect 184336 80489 184342 80501
rect 162410 80461 184342 80489
rect 162410 80449 162416 80461
rect 184336 80449 184342 80461
rect 184394 80449 184400 80501
rect 180016 80375 180022 80427
rect 180074 80415 180080 80427
rect 184624 80415 184630 80427
rect 180074 80387 184630 80415
rect 180074 80375 180080 80387
rect 184624 80375 184630 80387
rect 184682 80375 184688 80427
rect 149200 77711 149206 77763
rect 149258 77751 149264 77763
rect 184336 77751 184342 77763
rect 149258 77723 184342 77751
rect 149258 77711 149264 77723
rect 184336 77711 184342 77723
rect 184394 77711 184400 77763
rect 646960 77711 646966 77763
rect 647018 77751 647024 77763
rect 658288 77751 658294 77763
rect 647018 77723 658294 77751
rect 647018 77711 647024 77723
rect 658288 77711 658294 77723
rect 658346 77711 658352 77763
rect 149296 77637 149302 77689
rect 149354 77677 149360 77689
rect 184432 77677 184438 77689
rect 149354 77649 184438 77677
rect 149354 77637 149360 77649
rect 184432 77637 184438 77649
rect 184490 77637 184496 77689
rect 646576 77637 646582 77689
rect 646634 77677 646640 77689
rect 659440 77677 659446 77689
rect 646634 77649 659446 77677
rect 646634 77637 646640 77649
rect 659440 77637 659446 77649
rect 659498 77637 659504 77689
rect 149392 77563 149398 77615
rect 149450 77603 149456 77615
rect 184528 77603 184534 77615
rect 149450 77575 184534 77603
rect 149450 77563 149456 77575
rect 184528 77563 184534 77575
rect 184586 77563 184592 77615
rect 646672 77563 646678 77615
rect 646730 77603 646736 77615
rect 661744 77603 661750 77615
rect 646730 77575 661750 77603
rect 646730 77563 646736 77575
rect 661744 77563 661750 77575
rect 661802 77563 661808 77615
rect 156400 77489 156406 77541
rect 156458 77529 156464 77541
rect 184624 77529 184630 77541
rect 156458 77501 184630 77529
rect 156458 77489 156464 77501
rect 184624 77489 184630 77501
rect 184682 77489 184688 77541
rect 647920 77489 647926 77541
rect 647978 77529 647984 77541
rect 656944 77529 656950 77541
rect 647978 77501 656950 77529
rect 647978 77489 647984 77501
rect 656944 77489 656950 77501
rect 657002 77489 657008 77541
rect 646000 76083 646006 76135
rect 646058 76123 646064 76135
rect 657520 76123 657526 76135
rect 646058 76095 657526 76123
rect 646058 76083 646064 76095
rect 657520 76083 657526 76095
rect 657578 76083 657584 76135
rect 647056 74899 647062 74951
rect 647114 74939 647120 74951
rect 660112 74939 660118 74951
rect 647114 74911 660118 74939
rect 647114 74899 647120 74911
rect 660112 74899 660118 74911
rect 660170 74899 660176 74951
rect 148432 74825 148438 74877
rect 148490 74865 148496 74877
rect 184528 74865 184534 74877
rect 148490 74837 184534 74865
rect 148490 74825 148496 74837
rect 184528 74825 184534 74837
rect 184586 74825 184592 74877
rect 149104 74751 149110 74803
rect 149162 74791 149168 74803
rect 184624 74791 184630 74803
rect 149162 74763 184630 74791
rect 149162 74751 149168 74763
rect 184624 74751 184630 74763
rect 184682 74751 184688 74803
rect 151120 74677 151126 74729
rect 151178 74717 151184 74729
rect 184432 74717 184438 74729
rect 151178 74689 184438 74717
rect 151178 74677 151184 74689
rect 184432 74677 184438 74689
rect 184490 74677 184496 74729
rect 154096 74603 154102 74655
rect 154154 74643 154160 74655
rect 184336 74643 184342 74655
rect 154154 74615 184342 74643
rect 154154 74603 154160 74615
rect 184336 74603 184342 74615
rect 184394 74603 184400 74655
rect 647920 72087 647926 72139
rect 647978 72127 647984 72139
rect 660688 72127 660694 72139
rect 647978 72099 660694 72127
rect 647978 72087 647984 72099
rect 660688 72087 660694 72099
rect 660746 72087 660752 72139
rect 148240 71939 148246 71991
rect 148298 71979 148304 71991
rect 184432 71979 184438 71991
rect 148298 71951 184438 71979
rect 148298 71939 148304 71951
rect 184432 71939 184438 71951
rect 184490 71939 184496 71991
rect 149680 71865 149686 71917
rect 149738 71905 149744 71917
rect 184528 71905 184534 71917
rect 149738 71877 184534 71905
rect 149738 71865 149744 71877
rect 184528 71865 184534 71877
rect 184586 71865 184592 71917
rect 149584 71791 149590 71843
rect 149642 71831 149648 71843
rect 184336 71831 184342 71843
rect 149642 71803 184342 71831
rect 149642 71791 149648 71803
rect 184336 71791 184342 71803
rect 184394 71791 184400 71843
rect 647920 69423 647926 69475
rect 647978 69463 647984 69475
rect 661456 69463 661462 69475
rect 647978 69435 661462 69463
rect 647978 69423 647984 69435
rect 661456 69423 661462 69435
rect 661514 69423 661520 69475
rect 148816 69053 148822 69105
rect 148874 69093 148880 69105
rect 184336 69093 184342 69105
rect 148874 69065 184342 69093
rect 148874 69053 148880 69065
rect 184336 69053 184342 69065
rect 184394 69053 184400 69105
rect 149200 68979 149206 69031
rect 149258 69019 149264 69031
rect 184432 69019 184438 69031
rect 149258 68991 184438 69019
rect 149258 68979 149264 68991
rect 184432 68979 184438 68991
rect 184490 68979 184496 69031
rect 149584 68905 149590 68957
rect 149642 68945 149648 68957
rect 184336 68945 184342 68957
rect 149642 68917 184342 68945
rect 149642 68905 149648 68917
rect 184336 68905 184342 68917
rect 184394 68905 184400 68957
rect 149296 68831 149302 68883
rect 149354 68871 149360 68883
rect 184528 68871 184534 68883
rect 149354 68843 184534 68871
rect 149354 68831 149360 68843
rect 184528 68831 184534 68843
rect 184586 68831 184592 68883
rect 149104 66167 149110 66219
rect 149162 66207 149168 66219
rect 184528 66207 184534 66219
rect 149162 66179 184534 66207
rect 149162 66167 149168 66179
rect 184528 66167 184534 66179
rect 184586 66167 184592 66219
rect 646000 66167 646006 66219
rect 646058 66207 646064 66219
rect 652336 66207 652342 66219
rect 646058 66179 652342 66207
rect 646058 66167 646064 66179
rect 652336 66167 652342 66179
rect 652394 66167 652400 66219
rect 149392 66093 149398 66145
rect 149450 66133 149456 66145
rect 184624 66133 184630 66145
rect 149450 66105 184630 66133
rect 149450 66093 149456 66105
rect 184624 66093 184630 66105
rect 184682 66093 184688 66145
rect 149488 66019 149494 66071
rect 149546 66059 149552 66071
rect 184432 66059 184438 66071
rect 149546 66031 184438 66059
rect 149546 66019 149552 66031
rect 184432 66019 184438 66031
rect 184490 66019 184496 66071
rect 149008 65945 149014 65997
rect 149066 65985 149072 65997
rect 184336 65985 184342 65997
rect 149066 65957 184342 65985
rect 149066 65945 149072 65957
rect 184336 65945 184342 65957
rect 184394 65945 184400 65997
rect 647920 63577 647926 63629
rect 647978 63617 647984 63629
rect 663184 63617 663190 63629
rect 647978 63589 663190 63617
rect 647978 63577 647984 63589
rect 663184 63577 663190 63589
rect 663242 63577 663248 63629
rect 149392 63281 149398 63333
rect 149450 63321 149456 63333
rect 184624 63321 184630 63333
rect 149450 63293 184630 63321
rect 149450 63281 149456 63293
rect 184624 63281 184630 63293
rect 184682 63281 184688 63333
rect 149584 63207 149590 63259
rect 149642 63247 149648 63259
rect 184528 63247 184534 63259
rect 149642 63219 184534 63247
rect 149642 63207 149648 63219
rect 184528 63207 184534 63219
rect 184586 63207 184592 63259
rect 149200 63133 149206 63185
rect 149258 63173 149264 63185
rect 184336 63173 184342 63185
rect 149258 63145 184342 63173
rect 149258 63133 149264 63145
rect 184336 63133 184342 63145
rect 184394 63133 184400 63185
rect 149296 63059 149302 63111
rect 149354 63099 149360 63111
rect 184432 63099 184438 63111
rect 149354 63071 184438 63099
rect 149354 63059 149360 63071
rect 184432 63059 184438 63071
rect 184490 63059 184496 63111
rect 647920 60987 647926 61039
rect 647978 61027 647984 61039
rect 663472 61027 663478 61039
rect 647978 60999 663478 61027
rect 647978 60987 647984 60999
rect 663472 60987 663478 60999
rect 663530 60987 663536 61039
rect 149392 60395 149398 60447
rect 149450 60435 149456 60447
rect 184432 60435 184438 60447
rect 149450 60407 184438 60435
rect 149450 60395 149456 60407
rect 184432 60395 184438 60407
rect 184490 60395 184496 60447
rect 149488 60321 149494 60373
rect 149546 60361 149552 60373
rect 184336 60361 184342 60373
rect 149546 60333 184342 60361
rect 149546 60321 149552 60333
rect 184336 60321 184342 60333
rect 184394 60321 184400 60373
rect 149296 60247 149302 60299
rect 149354 60287 149360 60299
rect 184528 60287 184534 60299
rect 149354 60259 184534 60287
rect 149354 60247 149360 60259
rect 184528 60247 184534 60259
rect 184586 60247 184592 60299
rect 646000 59063 646006 59115
rect 646058 59103 646064 59115
rect 652240 59103 652246 59115
rect 646058 59075 652246 59103
rect 646058 59063 646064 59075
rect 652240 59063 652246 59075
rect 652298 59063 652304 59115
rect 149392 58989 149398 59041
rect 149450 59029 149456 59041
rect 184336 59029 184342 59041
rect 149450 59001 184342 59029
rect 149450 58989 149456 59001
rect 184336 58989 184342 59001
rect 184394 58989 184400 59041
rect 149392 57509 149398 57561
rect 149450 57549 149456 57561
rect 184336 57549 184342 57561
rect 149450 57521 184342 57549
rect 149450 57509 149456 57521
rect 184336 57509 184342 57521
rect 184394 57509 184400 57561
rect 149392 56177 149398 56229
rect 149450 56217 149456 56229
rect 184432 56217 184438 56229
rect 149450 56189 184438 56217
rect 149450 56177 149456 56189
rect 184432 56177 184438 56189
rect 184490 56177 184496 56229
rect 149488 56103 149494 56155
rect 149546 56143 149552 56155
rect 184336 56143 184342 56155
rect 149546 56115 184342 56143
rect 149546 56103 149552 56115
rect 184336 56103 184342 56115
rect 184394 56103 184400 56155
rect 149680 54623 149686 54675
rect 149738 54663 149744 54675
rect 184336 54663 184342 54675
rect 149738 54635 184342 54663
rect 149738 54623 149744 54635
rect 184336 54623 184342 54635
rect 184394 54623 184400 54675
rect 149392 53217 149398 53269
rect 149450 53257 149456 53269
rect 184336 53257 184342 53269
rect 149450 53229 184342 53257
rect 149450 53217 149456 53229
rect 184336 53217 184342 53229
rect 184394 53217 184400 53269
rect 434896 48111 434902 48163
rect 434954 48151 434960 48163
rect 475696 48151 475702 48163
rect 434954 48123 475702 48151
rect 434954 48111 434960 48123
rect 475696 48111 475702 48123
rect 475754 48111 475760 48163
rect 460336 48037 460342 48089
rect 460394 48077 460400 48089
rect 510352 48077 510358 48089
rect 460394 48049 510358 48077
rect 460394 48037 460400 48049
rect 510352 48037 510358 48049
rect 510410 48037 510416 48089
rect 394576 47963 394582 48015
rect 394634 48003 394640 48015
rect 406768 48003 406774 48015
rect 394634 47975 406774 48003
rect 394634 47963 394640 47975
rect 406768 47963 406774 47975
rect 406826 47963 406832 48015
rect 411856 47963 411862 48015
rect 411914 48003 411920 48015
rect 424048 48003 424054 48015
rect 411914 47975 424054 48003
rect 411914 47963 411920 47975
rect 424048 47963 424054 47975
rect 424106 47963 424112 48015
rect 426160 47963 426166 48015
rect 426218 48003 426224 48015
rect 492976 48003 492982 48015
rect 426218 47975 492982 48003
rect 426218 47963 426224 47975
rect 492976 47963 492982 47975
rect 493034 47963 493040 48015
rect 311056 47889 311062 47941
rect 311114 47929 311120 47941
rect 371920 47929 371926 47941
rect 311114 47901 371926 47929
rect 311114 47889 311120 47901
rect 371920 47889 371926 47901
rect 371978 47889 371984 47941
rect 405520 47889 405526 47941
rect 405578 47929 405584 47941
rect 441328 47929 441334 47941
rect 405578 47901 441334 47929
rect 405578 47889 405584 47901
rect 441328 47889 441334 47901
rect 441386 47889 441392 47941
rect 472240 47889 472246 47941
rect 472298 47929 472304 47941
rect 562480 47929 562486 47941
rect 472298 47901 562486 47929
rect 472298 47889 472304 47901
rect 562480 47889 562486 47901
rect 562538 47889 562544 47941
rect 320176 47815 320182 47867
rect 320234 47855 320240 47867
rect 529264 47855 529270 47867
rect 320234 47827 529270 47855
rect 320234 47815 320240 47827
rect 529264 47815 529270 47827
rect 529322 47815 529328 47867
rect 302896 47741 302902 47793
rect 302954 47781 302960 47793
rect 523888 47781 523894 47793
rect 302954 47753 523894 47781
rect 302954 47741 302960 47753
rect 523888 47741 523894 47753
rect 523946 47741 523952 47793
rect 233680 47667 233686 47719
rect 233738 47707 233744 47719
rect 475504 47707 475510 47719
rect 233738 47679 475510 47707
rect 233738 47667 233744 47679
rect 475504 47667 475510 47679
rect 475562 47667 475568 47719
rect 505360 47667 505366 47719
rect 505418 47707 505424 47719
rect 527920 47707 527926 47719
rect 505418 47679 527926 47707
rect 505418 47667 505424 47679
rect 527920 47667 527926 47679
rect 527978 47667 527984 47719
rect 268528 47593 268534 47645
rect 268586 47633 268592 47645
rect 517360 47633 517366 47645
rect 268586 47605 517366 47633
rect 268586 47593 268592 47605
rect 517360 47593 517366 47605
rect 517418 47593 517424 47645
rect 250960 47519 250966 47571
rect 251018 47559 251024 47571
rect 521200 47559 521206 47571
rect 251018 47531 521206 47559
rect 251018 47519 251024 47531
rect 521200 47519 521206 47531
rect 521258 47519 521264 47571
rect 145360 47075 145366 47127
rect 145418 47115 145424 47127
rect 199120 47115 199126 47127
rect 145418 47087 199126 47115
rect 145418 47075 145424 47087
rect 199120 47075 199126 47087
rect 199178 47075 199184 47127
rect 324304 46261 324310 46313
rect 324362 46301 324368 46313
rect 337456 46301 337462 46313
rect 324362 46273 337462 46301
rect 324362 46261 324368 46273
rect 337456 46261 337462 46273
rect 337514 46261 337520 46313
rect 345616 46261 345622 46313
rect 345674 46301 345680 46313
rect 354832 46301 354838 46313
rect 345674 46273 354838 46301
rect 345674 46261 345680 46273
rect 354832 46261 354838 46273
rect 354890 46261 354896 46313
rect 224560 44633 224566 44685
rect 224618 44673 224624 44685
rect 660880 44673 660886 44685
rect 224618 44645 660886 44673
rect 224618 44633 224624 44645
rect 660880 44633 660886 44645
rect 660938 44633 660944 44685
rect 523888 43967 523894 44019
rect 523946 44007 523952 44019
rect 525904 44007 525910 44019
rect 523946 43979 525910 44007
rect 523946 43967 523952 43979
rect 525904 43967 525910 43979
rect 525962 43967 525968 44019
rect 285808 43227 285814 43279
rect 285866 43267 285872 43279
rect 518704 43267 518710 43279
rect 285866 43239 518710 43267
rect 285866 43227 285872 43239
rect 518704 43227 518710 43239
rect 518762 43227 518768 43279
rect 399856 42339 399862 42391
rect 399914 42379 399920 42391
rect 411856 42379 411862 42391
rect 399914 42351 411862 42379
rect 399914 42339 399920 42351
rect 411856 42339 411862 42351
rect 411914 42339 411920 42391
rect 307216 41969 307222 42021
rect 307274 42009 307280 42021
rect 311056 42009 311062 42021
rect 307274 41981 311062 42009
rect 307274 41969 307280 41981
rect 311056 41969 311062 41981
rect 311114 41969 311120 42021
rect 362032 41969 362038 42021
rect 362090 42009 362096 42021
rect 365968 42009 365974 42021
rect 362090 41981 365974 42009
rect 362090 41969 362096 41981
rect 365968 41969 365974 41981
rect 366026 41969 366032 42021
rect 514000 41747 514006 41799
rect 514058 41787 514064 41799
rect 514864 41787 514870 41799
rect 514058 41759 514870 41787
rect 514058 41747 514064 41759
rect 514864 41747 514870 41759
rect 514922 41747 514928 41799
rect 365872 37381 365878 37433
rect 365930 37421 365936 37433
rect 399856 37421 399862 37433
rect 365930 37393 399862 37421
rect 365930 37381 365936 37393
rect 399856 37381 399862 37393
rect 399914 37381 399920 37433
rect 475504 37381 475510 37433
rect 475562 37421 475568 37433
rect 514000 37421 514006 37433
rect 475562 37393 514006 37421
rect 475562 37381 475568 37393
rect 514000 37381 514006 37393
rect 514058 37381 514064 37433
rect 365968 37307 365974 37359
rect 366026 37347 366032 37359
rect 389200 37347 389206 37359
rect 366026 37319 389206 37347
rect 366026 37307 366032 37319
rect 389200 37307 389206 37319
rect 389258 37307 389264 37359
<< via1 >>
rect 80566 1002267 80618 1002319
rect 82294 1002267 82346 1002319
rect 483670 1002267 483722 1002319
rect 486742 1002267 486794 1002319
rect 535702 991463 535754 991515
rect 538582 991463 538634 991515
rect 388630 990723 388682 990775
rect 389590 990723 389642 990775
rect 240886 982953 240938 983005
rect 241942 982953 241994 983005
rect 292534 982953 292586 983005
rect 296662 982953 296714 983005
rect 40150 961863 40202 961915
rect 60022 961863 60074 961915
rect 653782 960457 653834 960509
rect 679702 960457 679754 960509
rect 655414 892969 655466 893021
rect 676246 892969 676298 893021
rect 655222 892895 655274 892947
rect 676150 892895 676202 892947
rect 655126 892821 655178 892873
rect 676054 892821 676106 892873
rect 673366 892377 673418 892429
rect 676054 892377 676106 892429
rect 670966 891415 671018 891467
rect 676054 891415 676106 891467
rect 670870 890379 670922 890431
rect 676054 890379 676106 890431
rect 674230 887493 674282 887545
rect 676054 887493 676106 887545
rect 675094 887123 675146 887175
rect 676246 887123 676298 887175
rect 675190 887049 675242 887101
rect 676054 887049 676106 887101
rect 674038 885051 674090 885103
rect 676054 885051 676106 885103
rect 674902 884385 674954 884437
rect 676054 884385 676106 884437
rect 674902 884163 674954 884215
rect 676246 884163 676298 884215
rect 674614 883571 674666 883623
rect 676054 883571 676106 883623
rect 675286 882831 675338 882883
rect 679702 882831 679754 882883
rect 675766 882239 675818 882291
rect 680086 882239 680138 882291
rect 674422 881943 674474 881995
rect 676054 881943 676106 881995
rect 674326 881647 674378 881699
rect 680278 881647 680330 881699
rect 649462 881425 649514 881477
rect 679798 881425 679850 881477
rect 655318 881351 655370 881403
rect 675478 881351 675530 881403
rect 674134 880981 674186 881033
rect 674422 880981 674474 881033
rect 674422 880833 674474 880885
rect 675094 880833 675146 880885
rect 675094 880685 675146 880737
rect 680182 880685 680234 880737
rect 674998 879501 675050 879553
rect 679990 879501 680042 879553
rect 674518 878613 674570 878665
rect 675190 878613 675242 878665
rect 675190 878465 675242 878517
rect 679894 878465 679946 878517
rect 675766 878317 675818 878369
rect 675766 877799 675818 877851
rect 674326 876689 674378 876741
rect 675286 876689 675338 876741
rect 675094 874913 675146 874965
rect 675478 874913 675530 874965
rect 675190 874247 675242 874299
rect 675478 874247 675530 874299
rect 674998 873507 675050 873559
rect 675382 873507 675434 873559
rect 674902 872915 674954 872967
rect 675382 872915 675434 872967
rect 674038 872693 674090 872745
rect 674902 872693 674954 872745
rect 654166 872619 654218 872671
rect 675094 872619 675146 872671
rect 674230 870547 674282 870599
rect 675478 870547 675530 870599
rect 674614 869955 674666 870007
rect 675382 869955 675434 870007
rect 674518 869733 674570 869785
rect 674998 869733 675050 869785
rect 674134 868771 674186 868823
rect 675190 868771 675242 868823
rect 674902 867365 674954 867417
rect 675478 867365 675530 867417
rect 674422 865737 674474 865789
rect 675190 865737 675242 865789
rect 653782 863961 653834 864013
rect 675094 863961 675146 864013
rect 41782 816601 41834 816653
rect 47446 816601 47498 816653
rect 41782 816083 41834 816135
rect 44854 816083 44906 816135
rect 41590 815343 41642 815395
rect 44950 815343 45002 815395
rect 41782 814603 41834 814655
rect 43222 814603 43274 814655
rect 41590 813419 41642 813471
rect 44662 813419 44714 813471
rect 41782 812531 41834 812583
rect 44758 812531 44810 812583
rect 41590 810089 41642 810141
rect 42742 810089 42794 810141
rect 41590 808387 41642 808439
rect 42838 808387 42890 808439
rect 41782 807203 41834 807255
rect 43030 807203 43082 807255
rect 41590 806907 41642 806959
rect 42646 806907 42698 806959
rect 41782 803799 41834 803851
rect 43126 803799 43178 803851
rect 41494 803725 41546 803777
rect 44566 803725 44618 803777
rect 41590 803651 41642 803703
rect 42934 803651 42986 803703
rect 42742 800839 42794 800891
rect 43510 800839 43562 800891
rect 42838 800765 42890 800817
rect 43414 800765 43466 800817
rect 42742 800691 42794 800743
rect 57718 800691 57770 800743
rect 42838 800617 42890 800669
rect 57622 800617 57674 800669
rect 41398 800469 41450 800521
rect 43702 800469 43754 800521
rect 41878 800173 41930 800225
rect 42070 800173 42122 800225
rect 43318 800173 43370 800225
rect 41878 799951 41930 800003
rect 42646 797879 42698 797931
rect 42070 797435 42122 797487
rect 42742 797435 42794 797487
rect 42742 797287 42794 797339
rect 42166 796251 42218 796303
rect 43030 796251 43082 796303
rect 43030 796103 43082 796155
rect 43318 796103 43370 796155
rect 42070 795585 42122 795637
rect 42838 795585 42890 795637
rect 42166 794771 42218 794823
rect 42934 794771 42986 794823
rect 42934 794623 42986 794675
rect 43414 794623 43466 794675
rect 42070 794253 42122 794305
rect 42742 794253 42794 794305
rect 42166 793809 42218 793861
rect 43126 793809 43178 793861
rect 43126 793661 43178 793713
rect 43510 793661 43562 793713
rect 42262 792107 42314 792159
rect 43030 792107 43082 792159
rect 655222 792033 655274 792085
rect 675382 792033 675434 792085
rect 42262 790109 42314 790161
rect 43126 790109 43178 790161
rect 43126 789961 43178 790013
rect 43702 789961 43754 790013
rect 42166 789887 42218 789939
rect 42742 789887 42794 789939
rect 42166 789443 42218 789495
rect 43030 789443 43082 789495
rect 42742 789147 42794 789199
rect 58198 789147 58250 789199
rect 44950 789073 45002 789125
rect 58390 789073 58442 789125
rect 42166 786853 42218 786905
rect 43126 786853 43178 786905
rect 42166 786409 42218 786461
rect 42838 786409 42890 786461
rect 42070 785595 42122 785647
rect 42934 785595 42986 785647
rect 44854 785521 44906 785573
rect 59158 785521 59210 785573
rect 47446 785373 47498 785425
rect 59638 785373 59690 785425
rect 42166 785151 42218 785203
rect 42742 785151 42794 785203
rect 655030 783449 655082 783501
rect 674998 783449 675050 783501
rect 673270 782931 673322 782983
rect 675382 782931 675434 782983
rect 654358 780489 654410 780541
rect 675286 780489 675338 780541
rect 674998 778861 675050 778913
rect 675382 778861 675434 778913
rect 673174 778713 673226 778765
rect 675478 778713 675530 778765
rect 674614 773607 674666 773659
rect 675286 773607 675338 773659
rect 41782 773459 41834 773511
rect 47446 773459 47498 773511
rect 41782 772867 41834 772919
rect 44950 772867 45002 772919
rect 41782 772275 41834 772327
rect 45046 772275 45098 772327
rect 41590 772127 41642 772179
rect 61846 772127 61898 772179
rect 41782 771979 41834 772031
rect 43222 771979 43274 772031
rect 41494 771905 41546 771957
rect 62038 771905 62090 771957
rect 41782 771387 41834 771439
rect 43222 771387 43274 771439
rect 41590 767391 41642 767443
rect 43030 767391 43082 767443
rect 41590 766281 41642 766333
rect 42934 766281 42986 766333
rect 41782 765393 41834 765445
rect 43126 765393 43178 765445
rect 41782 763395 41834 763447
rect 42838 763395 42890 763447
rect 41590 760731 41642 760783
rect 44854 760731 44906 760783
rect 42838 757475 42890 757527
rect 58678 757475 58730 757527
rect 41302 757401 41354 757453
rect 43414 757401 43466 757453
rect 40342 757327 40394 757379
rect 41686 757327 41738 757379
rect 42742 757327 42794 757379
rect 43030 757327 43082 757379
rect 43606 757327 43658 757379
rect 42934 757253 42986 757305
rect 43510 757253 43562 757305
rect 42166 757179 42218 757231
rect 43318 757179 43370 757231
rect 42070 757105 42122 757157
rect 43126 757105 43178 757157
rect 41782 757031 41834 757083
rect 43030 757031 43082 757083
rect 41878 756957 41930 757009
rect 42934 756957 42986 757009
rect 41782 756735 41834 756787
rect 42070 754885 42122 754937
rect 42742 754885 42794 754937
rect 42166 754071 42218 754123
rect 42838 754071 42890 754123
rect 42838 753923 42890 753975
rect 43318 753923 43370 753975
rect 42070 753035 42122 753087
rect 42934 753035 42986 753087
rect 42934 752887 42986 752939
rect 43414 752887 43466 752939
rect 42166 751999 42218 752051
rect 43318 751999 43370 752051
rect 42070 751777 42122 751829
rect 43030 751777 43082 751829
rect 42070 751111 42122 751163
rect 43126 751111 43178 751163
rect 43126 750963 43178 751015
rect 43510 750963 43562 751015
rect 42166 750593 42218 750645
rect 42838 750593 42890 750645
rect 42070 749779 42122 749831
rect 42742 749779 42794 749831
rect 655702 748817 655754 748869
rect 675382 748817 675434 748869
rect 42166 747411 42218 747463
rect 43126 747411 43178 747463
rect 42838 747263 42890 747315
rect 43126 747263 43178 747315
rect 42166 746893 42218 746945
rect 42934 746893 42986 746945
rect 42934 746745 42986 746797
rect 43606 746745 43658 746797
rect 42070 746079 42122 746131
rect 43030 746079 43082 746131
rect 42358 745931 42410 745983
rect 54646 745931 54698 745983
rect 54742 745931 54794 745983
rect 57622 745931 57674 745983
rect 43318 745561 43370 745613
rect 59638 745561 59690 745613
rect 42166 745487 42218 745539
rect 42934 745487 42986 745539
rect 45046 745339 45098 745391
rect 58486 745339 58538 745391
rect 42166 743785 42218 743837
rect 43126 743785 43178 743837
rect 42070 743193 42122 743245
rect 42838 743193 42890 743245
rect 47446 742971 47498 743023
rect 59638 742971 59690 743023
rect 44950 742897 45002 742949
rect 59734 742897 59786 742949
rect 674422 742749 674474 742801
rect 675190 742749 675242 742801
rect 42166 742601 42218 742653
rect 42742 742601 42794 742653
rect 42166 741935 42218 741987
rect 42358 741935 42410 741987
rect 674902 741417 674954 741469
rect 675190 741417 675242 741469
rect 670774 737495 670826 737547
rect 675286 737495 675338 737547
rect 654070 737421 654122 737473
rect 674518 737421 674570 737473
rect 654166 737347 654218 737399
rect 675286 737347 675338 737399
rect 672598 734905 672650 734957
rect 675382 734905 675434 734957
rect 672982 734387 673034 734439
rect 675382 734387 675434 734439
rect 673078 734165 673130 734217
rect 675382 734165 675434 734217
rect 675190 733869 675242 733921
rect 675478 733869 675530 733921
rect 672886 732315 672938 732367
rect 675478 732315 675530 732367
rect 674518 732019 674570 732071
rect 675382 732019 675434 732071
rect 674422 730465 674474 730517
rect 675478 730465 675530 730517
rect 41782 730391 41834 730443
rect 47542 730391 47594 730443
rect 41782 729873 41834 729925
rect 44950 729873 45002 729925
rect 41782 729355 41834 729407
rect 45046 729355 45098 729407
rect 41782 728985 41834 729037
rect 43222 728985 43274 729037
rect 41590 728911 41642 728963
rect 62230 728911 62282 728963
rect 41686 728689 41738 728741
rect 62422 728689 62474 728741
rect 674134 728615 674186 728667
rect 675478 728615 675530 728667
rect 41782 728319 41834 728371
rect 43318 728319 43370 728371
rect 41782 727875 41834 727927
rect 43414 727875 43466 727927
rect 41782 726839 41834 726891
rect 43222 726839 43274 726891
rect 41782 725951 41834 726003
rect 42934 725951 42986 726003
rect 41590 720993 41642 721045
rect 43030 720993 43082 721045
rect 41590 720623 41642 720675
rect 43126 720623 43178 720675
rect 42262 719735 42314 719787
rect 42838 719735 42890 719787
rect 42166 719439 42218 719491
rect 43126 719439 43178 719491
rect 41590 719291 41642 719343
rect 43126 719291 43178 719343
rect 41494 717663 41546 717715
rect 47446 717663 47498 717715
rect 41590 717515 41642 717567
rect 42934 717515 42986 717567
rect 41878 715591 41930 715643
rect 42742 715591 42794 715643
rect 655606 714703 655658 714755
rect 676246 714703 676298 714755
rect 655414 714555 655466 714607
rect 676150 714555 676202 714607
rect 655126 714407 655178 714459
rect 676342 714407 676394 714459
rect 42838 714259 42890 714311
rect 59638 714259 59690 714311
rect 43030 714185 43082 714237
rect 43510 714185 43562 714237
rect 673366 714185 673418 714237
rect 676054 714185 676106 714237
rect 41686 714037 41738 714089
rect 43030 714037 43082 714089
rect 41782 713815 41834 713867
rect 42262 713741 42314 713793
rect 43606 713741 43658 713793
rect 41782 713519 41834 713571
rect 672790 713371 672842 713423
rect 676246 713371 676298 713423
rect 669718 713075 669770 713127
rect 670966 713075 671018 713127
rect 676054 713075 676106 713127
rect 670678 712631 670730 712683
rect 676054 712631 676106 712683
rect 669526 711891 669578 711943
rect 670870 711891 670922 711943
rect 676246 711891 676298 711943
rect 42070 711669 42122 711721
rect 42742 711669 42794 711721
rect 42742 711521 42794 711573
rect 43510 711521 43562 711573
rect 670582 711521 670634 711573
rect 676054 711521 676106 711573
rect 43030 711299 43082 711351
rect 674614 711299 674666 711351
rect 676054 711299 676106 711351
rect 42166 710855 42218 710907
rect 42838 710855 42890 710907
rect 42166 709893 42218 709945
rect 42742 709893 42794 709945
rect 42742 709745 42794 709797
rect 42070 708487 42122 708539
rect 43510 708487 43562 708539
rect 674998 708413 675050 708465
rect 676054 708413 676106 708465
rect 42070 708339 42122 708391
rect 43030 708339 43082 708391
rect 42166 707377 42218 707429
rect 43126 707377 43178 707429
rect 42166 706563 42218 706615
rect 42742 706563 42794 706615
rect 673270 705527 673322 705579
rect 676054 705527 676106 705579
rect 673174 704861 673226 704913
rect 676246 704861 676298 704913
rect 42358 704787 42410 704839
rect 43606 704787 43658 704839
rect 42166 704269 42218 704321
rect 42934 704269 42986 704321
rect 42070 703529 42122 703581
rect 43030 703529 43082 703581
rect 42166 702863 42218 702915
rect 42358 702863 42410 702915
rect 654358 702789 654410 702841
rect 675382 702789 675434 702841
rect 649462 702715 649514 702767
rect 679990 702715 680042 702767
rect 43510 702641 43562 702693
rect 58774 702641 58826 702693
rect 45046 702567 45098 702619
rect 58678 702567 58730 702619
rect 42166 702419 42218 702471
rect 42838 702419 42890 702471
rect 42070 700495 42122 700547
rect 43126 700495 43178 700547
rect 42166 700051 42218 700103
rect 42934 700051 42986 700103
rect 47542 699755 47594 699807
rect 59254 699755 59306 699807
rect 44950 699681 45002 699733
rect 58870 699681 58922 699733
rect 42166 699385 42218 699437
rect 42742 699385 42794 699437
rect 42070 698423 42122 698475
rect 43798 698423 43850 698475
rect 654166 694279 654218 694331
rect 674998 694279 675050 694331
rect 670966 693613 671018 693665
rect 675478 693613 675530 693665
rect 674902 692873 674954 692925
rect 675382 692873 675434 692925
rect 654070 691319 654122 691371
rect 675190 691319 675242 691371
rect 674614 690431 674666 690483
rect 675478 690431 675530 690483
rect 673174 689765 673226 689817
rect 675382 689765 675434 689817
rect 673366 689321 673418 689373
rect 675382 689321 675434 689373
rect 673270 689099 673322 689151
rect 675382 689099 675434 689151
rect 674998 688877 675050 688929
rect 675478 688877 675530 688929
rect 672694 687323 672746 687375
rect 675478 687323 675530 687375
rect 675190 687027 675242 687079
rect 675478 687027 675530 687079
rect 41782 686805 41834 686857
rect 50326 686805 50378 686857
rect 41782 686287 41834 686339
rect 47638 686287 47690 686339
rect 41590 685547 41642 685599
rect 47734 685547 47786 685599
rect 674326 685473 674378 685525
rect 675478 685473 675530 685525
rect 41782 685325 41834 685377
rect 43318 685325 43370 685377
rect 41782 684807 41834 684859
rect 43606 684807 43658 684859
rect 41782 683845 41834 683897
rect 43414 683845 43466 683897
rect 44950 683845 45002 683897
rect 674230 683623 674282 683675
rect 675478 683623 675530 683675
rect 41590 682957 41642 683009
rect 43222 682957 43274 683009
rect 45142 682957 45194 683009
rect 41782 680663 41834 680715
rect 43030 680663 43082 680715
rect 41590 676075 41642 676127
rect 43126 676075 43178 676127
rect 41590 674299 41642 674351
rect 42934 674299 42986 674351
rect 41590 674003 41642 674055
rect 47542 674003 47594 674055
rect 39766 673855 39818 673907
rect 41494 673855 41546 673907
rect 34486 672523 34538 672575
rect 42166 672523 42218 672575
rect 41974 671339 42026 671391
rect 43126 671339 43178 671391
rect 37366 671265 37418 671317
rect 43702 671265 43754 671317
rect 41494 671191 41546 671243
rect 43510 671191 43562 671243
rect 42166 671117 42218 671169
rect 43318 671117 43370 671169
rect 42838 671043 42890 671095
rect 59638 671043 59690 671095
rect 41782 670599 41834 670651
rect 42262 670599 42314 670651
rect 43414 670599 43466 670651
rect 41782 670303 41834 670355
rect 42166 668527 42218 668579
rect 43030 668527 43082 668579
rect 43126 668453 43178 668505
rect 655510 668379 655562 668431
rect 676246 668379 676298 668431
rect 43126 668157 43178 668209
rect 655318 668157 655370 668209
rect 676246 668157 676298 668209
rect 42166 667861 42218 667913
rect 42838 667861 42890 667913
rect 42838 667713 42890 667765
rect 43318 667713 43370 667765
rect 672790 667565 672842 667617
rect 675958 667565 676010 667617
rect 652246 666751 652298 666803
rect 668758 666751 668810 666803
rect 672790 666751 672842 666803
rect 676246 666751 676298 666803
rect 649750 666677 649802 666729
rect 670678 666677 670730 666729
rect 676150 666677 676202 666729
rect 670390 666011 670442 666063
rect 675958 666011 676010 666063
rect 668758 665493 668810 665545
rect 670582 665493 670634 665545
rect 675958 665493 676010 665545
rect 655222 665419 655274 665471
rect 676054 665419 676106 665471
rect 42166 665345 42218 665397
rect 42934 665345 42986 665397
rect 42070 665271 42122 665323
rect 45046 665271 45098 665323
rect 42934 665197 42986 665249
rect 43414 665197 43466 665249
rect 674422 665197 674474 665249
rect 676054 665197 676106 665249
rect 670678 664975 670730 665027
rect 675958 664975 676010 665027
rect 42070 663939 42122 663991
rect 43030 663939 43082 663991
rect 43126 663495 43178 663547
rect 42166 663347 42218 663399
rect 43126 663273 43178 663325
rect 43702 663273 43754 663325
rect 674134 662311 674186 662363
rect 676054 662311 676106 662363
rect 670774 660461 670826 660513
rect 676054 660461 676106 660513
rect 42070 660387 42122 660439
rect 42934 660387 42986 660439
rect 672886 660091 672938 660143
rect 676054 660091 676106 660143
rect 42166 659869 42218 659921
rect 42838 659869 42890 659921
rect 672982 659721 673034 659773
rect 676246 659721 676298 659773
rect 47734 659425 47786 659477
rect 59158 659425 59210 659477
rect 45046 659351 45098 659403
rect 58774 659351 58826 659403
rect 42070 659055 42122 659107
rect 43126 659055 43178 659107
rect 672598 658611 672650 658663
rect 676054 658611 676106 658663
rect 673078 658241 673130 658293
rect 676246 658241 676298 658293
rect 42070 657353 42122 657405
rect 43030 657353 43082 657405
rect 42166 656835 42218 656887
rect 42838 656835 42890 656887
rect 654166 656687 654218 656739
rect 675382 656687 675434 656739
rect 50326 656613 50378 656665
rect 58198 656613 58250 656665
rect 47638 656539 47690 656591
rect 58390 656539 58442 656591
rect 42166 656169 42218 656221
rect 42934 656169 42986 656221
rect 42166 655503 42218 655555
rect 45910 655503 45962 655555
rect 649558 654023 649610 654075
rect 679990 654097 680042 654149
rect 670870 648917 670922 648969
rect 675190 648917 675242 648969
rect 670774 648325 670826 648377
rect 675190 648325 675242 648377
rect 655798 648251 655850 648303
rect 674998 648251 675050 648303
rect 673846 648029 673898 648081
rect 675190 648029 675242 648081
rect 655990 645143 656042 645195
rect 675286 645143 675338 645195
rect 672982 644551 673034 644603
rect 675382 644551 675434 644603
rect 670582 644033 670634 644085
rect 675478 644033 675530 644085
rect 41782 643663 41834 643715
rect 50326 643663 50378 643715
rect 674998 643663 675050 643715
rect 675382 643663 675434 643715
rect 672886 643589 672938 643641
rect 675478 643589 675530 643641
rect 41782 643071 41834 643123
rect 47734 643071 47786 643123
rect 41494 642553 41546 642605
rect 61942 642553 61994 642605
rect 41686 642479 41738 642531
rect 62134 642479 62186 642531
rect 41590 642331 41642 642383
rect 47830 642331 47882 642383
rect 670486 642257 670538 642309
rect 675478 642257 675530 642309
rect 41782 642183 41834 642235
rect 43510 642183 43562 642235
rect 41782 641591 41834 641643
rect 43606 641591 43658 641643
rect 41782 640111 41834 640163
rect 43414 640111 43466 640163
rect 41590 633895 41642 633947
rect 43126 633895 43178 633947
rect 41878 631083 41930 631135
rect 43030 631083 43082 631135
rect 41590 630787 41642 630839
rect 47638 630787 47690 630839
rect 43126 628123 43178 628175
rect 43510 628123 43562 628175
rect 37366 627975 37418 628027
rect 43894 627975 43946 628027
rect 34486 627901 34538 627953
rect 43798 627901 43850 627953
rect 40150 627827 40202 627879
rect 43702 627827 43754 627879
rect 41494 627679 41546 627731
rect 43126 627679 43178 627731
rect 43222 627679 43274 627731
rect 42262 627605 42314 627657
rect 43030 627605 43082 627657
rect 42166 627531 42218 627583
rect 43222 627531 43274 627583
rect 43414 627457 43466 627509
rect 41782 627383 41834 627435
rect 41782 627161 41834 627213
rect 42838 625163 42890 625215
rect 43222 625163 43274 625215
rect 655414 624941 655466 624993
rect 676246 624941 676298 624993
rect 42166 624275 42218 624327
rect 58966 624275 59018 624327
rect 672790 623979 672842 624031
rect 676054 623979 676106 624031
rect 42166 623461 42218 623513
rect 42934 623461 42986 623513
rect 672598 623387 672650 623439
rect 676054 623387 676106 623439
rect 42934 623313 42986 623365
rect 43414 623313 43466 623365
rect 669622 623165 669674 623217
rect 670390 623165 670442 623217
rect 676342 623165 676394 623217
rect 670198 622425 670250 622477
rect 676054 622425 676106 622477
rect 655606 622351 655658 622403
rect 676246 622351 676298 622403
rect 655126 622203 655178 622255
rect 676150 622203 676202 622255
rect 42166 622055 42218 622107
rect 47926 622055 47978 622107
rect 674326 621981 674378 622033
rect 676246 621981 676298 622033
rect 42166 621907 42218 621959
rect 43030 621907 43082 621959
rect 670678 621907 670730 621959
rect 676054 621907 676106 621959
rect 43030 621759 43082 621811
rect 43702 621759 43754 621811
rect 42166 621611 42218 621663
rect 43510 621611 43562 621663
rect 670294 621315 670346 621367
rect 676054 621315 676106 621367
rect 42934 620945 42986 620997
rect 42070 620871 42122 620923
rect 42934 620797 42986 620849
rect 43798 620797 43850 620849
rect 43222 620649 43274 620701
rect 43606 620649 43658 620701
rect 42166 620353 42218 620405
rect 43126 620353 43178 620405
rect 43126 620205 43178 620257
rect 43894 620205 43946 620257
rect 669814 619835 669866 619887
rect 670678 619835 670730 619887
rect 674614 619021 674666 619073
rect 676054 619021 676106 619073
rect 674230 618799 674282 618851
rect 676246 618799 676298 618851
rect 42070 617837 42122 617889
rect 42838 617837 42890 617889
rect 42742 617319 42794 617371
rect 42166 617171 42218 617223
rect 670966 617097 671018 617149
rect 676246 617097 676298 617149
rect 42166 616653 42218 616705
rect 42934 616653 42986 616705
rect 672694 616505 672746 616557
rect 676054 616505 676106 616557
rect 47830 616283 47882 616335
rect 58966 616283 59018 616335
rect 47926 616209 47978 616261
rect 59638 616209 59690 616261
rect 42166 615987 42218 616039
rect 43030 615987 43082 616039
rect 673366 615913 673418 615965
rect 676054 615913 676106 615965
rect 673174 615173 673226 615225
rect 676246 615173 676298 615225
rect 673270 614433 673322 614485
rect 676054 614433 676106 614485
rect 42166 614137 42218 614189
rect 43126 614137 43178 614189
rect 42166 613619 42218 613671
rect 42838 613619 42890 613671
rect 655126 613471 655178 613523
rect 675382 613471 675434 613523
rect 50326 613397 50378 613449
rect 59638 613397 59690 613449
rect 47734 613323 47786 613375
rect 59542 613323 59594 613375
rect 42070 612953 42122 613005
rect 42742 612953 42794 613005
rect 42166 612361 42218 612413
rect 45910 612361 45962 612413
rect 649654 610659 649706 610711
rect 679990 610659 680042 610711
rect 673270 606885 673322 606937
rect 675190 606885 675242 606937
rect 670966 603259 671018 603311
rect 675382 603259 675434 603311
rect 673366 603037 673418 603089
rect 675382 603037 675434 603089
rect 655798 602075 655850 602127
rect 674998 602075 675050 602127
rect 653782 602001 653834 602053
rect 674902 602001 674954 602053
rect 673078 601927 673130 601979
rect 675286 601927 675338 601979
rect 41782 600447 41834 600499
rect 50326 600447 50378 600499
rect 41590 599707 41642 599759
rect 47830 599707 47882 599759
rect 673174 599559 673226 599611
rect 675382 599559 675434 599611
rect 41782 599337 41834 599389
rect 47926 599337 47978 599389
rect 670678 599263 670730 599315
rect 675382 599263 675434 599315
rect 41782 598967 41834 599019
rect 43222 598967 43274 599019
rect 672790 598893 672842 598945
rect 675382 598893 675434 598945
rect 674998 598671 675050 598723
rect 675478 598671 675530 598723
rect 41590 598227 41642 598279
rect 43510 598227 43562 598279
rect 672694 597117 672746 597169
rect 675478 597117 675530 597169
rect 674902 596821 674954 596873
rect 675382 596821 675434 596873
rect 41590 596155 41642 596207
rect 43318 596155 43370 596207
rect 45046 596155 45098 596207
rect 41782 593491 41834 593543
rect 43030 593491 43082 593543
rect 41878 590901 41930 590953
rect 43126 590901 43178 590953
rect 41590 590531 41642 590583
rect 42838 590531 42890 590583
rect 41974 589495 42026 589547
rect 43126 589495 43178 589547
rect 41590 589347 41642 589399
rect 43126 589347 43178 589399
rect 41590 587867 41642 587919
rect 42838 587867 42890 587919
rect 41590 587571 41642 587623
rect 47734 587571 47786 587623
rect 42358 584611 42410 584663
rect 43414 584611 43466 584663
rect 42070 584537 42122 584589
rect 43318 584537 43370 584589
rect 42166 584463 42218 584515
rect 43222 584463 43274 584515
rect 41782 584167 41834 584219
rect 41782 583945 41834 583997
rect 42166 582095 42218 582147
rect 43030 582095 43082 582147
rect 43030 581947 43082 581999
rect 43222 581947 43274 581999
rect 42166 580837 42218 580889
rect 58966 580837 59018 580889
rect 42070 580245 42122 580297
rect 42934 580245 42986 580297
rect 42934 580097 42986 580149
rect 43318 580097 43370 580149
rect 655702 579283 655754 579335
rect 676246 579283 676298 579335
rect 655510 579135 655562 579187
rect 676342 579135 676394 579187
rect 655318 578987 655370 579039
rect 676150 578987 676202 579039
rect 42166 578913 42218 578965
rect 48022 578913 48074 578965
rect 42166 578765 42218 578817
rect 42838 578765 42890 578817
rect 672598 578765 672650 578817
rect 676246 578765 676298 578817
rect 42166 577803 42218 577855
rect 43126 577803 43178 577855
rect 672502 577803 672554 577855
rect 676246 577803 676298 577855
rect 670102 577433 670154 577485
rect 676054 577433 676106 577485
rect 672598 577063 672650 577115
rect 676054 577063 676106 577115
rect 42070 576915 42122 576967
rect 43030 576915 43082 576967
rect 670294 576545 670346 576597
rect 676054 576545 676106 576597
rect 669910 576027 669962 576079
rect 670294 576027 670346 576079
rect 670390 575879 670442 575931
rect 676054 575879 676106 575931
rect 42166 574547 42218 574599
rect 43126 574547 43178 574599
rect 42166 574103 42218 574155
rect 42934 574103 42986 574155
rect 47926 573067 47978 573119
rect 58966 573067 59018 573119
rect 48022 572993 48074 573045
rect 59638 572993 59690 573045
rect 42166 572623 42218 572675
rect 42838 572623 42890 572675
rect 670870 572253 670922 572305
rect 676246 572253 676298 572305
rect 670774 571513 670826 571565
rect 676054 571513 676106 571565
rect 670486 571069 670538 571121
rect 676054 571069 676106 571121
rect 670582 570551 670634 570603
rect 676054 570551 676106 570603
rect 42070 570403 42122 570455
rect 43030 570403 43082 570455
rect 42166 570329 42218 570381
rect 42934 570329 42986 570381
rect 50326 570181 50378 570233
rect 59350 570181 59402 570233
rect 673846 570181 673898 570233
rect 676246 570181 676298 570233
rect 47830 570107 47882 570159
rect 59542 570107 59594 570159
rect 42070 569663 42122 569715
rect 42934 569663 42986 569715
rect 672982 569589 673034 569641
rect 676054 569589 676106 569641
rect 42166 569145 42218 569197
rect 46198 569145 46250 569197
rect 672886 569071 672938 569123
rect 676054 569071 676106 569123
rect 655702 567443 655754 567495
rect 675382 567443 675434 567495
rect 649846 567369 649898 567421
rect 679990 567369 680042 567421
rect 674422 559525 674474 559577
rect 675382 559525 675434 559577
rect 656566 558785 656618 558837
rect 674998 558785 675050 558837
rect 674614 558045 674666 558097
rect 675382 558045 675434 558097
rect 673846 555973 673898 556025
rect 675286 555973 675338 556025
rect 654166 555825 654218 555877
rect 675286 555825 675338 555877
rect 674902 555011 674954 555063
rect 675478 555011 675530 555063
rect 673750 554345 673802 554397
rect 675382 554345 675434 554397
rect 672886 553901 672938 553953
rect 675478 553901 675530 553953
rect 674998 553457 675050 553509
rect 675382 553457 675434 553509
rect 673654 553309 673706 553361
rect 675478 553309 675530 553361
rect 670870 551903 670922 551955
rect 675478 551903 675530 551955
rect 674326 548869 674378 548921
rect 675286 548869 675338 548921
rect 674230 548203 674282 548255
rect 675286 548203 675338 548255
rect 41590 543023 41642 543075
rect 50518 543023 50570 543075
rect 41782 542653 41834 542705
rect 48790 542653 48842 542705
rect 41782 542135 41834 542187
rect 48886 542135 48938 542187
rect 41782 541765 41834 541817
rect 43222 541765 43274 541817
rect 42742 541543 42794 541595
rect 57718 541543 57770 541595
rect 42838 541469 42890 541521
rect 57622 541469 57674 541521
rect 42166 539693 42218 539745
rect 42934 539693 42986 539745
rect 42166 538139 42218 538191
rect 42742 538139 42794 538191
rect 42166 536437 42218 536489
rect 42838 536437 42890 536489
rect 672502 533773 672554 533825
rect 675958 533773 676010 533825
rect 42070 533699 42122 533751
rect 42742 533699 42794 533751
rect 655606 533255 655658 533307
rect 676054 533255 676106 533307
rect 655414 533107 655466 533159
rect 676150 533107 676202 533159
rect 655222 532959 655274 533011
rect 676246 532959 676298 533011
rect 672406 532663 672458 532715
rect 672598 532663 672650 532715
rect 676054 532663 676106 532715
rect 42166 531479 42218 531531
rect 42742 531479 42794 531531
rect 670294 531479 670346 531531
rect 676246 531479 676298 531531
rect 42166 530887 42218 530939
rect 42838 530887 42890 530939
rect 42166 529407 42218 529459
rect 43030 529407 43082 529459
rect 673270 528001 673322 528053
rect 676246 528001 676298 528053
rect 42166 527779 42218 527831
rect 43126 527779 43178 527831
rect 48886 527483 48938 527535
rect 59638 527483 59690 527535
rect 673078 527409 673130 527461
rect 676246 527409 676298 527461
rect 42070 527187 42122 527239
rect 42838 527187 42890 527239
rect 670966 526669 671018 526721
rect 676054 526669 676106 526721
rect 42166 526447 42218 526499
rect 42934 526447 42986 526499
rect 672694 526299 672746 526351
rect 676054 526299 676106 526351
rect 42070 525929 42122 525981
rect 46678 525929 46730 525981
rect 670678 525929 670730 525981
rect 676246 525929 676298 525981
rect 673366 525189 673418 525241
rect 676054 525189 676106 525241
rect 48790 524967 48842 525019
rect 59638 524967 59690 525019
rect 673174 524819 673226 524871
rect 676054 524819 676106 524871
rect 50518 524671 50570 524723
rect 59350 524671 59402 524723
rect 672790 524449 672842 524501
rect 676246 524449 676298 524501
rect 42358 524227 42410 524279
rect 47830 524227 47882 524279
rect 649942 521267 649994 521319
rect 679798 521267 679850 521319
rect 43414 519935 43466 519987
rect 43414 519713 43466 519765
rect 43318 514089 43370 514141
rect 43510 514089 43562 514141
rect 655510 490039 655562 490091
rect 676246 490039 676298 490091
rect 655318 489891 655370 489943
rect 676150 489891 676202 489943
rect 655126 489743 655178 489795
rect 676342 489743 676394 489795
rect 670006 488115 670058 488167
rect 676054 488115 676106 488167
rect 676630 488115 676682 488167
rect 670198 487079 670250 487131
rect 676246 487079 676298 487131
rect 676534 487079 676586 487131
rect 674902 486635 674954 486687
rect 676054 486635 676106 486687
rect 674326 486561 674378 486613
rect 675958 486561 676010 486613
rect 674422 486487 674474 486539
rect 676246 486487 676298 486539
rect 674614 483749 674666 483801
rect 676054 483749 676106 483801
rect 674230 483675 674282 483727
rect 675958 483675 676010 483727
rect 670870 481899 670922 481951
rect 676054 481899 676106 481951
rect 672886 481529 672938 481581
rect 676246 481529 676298 481581
rect 673846 480789 673898 480841
rect 676054 480789 676106 480841
rect 673750 480419 673802 480471
rect 676054 480419 676106 480471
rect 673654 480049 673706 480101
rect 676246 480049 676298 480101
rect 676630 479235 676682 479287
rect 679702 479235 679754 479287
rect 650038 478125 650090 478177
rect 679894 478125 679946 478177
rect 41590 429211 41642 429263
rect 53206 429211 53258 429263
rect 673846 429137 673898 429189
rect 675286 429137 675338 429189
rect 41782 428915 41834 428967
rect 50326 428915 50378 428967
rect 41782 428323 41834 428375
rect 48022 428323 48074 428375
rect 41782 427953 41834 428005
rect 43318 427953 43370 428005
rect 41782 427361 41834 427413
rect 43414 427361 43466 427413
rect 41686 427213 41738 427265
rect 45334 427213 45386 427265
rect 41782 426843 41834 426895
rect 43318 426843 43370 426895
rect 41782 420405 41834 420457
rect 45526 420405 45578 420457
rect 41782 419073 41834 419125
rect 42838 419073 42890 419125
rect 41782 418555 41834 418607
rect 43126 418555 43178 418607
rect 41590 417815 41642 417867
rect 42934 417815 42986 417867
rect 41782 417741 41834 417793
rect 43030 417741 43082 417793
rect 41782 416927 41834 416979
rect 47926 416927 47978 416979
rect 41782 413375 41834 413427
rect 41782 413153 41834 413205
rect 42838 409823 42890 409875
rect 43222 409823 43274 409875
rect 42166 409675 42218 409727
rect 42838 409675 42890 409727
rect 42166 409453 42218 409505
rect 42934 409453 42986 409505
rect 42934 409305 42986 409357
rect 43126 409305 43178 409357
rect 43222 409009 43274 409061
rect 43414 409009 43466 409061
rect 42070 408047 42122 408099
rect 43030 408047 43082 408099
rect 42166 407973 42218 408025
rect 42934 407825 42986 407877
rect 42070 407455 42122 407507
rect 43126 407455 43178 407507
rect 42166 406863 42218 406915
rect 43030 406863 43082 406915
rect 42838 406049 42890 406101
rect 58486 406049 58538 406101
rect 42934 402571 42986 402623
rect 59350 402571 59402 402623
rect 655126 400573 655178 400625
rect 676150 400573 676202 400625
rect 655510 400499 655562 400551
rect 676246 400499 676298 400551
rect 655318 400425 655370 400477
rect 676054 400425 676106 400477
rect 673366 400351 673418 400403
rect 676246 400351 676298 400403
rect 53206 400277 53258 400329
rect 59734 400277 59786 400329
rect 50326 400203 50378 400255
rect 59542 400203 59594 400255
rect 48022 400129 48074 400181
rect 59638 400129 59690 400181
rect 672502 400129 672554 400181
rect 673846 400129 673898 400181
rect 676054 400129 676106 400181
rect 673078 397983 673130 398035
rect 675958 397983 676010 398035
rect 675190 397909 675242 397961
rect 676630 397909 676682 397961
rect 674518 397687 674570 397739
rect 676054 397687 676106 397739
rect 673174 395541 673226 395593
rect 676054 395541 676106 395593
rect 42070 394505 42122 394557
rect 57718 394505 57770 394557
rect 650134 388807 650186 388859
rect 679798 388807 679850 388859
rect 41782 386439 41834 386491
rect 53206 386439 53258 386491
rect 673270 385847 673322 385899
rect 674518 385847 674570 385899
rect 41590 385699 41642 385751
rect 50326 385699 50378 385751
rect 41782 385329 41834 385381
rect 48118 385329 48170 385381
rect 41590 385181 41642 385233
rect 43222 385181 43274 385233
rect 41782 384367 41834 384419
rect 43510 384367 43562 384419
rect 41782 383479 41834 383531
rect 43318 383479 43370 383531
rect 45430 383479 45482 383531
rect 653782 381629 653834 381681
rect 675094 381629 675146 381681
rect 34486 381555 34538 381607
rect 43318 381555 43370 381607
rect 652342 381555 652394 381607
rect 674998 381555 675050 381607
rect 40246 377189 40298 377241
rect 45622 377189 45674 377241
rect 41782 376893 41834 376945
rect 42934 376893 42986 376945
rect 41782 374747 41834 374799
rect 43030 374747 43082 374799
rect 41590 374599 41642 374651
rect 42838 374599 42890 374651
rect 39286 374303 39338 374355
rect 41782 374303 41834 374355
rect 39670 374229 39722 374281
rect 43126 374229 43178 374281
rect 41878 373859 41930 373911
rect 48022 373859 48074 373911
rect 673174 372083 673226 372135
rect 675382 372083 675434 372135
rect 41782 370159 41834 370211
rect 41782 369937 41834 369989
rect 42934 366681 42986 366733
rect 43222 366681 43274 366733
rect 42166 366533 42218 366585
rect 42934 366533 42986 366585
rect 42070 366237 42122 366289
rect 43126 366237 43178 366289
rect 42166 364979 42218 365031
rect 42838 364979 42890 365031
rect 42070 364683 42122 364735
rect 42838 364683 42890 364735
rect 42070 364239 42122 364291
rect 43126 364239 43178 364291
rect 42166 363795 42218 363847
rect 43030 363795 43082 363847
rect 42934 361427 42986 361479
rect 58486 361427 58538 361479
rect 42838 359947 42890 359999
rect 59158 359947 59210 359999
rect 655126 357135 655178 357187
rect 676246 357135 676298 357187
rect 53206 357061 53258 357113
rect 58390 357061 58442 357113
rect 50326 356987 50378 357039
rect 58486 356987 58538 357039
rect 48118 356913 48170 356965
rect 59638 356913 59690 356965
rect 673366 356173 673418 356225
rect 676246 356173 676298 356225
rect 673270 354767 673322 354819
rect 675958 354767 676010 354819
rect 672598 354397 672650 354449
rect 673270 354397 673322 354449
rect 655318 354323 655370 354375
rect 676054 354323 676106 354375
rect 655222 354249 655274 354301
rect 676150 354249 676202 354301
rect 672790 353879 672842 353931
rect 676054 353879 676106 353931
rect 42166 351289 42218 351341
rect 57718 351289 57770 351341
rect 674422 348625 674474 348677
rect 675958 348625 676010 348677
rect 675286 348551 675338 348603
rect 676246 348551 676298 348603
rect 675190 348477 675242 348529
rect 676054 348477 676106 348529
rect 674806 347515 674858 347567
rect 676054 347515 676106 347567
rect 674902 345739 674954 345791
rect 676150 345739 676202 345791
rect 674998 345665 675050 345717
rect 676246 345665 676298 345717
rect 675094 345591 675146 345643
rect 676054 345591 676106 345643
rect 41590 343223 41642 343275
rect 53206 343223 53258 343275
rect 41782 342853 41834 342905
rect 50326 342853 50378 342905
rect 650230 342705 650282 342757
rect 679702 342705 679754 342757
rect 41782 342335 41834 342387
rect 48118 342335 48170 342387
rect 41782 341965 41834 342017
rect 43510 341965 43562 342017
rect 41782 341373 41834 341425
rect 43222 341373 43274 341425
rect 675766 341373 675818 341425
rect 41782 340855 41834 340907
rect 43414 340855 43466 340907
rect 675766 340707 675818 340759
rect 666646 340633 666698 340685
rect 675478 340633 675530 340685
rect 41782 340485 41834 340537
rect 43318 340485 43370 340537
rect 45718 340485 45770 340537
rect 41782 339819 41834 339871
rect 43606 339819 43658 339871
rect 41590 339745 41642 339797
rect 45622 339893 45674 339945
rect 62614 339893 62666 339945
rect 675190 337229 675242 337281
rect 675478 337229 675530 337281
rect 674422 336563 674474 336615
rect 675382 336563 675434 336615
rect 675094 336045 675146 336097
rect 675382 336045 675434 336097
rect 41782 333085 41834 333137
rect 42742 333085 42794 333137
rect 674998 332715 675050 332767
rect 675382 332715 675434 332767
rect 674806 332197 674858 332249
rect 675478 332197 675530 332249
rect 674902 331753 674954 331805
rect 675382 331753 675434 331805
rect 41782 331531 41834 331583
rect 42934 331531 42986 331583
rect 41878 330939 41930 330991
rect 48214 330939 48266 330991
rect 41590 328719 41642 328771
rect 43030 328719 43082 328771
rect 654166 328275 654218 328327
rect 666646 328275 666698 328327
rect 41782 327017 41834 327069
rect 41782 326573 41834 326625
rect 42934 325759 42986 325811
rect 43126 325759 43178 325811
rect 42070 323317 42122 323369
rect 42454 323317 42506 323369
rect 42166 323095 42218 323147
rect 43030 323095 43082 323147
rect 41974 321615 42026 321667
rect 43126 321615 43178 321667
rect 42166 321467 42218 321519
rect 43126 321467 43178 321519
rect 42166 321245 42218 321297
rect 43030 321245 43082 321297
rect 42454 319617 42506 319669
rect 58486 319617 58538 319669
rect 43126 316731 43178 316783
rect 59158 316731 59210 316783
rect 53206 313845 53258 313897
rect 59734 313845 59786 313897
rect 50326 313771 50378 313823
rect 59542 313771 59594 313823
rect 48118 313697 48170 313749
rect 59638 313697 59690 313749
rect 654262 311181 654314 311233
rect 676246 311181 676298 311233
rect 654166 311107 654218 311159
rect 676150 311107 676202 311159
rect 654070 311033 654122 311085
rect 676342 311033 676394 311085
rect 42166 308073 42218 308125
rect 59062 308073 59114 308125
rect 45526 307777 45578 307829
rect 46102 307777 46154 307829
rect 674614 305335 674666 305387
rect 676054 305335 676106 305387
rect 675094 305261 675146 305313
rect 676246 305261 676298 305313
rect 674230 302597 674282 302649
rect 675958 302597 676010 302649
rect 674422 302523 674474 302575
rect 676054 302523 676106 302575
rect 674710 302449 674762 302501
rect 676246 302449 676298 302501
rect 674902 302375 674954 302427
rect 676054 302375 676106 302427
rect 46102 302301 46154 302353
rect 54646 302301 54698 302353
rect 43414 300895 43466 300947
rect 44278 300895 44330 300947
rect 62902 300895 62954 300947
rect 41782 299711 41834 299763
rect 50710 299711 50762 299763
rect 650326 299711 650378 299763
rect 679990 299711 680042 299763
rect 41878 299637 41930 299689
rect 44278 299637 44330 299689
rect 674326 299637 674378 299689
rect 676054 299637 676106 299689
rect 41590 299563 41642 299615
rect 60214 299563 60266 299615
rect 674998 299563 675050 299615
rect 676246 299563 676298 299615
rect 41782 298749 41834 298801
rect 43222 298749 43274 298801
rect 41782 298157 41834 298209
rect 43414 298157 43466 298209
rect 43606 298083 43658 298135
rect 62998 298083 63050 298135
rect 41782 297639 41834 297691
rect 43222 297639 43274 297691
rect 39862 296751 39914 296803
rect 43606 296751 43658 296803
rect 41782 296677 41834 296729
rect 43318 296677 43370 296729
rect 674710 295419 674762 295471
rect 675094 295419 675146 295471
rect 674614 294753 674666 294805
rect 675094 294753 675146 294805
rect 53302 293865 53354 293917
rect 59254 293865 59306 293917
rect 56182 293791 56234 293843
rect 60310 293791 60362 293843
rect 39670 293717 39722 293769
rect 58198 293717 58250 293769
rect 674422 292237 674474 292289
rect 675478 292237 675530 292289
rect 674230 291571 674282 291623
rect 675382 291571 675434 291623
rect 674902 291053 674954 291105
rect 675382 291053 675434 291105
rect 48310 290979 48362 291031
rect 59638 290979 59690 291031
rect 54646 290905 54698 290957
rect 58774 290831 58826 290883
rect 41782 289351 41834 289403
rect 43126 289351 43178 289403
rect 50710 288907 50762 288959
rect 59542 288907 59594 288959
rect 41782 288167 41834 288219
rect 42934 288167 42986 288219
rect 50326 288019 50378 288071
rect 59158 288019 59210 288071
rect 41878 287723 41930 287775
rect 45814 287723 45866 287775
rect 674326 287723 674378 287775
rect 675382 287723 675434 287775
rect 674998 286761 675050 286813
rect 675382 286761 675434 286813
rect 41590 285133 41642 285185
rect 42934 285133 42986 285185
rect 53206 285133 53258 285185
rect 59254 285133 59306 285185
rect 653782 284097 653834 284149
rect 658006 284097 658058 284149
rect 41782 283801 41834 283853
rect 41782 283505 41834 283557
rect 45334 282395 45386 282447
rect 53014 282395 53066 282447
rect 56086 282395 56138 282447
rect 57622 282395 57674 282447
rect 45526 282321 45578 282373
rect 59638 282321 59690 282373
rect 48118 282247 48170 282299
rect 58582 282247 58634 282299
rect 58774 282247 58826 282299
rect 63382 282173 63434 282225
rect 42070 280101 42122 280153
rect 42838 280101 42890 280153
rect 42166 279879 42218 279931
rect 42934 279879 42986 279931
rect 45334 279435 45386 279487
rect 58390 279435 58442 279487
rect 654262 279435 654314 279487
rect 663766 279435 663818 279487
rect 45622 279361 45674 279413
rect 58582 279361 58634 279413
rect 42166 278547 42218 278599
rect 43030 278547 43082 278599
rect 42070 278473 42122 278525
rect 42934 278473 42986 278525
rect 314902 278325 314954 278377
rect 408310 278325 408362 278377
rect 381046 278251 381098 278303
rect 571414 278251 571466 278303
rect 319510 278177 319562 278229
rect 418966 278177 419018 278229
rect 320950 278103 321002 278155
rect 422518 278103 422570 278155
rect 386518 278029 386570 278081
rect 585622 278029 585674 278081
rect 53014 277955 53066 278007
rect 138262 277955 138314 278007
rect 323830 277955 323882 278007
rect 429622 277955 429674 278007
rect 63382 277881 63434 277933
rect 382390 277881 382442 277933
rect 408886 277881 408938 277933
rect 672502 277881 672554 277933
rect 326422 277807 326474 277859
rect 437014 277807 437066 277859
rect 317878 277733 317930 277785
rect 415702 277733 415754 277785
rect 329302 277659 329354 277711
rect 444118 277659 444170 277711
rect 332374 277585 332426 277637
rect 451222 277585 451274 277637
rect 334966 277511 335018 277563
rect 458230 277511 458282 277563
rect 337846 277437 337898 277489
rect 465334 277437 465386 277489
rect 341014 277363 341066 277415
rect 472438 277363 472490 277415
rect 343894 277289 343946 277341
rect 479542 277289 479594 277341
rect 42070 277215 42122 277267
rect 43126 277215 43178 277267
rect 373846 277215 373898 277267
rect 554038 277215 554090 277267
rect 375094 277141 375146 277193
rect 557590 277141 557642 277193
rect 376822 277067 376874 277119
rect 561142 277067 561194 277119
rect 377974 276993 378026 277045
rect 564694 276993 564746 277045
rect 379414 276919 379466 276971
rect 568246 276919 568298 276971
rect 316630 276845 316682 276897
rect 412150 276845 412202 276897
rect 382294 276771 382346 276823
rect 575254 276771 575306 276823
rect 383638 276697 383690 276749
rect 578806 276697 578858 276749
rect 385366 276623 385418 276675
rect 582358 276623 582410 276675
rect 675766 276623 675818 276675
rect 679798 276623 679850 276675
rect 322102 276549 322154 276601
rect 426358 276549 426410 276601
rect 387958 276475 388010 276527
rect 589462 276475 589514 276527
rect 675286 276475 675338 276527
rect 679702 276475 679754 276527
rect 42838 276401 42890 276453
rect 53302 276401 53354 276453
rect 286102 276401 286154 276453
rect 336502 276401 336554 276453
rect 356182 276401 356234 276453
rect 510262 276401 510314 276453
rect 284470 276327 284522 276379
rect 332950 276327 333002 276379
rect 359158 276327 359210 276379
rect 517366 276327 517418 276379
rect 287350 276253 287402 276305
rect 340054 276253 340106 276305
rect 361750 276253 361802 276305
rect 524470 276253 524522 276305
rect 288694 276179 288746 276231
rect 343606 276179 343658 276231
rect 364630 276179 364682 276231
rect 531574 276179 531626 276231
rect 291862 276105 291914 276157
rect 350710 276105 350762 276157
rect 367702 276105 367754 276157
rect 538678 276105 538730 276157
rect 290326 276031 290378 276083
rect 347158 276031 347210 276083
rect 371926 276031 371978 276083
rect 549334 276031 549386 276083
rect 293014 275957 293066 276009
rect 354262 275957 354314 276009
rect 371062 275957 371114 276009
rect 546934 275957 546986 276009
rect 294646 275883 294698 275935
rect 357814 275883 357866 275935
rect 370294 275883 370346 275935
rect 545782 275883 545834 275935
rect 296470 275809 296522 275861
rect 362518 275809 362570 275861
rect 373462 275809 373514 275861
rect 552790 275809 552842 275861
rect 297334 275735 297386 275787
rect 364918 275735 364970 275787
rect 374614 275735 374666 275787
rect 556342 275735 556394 275787
rect 295894 275661 295946 275713
rect 361366 275661 361418 275713
rect 377494 275661 377546 275713
rect 563446 275661 563498 275713
rect 298966 275587 299018 275639
rect 368470 275587 368522 275639
rect 376246 275587 376298 275639
rect 559894 275587 559946 275639
rect 297814 275513 297866 275565
rect 366070 275513 366122 275565
rect 380566 275513 380618 275565
rect 570550 275513 570602 275565
rect 300214 275439 300266 275491
rect 372022 275439 372074 275491
rect 381814 275439 381866 275491
rect 574102 275439 574154 275491
rect 299158 275365 299210 275417
rect 369622 275365 369674 275417
rect 388918 275365 388970 275417
rect 591862 275365 591914 275417
rect 303286 275291 303338 275343
rect 379126 275291 379178 275343
rect 389590 275291 389642 275343
rect 593014 275291 593066 275343
rect 304438 275217 304490 275269
rect 382582 275217 382634 275269
rect 391990 275217 392042 275269
rect 598966 275217 599018 275269
rect 307318 275143 307370 275195
rect 389686 275143 389738 275195
rect 396310 275143 396362 275195
rect 609526 275143 609578 275195
rect 310390 275069 310442 275121
rect 396790 275069 396842 275121
rect 401782 275069 401834 275121
rect 623734 275069 623786 275121
rect 311638 274995 311690 275047
rect 400342 274995 400394 275047
rect 404950 274995 405002 275047
rect 630838 274995 630890 275047
rect 283030 274921 283082 274973
rect 329398 274921 329450 274973
rect 344566 274921 344618 274973
rect 481942 274921 481994 274973
rect 281782 274847 281834 274899
rect 325846 274847 325898 274899
rect 339094 274847 339146 274899
rect 467734 274847 467786 274899
rect 336022 274773 336074 274825
rect 460630 274773 460682 274825
rect 333142 274699 333194 274751
rect 453526 274699 453578 274751
rect 330454 274625 330506 274677
rect 446422 274625 446474 274677
rect 328822 274551 328874 274603
rect 442870 274551 442922 274603
rect 325942 274477 325994 274529
rect 435862 274477 435914 274529
rect 323350 274403 323402 274455
rect 428758 274403 428810 274455
rect 320182 274329 320234 274381
rect 421654 274329 421706 274381
rect 315958 274255 316010 274307
rect 410998 274255 411050 274307
rect 317302 274181 317354 274233
rect 414550 274181 414602 274233
rect 314710 274107 314762 274159
rect 407446 274107 407498 274159
rect 348502 274033 348554 274085
rect 401494 274033 401546 274085
rect 341206 273959 341258 274011
rect 387382 273959 387434 274011
rect 326806 273885 326858 273937
rect 373174 273885 373226 273937
rect 334294 273811 334346 273863
rect 380278 273811 380330 273863
rect 347062 273737 347114 273789
rect 394486 273737 394538 273789
rect 331222 273663 331274 273715
rect 376726 273663 376778 273715
rect 42934 273515 42986 273567
rect 56182 273515 56234 273567
rect 160438 273515 160490 273567
rect 207478 273515 207530 273567
rect 230134 273515 230186 273567
rect 242902 273515 242954 273567
rect 270262 273515 270314 273567
rect 297526 273515 297578 273567
rect 299350 273515 299402 273567
rect 305302 273515 305354 273567
rect 306934 273515 306986 273567
rect 406582 273589 406634 273641
rect 327094 273515 327146 273567
rect 349462 273515 349514 273567
rect 493750 273515 493802 273567
rect 635542 273515 635594 273567
rect 130870 273441 130922 273493
rect 192982 273441 193034 273493
rect 195862 273441 195914 273493
rect 221494 273441 221546 273493
rect 275350 273441 275402 273493
rect 310486 273441 310538 273493
rect 310582 273441 310634 273493
rect 344758 273441 344810 273493
rect 350038 273441 350090 273493
rect 494902 273441 494954 273493
rect 526966 273441 527018 273493
rect 624982 273441 625034 273493
rect 142678 273367 142730 273419
rect 208150 273367 208202 273419
rect 219574 273367 219626 273419
rect 238678 273367 238730 273419
rect 277078 273367 277130 273419
rect 314038 273367 314090 273419
rect 352438 273367 352490 273419
rect 500854 273367 500906 273419
rect 133270 273293 133322 273345
rect 135286 273293 135338 273345
rect 135574 273293 135626 273345
rect 209782 273293 209834 273345
rect 279670 273293 279722 273345
rect 321142 273293 321194 273345
rect 352630 273293 352682 273345
rect 502006 273293 502058 273345
rect 68278 273219 68330 273271
rect 142582 273219 142634 273271
rect 153334 273219 153386 273271
rect 207382 273219 207434 273271
rect 278230 273219 278282 273271
rect 317590 273219 317642 273271
rect 355510 273219 355562 273271
rect 509110 273219 509162 273271
rect 132022 273145 132074 273197
rect 209878 273145 209930 273197
rect 218326 273145 218378 273197
rect 238102 273145 238154 273197
rect 285622 273145 285674 273197
rect 335350 273145 335402 273197
rect 355030 273145 355082 273197
rect 507958 273145 508010 273197
rect 508246 273145 508298 273197
rect 555190 273145 555242 273197
rect 127318 273071 127370 273123
rect 209974 273071 210026 273123
rect 216022 273071 216074 273123
rect 236950 273071 237002 273123
rect 286774 273071 286826 273123
rect 128470 272997 128522 273049
rect 210166 272997 210218 273049
rect 220726 272997 220778 273049
rect 239158 272997 239210 273049
rect 289942 272997 289994 273049
rect 306646 273071 306698 273123
rect 334198 273071 334250 273123
rect 358582 273071 358634 273123
rect 123766 272923 123818 272975
rect 209014 272923 209066 272975
rect 217174 272923 217226 272975
rect 237622 272923 237674 272975
rect 274198 272923 274250 272975
rect 305302 272923 305354 272975
rect 338902 272997 338954 273049
rect 360982 272997 361034 273049
rect 375190 273071 375242 273123
rect 514966 273071 515018 273123
rect 116662 272849 116714 272901
rect 207094 272849 207146 272901
rect 213622 272849 213674 272901
rect 236278 272849 236330 272901
rect 292246 272849 292298 272901
rect 306838 272923 306890 272975
rect 358966 272923 359018 272975
rect 361270 272923 361322 272975
rect 516214 272997 516266 273049
rect 120214 272775 120266 272827
rect 207862 272775 207914 272827
rect 212470 272775 212522 272827
rect 235702 272775 235754 272827
rect 292726 272775 292778 272827
rect 346006 272849 346058 272901
rect 363574 272849 363626 272901
rect 522070 272923 522122 272975
rect 113110 272701 113162 272753
rect 206230 272701 206282 272753
rect 211222 272701 211274 272753
rect 235030 272701 235082 272753
rect 295414 272701 295466 272753
rect 110806 272627 110858 272679
rect 205462 272627 205514 272679
rect 214774 272627 214826 272679
rect 236470 272627 236522 272679
rect 298294 272701 298346 272753
rect 351862 272775 351914 272827
rect 364150 272775 364202 272827
rect 523318 272849 523370 272901
rect 523990 272849 524042 272901
rect 639094 272849 639146 272901
rect 302038 272627 302090 272679
rect 106102 272553 106154 272605
rect 204022 272553 204074 272605
rect 208918 272553 208970 272605
rect 234358 272553 234410 272605
rect 270550 272553 270602 272605
rect 298678 272553 298730 272605
rect 301366 272553 301418 272605
rect 353110 272701 353162 272753
rect 366550 272701 366602 272753
rect 374518 272701 374570 272753
rect 529174 272775 529226 272827
rect 530422 272701 530474 272753
rect 532822 272701 532874 272753
rect 611926 272701 611978 272753
rect 302326 272627 302378 272679
rect 360214 272627 360266 272679
rect 367126 272627 367178 272679
rect 537430 272627 537482 272679
rect 103702 272479 103754 272531
rect 203542 272479 203594 272531
rect 210070 272479 210122 272531
rect 234550 272479 234602 272531
rect 234934 272479 234986 272531
rect 244822 272479 244874 272531
rect 272278 272479 272330 272531
rect 301942 272479 301994 272531
rect 367222 272553 367274 272605
rect 372694 272553 372746 272605
rect 374326 272479 374378 272531
rect 374518 272553 374570 272605
rect 536278 272553 536330 272605
rect 551638 272479 551690 272531
rect 98998 272405 99050 272457
rect 199126 272405 199178 272457
rect 232534 272405 232586 272457
rect 243670 272405 243722 272457
rect 272758 272405 272810 272457
rect 303478 272405 303530 272457
rect 307126 272405 307178 272457
rect 96598 272331 96650 272383
rect 201622 272331 201674 272383
rect 207670 272331 207722 272383
rect 233878 272331 233930 272383
rect 236086 272331 236138 272383
rect 245302 272331 245354 272383
rect 273430 272331 273482 272383
rect 305782 272331 305834 272383
rect 309910 272331 309962 272383
rect 326902 272405 326954 272457
rect 381430 272405 381482 272457
rect 381526 272405 381578 272457
rect 572950 272405 573002 272457
rect 84790 272257 84842 272309
rect 86326 272257 86378 272309
rect 104854 272257 104906 272309
rect 106486 272257 106538 272309
rect 198262 272257 198314 272309
rect 224374 272257 224426 272309
rect 227830 272257 227882 272309
rect 242134 272257 242186 272309
rect 275158 272257 275210 272309
rect 309334 272257 309386 272309
rect 312790 272257 312842 272309
rect 388534 272331 388586 272383
rect 407446 272331 407498 272383
rect 587158 272331 587210 272383
rect 165142 272183 165194 272235
rect 166966 272183 167018 272235
rect 65878 272109 65930 272161
rect 192406 272183 192458 272235
rect 194710 272183 194762 272235
rect 224470 272183 224522 272235
rect 276310 272183 276362 272235
rect 312886 272183 312938 272235
rect 191158 272109 191210 272161
rect 227158 272109 227210 272161
rect 228982 272109 229034 272161
rect 242422 272109 242474 272161
rect 277750 272109 277802 272161
rect 316438 272183 316490 272235
rect 395638 272257 395690 272309
rect 395926 272257 395978 272309
rect 608374 272257 608426 272309
rect 402742 272183 402794 272235
rect 402934 272183 402986 272235
rect 622582 272183 622634 272235
rect 315478 272109 315530 272161
rect 409846 272109 409898 272161
rect 413686 272109 413738 272161
rect 643894 272109 643946 272161
rect 167542 272035 167594 272087
rect 210646 272035 210698 272087
rect 271030 272035 271082 272087
rect 299926 272035 299978 272087
rect 174646 271961 174698 272013
rect 210550 271961 210602 272013
rect 231382 271961 231434 272013
rect 243094 271961 243146 272013
rect 299446 271961 299498 272013
rect 328246 272035 328298 272087
rect 346966 272035 347018 272087
rect 487798 272035 487850 272087
rect 302326 271961 302378 272013
rect 324694 271961 324746 272013
rect 346486 271961 346538 272013
rect 486646 271961 486698 272013
rect 159286 271887 159338 271939
rect 198646 271887 198698 271939
rect 201814 271887 201866 271939
rect 223702 271887 223754 271939
rect 233686 271887 233738 271939
rect 244054 271887 244106 271939
rect 303958 271887 304010 271939
rect 326902 271887 326954 271939
rect 344086 271887 344138 271939
rect 480694 271887 480746 271939
rect 147382 271813 147434 271865
rect 149686 271813 149738 271865
rect 166294 271813 166346 271865
rect 201526 271813 201578 271865
rect 205366 271813 205418 271865
rect 232630 271813 232682 271865
rect 284950 271813 285002 271865
rect 306646 271813 306698 271865
rect 351382 271813 351434 271865
rect 355414 271813 355466 271865
rect 101302 271739 101354 271791
rect 103606 271739 103658 271791
rect 173398 271739 173450 271791
rect 206038 271739 206090 271791
rect 341494 271739 341546 271791
rect 473686 271813 473738 271865
rect 355606 271739 355658 271791
rect 466582 271739 466634 271791
rect 115510 271665 115562 271717
rect 118006 271665 118058 271717
rect 192310 271665 192362 271717
rect 224566 271665 224618 271717
rect 335446 271665 335498 271717
rect 459478 271665 459530 271717
rect 75286 271591 75338 271643
rect 77686 271591 77738 271643
rect 129718 271591 129770 271643
rect 132406 271591 132458 271643
rect 150934 271591 150986 271643
rect 152374 271591 152426 271643
rect 181750 271591 181802 271643
rect 210454 271591 210506 271643
rect 332566 271591 332618 271643
rect 452374 271591 452426 271643
rect 89494 271517 89546 271569
rect 92086 271517 92138 271569
rect 180502 271517 180554 271569
rect 205846 271517 205898 271569
rect 329974 271517 330026 271569
rect 445270 271517 445322 271569
rect 185206 271443 185258 271495
rect 210358 271443 210410 271495
rect 326902 271443 326954 271495
rect 438166 271443 438218 271495
rect 193558 271369 193610 271421
rect 221686 271369 221738 271421
rect 324022 271369 324074 271421
rect 431062 271369 431114 271421
rect 161590 271295 161642 271347
rect 163894 271295 163946 271347
rect 188758 271295 188810 271347
rect 210262 271295 210314 271347
rect 321430 271295 321482 271347
rect 423958 271295 424010 271347
rect 184054 271221 184106 271273
rect 205750 271221 205802 271273
rect 237238 271221 237290 271273
rect 245590 271221 245642 271273
rect 318358 271221 318410 271273
rect 416950 271221 417002 271273
rect 76534 271147 76586 271199
rect 175798 271147 175850 271199
rect 178294 271147 178346 271199
rect 195670 271147 195722 271199
rect 199414 271147 199466 271199
rect 221590 271147 221642 271199
rect 238486 271147 238538 271199
rect 246070 271147 246122 271199
rect 338614 271147 338666 271199
rect 355606 271147 355658 271199
rect 357910 271147 357962 271199
rect 375190 271147 375242 271199
rect 387286 271147 387338 271199
rect 407446 271147 407498 271199
rect 187606 271073 187658 271125
rect 205942 271073 205994 271125
rect 240790 271073 240842 271125
rect 247222 271073 247274 271125
rect 85942 270999 85994 271051
rect 198550 270999 198602 271051
rect 221878 270999 221930 271051
rect 239350 270999 239402 271051
rect 239542 270999 239594 271051
rect 241270 270999 241322 271051
rect 241942 270999 241994 271051
rect 247702 270999 247754 271051
rect 334102 270999 334154 271051
rect 337750 270999 337802 271051
rect 223030 270925 223082 270977
rect 240022 270925 240074 270977
rect 243190 270925 243242 270977
rect 247990 270925 248042 270977
rect 224278 270851 224330 270903
rect 240502 270851 240554 270903
rect 244342 270851 244394 270903
rect 248662 270851 248714 270903
rect 338710 270851 338762 270903
rect 341302 270851 341354 270903
rect 645238 270851 645290 270903
rect 652342 270851 652394 270903
rect 225430 270777 225482 270829
rect 241078 270777 241130 270829
rect 245494 270777 245546 270829
rect 249142 270777 249194 270829
rect 342742 270777 342794 270829
rect 348310 270777 348362 270829
rect 94198 270703 94250 270755
rect 94966 270703 95018 270755
rect 108406 270703 108458 270755
rect 109366 270703 109418 270755
rect 119062 270703 119114 270755
rect 120886 270703 120938 270755
rect 122614 270703 122666 270755
rect 123766 270703 123818 270755
rect 136822 270703 136874 270755
rect 138166 270703 138218 270755
rect 138262 270703 138314 270755
rect 151606 270703 151658 270755
rect 154486 270703 154538 270755
rect 155446 270703 155498 270755
rect 168694 270703 168746 270755
rect 169846 270703 169898 270755
rect 179350 270703 179402 270755
rect 181366 270703 181418 270755
rect 182902 270703 182954 270755
rect 184246 270703 184298 270755
rect 185494 270703 185546 270755
rect 186454 270703 186506 270755
rect 226582 270703 226634 270755
rect 239542 270703 239594 270755
rect 239638 270703 239690 270755
rect 246454 270703 246506 270755
rect 246742 270703 246794 270755
rect 249622 270703 249674 270755
rect 408982 270703 409034 270755
rect 413398 270703 413450 270755
rect 145078 270629 145130 270681
rect 214486 270629 214538 270681
rect 279286 270629 279338 270681
rect 293302 270629 293354 270681
rect 293398 270629 293450 270681
rect 318838 270629 318890 270681
rect 348118 270629 348170 270681
rect 490198 270629 490250 270681
rect 141526 270555 141578 270607
rect 213814 270555 213866 270607
rect 280150 270555 280202 270607
rect 322390 270555 322442 270607
rect 348406 270555 348458 270607
rect 491350 270555 491402 270607
rect 137974 270481 138026 270533
rect 212662 270481 212714 270533
rect 264694 270481 264746 270533
rect 283318 270481 283370 270533
rect 134422 270407 134474 270459
rect 211894 270407 211946 270459
rect 253942 270407 253994 270459
rect 257302 270407 257354 270459
rect 262006 270407 262058 270459
rect 277462 270407 277514 270459
rect 280630 270407 280682 270459
rect 323542 270481 323594 270533
rect 350710 270481 350762 270533
rect 497302 270481 497354 270533
rect 283702 270407 283754 270459
rect 125014 270333 125066 270385
rect 209494 270333 209546 270385
rect 262486 270333 262538 270385
rect 278614 270333 278666 270385
rect 284182 270333 284234 270385
rect 293302 270407 293354 270459
rect 319990 270407 320042 270459
rect 351286 270407 351338 270459
rect 498454 270407 498506 270459
rect 121462 270259 121514 270311
rect 208342 270259 208394 270311
rect 210550 270259 210602 270311
rect 222838 270259 222890 270311
rect 255286 270259 255338 270311
rect 260854 270259 260906 270311
rect 262966 270259 263018 270311
rect 279766 270259 279818 270311
rect 286294 270259 286346 270311
rect 330646 270333 330698 270385
rect 354070 270333 354122 270385
rect 505558 270333 505610 270385
rect 114358 270185 114410 270237
rect 206422 270185 206474 270237
rect 264886 270185 264938 270237
rect 284566 270185 284618 270237
rect 287926 270185 287978 270237
rect 292918 270185 292970 270237
rect 331798 270259 331850 270311
rect 353686 270259 353738 270311
rect 504406 270259 504458 270311
rect 334102 270185 334154 270237
rect 356758 270185 356810 270237
rect 511510 270185 511562 270237
rect 117910 270111 117962 270163
rect 207574 270111 207626 270163
rect 210454 270111 210506 270163
rect 224758 270111 224810 270163
rect 265366 270111 265418 270163
rect 109558 270037 109610 270089
rect 205270 270037 205322 270089
rect 210358 270037 210410 270089
rect 225526 270037 225578 270089
rect 266518 270037 266570 270089
rect 288502 270111 288554 270163
rect 342454 270111 342506 270163
rect 356950 270111 357002 270163
rect 512662 270111 512714 270163
rect 107254 269963 107306 270015
rect 204694 269963 204746 270015
rect 210262 269963 210314 270015
rect 226678 269963 226730 270015
rect 285718 270037 285770 270089
rect 288022 269963 288074 270015
rect 102550 269889 102602 269941
rect 203350 269889 203402 269941
rect 205846 269889 205898 269941
rect 224086 269889 224138 269941
rect 261814 269889 261866 269941
rect 276214 269889 276266 269941
rect 276406 269889 276458 269941
rect 292822 270037 292874 270089
rect 292918 270037 292970 270089
rect 338710 270037 338762 270089
rect 359830 270037 359882 270089
rect 519766 270037 519818 270089
rect 290614 269963 290666 270015
rect 342742 269963 342794 270015
rect 359350 269963 359402 270015
rect 518518 269963 518570 270015
rect 291094 269889 291146 269941
rect 349558 269889 349610 269941
rect 362710 269889 362762 269941
rect 526870 269889 526922 269941
rect 100150 269815 100202 269867
rect 202870 269815 202922 269867
rect 206038 269815 206090 269867
rect 222358 269815 222410 269867
rect 261238 269815 261290 269867
rect 275062 269815 275114 269867
rect 275254 269815 275306 269867
rect 289270 269815 289322 269867
rect 293974 269815 294026 269867
rect 356662 269815 356714 269867
rect 362230 269815 362282 269867
rect 525622 269815 525674 269867
rect 95446 269741 95498 269793
rect 201142 269741 201194 269793
rect 201526 269741 201578 269793
rect 220534 269741 220586 269793
rect 256246 269741 256298 269793
rect 263254 269741 263306 269793
rect 267766 269741 267818 269793
rect 291574 269741 291626 269793
rect 293494 269741 293546 269793
rect 351382 269741 351434 269793
rect 365302 269741 365354 269793
rect 532726 269741 532778 269793
rect 93046 269667 93098 269719
rect 200950 269667 201002 269719
rect 205942 269667 205994 269719
rect 226006 269667 226058 269719
rect 259894 269667 259946 269719
rect 271510 269667 271562 269719
rect 90646 269593 90698 269645
rect 199702 269593 199754 269645
rect 205750 269593 205802 269645
rect 225238 269593 225290 269645
rect 249046 269593 249098 269645
rect 250294 269593 250346 269645
rect 255766 269593 255818 269645
rect 262102 269593 262154 269645
rect 269686 269593 269738 269645
rect 296374 269667 296426 269719
rect 297046 269667 297098 269719
rect 363670 269667 363722 269719
rect 365494 269667 365546 269719
rect 533878 269667 533930 269719
rect 271702 269593 271754 269645
rect 293782 269593 293834 269645
rect 299638 269593 299690 269645
rect 370774 269593 370826 269645
rect 83638 269519 83690 269571
rect 198070 269519 198122 269571
rect 206518 269519 206570 269571
rect 233398 269519 233450 269571
rect 269206 269519 269258 269571
rect 295126 269519 295178 269571
rect 302614 269519 302666 269571
rect 377878 269519 377930 269571
rect 87190 269445 87242 269497
rect 199030 269445 199082 269497
rect 202966 269445 203018 269497
rect 231958 269445 232010 269497
rect 271510 269445 271562 269497
rect 301078 269445 301130 269497
rect 305686 269445 305738 269497
rect 379606 269445 379658 269497
rect 82390 269371 82442 269423
rect 197398 269371 197450 269423
rect 204118 269371 204170 269423
rect 232150 269371 232202 269423
rect 258646 269371 258698 269423
rect 269110 269371 269162 269423
rect 272950 269371 273002 269423
rect 304630 269371 304682 269423
rect 308278 269371 308330 269423
rect 385078 269593 385130 269645
rect 387382 269593 387434 269645
rect 399190 269593 399242 269645
rect 379894 269519 379946 269571
rect 569398 269519 569450 269571
rect 384118 269445 384170 269497
rect 580054 269445 580106 269497
rect 379798 269371 379850 269423
rect 384982 269371 385034 269423
rect 385078 269371 385130 269423
rect 392086 269371 392138 269423
rect 394390 269371 394442 269423
rect 604822 269371 604874 269423
rect 81238 269297 81290 269349
rect 196822 269297 196874 269349
rect 200662 269297 200714 269349
rect 230998 269297 231050 269349
rect 268630 269297 268682 269349
rect 271702 269297 271754 269349
rect 278902 269297 278954 269349
rect 293398 269297 293450 269349
rect 311158 269297 311210 269349
rect 387382 269297 387434 269349
rect 399958 269297 400010 269349
rect 619030 269297 619082 269349
rect 74134 269223 74186 269275
rect 194998 269223 195050 269275
rect 197110 269223 197162 269275
rect 229558 269223 229610 269275
rect 260566 269223 260618 269275
rect 273910 269223 273962 269275
rect 314230 269223 314282 269275
rect 406294 269223 406346 269275
rect 146230 269149 146282 269201
rect 214966 269149 215018 269201
rect 267094 269149 267146 269201
rect 275254 269149 275306 269201
rect 277558 269149 277610 269201
rect 315286 269149 315338 269201
rect 345430 269149 345482 269201
rect 484246 269149 484298 269201
rect 148630 269075 148682 269127
rect 215734 269075 215786 269127
rect 253366 269075 253418 269127
rect 256150 269075 256202 269127
rect 257014 269075 257066 269127
rect 264406 269075 264458 269127
rect 268438 269075 268490 269127
rect 276406 269075 276458 269127
rect 281302 269075 281354 269127
rect 302326 269075 302378 269127
rect 306358 269075 306410 269127
rect 341206 269075 341258 269127
rect 345238 269075 345290 269127
rect 483094 269075 483146 269127
rect 149782 269001 149834 269053
rect 216214 269001 216266 269053
rect 266038 269001 266090 269053
rect 286870 269001 286922 269053
rect 303766 269001 303818 269053
rect 334294 269001 334346 269053
rect 342646 269001 342698 269053
rect 477142 269001 477194 269053
rect 152182 268927 152234 268979
rect 216694 268927 216746 268979
rect 260086 268927 260138 268979
rect 272662 268927 272714 268979
rect 282070 268927 282122 268979
rect 299350 268927 299402 268979
rect 302038 268927 302090 268979
rect 331222 268927 331274 268979
rect 339766 268927 339818 268979
rect 470134 268927 470186 268979
rect 155734 268853 155786 268905
rect 217366 268853 217418 268905
rect 300694 268853 300746 268905
rect 326806 268853 326858 268905
rect 336886 268853 336938 268905
rect 463030 268853 463082 268905
rect 156886 268779 156938 268831
rect 218134 268779 218186 268831
rect 258166 268779 258218 268831
rect 267958 268779 268010 268831
rect 289174 268779 289226 268831
rect 310582 268779 310634 268831
rect 334294 268779 334346 268831
rect 455926 268779 455978 268831
rect 162838 268705 162890 268757
rect 219286 268705 219338 268757
rect 257686 268705 257738 268757
rect 266806 268705 266858 268757
rect 295222 268705 295274 268757
rect 306838 268705 306890 268757
rect 331222 268705 331274 268757
rect 448822 268705 448874 268757
rect 163990 268631 164042 268683
rect 219958 268631 220010 268683
rect 254614 268631 254666 268683
rect 258550 268631 258602 268683
rect 259414 268631 259466 268683
rect 270358 268631 270410 268683
rect 275830 268631 275882 268683
rect 311734 268631 311786 268683
rect 328342 268631 328394 268683
rect 441718 268631 441770 268683
rect 42166 268557 42218 268609
rect 48310 268557 48362 268609
rect 169750 268557 169802 268609
rect 221206 268557 221258 268609
rect 274678 268557 274730 268609
rect 308182 268557 308234 268609
rect 325750 268557 325802 268609
rect 434614 268557 434666 268609
rect 171094 268483 171146 268535
rect 221782 268483 221834 268535
rect 253174 268483 253226 268535
rect 254998 268483 255050 268535
rect 267286 268483 267338 268535
rect 290422 268483 290474 268535
rect 322582 268483 322634 268535
rect 427510 268483 427562 268535
rect 176950 268409 177002 268461
rect 223414 268409 223466 268461
rect 319702 268409 319754 268461
rect 420502 268409 420554 268461
rect 178198 268335 178250 268387
rect 223606 268335 223658 268387
rect 247894 268335 247946 268387
rect 249814 268335 249866 268387
rect 255094 268335 255146 268387
rect 259702 268335 259754 268387
rect 264118 268335 264170 268387
rect 282166 268335 282218 268387
rect 317110 268335 317162 268387
rect 408982 268335 409034 268387
rect 198646 268261 198698 268313
rect 218614 268261 218666 268313
rect 221494 268261 221546 268313
rect 229078 268261 229130 268313
rect 309238 268261 309290 268313
rect 347062 268261 347114 268313
rect 192982 268187 193034 268239
rect 210742 268187 210794 268239
rect 223702 268187 223754 268239
rect 231478 268187 231530 268239
rect 257494 268187 257546 268239
rect 265654 268187 265706 268239
rect 209782 268113 209834 268165
rect 212374 268113 212426 268165
rect 212470 268113 212522 268165
rect 218902 268113 218954 268165
rect 224374 268113 224426 268165
rect 230038 268113 230090 268165
rect 263638 268113 263690 268165
rect 281014 268187 281066 268239
rect 312310 268187 312362 268239
rect 348502 268187 348554 268239
rect 408502 268187 408554 268239
rect 640342 268187 640394 268239
rect 330742 268113 330794 268165
rect 343798 268113 343850 268165
rect 371254 268113 371306 268165
rect 548086 268113 548138 268165
rect 207382 268039 207434 268091
rect 216886 268039 216938 268091
rect 224470 268039 224522 268091
rect 228406 268039 228458 268091
rect 252694 268039 252746 268091
rect 253750 268039 253802 268091
rect 333622 268039 333674 268091
rect 351382 268039 351434 268091
rect 209878 267965 209930 268017
rect 211414 267965 211466 268017
rect 221590 267965 221642 268017
rect 230518 267965 230570 268017
rect 336694 267965 336746 268017
rect 357622 267965 357674 268017
rect 210646 267891 210698 267943
rect 221014 267891 221066 267943
rect 221686 267891 221738 267943
rect 227830 267891 227882 267943
rect 339286 267891 339338 267943
rect 362806 267891 362858 267943
rect 199126 267817 199178 267869
rect 202294 267817 202346 267869
rect 207478 267817 207530 267869
rect 212470 267817 212522 267869
rect 224566 267817 224618 267869
rect 227638 267817 227690 267869
rect 282550 267817 282602 267869
rect 299446 267817 299498 267869
rect 342166 267817 342218 267869
rect 365686 267817 365738 267869
rect 401302 267817 401354 267869
rect 402934 267817 402986 267869
rect 409942 267817 409994 267869
rect 413686 267817 413738 267869
rect 388726 267743 388778 267795
rect 645238 267743 645290 267795
rect 351958 267669 352010 267721
rect 499606 267669 499658 267721
rect 354838 267595 354890 267647
rect 506710 267595 506762 267647
rect 357430 267521 357482 267573
rect 513814 267521 513866 267573
rect 360310 267447 360362 267499
rect 520918 267447 520970 267499
rect 363382 267373 363434 267425
rect 528022 267373 528074 267425
rect 365974 267299 366026 267351
rect 535126 267299 535178 267351
rect 368950 267225 369002 267277
rect 542230 267225 542282 267277
rect 372502 267151 372554 267203
rect 550486 267151 550538 267203
rect 384886 267077 384938 267129
rect 581206 267077 581258 267129
rect 386038 267003 386090 267055
rect 584758 267003 584810 267055
rect 387766 266929 387818 266981
rect 588310 266929 588362 266981
rect 301846 266855 301898 266907
rect 375286 266855 375338 266907
rect 393238 266855 393290 266907
rect 602518 266855 602570 266907
rect 305014 266781 305066 266833
rect 383542 266781 383594 266833
rect 394678 266781 394730 266833
rect 606070 266781 606122 266833
rect 306166 266707 306218 266759
rect 386134 266707 386186 266759
rect 397558 266707 397610 266759
rect 613078 266707 613130 266759
rect 308086 266633 308138 266685
rect 390934 266633 390986 266685
rect 398230 266633 398282 266685
rect 614326 266633 614378 266685
rect 308758 266559 308810 266611
rect 392950 266559 393002 266611
rect 400630 266559 400682 266611
rect 620182 266559 620234 266611
rect 310678 266485 310730 266537
rect 398038 266485 398090 266537
rect 403222 266485 403274 266537
rect 627286 266485 627338 266537
rect 313078 266411 313130 266463
rect 403894 266411 403946 266463
rect 406102 266411 406154 266463
rect 634390 266411 634442 266463
rect 313558 266337 313610 266389
rect 405046 266337 405098 266389
rect 409174 266337 409226 266389
rect 641494 266337 641546 266389
rect 348886 266263 348938 266315
rect 492598 266263 492650 266315
rect 346006 266189 346058 266241
rect 485494 266189 485546 266241
rect 343318 266115 343370 266167
rect 478390 266115 478442 266167
rect 340246 266041 340298 266093
rect 471286 266041 471338 266093
rect 337366 265967 337418 266019
rect 464182 265967 464234 266019
rect 334774 265893 334826 265945
rect 457078 265893 457130 265945
rect 331894 265819 331946 265871
rect 449974 265819 450026 265871
rect 408022 265745 408074 265797
rect 523990 265745 524042 265797
rect 327574 265671 327626 265723
rect 439318 265671 439370 265723
rect 324502 265597 324554 265649
rect 432310 265597 432362 265649
rect 321622 265523 321674 265575
rect 425206 265523 425258 265575
rect 319030 265449 319082 265501
rect 418102 265449 418154 265501
rect 656566 265375 656618 265427
rect 676246 265375 676298 265427
rect 656470 265227 656522 265279
rect 676150 265227 676202 265279
rect 656086 265079 656138 265131
rect 676342 265079 676394 265131
rect 23158 265005 23210 265057
rect 43510 265005 43562 265057
rect 671830 265005 671882 265057
rect 673270 265005 673322 265057
rect 676246 265005 676298 265057
rect 43318 264931 43370 264983
rect 44278 264931 44330 264983
rect 669814 264931 669866 264983
rect 43222 264857 43274 264909
rect 44182 264857 44234 264909
rect 669622 264857 669674 264909
rect 365686 264783 365738 264835
rect 475990 264783 476042 264835
rect 325366 264709 325418 264761
rect 433462 264709 433514 264761
rect 362806 264635 362858 264687
rect 468886 264635 468938 264687
rect 357622 264561 357674 264613
rect 461782 264561 461834 264613
rect 328054 264487 328106 264539
rect 440566 264487 440618 264539
rect 343798 264413 343850 264465
rect 447670 264413 447722 264465
rect 351382 264339 351434 264391
rect 454774 264339 454826 264391
rect 399382 264043 399434 264095
rect 411670 264043 411722 264095
rect 390838 263969 390890 264021
rect 596566 263969 596618 264021
rect 392278 263895 392330 263947
rect 600118 263895 600170 263947
rect 395446 263821 395498 263873
rect 607222 263821 607274 263873
rect 401110 263747 401162 263799
rect 403990 263673 404042 263725
rect 411670 263747 411722 263799
rect 617878 263747 617930 263799
rect 23542 263599 23594 263651
rect 44182 263599 44234 263651
rect 405430 263599 405482 263651
rect 621430 263673 621482 263725
rect 23062 263525 23114 263577
rect 44278 263525 44330 263577
rect 409654 263525 409706 263577
rect 628438 263599 628490 263651
rect 631990 263525 632042 263577
rect 642646 263451 642698 263503
rect 23350 262119 23402 262171
rect 43318 262119 43370 262171
rect 420406 262119 420458 262171
rect 606166 262119 606218 262171
rect 675190 262119 675242 262171
rect 676246 262119 676298 262171
rect 674806 259899 674858 259951
rect 676246 259899 676298 259951
rect 673270 259529 673322 259581
rect 673462 259529 673514 259581
rect 674710 259307 674762 259359
rect 676054 259307 676106 259359
rect 420406 259233 420458 259285
rect 606262 259233 606314 259285
rect 675286 259233 675338 259285
rect 676246 259233 676298 259285
rect 151606 257753 151658 257805
rect 169750 257753 169802 257805
rect 187222 257753 187274 257805
rect 189718 257753 189770 257805
rect 41782 256421 41834 256473
rect 56086 256421 56138 256473
rect 674614 256421 674666 256473
rect 675958 256421 676010 256473
rect 41590 256347 41642 256399
rect 58966 256347 59018 256399
rect 420406 256347 420458 256399
rect 606358 256347 606410 256399
rect 674902 256347 674954 256399
rect 676054 256347 676106 256399
rect 41782 255977 41834 256029
rect 53206 255977 53258 256029
rect 41782 255533 41834 255585
rect 43414 255533 43466 255585
rect 41782 255015 41834 255067
rect 43414 255015 43466 255067
rect 47926 254941 47978 254993
rect 186070 254941 186122 254993
rect 48022 254867 48074 254919
rect 186262 254867 186314 254919
rect 420406 253461 420458 253513
rect 603286 253461 603338 253513
rect 646678 253461 646730 253513
rect 679798 253461 679850 253513
rect 141046 252499 141098 252551
rect 171382 252499 171434 252551
rect 106486 252425 106538 252477
rect 156886 252425 156938 252477
rect 97846 252351 97898 252403
rect 154006 252351 154058 252403
rect 103606 252277 103658 252329
rect 159766 252277 159818 252329
rect 109366 252203 109418 252255
rect 177046 252203 177098 252255
rect 86326 252129 86378 252181
rect 165526 252129 165578 252181
rect 94966 252055 95018 252107
rect 174166 252055 174218 252107
rect 92086 251981 92138 252033
rect 182806 251981 182858 252033
rect 670390 250649 670442 250701
rect 675382 250649 675434 250701
rect 420406 250575 420458 250627
rect 603382 250575 603434 250627
rect 120886 249835 120938 249887
rect 145558 249835 145610 249887
rect 132406 249761 132458 249813
rect 162742 249761 162794 249813
rect 135286 249687 135338 249739
rect 168502 249687 168554 249739
rect 118006 249613 118058 249665
rect 156982 249613 157034 249665
rect 138166 249539 138218 249591
rect 180022 249539 180074 249591
rect 126646 249465 126698 249517
rect 177238 249465 177290 249517
rect 123766 249391 123818 249443
rect 174454 249391 174506 249443
rect 80566 249317 80618 249369
rect 145462 249317 145514 249369
rect 77686 249243 77738 249295
rect 145366 249243 145418 249295
rect 48214 249169 48266 249221
rect 186742 249169 186794 249221
rect 47734 249095 47786 249147
rect 186454 249095 186506 249147
rect 674806 247911 674858 247963
rect 675382 247911 675434 247963
rect 420310 247763 420362 247815
rect 603478 247763 603530 247815
rect 420406 247689 420458 247741
rect 629206 247689 629258 247741
rect 655894 247615 655946 247667
rect 670390 247615 670442 247667
rect 674806 247023 674858 247075
rect 675478 247023 675530 247075
rect 112246 246653 112298 246705
rect 185782 246653 185834 246705
rect 47542 246579 47594 246631
rect 186358 246579 186410 246631
rect 47638 246505 47690 246557
rect 186646 246505 186698 246557
rect 47446 246431 47498 246483
rect 186550 246431 186602 246483
rect 45814 246357 45866 246409
rect 186934 246357 186986 246409
rect 44854 246283 44906 246335
rect 186166 246283 186218 246335
rect 44566 246209 44618 246261
rect 185974 246209 186026 246261
rect 674902 245839 674954 245891
rect 675382 245839 675434 245891
rect 41590 245469 41642 245521
rect 43030 245469 43082 245521
rect 41686 245395 41738 245447
rect 42838 245395 42890 245447
rect 41878 245025 41930 245077
rect 42934 245025 42986 245077
rect 44662 244951 44714 245003
rect 186838 244951 186890 245003
rect 41590 244877 41642 244929
rect 142486 244877 142538 244929
rect 41686 244803 41738 244855
rect 159958 244803 160010 244855
rect 420406 244803 420458 244855
rect 629302 244803 629354 244855
rect 41494 244655 41546 244707
rect 42742 244655 42794 244707
rect 169750 243027 169802 243079
rect 180118 243027 180170 243079
rect 44758 242805 44810 242857
rect 185686 242805 185738 242857
rect 44854 242731 44906 242783
rect 185878 242731 185930 242783
rect 674614 242731 674666 242783
rect 675382 242731 675434 242783
rect 44566 242657 44618 242709
rect 187030 242657 187082 242709
rect 41590 242583 41642 242635
rect 142678 242583 142730 242635
rect 420310 241917 420362 241969
rect 600406 241917 600458 241969
rect 41782 240585 41834 240637
rect 41782 240363 41834 240415
rect 368662 239919 368714 239971
rect 412054 239919 412106 239971
rect 413014 239919 413066 239971
rect 442198 239919 442250 239971
rect 409558 239845 409610 239897
rect 412150 239845 412202 239897
rect 350710 239771 350762 239823
rect 508630 239771 508682 239823
rect 360022 239697 360074 239749
rect 434614 239697 434666 239749
rect 366550 239623 366602 239675
rect 446710 239623 446762 239675
rect 396694 239549 396746 239601
rect 412246 239549 412298 239601
rect 412918 239549 412970 239601
rect 495766 239549 495818 239601
rect 383062 239475 383114 239527
rect 470902 239475 470954 239527
rect 371638 239401 371690 239453
rect 458806 239401 458858 239453
rect 406102 239327 406154 239379
rect 412342 239327 412394 239379
rect 412822 239327 412874 239379
rect 502582 239327 502634 239379
rect 378454 239253 378506 239305
rect 488278 239253 488330 239305
rect 398422 239179 398474 239231
rect 532822 239179 532874 239231
rect 411766 239105 411818 239157
rect 412630 239105 412682 239157
rect 420310 239105 420362 239157
rect 599062 239105 599114 239157
rect 380854 239031 380906 239083
rect 412438 239031 412490 239083
rect 324406 238957 324458 239009
rect 455158 238957 455210 239009
rect 323926 238883 323978 238935
rect 455062 238883 455114 238935
rect 326710 238809 326762 238861
rect 462550 238809 462602 238861
rect 328918 238735 328970 238787
rect 464758 238735 464810 238787
rect 329878 238661 329930 238713
rect 468598 238661 468650 238713
rect 332662 238587 332714 238639
rect 474646 238587 474698 238639
rect 335734 238513 335786 238565
rect 480694 238513 480746 238565
rect 336694 238439 336746 238491
rect 479158 238439 479210 238491
rect 338998 238365 339050 238417
rect 486742 238365 486794 238417
rect 341782 238291 341834 238343
rect 492790 238291 492842 238343
rect 345334 238217 345386 238269
rect 500278 238217 500330 238269
rect 346678 238143 346730 238195
rect 503350 238143 503402 238195
rect 349942 238069 349994 238121
rect 509398 238069 509450 238121
rect 353494 237995 353546 238047
rect 514678 237995 514730 238047
rect 352726 237921 352778 237973
rect 512758 237921 512810 237973
rect 355702 237847 355754 237899
rect 521494 237847 521546 237899
rect 358582 237773 358634 237825
rect 526006 237773 526058 237825
rect 363094 237699 363146 237751
rect 535126 237699 535178 237751
rect 275350 237625 275402 237677
rect 357718 237625 357770 237677
rect 361750 237625 361802 237677
rect 533494 237625 533546 237677
rect 277078 237551 277130 237603
rect 363670 237551 363722 237603
rect 364438 237551 364490 237603
rect 535798 237551 535850 237603
rect 320854 237477 320906 237529
rect 449302 237477 449354 237529
rect 317590 237403 317642 237455
rect 444502 237403 444554 237455
rect 317110 237329 317162 237381
rect 441430 237329 441482 237381
rect 314806 237255 314858 237307
rect 438358 237255 438410 237307
rect 311542 237181 311594 237233
rect 432406 237181 432458 237233
rect 308566 237107 308618 237159
rect 411478 237107 411530 237159
rect 411670 237107 411722 237159
rect 412726 237107 412778 237159
rect 310774 237033 310826 237085
rect 411190 237033 411242 237085
rect 411574 237033 411626 237085
rect 412822 237033 412874 237085
rect 305782 236959 305834 237011
rect 420310 236959 420362 237011
rect 300214 236885 300266 236937
rect 407158 236885 407210 236937
rect 408982 236885 409034 236937
rect 413974 236885 414026 236937
rect 279862 236811 279914 236863
rect 368854 236811 368906 236863
rect 382582 236811 382634 236863
rect 388726 236811 388778 236863
rect 406006 236811 406058 236863
rect 409174 236811 409226 236863
rect 411478 236811 411530 236863
rect 426358 236811 426410 236863
rect 278422 236737 278474 236789
rect 366742 236737 366794 236789
rect 388342 236737 388394 236789
rect 389014 236737 389066 236789
rect 389398 236737 389450 236789
rect 409366 236737 409418 236789
rect 411190 236737 411242 236789
rect 428662 236737 428714 236789
rect 42166 236663 42218 236715
rect 42742 236663 42794 236715
rect 377782 236663 377834 236715
rect 388630 236663 388682 236715
rect 408694 236663 408746 236715
rect 413686 236663 413738 236715
rect 408790 236589 408842 236641
rect 413398 236589 413450 236641
rect 42742 236515 42794 236567
rect 43030 236515 43082 236567
rect 387958 236515 388010 236567
rect 388630 236515 388682 236567
rect 405910 236515 405962 236567
rect 412534 236515 412586 236567
rect 411478 236441 411530 236493
rect 412918 236441 412970 236493
rect 414550 236367 414602 236419
rect 430102 236367 430154 236419
rect 385942 236293 385994 236345
rect 492022 236293 492074 236345
rect 397366 236219 397418 236271
rect 505654 236219 505706 236271
rect 240214 236071 240266 236123
rect 263734 236071 263786 236123
rect 273046 236071 273098 236123
rect 305110 236071 305162 236123
rect 352150 236071 352202 236123
rect 511606 236145 511658 236197
rect 410038 236071 410090 236123
rect 528502 236071 528554 236123
rect 208438 235997 208490 236049
rect 223222 235997 223274 236049
rect 247990 235997 248042 236049
rect 273718 235997 273770 236049
rect 287062 235997 287114 236049
rect 318262 235997 318314 236049
rect 362518 235997 362570 236049
rect 392758 235997 392810 236049
rect 207478 235923 207530 235975
rect 223990 235923 224042 235975
rect 243286 235923 243338 235975
rect 270934 235923 270986 235975
rect 277558 235923 277610 235975
rect 313942 235923 313994 235975
rect 319894 235923 319946 235975
rect 366550 235923 366602 235975
rect 406006 235997 406058 236049
rect 406294 235997 406346 236049
rect 414646 235997 414698 236049
rect 209686 235849 209738 235901
rect 226198 235849 226250 235901
rect 234262 235849 234314 235901
rect 264694 235849 264746 235901
rect 276118 235849 276170 235901
rect 310102 235849 310154 235901
rect 313846 235849 313898 235901
rect 360022 235849 360074 235901
rect 208918 235775 208970 235827
rect 226966 235775 227018 235827
rect 237526 235775 237578 235827
rect 267958 235775 268010 235827
rect 279286 235775 279338 235827
rect 318358 235775 318410 235827
rect 326134 235775 326186 235827
rect 371638 235849 371690 235901
rect 211222 235701 211274 235753
rect 229270 235701 229322 235753
rect 231190 235701 231242 235753
rect 259030 235701 259082 235753
rect 262870 235701 262922 235753
rect 305014 235701 305066 235753
rect 364054 235701 364106 235753
rect 371830 235849 371882 235901
rect 392566 235849 392618 235901
rect 386710 235775 386762 235827
rect 411670 235923 411722 235975
rect 401206 235849 401258 235901
rect 411766 235849 411818 235901
rect 393142 235775 393194 235827
rect 406102 235775 406154 235827
rect 410902 235775 410954 235827
rect 413014 235775 413066 235827
rect 378838 235701 378890 235753
rect 392854 235701 392906 235753
rect 392950 235701 393002 235753
rect 398422 235701 398474 235753
rect 398614 235701 398666 235753
rect 528406 235701 528458 235753
rect 210646 235627 210698 235679
rect 230038 235627 230090 235679
rect 285142 235627 285194 235679
rect 323350 235627 323402 235679
rect 326230 235627 326282 235679
rect 460246 235627 460298 235679
rect 210070 235553 210122 235605
rect 227830 235553 227882 235605
rect 236470 235553 236522 235605
rect 282934 235553 282986 235605
rect 286678 235553 286730 235605
rect 326806 235553 326858 235605
rect 332566 235553 332618 235605
rect 472342 235553 472394 235605
rect 212950 235479 213002 235531
rect 232342 235479 232394 235531
rect 238006 235479 238058 235531
rect 285910 235479 285962 235531
rect 290326 235479 290378 235531
rect 334294 235479 334346 235531
rect 348886 235479 348938 235531
rect 397366 235479 397418 235531
rect 42166 235405 42218 235457
rect 42838 235405 42890 235457
rect 211990 235405 212042 235457
rect 233014 235405 233066 235457
rect 242134 235405 242186 235457
rect 293398 235405 293450 235457
rect 295222 235405 295274 235457
rect 348694 235405 348746 235457
rect 392854 235405 392906 235457
rect 396694 235405 396746 235457
rect 396790 235405 396842 235457
rect 588982 235479 589034 235531
rect 403030 235405 403082 235457
rect 588694 235405 588746 235457
rect 206998 235331 207050 235383
rect 221782 235331 221834 235383
rect 223894 235331 223946 235383
rect 244726 235331 244778 235383
rect 254230 235331 254282 235383
rect 306742 235331 306794 235383
rect 339478 235331 339530 235383
rect 395254 235331 395306 235383
rect 398518 235331 398570 235383
rect 590422 235331 590474 235383
rect 214198 235257 214250 235309
rect 235318 235257 235370 235309
rect 239350 235257 239402 235309
rect 287350 235257 287402 235309
rect 288886 235257 288938 235309
rect 345718 235257 345770 235309
rect 396310 235257 396362 235309
rect 588886 235257 588938 235309
rect 220630 235183 220682 235235
rect 241846 235183 241898 235235
rect 249718 235183 249770 235235
rect 302326 235183 302378 235235
rect 305206 235183 305258 235235
rect 365686 235183 365738 235235
rect 374518 235183 374570 235235
rect 381622 235183 381674 235235
rect 394966 235183 395018 235235
rect 403030 235183 403082 235235
rect 403126 235183 403178 235235
rect 587926 235183 587978 235235
rect 206134 235109 206186 235161
rect 215926 235109 215978 235161
rect 232918 235109 232970 235161
rect 262006 235109 262058 235161
rect 266134 235109 266186 235161
rect 324502 235109 324554 235161
rect 327670 235109 327722 235161
rect 390358 235109 390410 235161
rect 392182 235109 392234 235161
rect 592342 235109 592394 235161
rect 203254 235035 203306 235087
rect 211510 235035 211562 235087
rect 213430 235035 213482 235087
rect 233398 235035 233450 235087
rect 235702 235035 235754 235087
rect 265270 235035 265322 235087
rect 268918 235035 268970 235087
rect 331414 235035 331466 235087
rect 334966 235035 335018 235087
rect 393526 235035 393578 235087
rect 394582 235035 394634 235087
rect 597718 235035 597770 235087
rect 208822 234961 208874 235013
rect 224758 234961 224810 235013
rect 225526 234961 225578 235013
rect 260182 234961 260234 235013
rect 260278 234961 260330 235013
rect 323254 234961 323306 235013
rect 333430 234961 333482 235013
rect 211030 234887 211082 234939
rect 231574 234887 231626 234939
rect 243862 234887 243914 234939
rect 296470 234887 296522 234939
rect 296566 234887 296618 234939
rect 361942 234887 361994 234939
rect 209302 234813 209354 234865
rect 228502 234813 228554 234865
rect 229750 234813 229802 234865
rect 253558 234813 253610 234865
rect 257494 234813 257546 234865
rect 308182 234813 308234 234865
rect 321622 234813 321674 234865
rect 378550 234813 378602 234865
rect 389878 234961 389930 235013
rect 403126 234961 403178 235013
rect 403606 234961 403658 235013
rect 615862 234961 615914 235013
rect 381622 234887 381674 234939
rect 398806 234887 398858 234939
rect 406678 234887 406730 234939
rect 621814 234887 621866 234939
rect 395734 234813 395786 234865
rect 398230 234813 398282 234865
rect 405046 234813 405098 234865
rect 407926 234813 407978 234865
rect 408790 234813 408842 234865
rect 409942 234813 409994 234865
rect 627862 234813 627914 234865
rect 202870 234739 202922 234791
rect 214774 234739 214826 234791
rect 225142 234739 225194 234791
rect 247702 234739 247754 234791
rect 251158 234739 251210 234791
rect 304150 234739 304202 234791
rect 315286 234739 315338 234791
rect 396406 234739 396458 234791
rect 396502 234739 396554 234791
rect 406870 234739 406922 234791
rect 412150 234739 412202 234791
rect 632374 234739 632426 234791
rect 204790 234665 204842 234717
rect 214870 234665 214922 234717
rect 222358 234665 222410 234717
rect 243958 234665 244010 234717
rect 246646 234665 246698 234717
rect 299350 234665 299402 234717
rect 301750 234665 301802 234717
rect 398902 234665 398954 234717
rect 411286 234665 411338 234717
rect 630934 234665 630986 234717
rect 42166 234591 42218 234643
rect 42742 234591 42794 234643
rect 202006 234591 202058 234643
rect 213430 234591 213482 234643
rect 251062 234591 251114 234643
rect 273622 234591 273674 234643
rect 280630 234591 280682 234643
rect 321046 234591 321098 234643
rect 323542 234591 323594 234643
rect 434902 234591 434954 234643
rect 204214 234517 204266 234569
rect 215542 234517 215594 234569
rect 237046 234517 237098 234569
rect 258070 234517 258122 234569
rect 262486 234517 262538 234569
rect 290902 234517 290954 234569
rect 295702 234517 295754 234569
rect 341398 234517 341450 234569
rect 345910 234517 345962 234569
rect 400342 234517 400394 234569
rect 410806 234517 410858 234569
rect 522646 234517 522698 234569
rect 206518 234443 206570 234495
rect 204406 234369 204458 234421
rect 210166 234369 210218 234421
rect 201526 234295 201578 234347
rect 211894 234295 211946 234347
rect 250486 234443 250538 234495
rect 269398 234443 269450 234495
rect 271606 234443 271658 234495
rect 301270 234443 301322 234495
rect 306262 234443 306314 234495
rect 358390 234443 358442 234495
rect 383638 234443 383690 234495
rect 396502 234443 396554 234495
rect 396598 234443 396650 234495
rect 408022 234443 408074 234495
rect 409270 234443 409322 234495
rect 521206 234443 521258 234495
rect 215926 234369 215978 234421
rect 221014 234369 221066 234421
rect 235606 234369 235658 234421
rect 250582 234369 250634 234421
rect 255286 234369 255338 234421
rect 277078 234369 277130 234421
rect 283990 234369 284042 234421
rect 311350 234369 311402 234421
rect 314422 234369 314474 234421
rect 423382 234369 423434 234421
rect 222454 234295 222506 234347
rect 239830 234295 239882 234347
rect 260470 234295 260522 234347
rect 261238 234295 261290 234347
rect 288022 234295 288074 234347
rect 308470 234295 308522 234347
rect 416374 234295 416426 234347
rect 207862 234221 207914 234273
rect 200278 234147 200330 234199
rect 210358 234147 210410 234199
rect 214870 234221 214922 234273
rect 219382 234221 219434 234273
rect 244342 234221 244394 234273
rect 264886 234221 264938 234273
rect 268534 234221 268586 234273
rect 293782 234221 293834 234273
rect 312694 234221 312746 234273
rect 418294 234221 418346 234273
rect 225526 234147 225578 234199
rect 256534 234147 256586 234199
rect 279286 234147 279338 234199
rect 283894 234147 283946 234199
rect 320758 234147 320810 234199
rect 330454 234147 330506 234199
rect 374710 234147 374762 234199
rect 378550 234147 378602 234199
rect 385942 234147 385994 234199
rect 395830 234147 395882 234199
rect 403126 234147 403178 234199
rect 403222 234147 403274 234199
rect 498550 234147 498602 234199
rect 200182 234073 200234 234125
rect 208822 234073 208874 234125
rect 210166 234073 210218 234125
rect 217942 234073 217994 234125
rect 247414 234073 247466 234125
rect 266326 234073 266378 234125
rect 267094 234073 267146 234125
rect 290998 234073 291050 234125
rect 294838 234073 294890 234125
rect 339094 234073 339146 234125
rect 358006 234073 358058 234125
rect 394870 234073 394922 234125
rect 401782 234073 401834 234125
rect 486646 234073 486698 234125
rect 42070 233999 42122 234051
rect 42934 233999 42986 234051
rect 198742 233999 198794 234051
rect 207382 233999 207434 234051
rect 198358 233925 198410 233977
rect 205942 233925 205994 233977
rect 206902 233925 206954 233977
rect 220246 233999 220298 234051
rect 259798 233999 259850 234051
rect 281878 233999 281930 234051
rect 299830 233999 299882 234051
rect 344662 233999 344714 234051
rect 365878 233999 365930 234051
rect 382774 233999 382826 234051
rect 399094 233999 399146 234051
rect 400150 233999 400202 234051
rect 400246 233999 400298 234051
rect 211510 233925 211562 233977
rect 216502 233925 216554 233977
rect 296086 233925 296138 233977
rect 339766 233925 339818 233977
rect 341206 233925 341258 233977
rect 378454 233925 378506 233977
rect 382102 233925 382154 233977
rect 400726 233925 400778 233977
rect 408022 233999 408074 234051
rect 475222 233999 475274 234051
rect 479254 233925 479306 233977
rect 197494 233851 197546 233903
rect 204310 233851 204362 233903
rect 196918 233777 196970 233829
rect 202870 233777 202922 233829
rect 205174 233777 205226 233829
rect 214486 233851 214538 233903
rect 253462 233851 253514 233903
rect 270838 233851 270890 233903
rect 294454 233851 294506 233903
rect 331222 233851 331274 233903
rect 339862 233851 339914 233903
rect 351382 233851 351434 233903
rect 361270 233851 361322 233903
rect 211606 233777 211658 233829
rect 230710 233777 230762 233829
rect 242902 233777 242954 233829
rect 260854 233777 260906 233829
rect 267478 233777 267530 233829
rect 285046 233777 285098 233829
rect 297238 233777 297290 233829
rect 328342 233777 328394 233829
rect 332182 233777 332234 233829
rect 383062 233777 383114 233829
rect 432022 233851 432074 233903
rect 400726 233777 400778 233829
rect 411766 233777 411818 233829
rect 197974 233703 198026 233755
rect 203638 233703 203690 233755
rect 203926 233703 203978 233755
rect 214198 233703 214250 233755
rect 195670 233629 195722 233681
rect 201334 233629 201386 233681
rect 202486 233629 202538 233681
rect 212566 233629 212618 233681
rect 192886 233555 192938 233607
rect 195286 233555 195338 233607
rect 195574 233555 195626 233607
rect 199798 233555 199850 233607
rect 201046 233555 201098 233607
rect 209686 233555 209738 233607
rect 194230 233481 194282 233533
rect 198358 233481 198410 233533
rect 199126 233481 199178 233533
rect 205078 233481 205130 233533
rect 205558 233481 205610 233533
rect 218710 233703 218762 233755
rect 258358 233703 258410 233755
rect 278230 233703 278282 233755
rect 304822 233703 304874 233755
rect 334102 233703 334154 233755
rect 338614 233703 338666 233755
rect 464566 233703 464618 233755
rect 214486 233629 214538 233681
rect 217174 233629 217226 233681
rect 287446 233629 287498 233681
rect 311254 233629 311306 233681
rect 324790 233629 324842 233681
rect 342646 233629 342698 233681
rect 343510 233629 343562 233681
rect 411478 233629 411530 233681
rect 259894 233555 259946 233607
rect 267766 233555 267818 233607
rect 288406 233555 288458 233607
rect 313846 233555 313898 233607
rect 329302 233555 329354 233607
rect 449302 233555 449354 233607
rect 240598 233481 240650 233533
rect 290422 233481 290474 233533
rect 297142 233481 297194 233533
rect 319606 233481 319658 233533
rect 335350 233481 335402 233533
rect 463606 233481 463658 233533
rect 194614 233407 194666 233459
rect 196054 233407 196106 233459
rect 196534 233407 196586 233459
rect 200566 233407 200618 233459
rect 200662 233407 200714 233459
rect 208150 233407 208202 233459
rect 233398 233407 233450 233459
rect 235990 233407 236042 233459
rect 264406 233407 264458 233459
rect 271894 233407 271946 233459
rect 292918 233407 292970 233459
rect 311062 233407 311114 233459
rect 317206 233407 317258 233459
rect 410902 233407 410954 233459
rect 192406 233333 192458 233385
rect 193750 233333 193802 233385
rect 193846 233333 193898 233385
rect 196822 233333 196874 233385
rect 197878 233333 197930 233385
rect 202102 233333 202154 233385
rect 202390 233333 202442 233385
rect 211126 233333 211178 233385
rect 228406 233333 228458 233385
rect 236374 233333 236426 233385
rect 261622 233333 261674 233385
rect 269014 233333 269066 233385
rect 270550 233333 270602 233385
rect 274678 233333 274730 233385
rect 311158 233333 311210 233385
rect 414550 233333 414602 233385
rect 193462 233259 193514 233311
rect 194614 233259 194666 233311
rect 195190 233259 195242 233311
rect 195862 233259 195914 233311
rect 196150 233259 196202 233311
rect 199126 233259 199178 233311
rect 199702 233259 199754 233311
rect 206614 233259 206666 233311
rect 226678 233259 226730 233311
rect 238966 233259 239018 233311
rect 257974 233259 258026 233311
rect 269110 233259 269162 233311
rect 270262 233259 270314 233311
rect 273526 233259 273578 233311
rect 320278 233259 320330 233311
rect 448246 233259 448298 233311
rect 262102 233185 262154 233237
rect 334198 233185 334250 233237
rect 340822 233185 340874 233237
rect 491254 233185 491306 233237
rect 495382 233185 495434 233237
rect 622678 233185 622730 233237
rect 260662 233111 260714 233163
rect 331318 233111 331370 233163
rect 347062 233111 347114 233163
rect 501046 233111 501098 233163
rect 265750 233037 265802 233089
rect 338038 233037 338090 233089
rect 350326 233037 350378 233089
rect 507094 233037 507146 233089
rect 290806 232963 290858 233015
rect 374614 232963 374666 233015
rect 398806 232963 398858 233015
rect 557014 232963 557066 233015
rect 263926 232889 263978 232941
rect 337270 232889 337322 232941
rect 353110 232889 353162 232941
rect 513142 232889 513194 232941
rect 513238 232889 513290 232941
rect 519190 232889 519242 232941
rect 237622 232815 237674 232867
rect 284374 232815 284426 232867
rect 289942 232815 289994 232867
rect 382870 232815 382922 232867
rect 411766 232815 411818 232867
rect 265174 232741 265226 232793
rect 340246 232741 340298 232793
rect 216598 232667 216650 232719
rect 242134 232667 242186 232719
rect 266614 232667 266666 232719
rect 343222 232667 343274 232719
rect 219766 232593 219818 232645
rect 248086 232593 248138 232645
rect 268438 232593 268490 232645
rect 346294 232741 346346 232793
rect 356278 232741 356330 232793
rect 513046 232741 513098 232793
rect 572086 232815 572138 232867
rect 521206 232741 521258 232793
rect 626422 232741 626474 232793
rect 218038 232519 218090 232571
rect 245110 232519 245162 232571
rect 274870 232519 274922 232571
rect 346966 232667 347018 232719
rect 361366 232667 361418 232719
rect 362134 232667 362186 232719
rect 531286 232667 531338 232719
rect 356086 232593 356138 232645
rect 365398 232593 365450 232645
rect 537238 232593 537290 232645
rect 343894 232519 343946 232571
rect 355318 232519 355370 232571
rect 365014 232519 365066 232571
rect 539542 232519 539594 232571
rect 222550 232445 222602 232497
rect 254230 232445 254282 232497
rect 269686 232445 269738 232497
rect 349366 232445 349418 232497
rect 368182 232445 368234 232497
rect 543382 232445 543434 232497
rect 221110 232371 221162 232423
rect 251158 232371 251210 232423
rect 271222 232371 271274 232423
rect 352342 232371 352394 232423
rect 366262 232371 366314 232423
rect 542614 232371 542666 232423
rect 222934 232297 222986 232349
rect 255670 232297 255722 232349
rect 272950 232297 273002 232349
rect 343894 232297 343946 232349
rect 343990 232297 344042 232349
rect 350518 232297 350570 232349
rect 371158 232297 371210 232349
rect 549430 232297 549482 232349
rect 226294 232223 226346 232275
rect 261718 232223 261770 232275
rect 274198 232223 274250 232275
rect 358294 232223 358346 232275
rect 372694 232223 372746 232275
rect 552406 232223 552458 232275
rect 224278 232149 224330 232201
rect 257206 232149 257258 232201
rect 277462 232149 277514 232201
rect 364438 232149 364490 232201
rect 368086 232149 368138 232201
rect 545590 232149 545642 232201
rect 227062 232075 227114 232127
rect 263254 232075 263306 232127
rect 275734 232075 275786 232127
rect 346966 232075 347018 232127
rect 350518 232075 350570 232127
rect 367126 232075 367178 232127
rect 369526 232075 369578 232127
rect 548566 232075 548618 232127
rect 147670 232001 147722 232053
rect 154102 232001 154154 232053
rect 233878 232001 233930 232053
rect 274486 232001 274538 232053
rect 280246 232001 280298 232053
rect 370390 232001 370442 232053
rect 375766 232001 375818 232053
rect 558454 232001 558506 232053
rect 234838 231927 234890 231979
rect 278326 231927 278378 231979
rect 278998 231927 279050 231979
rect 367414 231927 367466 231979
rect 372310 231927 372362 231979
rect 554710 231927 554762 231979
rect 233206 231853 233258 231905
rect 275350 231853 275402 231905
rect 281974 231853 282026 231905
rect 373462 231853 373514 231905
rect 374038 231853 374090 231905
rect 557590 231853 557642 231905
rect 236086 231779 236138 231831
rect 281302 231779 281354 231831
rect 295318 231779 295370 231831
rect 400246 231779 400298 231831
rect 405046 231779 405098 231831
rect 604534 231779 604586 231831
rect 259126 231705 259178 231757
rect 328150 231705 328202 231757
rect 346966 231705 347018 231757
rect 362134 231705 362186 231757
rect 367126 231705 367178 231757
rect 495094 231705 495146 231757
rect 498550 231705 498602 231757
rect 614998 231705 615050 231757
rect 258742 231631 258794 231683
rect 326710 231631 326762 231683
rect 337558 231631 337610 231683
rect 485206 231631 485258 231683
rect 255766 231557 255818 231609
rect 320662 231557 320714 231609
rect 327094 231557 327146 231609
rect 464086 231557 464138 231609
rect 248374 231483 248426 231535
rect 305494 231483 305546 231535
rect 312214 231483 312266 231535
rect 433846 231483 433898 231535
rect 292534 231409 292586 231461
rect 379990 231409 380042 231461
rect 400438 231409 400490 231461
rect 520726 231409 520778 231461
rect 293110 231335 293162 231387
rect 371638 231335 371690 231387
rect 400342 231335 400394 231387
rect 499606 231335 499658 231387
rect 281206 231261 281258 231313
rect 289270 231261 289322 231313
rect 293494 231261 293546 231313
rect 364246 231261 364298 231313
rect 395254 231261 395306 231313
rect 485974 231261 486026 231313
rect 257590 231187 257642 231239
rect 325174 231187 325226 231239
rect 334102 231187 334154 231239
rect 416470 231187 416522 231239
rect 256150 231113 256202 231165
rect 322102 231113 322154 231165
rect 331222 231113 331274 231165
rect 395350 231113 395402 231165
rect 395734 231113 395786 231165
rect 473878 231113 473930 231165
rect 149398 231039 149450 231091
rect 159862 231039 159914 231091
rect 252982 231039 253034 231091
rect 314518 231039 314570 231091
rect 328342 231039 328394 231091
rect 368758 231039 368810 231091
rect 245206 230965 245258 231017
rect 299446 230965 299498 231017
rect 308182 230965 308234 231017
rect 323638 230965 323690 231017
rect 344662 230965 344714 231017
rect 409654 230965 409706 231017
rect 416374 230965 416426 231017
rect 424054 230965 424106 231017
rect 326806 230891 326858 230943
rect 380278 230891 380330 230943
rect 385942 230891 385994 230943
rect 449686 230891 449738 230943
rect 290710 230817 290762 230869
rect 297430 230817 297482 230869
rect 313942 230817 313994 230869
rect 346966 230817 347018 230869
rect 358390 230817 358442 230869
rect 419542 230817 419594 230869
rect 323350 230743 323402 230795
rect 377110 230743 377162 230795
rect 320758 230669 320810 230721
rect 368566 230669 368618 230721
rect 368758 230669 368810 230721
rect 401398 230669 401450 230721
rect 302326 230595 302378 230647
rect 308566 230595 308618 230647
rect 323254 230595 323306 230647
rect 329590 230595 329642 230647
rect 354262 230595 354314 230647
rect 306742 230521 306794 230573
rect 317590 230521 317642 230573
rect 321046 230521 321098 230573
rect 368182 230521 368234 230573
rect 404470 230595 404522 230647
rect 299350 230447 299402 230499
rect 302518 230447 302570 230499
rect 304150 230447 304202 230499
rect 311638 230447 311690 230499
rect 318358 230447 318410 230499
rect 365110 230447 365162 230499
rect 398902 230447 398954 230499
rect 410518 230447 410570 230499
rect 423382 230447 423434 230499
rect 436150 230447 436202 230499
rect 248950 230373 249002 230425
rect 304822 230373 304874 230425
rect 321238 230373 321290 230425
rect 451990 230373 452042 230425
rect 228886 230299 228938 230351
rect 267862 230299 267914 230351
rect 269110 230299 269162 230351
rect 322966 230299 323018 230351
rect 325750 230299 325802 230351
rect 461014 230299 461066 230351
rect 463606 230299 463658 230351
rect 478390 230299 478442 230351
rect 247030 230225 247082 230277
rect 303958 230225 304010 230277
rect 305110 230225 305162 230277
rect 326806 230225 326858 230277
rect 248758 230151 248810 230203
rect 307030 230151 307082 230203
rect 324022 230151 324074 230203
rect 458038 230225 458090 230277
rect 464566 230225 464618 230277
rect 484438 230225 484490 230277
rect 328534 230151 328586 230203
rect 467062 230151 467114 230203
rect 475222 230151 475274 230203
rect 601462 230151 601514 230203
rect 251926 230077 251978 230129
rect 310774 230077 310826 230129
rect 331606 230077 331658 230129
rect 473110 230077 473162 230129
rect 479254 230077 479306 230129
rect 609046 230077 609098 230129
rect 251542 230003 251594 230055
rect 313078 230003 313130 230055
rect 336310 230003 336362 230055
rect 482134 230003 482186 230055
rect 486646 230003 486698 230055
rect 612118 230003 612170 230055
rect 227446 229929 227498 229981
rect 264790 229929 264842 229981
rect 290902 229929 290954 229981
rect 331894 229929 331946 229981
rect 348502 229929 348554 229981
rect 504022 229929 504074 229981
rect 253078 229855 253130 229907
rect 316150 229855 316202 229907
rect 351766 229855 351818 229907
rect 510166 229855 510218 229907
rect 512182 229855 512234 229907
rect 625558 229855 625610 229907
rect 146902 229781 146954 229833
rect 151222 229781 151274 229833
rect 239734 229781 239786 229833
rect 288886 229781 288938 229833
rect 291190 229781 291242 229833
rect 382966 229781 383018 229833
rect 389110 229781 389162 229833
rect 396982 229781 397034 229833
rect 406966 229781 407018 229833
rect 565942 229781 565994 229833
rect 220150 229707 220202 229759
rect 249718 229707 249770 229759
rect 255190 229707 255242 229759
rect 316822 229707 316874 229759
rect 354838 229707 354890 229759
rect 516118 229707 516170 229759
rect 528406 229707 528458 229759
rect 605974 229707 606026 229759
rect 221590 229633 221642 229685
rect 252598 229633 252650 229685
rect 254806 229633 254858 229685
rect 319126 229633 319178 229685
rect 360886 229633 360938 229685
rect 241078 229559 241130 229611
rect 291958 229559 292010 229611
rect 298102 229559 298154 229611
rect 362806 229559 362858 229611
rect 369910 229633 369962 229685
rect 378550 229633 378602 229685
rect 378646 229633 378698 229685
rect 522166 229633 522218 229685
rect 522646 229633 522698 229685
rect 630166 229633 630218 229685
rect 528310 229559 528362 229611
rect 528502 229559 528554 229611
rect 628630 229559 628682 229611
rect 215254 229485 215306 229537
rect 239062 229485 239114 229537
rect 244246 229485 244298 229537
rect 298006 229485 298058 229537
rect 298390 229485 298442 229537
rect 406774 229485 406826 229537
rect 406870 229485 406922 229537
rect 575062 229485 575114 229537
rect 264310 229411 264362 229463
rect 334966 229411 335018 229463
rect 366646 229411 366698 229463
rect 540310 229411 540362 229463
rect 231862 229337 231914 229389
rect 272278 229337 272330 229389
rect 273526 229337 273578 229389
rect 347062 229337 347114 229389
rect 357622 229337 357674 229389
rect 378646 229337 378698 229389
rect 378742 229337 378794 229389
rect 546358 229337 546410 229389
rect 230806 229263 230858 229315
rect 270742 229263 270794 229315
rect 283510 229263 283562 229315
rect 367510 229263 367562 229315
rect 374134 229263 374186 229315
rect 555382 229263 555434 229315
rect 233494 229189 233546 229241
rect 276790 229189 276842 229241
rect 282166 229189 282218 229241
rect 371254 229189 371306 229241
rect 377206 229189 377258 229241
rect 561430 229189 561482 229241
rect 231958 229115 232010 229167
rect 273814 229115 273866 229167
rect 284758 229115 284810 229167
rect 371542 229115 371594 229167
rect 376822 229115 376874 229167
rect 563638 229115 563690 229167
rect 235222 229041 235274 229093
rect 279862 229041 279914 229093
rect 286294 229041 286346 229093
rect 374518 229041 374570 229093
rect 380470 229041 380522 229093
rect 567478 229041 567530 229093
rect 238390 228967 238442 229019
rect 283606 228967 283658 229019
rect 287926 228967 287978 229019
rect 374422 228967 374474 229019
rect 379894 228967 379946 229019
rect 569782 228967 569834 229019
rect 245782 228893 245834 228945
rect 300982 228893 301034 228945
rect 317974 228893 318026 228945
rect 445942 228893 445994 228945
rect 449302 228893 449354 228945
rect 466390 228893 466442 228945
rect 246166 228819 246218 228871
rect 298678 228819 298730 228871
rect 314902 228819 314954 228871
rect 439990 228819 440042 228871
rect 242518 228745 242570 228797
rect 294934 228745 294986 228797
rect 308950 228745 309002 228797
rect 427798 228745 427850 228797
rect 428278 228745 428330 228797
rect 547894 228745 547946 228797
rect 241654 228671 241706 228723
rect 289750 228671 289802 228723
rect 306166 228671 306218 228723
rect 230326 228597 230378 228649
rect 269302 228597 269354 228649
rect 269398 228597 269450 228649
rect 307702 228597 307754 228649
rect 309334 228671 309386 228723
rect 425590 228671 425642 228723
rect 432022 228671 432074 228723
rect 529750 228671 529802 228723
rect 421846 228597 421898 228649
rect 434902 228597 434954 228649
rect 454294 228597 454346 228649
rect 190198 228523 190250 228575
rect 192310 228523 192362 228575
rect 228790 228523 228842 228575
rect 266230 228523 266282 228575
rect 266326 228523 266378 228575
rect 301750 228523 301802 228575
rect 304438 228523 304490 228575
rect 418774 228523 418826 228575
rect 455062 228523 455114 228575
rect 456502 228523 456554 228575
rect 535798 228523 535850 228575
rect 538006 228523 538058 228575
rect 544342 228523 544394 228575
rect 547126 228523 547178 228575
rect 556150 228523 556202 228575
rect 557686 228523 557738 228575
rect 567382 228523 567434 228575
rect 569014 228523 569066 228575
rect 224374 228449 224426 228501
rect 258742 228449 258794 228501
rect 260470 228449 260522 228501
rect 286678 228449 286730 228501
rect 289366 228449 289418 228501
rect 380086 228449 380138 228501
rect 403318 228449 403370 228501
rect 517654 228449 517706 228501
rect 264886 228375 264938 228427
rect 295702 228375 295754 228427
rect 303478 228375 303530 228427
rect 413494 228375 413546 228427
rect 535798 228375 535850 228427
rect 537910 228375 537962 228427
rect 260854 228301 260906 228353
rect 292630 228301 292682 228353
rect 293878 228301 293930 228353
rect 381718 228301 381770 228353
rect 393526 228301 393578 228353
rect 476950 228301 477002 228353
rect 250582 228227 250634 228279
rect 276502 228227 276554 228279
rect 288022 228227 288074 228279
rect 328918 228227 328970 228279
rect 357718 228227 357770 228279
rect 359926 228227 359978 228279
rect 270838 228153 270890 228205
rect 313846 228153 313898 228205
rect 258070 228079 258122 228131
rect 280630 228079 280682 228131
rect 311062 228079 311114 228131
rect 392374 228153 392426 228205
rect 396406 228153 396458 228205
rect 437686 228153 437738 228205
rect 314038 228079 314090 228131
rect 383254 228079 383306 228131
rect 390358 228079 390410 228131
rect 461878 228079 461930 228131
rect 290998 228005 291050 228057
rect 341014 228005 341066 228057
rect 344182 228005 344234 228057
rect 412726 228005 412778 228057
rect 281878 227931 281930 227983
rect 325846 227931 325898 227983
rect 341398 227931 341450 227983
rect 398326 227931 398378 227983
rect 250198 227857 250250 227909
rect 310006 227857 310058 227909
rect 310102 227857 310154 227909
rect 359158 227857 359210 227909
rect 293782 227783 293834 227835
rect 343990 227783 344042 227835
rect 301270 227709 301322 227761
rect 350038 227709 350090 227761
rect 319606 227635 319658 227687
rect 149398 227561 149450 227613
rect 182902 227561 182954 227613
rect 279286 227561 279338 227613
rect 319894 227561 319946 227613
rect 326806 227635 326858 227687
rect 353110 227635 353162 227687
rect 403702 227561 403754 227613
rect 418294 227561 418346 227613
rect 433174 227561 433226 227613
rect 187126 227487 187178 227539
rect 190774 227487 190826 227539
rect 213814 227487 213866 227539
rect 237526 227487 237578 227539
rect 249334 227487 249386 227539
rect 306262 227487 306314 227539
rect 311350 227487 311402 227539
rect 375766 227487 375818 227539
rect 390070 227487 390122 227539
rect 588598 227487 588650 227539
rect 596182 227487 596234 227539
rect 616630 227487 616682 227539
rect 629302 227487 629354 227539
rect 634006 227487 634058 227539
rect 216118 227413 216170 227465
rect 239830 227413 239882 227465
rect 253846 227413 253898 227465
rect 315382 227413 315434 227465
rect 318262 227413 318314 227465
rect 381814 227413 381866 227465
rect 390838 227413 390890 227465
rect 590134 227413 590186 227465
rect 593014 227413 593066 227465
rect 611254 227413 611306 227465
rect 215734 227339 215786 227391
rect 238390 227339 238442 227391
rect 284662 227339 284714 227391
rect 306646 227339 306698 227391
rect 311254 227339 311306 227391
rect 384022 227339 384074 227391
rect 388246 227339 388298 227391
rect 585622 227339 585674 227391
rect 595894 227339 595946 227391
rect 614326 227339 614378 227391
rect 274678 227265 274730 227317
rect 348598 227265 348650 227317
rect 392278 227265 392330 227317
rect 593110 227265 593162 227317
rect 597430 227265 597482 227317
rect 619606 227265 619658 227317
rect 220342 227191 220394 227243
rect 247414 227191 247466 227243
rect 247702 227191 247754 227243
rect 257974 227191 258026 227243
rect 271990 227191 272042 227243
rect 351574 227191 351626 227243
rect 603478 227191 603530 227243
rect 636214 227191 636266 227243
rect 219478 227117 219530 227169
rect 245878 227117 245930 227169
rect 263734 227117 263786 227169
rect 288118 227117 288170 227169
rect 289270 227117 289322 227169
rect 369622 227117 369674 227169
rect 388150 227117 388202 227169
rect 584854 227117 584906 227169
rect 606358 227117 606410 227169
rect 638518 227117 638570 227169
rect 238774 227043 238826 227095
rect 254902 227043 254954 227095
rect 259030 227043 259082 227095
rect 269974 227043 270026 227095
rect 275254 227043 275306 227095
rect 357622 227043 357674 227095
rect 392662 227043 392714 227095
rect 593974 227043 594026 227095
rect 599062 227043 599114 227095
rect 633142 227043 633194 227095
rect 212374 226969 212426 227021
rect 234550 226969 234602 227021
rect 236374 226969 236426 227021
rect 264022 226969 264074 227021
rect 276694 226969 276746 227021
rect 360598 226969 360650 227021
rect 391222 226969 391274 227021
rect 590902 226969 590954 227021
rect 221686 226895 221738 226947
rect 250390 226895 250442 226947
rect 253558 226895 253610 226947
rect 266998 226895 267050 226947
rect 273430 226895 273482 226947
rect 354550 226895 354602 226947
rect 359830 226895 359882 226947
rect 393142 226895 393194 226947
rect 395542 226895 395594 226947
rect 224854 226821 224906 226873
rect 256438 226821 256490 226873
rect 277942 226821 277994 226873
rect 363766 226821 363818 226873
rect 364246 226821 364298 226873
rect 396118 226821 396170 226873
rect 397654 226895 397706 226947
rect 603670 226969 603722 227021
rect 606262 226969 606314 227021
rect 639190 226969 639242 227021
rect 603382 226895 603434 226947
rect 636886 226895 636938 226947
rect 599158 226821 599210 226873
rect 600406 226821 600458 226873
rect 634678 226821 634730 226873
rect 223318 226747 223370 226799
rect 253462 226747 253514 226799
rect 279766 226747 279818 226799
rect 366742 226747 366794 226799
rect 374614 226747 374666 226799
rect 391510 226747 391562 226799
rect 397174 226747 397226 226799
rect 602998 226747 603050 226799
rect 603286 226747 603338 226799
rect 637750 226747 637802 226799
rect 226582 226673 226634 226725
rect 259414 226673 259466 226725
rect 271894 226673 271946 226725
rect 336406 226673 336458 226725
rect 371638 226673 371690 226725
rect 393814 226673 393866 226725
rect 400822 226673 400874 226725
rect 609814 226673 609866 226725
rect 227926 226599 227978 226651
rect 262486 226599 262538 226651
rect 264694 226599 264746 226651
rect 276118 226599 276170 226651
rect 285718 226599 285770 226651
rect 378742 226599 378794 226651
rect 381718 226599 381770 226651
rect 397654 226599 397706 226651
rect 588886 226599 588938 226651
rect 600790 226599 600842 226651
rect 606166 226599 606218 226651
rect 639958 226599 640010 226651
rect 231094 226525 231146 226577
rect 268534 226525 268586 226577
rect 270934 226525 270986 226577
rect 294262 226525 294314 226577
rect 297430 226525 297482 226577
rect 390070 226525 390122 226577
rect 402166 226525 402218 226577
rect 612790 226525 612842 226577
rect 229558 226451 229610 226503
rect 265558 226451 265610 226503
rect 288502 226451 288554 226503
rect 384790 226451 384842 226503
rect 385750 226451 385802 226503
rect 392086 226451 392138 226503
rect 404374 226451 404426 226503
rect 617302 226451 617354 226503
rect 232534 226377 232586 226429
rect 271606 226377 271658 226429
rect 291574 226377 291626 226429
rect 214582 226303 214634 226355
rect 236854 226303 236906 226355
rect 241750 226303 241802 226355
rect 217846 226229 217898 226281
rect 242902 226229 242954 226281
rect 215638 226155 215690 226207
rect 240598 226155 240650 226207
rect 246550 226155 246602 226207
rect 254902 226303 254954 226355
rect 285142 226303 285194 226355
rect 306646 226377 306698 226429
rect 378070 226377 378122 226429
rect 379990 226377 380042 226429
rect 394582 226377 394634 226429
rect 402646 226377 402698 226429
rect 613558 226377 613610 226429
rect 629206 226377 629258 226429
rect 635446 226377 635498 226429
rect 390838 226303 390890 226355
rect 404950 226303 405002 226355
rect 618070 226303 618122 226355
rect 254998 226229 255050 226281
rect 297238 226229 297290 226281
rect 297622 226229 297674 226281
rect 402838 226229 402890 226281
rect 407734 226229 407786 226281
rect 624118 226229 624170 226281
rect 151126 226081 151178 226133
rect 187126 226081 187178 226133
rect 218326 226081 218378 226133
rect 246646 226081 246698 226133
rect 291190 226155 291242 226207
rect 300694 226155 300746 226207
rect 408982 226155 409034 226207
rect 300214 226081 300266 226133
rect 301366 226081 301418 226133
rect 411286 226081 411338 226133
rect 411382 226081 411434 226133
rect 631702 226081 631754 226133
rect 213046 226007 213098 226059
rect 233782 226007 233834 226059
rect 238966 226007 239018 226059
rect 217462 225933 217514 225985
rect 241270 225933 241322 225985
rect 244822 226007 244874 226059
rect 254998 226007 255050 226059
rect 257110 226007 257162 226059
rect 261046 225933 261098 225985
rect 324502 226007 324554 226059
rect 339478 226007 339530 226059
rect 321334 225933 321386 225985
rect 334294 225933 334346 225985
rect 345718 225933 345770 225985
rect 386998 225933 387050 225985
rect 387286 226007 387338 226059
rect 582646 226007 582698 226059
rect 591478 226007 591530 226059
rect 608278 226007 608330 226059
rect 387766 225933 387818 225985
rect 388054 225933 388106 225985
rect 584086 225933 584138 225985
rect 590422 225933 590474 225985
rect 218806 225859 218858 225911
rect 244342 225859 244394 225911
rect 244726 225859 244778 225911
rect 254902 225859 254954 225911
rect 269014 225859 269066 225911
rect 330454 225859 330506 225911
rect 331414 225859 331466 225911
rect 345526 225859 345578 225911
rect 365686 225859 365738 225911
rect 382678 225859 382730 225911
rect 382966 225859 383018 225911
rect 388726 225859 388778 225911
rect 389494 225859 389546 225911
rect 587158 225859 587210 225911
rect 588694 225859 588746 225911
rect 598486 225859 598538 225911
rect 605302 225859 605354 225911
rect 217078 225785 217130 225837
rect 243574 225785 243626 225837
rect 267766 225785 267818 225837
rect 327382 225785 327434 225837
rect 368566 225785 368618 225837
rect 374230 225785 374282 225837
rect 374422 225785 374474 225837
rect 385558 225785 385610 225837
rect 386614 225785 386666 225837
rect 285046 225711 285098 225763
rect 342550 225711 342602 225763
rect 371350 225711 371402 225763
rect 376438 225711 376490 225763
rect 380086 225711 380138 225763
rect 388630 225711 388682 225763
rect 388726 225711 388778 225763
rect 389302 225711 389354 225763
rect 392086 225785 392138 225837
rect 579574 225785 579626 225837
rect 581110 225711 581162 225763
rect 588982 225711 589034 225763
rect 602230 225711 602282 225763
rect 278230 225637 278282 225689
rect 324406 225637 324458 225689
rect 339094 225637 339146 225689
rect 396886 225637 396938 225689
rect 396982 225637 397034 225689
rect 586390 225637 586442 225689
rect 273622 225563 273674 225615
rect 309334 225563 309386 225615
rect 315766 225563 315818 225615
rect 439126 225563 439178 225615
rect 265270 225489 265322 225541
rect 279094 225489 279146 225541
rect 243958 225415 244010 225467
rect 251926 225415 251978 225467
rect 262006 225415 262058 225467
rect 273046 225415 273098 225467
rect 273718 225415 273770 225467
rect 303190 225489 303242 225541
rect 309910 225489 309962 225541
rect 427030 225489 427082 225541
rect 306742 225415 306794 225467
rect 420982 225415 421034 225467
rect 241846 225341 241898 225393
rect 248854 225341 248906 225393
rect 303862 225341 303914 225393
rect 415030 225341 415082 225393
rect 302134 225267 302186 225319
rect 411958 225267 412010 225319
rect 277078 225193 277130 225245
rect 318358 225193 318410 225245
rect 339766 225193 339818 225245
rect 399958 225193 400010 225245
rect 400150 225193 400202 225245
rect 606742 225193 606794 225245
rect 305014 225119 305066 225171
rect 333526 225119 333578 225171
rect 349750 225119 349802 225171
rect 405910 225119 405962 225171
rect 410422 225119 410474 225171
rect 629398 225119 629450 225171
rect 252694 225045 252746 225097
rect 312310 225045 312362 225097
rect 367510 225045 367562 225097
rect 371350 225045 371402 225097
rect 371446 225045 371498 225097
rect 372694 225045 372746 225097
rect 374518 225045 374570 225097
rect 382582 225045 382634 225097
rect 382678 225045 382730 225097
rect 418006 225045 418058 225097
rect 354358 224971 354410 225023
rect 408214 224971 408266 225023
rect 348694 224897 348746 224949
rect 399094 224897 399146 224949
rect 149302 224823 149354 224875
rect 165622 224823 165674 224875
rect 362806 224823 362858 224875
rect 405142 224823 405194 224875
rect 149398 224749 149450 224801
rect 171286 224749 171338 224801
rect 361942 224749 361994 224801
rect 402166 224749 402218 224801
rect 149494 224675 149546 224727
rect 174262 224675 174314 224727
rect 267958 224675 268010 224727
rect 282070 224675 282122 224727
rect 282550 224675 282602 224727
rect 371446 224675 371498 224727
rect 371542 224675 371594 224727
rect 379510 224675 379562 224727
rect 382870 224675 382922 224727
rect 386326 224675 386378 224727
rect 390454 224675 390506 224727
rect 589366 224675 589418 224727
rect 323158 224601 323210 224653
rect 452758 224601 452810 224653
rect 319414 224527 319466 224579
rect 447478 224527 447530 224579
rect 322294 224453 322346 224505
rect 453430 224453 453482 224505
rect 325078 224379 325130 224431
rect 459574 224379 459626 224431
rect 328246 224305 328298 224357
rect 465622 224305 465674 224357
rect 331510 224231 331562 224283
rect 471574 224231 471626 224283
rect 276502 224157 276554 224209
rect 277558 224157 277610 224209
rect 338134 224157 338186 224209
rect 482902 224157 482954 224209
rect 334486 224083 334538 224135
rect 477622 224083 477674 224135
rect 337174 224009 337226 224061
rect 483766 224009 483818 224061
rect 340438 223935 340490 223987
rect 489718 223935 489770 223987
rect 343606 223861 343658 223913
rect 497302 223861 497354 223913
rect 263542 223787 263594 223839
rect 335734 223787 335786 223839
rect 346582 223787 346634 223839
rect 501814 223787 501866 223839
rect 261910 223713 261962 223765
rect 332662 223713 332714 223765
rect 348022 223713 348074 223765
rect 504790 223713 504842 223765
rect 266518 223639 266570 223691
rect 341782 223639 341834 223691
rect 349558 223639 349610 223691
rect 507862 223639 507914 223691
rect 268054 223565 268106 223617
rect 344854 223565 344906 223617
rect 350806 223565 350858 223617
rect 510838 223565 510890 223617
rect 264598 223491 264650 223543
rect 338710 223491 338762 223543
rect 348118 223491 348170 223543
rect 506326 223491 506378 223543
rect 269494 223417 269546 223469
rect 347734 223417 347786 223469
rect 351190 223417 351242 223469
rect 512374 223417 512426 223469
rect 271126 223343 271178 223395
rect 350806 223343 350858 223395
rect 352534 223343 352586 223395
rect 513910 223343 513962 223395
rect 354070 223269 354122 223321
rect 516982 223269 517034 223321
rect 272566 223195 272618 223247
rect 353878 223195 353930 223247
rect 355606 223195 355658 223247
rect 519862 223195 519914 223247
rect 286198 223121 286250 223173
rect 381046 223121 381098 223173
rect 394870 223121 394922 223173
rect 523798 223121 523850 223173
rect 316342 223047 316394 223099
rect 441430 223047 441482 223099
rect 318550 222973 318602 223025
rect 443734 222973 443786 223025
rect 313366 222899 313418 222951
rect 435382 222899 435434 222951
rect 310294 222825 310346 222877
rect 429334 222825 429386 222877
rect 307990 222751 308042 222803
rect 422518 222751 422570 222803
rect 312598 222677 312650 222729
rect 431542 222677 431594 222729
rect 307222 222603 307274 222655
rect 423286 222603 423338 222655
rect 304246 222529 304298 222581
rect 417238 222529 417290 222581
rect 302806 222455 302858 222507
rect 414262 222455 414314 222507
rect 283126 222381 283178 222433
rect 374998 222381 375050 222433
rect 391798 222381 391850 222433
rect 496534 222381 496586 222433
rect 281590 222307 281642 222359
rect 371926 222307 371978 222359
rect 374710 222307 374762 222359
rect 467830 222307 467882 222359
rect 274102 222233 274154 222285
rect 356854 222233 356906 222285
rect 656182 222011 656234 222063
rect 676246 222011 676298 222063
rect 149494 221863 149546 221915
rect 162646 221863 162698 221915
rect 655990 221863 656042 221915
rect 676246 221863 676298 221915
rect 149398 221789 149450 221841
rect 168406 221789 168458 221841
rect 42070 221715 42122 221767
rect 50326 221715 50378 221767
rect 159958 221715 160010 221767
rect 184342 221715 184394 221767
rect 195766 221715 195818 221767
rect 197542 221715 197594 221767
rect 512758 221715 512810 221767
rect 515398 221715 515450 221767
rect 673462 219865 673514 219917
rect 676246 219865 676298 219917
rect 147670 219051 147722 219103
rect 174358 219051 174410 219103
rect 655798 219051 655850 219103
rect 676054 219051 676106 219103
rect 149398 218977 149450 219029
rect 177142 218977 177194 219029
rect 149494 218903 149546 218955
rect 179926 218903 179978 218955
rect 143062 218829 143114 218881
rect 184342 218829 184394 218881
rect 673366 218755 673418 218807
rect 676054 218755 676106 218807
rect 147286 217719 147338 217771
rect 151798 217719 151850 217771
rect 149398 216387 149450 216439
rect 159958 216387 160010 216439
rect 41782 213649 41834 213701
rect 45334 213649 45386 213701
rect 147574 213279 147626 213331
rect 151702 213279 151754 213331
rect 674806 213205 674858 213257
rect 676054 213205 676106 213257
rect 41782 213131 41834 213183
rect 45622 213131 45674 213183
rect 147382 213131 147434 213183
rect 151510 213131 151562 213183
rect 675094 213131 675146 213183
rect 676246 213131 676298 213183
rect 146902 212835 146954 212887
rect 152086 212835 152138 212887
rect 180118 212835 180170 212887
rect 187030 212835 187082 212887
rect 41590 212761 41642 212813
rect 45526 212761 45578 212813
rect 41782 212169 41834 212221
rect 43414 212169 43466 212221
rect 674614 211873 674666 211925
rect 676054 211873 676106 211925
rect 41782 211651 41834 211703
rect 44854 211651 44906 211703
rect 41590 211281 41642 211333
rect 50614 211281 50666 211333
rect 41782 210689 41834 210741
rect 43318 210689 43370 210741
rect 147382 210467 147434 210519
rect 151606 210467 151658 210519
rect 674710 210393 674762 210445
rect 675958 210393 676010 210445
rect 147382 210319 147434 210371
rect 151414 210319 151466 210371
rect 674902 210319 674954 210371
rect 676054 210319 676106 210371
rect 674998 210245 675050 210297
rect 676246 210245 676298 210297
rect 41782 210097 41834 210149
rect 50422 210097 50474 210149
rect 41590 209801 41642 209853
rect 43510 209801 43562 209853
rect 146902 208321 146954 208373
rect 151990 208321 152042 208373
rect 146998 207359 147050 207411
rect 151318 207359 151370 207411
rect 646774 207359 646826 207411
rect 679990 207359 680042 207411
rect 147094 206249 147146 206301
rect 151894 206249 151946 206301
rect 675766 206101 675818 206153
rect 675094 205657 675146 205709
rect 675478 205657 675530 205709
rect 675766 205583 675818 205635
rect 149398 204547 149450 204599
rect 157078 204547 157130 204599
rect 147670 204029 147722 204081
rect 154198 204029 154250 204081
rect 41782 203289 41834 203341
rect 43030 203289 43082 203341
rect 41782 202771 41834 202823
rect 42934 202771 42986 202823
rect 41974 202105 42026 202157
rect 44662 202105 44714 202157
rect 675190 201883 675242 201935
rect 675478 201883 675530 201935
rect 41974 201661 42026 201713
rect 44758 201661 44810 201713
rect 149494 201661 149546 201713
rect 180118 201661 180170 201713
rect 41782 201587 41834 201639
rect 42742 201587 42794 201639
rect 149398 201587 149450 201639
rect 182998 201587 183050 201639
rect 143062 201513 143114 201565
rect 184342 201513 184394 201565
rect 655606 201513 655658 201565
rect 675094 201513 675146 201565
rect 674806 201291 674858 201343
rect 675382 201291 675434 201343
rect 41782 201217 41834 201269
rect 44566 201217 44618 201269
rect 674998 200847 675050 200899
rect 675382 200847 675434 200899
rect 41590 198849 41642 198901
rect 42838 198849 42890 198901
rect 147478 198775 147530 198827
rect 152182 198775 152234 198827
rect 149398 198701 149450 198753
rect 165718 198701 165770 198753
rect 181366 198627 181418 198679
rect 184438 198627 184490 198679
rect 178294 198553 178346 198605
rect 184342 198553 184394 198605
rect 674902 197739 674954 197791
rect 675382 197739 675434 197791
rect 41878 197369 41930 197421
rect 41878 197147 41930 197199
rect 674614 196999 674666 197051
rect 675478 196999 675530 197051
rect 674710 196555 674762 196607
rect 675382 196555 675434 196607
rect 147286 195963 147338 196015
rect 168598 195963 168650 196015
rect 149398 195889 149450 195941
rect 171478 195889 171530 195941
rect 149302 195815 149354 195867
rect 177334 195815 177386 195867
rect 166966 195741 167018 195793
rect 184534 195741 184586 195793
rect 169846 195667 169898 195719
rect 184438 195667 184490 195719
rect 172726 195593 172778 195645
rect 184342 195593 184394 195645
rect 42070 193447 42122 193499
rect 42838 193447 42890 193499
rect 149398 193151 149450 193203
rect 160054 193151 160106 193203
rect 149494 193003 149546 193055
rect 162838 193003 162890 193055
rect 152374 192929 152426 192981
rect 184630 192929 184682 192981
rect 155446 192855 155498 192907
rect 184534 192855 184586 192907
rect 158134 192781 158186 192833
rect 184342 192781 184394 192833
rect 163894 192707 163946 192759
rect 184438 192707 184490 192759
rect 42166 192189 42218 192241
rect 42742 192189 42794 192241
rect 42070 191449 42122 191501
rect 43030 191449 43082 191501
rect 149398 191079 149450 191131
rect 157174 191079 157226 191131
rect 42166 191005 42218 191057
rect 42934 191005 42986 191057
rect 147286 190117 147338 190169
rect 154294 190117 154346 190169
rect 143926 190043 143978 190095
rect 184534 190043 184586 190095
rect 149686 189969 149738 190021
rect 184342 189969 184394 190021
rect 171382 189895 171434 189947
rect 184438 189895 184490 189947
rect 180022 189821 180074 189873
rect 184342 189821 184394 189873
rect 162742 187157 162794 187209
rect 184438 187157 184490 187209
rect 168502 187083 168554 187135
rect 184342 187083 184394 187135
rect 174454 187009 174506 187061
rect 184534 187009 184586 187061
rect 177238 186935 177290 186987
rect 184630 186935 184682 186987
rect 149398 185751 149450 185803
rect 186070 185751 186122 185803
rect 145558 184271 145610 184323
rect 184342 184271 184394 184323
rect 156982 184197 157034 184249
rect 184438 184197 184490 184249
rect 177046 184123 177098 184175
rect 184534 184123 184586 184175
rect 645142 183087 645194 183139
rect 649366 183087 649418 183139
rect 149302 182939 149354 182991
rect 185974 182939 186026 182991
rect 149590 182865 149642 182917
rect 186166 182865 186218 182917
rect 42166 182199 42218 182251
rect 48118 182199 48170 182251
rect 149398 181533 149450 181585
rect 165814 181533 165866 181585
rect 149494 181459 149546 181511
rect 174454 181459 174506 181511
rect 154006 181385 154058 181437
rect 184630 181385 184682 181437
rect 156886 181311 156938 181363
rect 184342 181311 184394 181363
rect 159766 181237 159818 181289
rect 184438 181237 184490 181289
rect 174166 181163 174218 181215
rect 184534 181163 184586 181215
rect 149206 179979 149258 180031
rect 185494 179979 185546 180031
rect 645142 179387 645194 179439
rect 649462 179387 649514 179439
rect 149494 178721 149546 178773
rect 162742 178721 162794 178773
rect 149398 178647 149450 178699
rect 171382 178647 171434 178699
rect 149302 178573 149354 178625
rect 183094 178573 183146 178625
rect 145462 178499 145514 178551
rect 184438 178499 184490 178551
rect 165526 178425 165578 178477
rect 184342 178425 184394 178477
rect 182806 178351 182858 178403
rect 186742 178351 186794 178403
rect 655702 176131 655754 176183
rect 676150 176131 676202 176183
rect 655510 175983 655562 176035
rect 676246 175983 676298 176035
rect 655414 175835 655466 175887
rect 676342 175835 676394 175887
rect 149398 175761 149450 175813
rect 156886 175761 156938 175813
rect 149494 175687 149546 175739
rect 168502 175687 168554 175739
rect 143062 175613 143114 175665
rect 184438 175613 184490 175665
rect 145366 175539 145418 175591
rect 184342 175539 184394 175591
rect 147670 175021 147722 175073
rect 154006 175021 154058 175073
rect 645142 174873 645194 174925
rect 649558 174873 649610 174925
rect 149206 174207 149258 174259
rect 186262 174207 186314 174259
rect 148918 174059 148970 174111
rect 149398 174059 149450 174111
rect 148534 172727 148586 172779
rect 184534 172727 184586 172779
rect 148726 172653 148778 172705
rect 184630 172653 184682 172705
rect 148342 172579 148394 172631
rect 184342 172579 184394 172631
rect 149014 172505 149066 172557
rect 184438 172505 184490 172557
rect 645142 171025 645194 171077
rect 649654 171025 649706 171077
rect 674806 170285 674858 170337
rect 676054 170285 676106 170337
rect 675286 169915 675338 169967
rect 676054 169915 676106 169967
rect 148630 169841 148682 169893
rect 184630 169841 184682 169893
rect 148822 169767 148874 169819
rect 184438 169767 184490 169819
rect 148246 169693 148298 169745
rect 184342 169693 184394 169745
rect 149302 169619 149354 169671
rect 184534 169619 184586 169671
rect 645142 168213 645194 168265
rect 649846 168213 649898 168265
rect 674902 167695 674954 167747
rect 676054 167695 676106 167747
rect 675190 167103 675242 167155
rect 676246 167103 676298 167155
rect 674998 167029 675050 167081
rect 676054 167029 676106 167081
rect 148438 166955 148490 167007
rect 184342 166955 184394 167007
rect 149398 166881 149450 166933
rect 184438 166881 184490 166933
rect 154102 166807 154154 166859
rect 184534 166807 184586 166859
rect 148726 166659 148778 166711
rect 149110 166659 149162 166711
rect 674710 166215 674762 166267
rect 676054 166215 676106 166267
rect 646870 164365 646922 164417
rect 676054 164365 676106 164417
rect 647062 164291 647114 164343
rect 676246 164291 676298 164343
rect 646966 164217 647018 164269
rect 676150 164217 676202 164269
rect 182902 164069 182954 164121
rect 185302 164069 185354 164121
rect 159862 163995 159914 164047
rect 184342 163995 184394 164047
rect 165622 163921 165674 163973
rect 184438 163921 184490 163973
rect 151222 163847 151274 163899
rect 184342 163847 184394 163899
rect 645142 163329 645194 163381
rect 649942 163329 649994 163381
rect 162646 161183 162698 161235
rect 184534 161183 184586 161235
rect 168406 161109 168458 161161
rect 184630 161109 184682 161161
rect 675670 161109 675722 161161
rect 171286 161035 171338 161087
rect 184342 161035 184394 161087
rect 174262 160961 174314 161013
rect 184438 160961 184490 161013
rect 675670 160591 675722 160643
rect 670390 160443 670442 160495
rect 675382 160443 675434 160495
rect 645142 159703 645194 159755
rect 650038 159703 650090 159755
rect 146902 159111 146954 159163
rect 151222 159111 151274 159163
rect 151798 158371 151850 158423
rect 184438 158371 184490 158423
rect 174358 158297 174410 158349
rect 184342 158297 184394 158349
rect 179926 158223 179978 158275
rect 184534 158223 184586 158275
rect 177142 158149 177194 158201
rect 184630 158149 184682 158201
rect 674806 157705 674858 157757
rect 675382 157705 675434 157757
rect 674902 157039 674954 157091
rect 675478 157039 675530 157091
rect 675190 156521 675242 156573
rect 675382 156521 675434 156573
rect 645142 156003 645194 156055
rect 650134 156003 650186 156055
rect 674998 155855 675050 155907
rect 675382 155855 675434 155907
rect 149302 155707 149354 155759
rect 174550 155707 174602 155759
rect 148822 155633 148874 155685
rect 180022 155633 180074 155685
rect 148918 155559 148970 155611
rect 149302 155559 149354 155611
rect 149686 155559 149738 155611
rect 182806 155559 182858 155611
rect 151702 155485 151754 155537
rect 184534 155485 184586 155537
rect 658006 155485 658058 155537
rect 670390 155485 670442 155537
rect 151510 155411 151562 155463
rect 184438 155411 184490 155463
rect 152086 155337 152138 155389
rect 184630 155337 184682 155389
rect 159958 155263 160010 155315
rect 184342 155263 184394 155315
rect 149206 152747 149258 152799
rect 177046 152747 177098 152799
rect 149686 152673 149738 152725
rect 177142 152673 177194 152725
rect 151414 152599 151466 152651
rect 184534 152599 184586 152651
rect 151606 152525 151658 152577
rect 184342 152525 184394 152577
rect 645142 152525 645194 152577
rect 650230 152525 650282 152577
rect 151990 152451 152042 152503
rect 184438 152451 184490 152503
rect 149206 151785 149258 151837
rect 159958 151785 160010 151837
rect 674710 151415 674762 151467
rect 675382 151415 675434 151467
rect 149206 149861 149258 149913
rect 174166 149861 174218 149913
rect 149686 149787 149738 149839
rect 179926 149787 179978 149839
rect 151318 149713 151370 149765
rect 184342 149713 184394 149765
rect 151894 149639 151946 149691
rect 184438 149639 184490 149691
rect 154198 149565 154250 149617
rect 184534 149565 184586 149617
rect 157078 149491 157130 149543
rect 184342 149491 184394 149543
rect 645142 148159 645194 148211
rect 650326 148159 650378 148211
rect 149206 146975 149258 147027
rect 168406 146975 168458 147027
rect 149686 146901 149738 146953
rect 171574 146901 171626 146953
rect 182998 146827 183050 146879
rect 186742 146827 186794 146879
rect 165718 146753 165770 146805
rect 184342 146753 184394 146805
rect 180118 146679 180170 146731
rect 185398 146679 185450 146731
rect 152182 146605 152234 146657
rect 184438 146605 184490 146657
rect 148630 145495 148682 145547
rect 147862 145421 147914 145473
rect 148342 145421 148394 145473
rect 148342 145273 148394 145325
rect 149206 144089 149258 144141
rect 162934 144089 162986 144141
rect 149686 144015 149738 144067
rect 165622 144015 165674 144067
rect 162838 143941 162890 143993
rect 184534 143941 184586 143993
rect 168598 143867 168650 143919
rect 184438 143867 184490 143919
rect 171478 143793 171530 143845
rect 184342 143793 184394 143845
rect 177334 143719 177386 143771
rect 184630 143719 184682 143771
rect 149686 142313 149738 142365
rect 159862 142313 159914 142365
rect 149206 142239 149258 142291
rect 156982 142239 157034 142291
rect 148822 141203 148874 141255
rect 154102 141203 154154 141255
rect 154294 141055 154346 141107
rect 184534 141055 184586 141107
rect 157174 140981 157226 141033
rect 184438 140981 184490 141033
rect 160054 140907 160106 140959
rect 184342 140907 184394 140959
rect 147094 140167 147146 140219
rect 151126 140167 151178 140219
rect 149206 138243 149258 138295
rect 165526 138243 165578 138295
rect 149206 135431 149258 135483
rect 159766 135431 159818 135483
rect 149686 135357 149738 135409
rect 162646 135357 162698 135409
rect 162742 135283 162794 135335
rect 184534 135283 184586 135335
rect 165814 135209 165866 135261
rect 184438 135209 184490 135261
rect 149494 135135 149546 135187
rect 149686 135135 149738 135187
rect 174454 135135 174506 135187
rect 184342 135135 184394 135187
rect 174550 133951 174602 134003
rect 185686 133951 185738 134003
rect 159958 133877 160010 133929
rect 185590 133877 185642 133929
rect 149398 132545 149450 132597
rect 171286 132545 171338 132597
rect 149494 132471 149546 132523
rect 174262 132471 174314 132523
rect 183094 132397 183146 132449
rect 184630 132397 184682 132449
rect 168502 132323 168554 132375
rect 184534 132323 184586 132375
rect 171382 132249 171434 132301
rect 184342 132249 184394 132301
rect 156886 132175 156938 132227
rect 184438 132175 184490 132227
rect 147190 130251 147242 130303
rect 151126 130251 151178 130303
rect 655318 130103 655370 130155
rect 676150 130103 676202 130155
rect 655222 129955 655274 130007
rect 676246 129955 676298 130007
rect 655126 129807 655178 129859
rect 676342 129807 676394 129859
rect 645718 129585 645770 129637
rect 676246 129585 676298 129637
rect 149302 129511 149354 129563
rect 184630 129511 184682 129563
rect 149206 129437 149258 129489
rect 184438 129437 184490 129489
rect 148246 129363 148298 129415
rect 148438 129363 148490 129415
rect 149590 129363 149642 129415
rect 184534 129363 184586 129415
rect 154006 129289 154058 129341
rect 184342 129289 184394 129341
rect 646486 126847 646538 126899
rect 676246 126847 676298 126899
rect 646582 126773 646634 126825
rect 676150 126773 676202 126825
rect 674134 126699 674186 126751
rect 676054 126699 676106 126751
rect 149014 126625 149066 126677
rect 184438 126625 184490 126677
rect 148726 126551 148778 126603
rect 184534 126551 184586 126603
rect 149686 126477 149738 126529
rect 184342 126477 184394 126529
rect 674230 124627 674282 124679
rect 676054 124627 676106 124679
rect 674038 124035 674090 124087
rect 675958 124035 676010 124087
rect 674614 123961 674666 124013
rect 676054 123961 676106 124013
rect 675190 123887 675242 123939
rect 676246 123887 676298 123939
rect 148630 123813 148682 123865
rect 184342 123813 184394 123865
rect 148438 123739 148490 123791
rect 184438 123739 184490 123791
rect 147862 123665 147914 123717
rect 184342 123665 184394 123717
rect 148342 123591 148394 123643
rect 184534 123591 184586 123643
rect 179926 123517 179978 123569
rect 186166 123517 186218 123569
rect 674422 122111 674474 122163
rect 676054 122111 676106 122163
rect 674710 121149 674762 121201
rect 676054 121149 676106 121201
rect 674326 121075 674378 121127
rect 676246 121075 676298 121127
rect 674806 121001 674858 121053
rect 676054 121001 676106 121053
rect 147958 120927 148010 120979
rect 184438 120927 184490 120979
rect 148246 120853 148298 120905
rect 184534 120853 184586 120905
rect 171574 120779 171626 120831
rect 184630 120779 184682 120831
rect 174166 120705 174218 120757
rect 184342 120705 184394 120757
rect 647830 118337 647882 118389
rect 676246 118337 676298 118389
rect 149398 118263 149450 118315
rect 168502 118263 168554 118315
rect 149494 118189 149546 118241
rect 174358 118189 174410 118241
rect 647926 118189 647978 118241
rect 676150 118189 676202 118241
rect 149398 118115 149450 118167
rect 182902 118115 182954 118167
rect 645238 118115 645290 118167
rect 676054 118115 676106 118167
rect 159862 118041 159914 118093
rect 184630 118041 184682 118093
rect 162934 117967 162986 118019
rect 184534 117967 184586 118019
rect 165622 117893 165674 117945
rect 184438 117893 184490 117945
rect 168406 117819 168458 117871
rect 184342 117819 184394 117871
rect 675094 115377 675146 115429
rect 675286 115377 675338 115429
rect 149398 115303 149450 115355
rect 165718 115303 165770 115355
rect 149494 115229 149546 115281
rect 179926 115229 179978 115281
rect 647926 115229 647978 115281
rect 665302 115229 665354 115281
rect 151222 115155 151274 115207
rect 184534 115155 184586 115207
rect 663766 115155 663818 115207
rect 665206 115155 665258 115207
rect 154102 115081 154154 115133
rect 184438 115081 184490 115133
rect 156982 115007 157034 115059
rect 184342 115007 184394 115059
rect 674614 114785 674666 114837
rect 675190 114785 675242 114837
rect 674134 114119 674186 114171
rect 675382 114119 675434 114171
rect 148726 113675 148778 113727
rect 149014 113675 149066 113727
rect 149014 113527 149066 113579
rect 149206 113527 149258 113579
rect 149398 112861 149450 112913
rect 159862 112861 159914 112913
rect 674230 112491 674282 112543
rect 675382 112491 675434 112543
rect 149494 112343 149546 112395
rect 162742 112343 162794 112395
rect 182806 112269 182858 112321
rect 184342 112269 184394 112321
rect 665206 112269 665258 112321
rect 675094 112269 675146 112321
rect 180022 112195 180074 112247
rect 184438 112195 184490 112247
rect 177142 112121 177194 112173
rect 184534 112121 184586 112173
rect 674038 111677 674090 111729
rect 675382 111677 675434 111729
rect 674422 111307 674474 111359
rect 675382 111307 675434 111359
rect 674710 110641 674762 110693
rect 675382 110641 675434 110693
rect 149398 109531 149450 109583
rect 156886 109531 156938 109583
rect 165526 109383 165578 109435
rect 184342 109383 184394 109435
rect 177046 109309 177098 109361
rect 184438 109309 184490 109361
rect 147670 108347 147722 108399
rect 154006 108347 154058 108399
rect 674326 107311 674378 107363
rect 675382 107311 675434 107363
rect 146998 106571 147050 106623
rect 151222 106571 151274 106623
rect 159766 106497 159818 106549
rect 184534 106497 184586 106549
rect 162646 106423 162698 106475
rect 184342 106423 184394 106475
rect 171286 106349 171338 106401
rect 184630 106349 184682 106401
rect 674806 106349 674858 106401
rect 675382 106349 675434 106401
rect 174262 106275 174314 106327
rect 184438 106275 184490 106327
rect 151126 105091 151178 105143
rect 184726 105091 184778 105143
rect 647926 103759 647978 103811
rect 661174 103759 661226 103811
rect 645718 103685 645770 103737
rect 657526 103685 657578 103737
rect 148918 103611 148970 103663
rect 184438 103611 184490 103663
rect 148822 103537 148874 103589
rect 184342 103537 184394 103589
rect 149302 103463 149354 103515
rect 184534 103463 184586 103515
rect 645142 102057 645194 102109
rect 652438 102057 652490 102109
rect 149398 100799 149450 100851
rect 168406 100799 168458 100851
rect 148150 100725 148202 100777
rect 184534 100725 184586 100777
rect 149206 100651 149258 100703
rect 184630 100651 184682 100703
rect 149110 100577 149162 100629
rect 184342 100577 184394 100629
rect 149686 100503 149738 100555
rect 184438 100503 184490 100555
rect 149398 97987 149450 98039
rect 184246 97987 184298 98039
rect 149494 97913 149546 97965
rect 186166 97913 186218 97965
rect 647926 97913 647978 97965
rect 662518 97913 662570 97965
rect 148726 97839 148778 97891
rect 184342 97839 184394 97891
rect 149014 97765 149066 97817
rect 184438 97765 184490 97817
rect 168502 97691 168554 97743
rect 184534 97691 184586 97743
rect 645430 95915 645482 95967
rect 653686 95915 653738 95967
rect 149494 95101 149546 95153
rect 165526 95101 165578 95153
rect 149398 95027 149450 95079
rect 180022 95027 180074 95079
rect 174358 94879 174410 94931
rect 184342 94879 184394 94931
rect 165718 94731 165770 94783
rect 184342 94731 184394 94783
rect 182902 94657 182954 94709
rect 186262 94657 186314 94709
rect 179926 94583 179978 94635
rect 184630 94583 184682 94635
rect 646774 92659 646826 92711
rect 663094 92659 663146 92711
rect 149398 92363 149450 92415
rect 159574 92363 159626 92415
rect 645526 92363 645578 92415
rect 661750 92363 661802 92415
rect 646486 92289 646538 92341
rect 660694 92289 660746 92341
rect 646870 92215 646922 92267
rect 659830 92215 659882 92267
rect 149494 92141 149546 92193
rect 162358 92141 162410 92193
rect 647158 92141 647210 92193
rect 658870 92141 658922 92193
rect 148438 92067 148490 92119
rect 184630 92067 184682 92119
rect 148246 91993 148298 92045
rect 184534 91993 184586 92045
rect 159862 91919 159914 91971
rect 184438 91919 184490 91971
rect 162742 91845 162794 91897
rect 184342 91845 184394 91897
rect 148534 89181 148586 89233
rect 184630 89181 184682 89233
rect 151222 89107 151274 89159
rect 184534 89107 184586 89159
rect 154006 89033 154058 89085
rect 184438 89033 184490 89085
rect 156886 88959 156938 89011
rect 184342 88959 184394 89011
rect 645910 87479 645962 87531
rect 650902 87479 650954 87531
rect 647926 87257 647978 87309
rect 658006 87257 658058 87309
rect 149494 87035 149546 87087
rect 156406 87035 156458 87087
rect 647062 87035 647114 87087
rect 663286 87035 663338 87087
rect 148726 86443 148778 86495
rect 154102 86443 154154 86495
rect 148342 86369 148394 86421
rect 184438 86369 184490 86421
rect 148630 86295 148682 86347
rect 184534 86295 184586 86347
rect 149590 86221 149642 86273
rect 184342 86221 184394 86273
rect 645910 84149 645962 84201
rect 657046 84149 657098 84201
rect 147094 83557 147146 83609
rect 151126 83557 151178 83609
rect 646774 83557 646826 83609
rect 651766 83557 651818 83609
rect 165526 83483 165578 83535
rect 184438 83483 184490 83535
rect 168406 83409 168458 83461
rect 184342 83409 184394 83461
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 647830 81781 647882 81833
rect 663382 81781 663434 81833
rect 657046 81633 657098 81685
rect 658582 81633 658634 81685
rect 647734 81559 647786 81611
rect 662422 81559 662474 81611
rect 660886 80967 660938 81019
rect 668374 80967 668426 81019
rect 647926 80745 647978 80797
rect 662518 80745 662570 80797
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 149686 80597 149738 80649
rect 184438 80597 184490 80649
rect 159574 80523 159626 80575
rect 184534 80523 184586 80575
rect 162358 80449 162410 80501
rect 184342 80449 184394 80501
rect 180022 80375 180074 80427
rect 184630 80375 184682 80427
rect 149206 77711 149258 77763
rect 184342 77711 184394 77763
rect 646966 77711 647018 77763
rect 658294 77711 658346 77763
rect 149302 77637 149354 77689
rect 184438 77637 184490 77689
rect 646582 77637 646634 77689
rect 659446 77637 659498 77689
rect 149398 77563 149450 77615
rect 184534 77563 184586 77615
rect 646678 77563 646730 77615
rect 661750 77563 661802 77615
rect 156406 77489 156458 77541
rect 184630 77489 184682 77541
rect 647926 77489 647978 77541
rect 656950 77489 657002 77541
rect 646006 76083 646058 76135
rect 657526 76083 657578 76135
rect 647062 74899 647114 74951
rect 660118 74899 660170 74951
rect 148438 74825 148490 74877
rect 184534 74825 184586 74877
rect 149110 74751 149162 74803
rect 184630 74751 184682 74803
rect 151126 74677 151178 74729
rect 184438 74677 184490 74729
rect 154102 74603 154154 74655
rect 184342 74603 184394 74655
rect 647926 72087 647978 72139
rect 660694 72087 660746 72139
rect 148246 71939 148298 71991
rect 184438 71939 184490 71991
rect 149686 71865 149738 71917
rect 184534 71865 184586 71917
rect 149590 71791 149642 71843
rect 184342 71791 184394 71843
rect 647926 69423 647978 69475
rect 661462 69423 661514 69475
rect 148822 69053 148874 69105
rect 184342 69053 184394 69105
rect 149206 68979 149258 69031
rect 184438 68979 184490 69031
rect 149590 68905 149642 68957
rect 184342 68905 184394 68957
rect 149302 68831 149354 68883
rect 184534 68831 184586 68883
rect 149110 66167 149162 66219
rect 184534 66167 184586 66219
rect 646006 66167 646058 66219
rect 652342 66167 652394 66219
rect 149398 66093 149450 66145
rect 184630 66093 184682 66145
rect 149494 66019 149546 66071
rect 184438 66019 184490 66071
rect 149014 65945 149066 65997
rect 184342 65945 184394 65997
rect 647926 63577 647978 63629
rect 663190 63577 663242 63629
rect 149398 63281 149450 63333
rect 184630 63281 184682 63333
rect 149590 63207 149642 63259
rect 184534 63207 184586 63259
rect 149206 63133 149258 63185
rect 184342 63133 184394 63185
rect 149302 63059 149354 63111
rect 184438 63059 184490 63111
rect 647926 60987 647978 61039
rect 663478 60987 663530 61039
rect 149398 60395 149450 60447
rect 184438 60395 184490 60447
rect 149494 60321 149546 60373
rect 184342 60321 184394 60373
rect 149302 60247 149354 60299
rect 184534 60247 184586 60299
rect 646006 59063 646058 59115
rect 652246 59063 652298 59115
rect 149398 58989 149450 59041
rect 184342 58989 184394 59041
rect 149398 57509 149450 57561
rect 184342 57509 184394 57561
rect 149398 56177 149450 56229
rect 184438 56177 184490 56229
rect 149494 56103 149546 56155
rect 184342 56103 184394 56155
rect 149686 54623 149738 54675
rect 184342 54623 184394 54675
rect 149398 53217 149450 53269
rect 184342 53217 184394 53269
rect 434902 48111 434954 48163
rect 475702 48111 475754 48163
rect 460342 48037 460394 48089
rect 510358 48037 510410 48089
rect 394582 47963 394634 48015
rect 406774 47963 406826 48015
rect 411862 47963 411914 48015
rect 424054 47963 424106 48015
rect 426166 47963 426218 48015
rect 492982 47963 493034 48015
rect 311062 47889 311114 47941
rect 371926 47889 371978 47941
rect 405526 47889 405578 47941
rect 441334 47889 441386 47941
rect 472246 47889 472298 47941
rect 562486 47889 562538 47941
rect 320182 47815 320234 47867
rect 529270 47815 529322 47867
rect 302902 47741 302954 47793
rect 523894 47741 523946 47793
rect 233686 47667 233738 47719
rect 475510 47667 475562 47719
rect 505366 47667 505418 47719
rect 527926 47667 527978 47719
rect 268534 47593 268586 47645
rect 517366 47593 517418 47645
rect 250966 47519 251018 47571
rect 521206 47519 521258 47571
rect 145366 47075 145418 47127
rect 199126 47075 199178 47127
rect 324310 46261 324362 46313
rect 337462 46261 337514 46313
rect 345622 46261 345674 46313
rect 354838 46261 354890 46313
rect 224566 44633 224618 44685
rect 660886 44633 660938 44685
rect 523894 43967 523946 44019
rect 525910 43967 525962 44019
rect 285814 43227 285866 43279
rect 518710 43227 518762 43279
rect 399862 42339 399914 42391
rect 411862 42339 411914 42391
rect 307222 41969 307274 42021
rect 311062 41969 311114 42021
rect 362038 41969 362090 42021
rect 365974 41969 366026 42021
rect 514006 41747 514058 41799
rect 514870 41747 514922 41799
rect 365878 37381 365930 37433
rect 399862 37381 399914 37433
rect 475510 37381 475562 37433
rect 514006 37381 514058 37433
rect 365974 37307 366026 37359
rect 389206 37307 389258 37359
<< metal2 >>
rect 82292 1002358 82348 1002367
rect 80566 1002319 80618 1002325
rect 82292 1002293 82294 1002302
rect 80566 1002261 80618 1002267
rect 82346 1002293 82348 1002302
rect 483668 1002358 483724 1002367
rect 483668 1002293 483670 1002302
rect 82294 1002261 82346 1002267
rect 483722 1002293 483724 1002302
rect 486742 1002319 486794 1002325
rect 483670 1002261 483722 1002267
rect 486742 1002261 486794 1002267
rect 80578 982979 80606 1002261
rect 132404 997770 132460 997779
rect 132404 997705 132460 997714
rect 184244 997770 184300 997779
rect 184244 997705 184300 997714
rect 132418 982979 132446 997705
rect 184258 982979 184286 997705
rect 233218 982979 233246 997742
rect 241172 997178 241228 997187
rect 241172 997113 241228 997122
rect 240886 983005 240938 983011
rect 80564 982970 80620 982979
rect 80564 982905 80620 982914
rect 132404 982970 132460 982979
rect 132404 982905 132460 982914
rect 184244 982970 184300 982979
rect 184244 982905 184300 982914
rect 233204 982970 233260 982979
rect 233204 982905 233260 982914
rect 240884 982970 240886 982979
rect 241186 982979 241214 997113
rect 241954 983011 241982 997742
rect 241942 983005 241994 983011
rect 240938 982970 240940 982979
rect 240884 982905 240940 982914
rect 241172 982970 241228 982979
rect 285058 982979 285086 997742
rect 293108 997178 293164 997187
rect 293108 997113 293164 997122
rect 292534 983005 292586 983011
rect 241942 982947 241994 982953
rect 285044 982970 285100 982979
rect 241172 982905 241228 982914
rect 285044 982905 285100 982914
rect 292532 982970 292534 982979
rect 293122 982979 293150 997113
rect 296674 983011 296702 997742
rect 388642 990781 388670 997742
rect 388630 990775 388682 990781
rect 388630 990717 388682 990723
rect 389590 990775 389642 990781
rect 389590 990717 389642 990723
rect 389602 983275 389630 990717
rect 389588 983266 389644 983275
rect 389588 983201 389644 983210
rect 296662 983005 296714 983011
rect 292586 982970 292588 982979
rect 292532 982905 292588 982914
rect 293108 982970 293164 982979
rect 394594 982979 394622 997742
rect 400340 997178 400396 997187
rect 400340 997113 400396 997122
rect 400354 982979 400382 997113
rect 486754 982979 486782 1002261
rect 535700 997770 535756 997779
rect 535700 997705 535756 997714
rect 639380 997770 639436 997779
rect 639380 997705 639436 997714
rect 535714 991521 535742 997705
rect 535702 991515 535754 991521
rect 535702 991457 535754 991463
rect 538582 991515 538634 991521
rect 538582 991457 538634 991463
rect 538594 982979 538622 991457
rect 639394 982979 639422 997705
rect 296662 982947 296714 982953
rect 394580 982970 394636 982979
rect 293108 982905 293164 982914
rect 394580 982905 394636 982914
rect 400340 982970 400396 982979
rect 400340 982905 400396 982914
rect 486740 982970 486796 982979
rect 486740 982905 486796 982914
rect 538580 982970 538636 982979
rect 538580 982905 538636 982914
rect 639380 982970 639436 982979
rect 639380 982905 639436 982914
rect 40148 961954 40204 961963
rect 40148 961889 40150 961898
rect 40202 961889 40204 961898
rect 60022 961915 60074 961921
rect 40150 961857 40202 961863
rect 60022 961857 60074 961863
rect 60034 961815 60062 961857
rect 60020 961806 60076 961815
rect 60020 961741 60076 961750
rect 653782 960509 653834 960515
rect 653780 960474 653782 960483
rect 679702 960509 679754 960515
rect 653834 960474 653836 960483
rect 679702 960451 679754 960457
rect 653780 960409 653836 960418
rect 679714 958559 679742 960451
rect 679700 958550 679756 958559
rect 679700 958485 679756 958494
rect 676148 894170 676204 894179
rect 676148 894105 676204 894114
rect 676052 893430 676108 893439
rect 676052 893365 676108 893374
rect 655414 893021 655466 893027
rect 655414 892963 655466 892969
rect 655222 892947 655274 892953
rect 655222 892889 655274 892895
rect 655126 892873 655178 892879
rect 655126 892815 655178 892821
rect 649462 881477 649514 881483
rect 649462 881419 649514 881425
rect 649474 861134 649502 881419
rect 654166 872671 654218 872677
rect 654166 872613 654218 872619
rect 653782 864013 653834 864019
rect 654178 863987 654206 872613
rect 655138 866503 655166 892815
rect 655234 867687 655262 892889
rect 655318 881403 655370 881409
rect 655318 881345 655370 881351
rect 655220 867678 655276 867687
rect 655220 867613 655276 867622
rect 655124 866494 655180 866503
rect 655124 866429 655180 866438
rect 655330 865319 655358 881345
rect 655426 868871 655454 892963
rect 676066 892879 676094 893365
rect 676162 892953 676190 894105
rect 676244 893578 676300 893587
rect 676244 893513 676300 893522
rect 676258 893027 676286 893513
rect 676246 893021 676298 893027
rect 676246 892963 676298 892969
rect 676150 892947 676202 892953
rect 676150 892889 676202 892895
rect 676054 892873 676106 892879
rect 676054 892815 676106 892821
rect 676052 892468 676108 892477
rect 673366 892429 673418 892435
rect 676052 892403 676054 892412
rect 673366 892371 673418 892377
rect 676106 892403 676108 892412
rect 676054 892371 676106 892377
rect 670966 891467 671018 891473
rect 670966 891409 671018 891415
rect 670870 890431 670922 890437
rect 670870 890373 670922 890379
rect 655412 868862 655468 868871
rect 655412 868797 655468 868806
rect 655316 865310 655372 865319
rect 655316 865245 655372 865254
rect 653782 863955 653834 863961
rect 654164 863978 654220 863987
rect 653794 862951 653822 863955
rect 654164 863913 654220 863922
rect 653780 862942 653836 862951
rect 653780 862877 653836 862886
rect 649378 861106 649502 861134
rect 41780 816692 41836 816701
rect 41780 816627 41782 816636
rect 41834 816627 41836 816636
rect 47446 816653 47498 816659
rect 41782 816595 41834 816601
rect 47446 816595 47498 816601
rect 41780 816174 41836 816183
rect 41780 816109 41782 816118
rect 41834 816109 41836 816118
rect 44854 816135 44906 816141
rect 41782 816077 41834 816083
rect 44854 816077 44906 816083
rect 41588 815434 41644 815443
rect 41588 815369 41590 815378
rect 41642 815369 41644 815378
rect 41590 815337 41642 815343
rect 41780 814694 41836 814703
rect 41780 814629 41782 814638
rect 41834 814629 41836 814638
rect 43222 814655 43274 814661
rect 41782 814597 41834 814603
rect 43222 814597 43274 814603
rect 41588 813510 41644 813519
rect 41588 813445 41590 813454
rect 41642 813445 41644 813454
rect 41590 813413 41642 813419
rect 41780 812622 41836 812631
rect 41780 812557 41782 812566
rect 41834 812557 41836 812566
rect 41782 812525 41834 812531
rect 41396 812030 41452 812039
rect 41396 811965 41452 811974
rect 40244 811290 40300 811299
rect 40244 811225 40300 811234
rect 28820 804482 28876 804491
rect 28820 804417 28876 804426
rect 28834 803899 28862 804417
rect 28820 803890 28876 803899
rect 28820 803825 28876 803834
rect 40258 801383 40286 811225
rect 40244 801374 40300 801383
rect 40244 801309 40300 801318
rect 41410 800527 41438 811965
rect 41972 811660 42028 811669
rect 41972 811595 42028 811604
rect 41588 810550 41644 810559
rect 41588 810485 41644 810494
rect 41602 810147 41630 810485
rect 41590 810141 41642 810147
rect 41590 810083 41642 810089
rect 41684 809958 41740 809967
rect 41684 809893 41740 809902
rect 41588 808478 41644 808487
rect 41588 808413 41590 808422
rect 41642 808413 41644 808422
rect 41590 808381 41642 808387
rect 41588 806998 41644 807007
rect 41588 806933 41590 806942
rect 41642 806933 41644 806942
rect 41590 806901 41642 806907
rect 41588 805518 41644 805527
rect 41588 805453 41644 805462
rect 41492 803890 41548 803899
rect 41492 803825 41548 803834
rect 41506 803783 41534 803825
rect 41494 803777 41546 803783
rect 41494 803719 41546 803725
rect 41602 803709 41630 805453
rect 41590 803703 41642 803709
rect 41590 803645 41642 803651
rect 41398 800521 41450 800527
rect 41698 800495 41726 809893
rect 41876 809662 41932 809671
rect 41876 809597 41932 809606
rect 41780 807738 41836 807747
rect 41780 807673 41836 807682
rect 41794 807261 41822 807673
rect 41782 807255 41834 807261
rect 41782 807197 41834 807203
rect 41780 806258 41836 806267
rect 41780 806193 41836 806202
rect 41794 803857 41822 806193
rect 41782 803851 41834 803857
rect 41782 803793 41834 803799
rect 41398 800463 41450 800469
rect 41684 800486 41740 800495
rect 41684 800421 41740 800430
rect 41890 800231 41918 809597
rect 41986 800347 42014 811595
rect 42742 810141 42794 810147
rect 42742 810083 42794 810089
rect 42164 808182 42220 808191
rect 42164 808117 42220 808126
rect 42068 806628 42124 806637
rect 42068 806563 42124 806572
rect 41972 800338 42028 800347
rect 41972 800273 42028 800282
rect 42082 800231 42110 806563
rect 42178 800347 42206 808117
rect 42646 806959 42698 806965
rect 42646 806901 42698 806907
rect 42164 800338 42220 800347
rect 42164 800273 42220 800282
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 42070 800225 42122 800231
rect 42070 800167 42122 800173
rect 41878 800003 41930 800009
rect 41878 799945 41930 799951
rect 41890 799422 41918 799945
rect 41972 798118 42028 798127
rect 41972 798053 42028 798062
rect 41986 797605 42014 798053
rect 42658 797937 42686 806901
rect 42754 800897 42782 810083
rect 42838 808439 42890 808445
rect 42838 808381 42890 808387
rect 42742 800891 42794 800897
rect 42742 800833 42794 800839
rect 42850 800823 42878 808381
rect 43030 807255 43082 807261
rect 43030 807197 43082 807203
rect 42934 803703 42986 803709
rect 42934 803645 42986 803651
rect 42838 800817 42890 800823
rect 42838 800759 42890 800765
rect 42742 800743 42794 800749
rect 42742 800685 42794 800691
rect 42646 797931 42698 797937
rect 42646 797873 42698 797879
rect 42754 797493 42782 800685
rect 42838 800669 42890 800675
rect 42838 800611 42890 800617
rect 42070 797487 42122 797493
rect 42070 797429 42122 797435
rect 42742 797487 42794 797493
rect 42742 797429 42794 797435
rect 42082 796980 42110 797429
rect 42742 797339 42794 797345
rect 42742 797281 42794 797287
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42178 795765 42206 796245
rect 42070 795637 42122 795643
rect 42070 795579 42122 795585
rect 42082 795130 42110 795579
rect 42166 794823 42218 794829
rect 42166 794765 42218 794771
rect 42178 794569 42206 794765
rect 42754 794311 42782 797281
rect 42850 795643 42878 800611
rect 42838 795637 42890 795643
rect 42838 795579 42890 795585
rect 42836 795454 42892 795463
rect 42836 795389 42892 795398
rect 42070 794305 42122 794311
rect 42070 794247 42122 794253
rect 42742 794305 42794 794311
rect 42742 794247 42794 794253
rect 42082 793946 42110 794247
rect 42166 793861 42218 793867
rect 42166 793803 42218 793809
rect 42178 793280 42206 793803
rect 41780 792938 41836 792947
rect 41780 792873 41836 792882
rect 41794 792729 41822 792873
rect 42262 792159 42314 792165
rect 42262 792101 42314 792107
rect 42274 790260 42302 792101
rect 42850 792014 42878 795389
rect 42946 794829 42974 803645
rect 43042 796309 43070 807197
rect 43126 803851 43178 803857
rect 43126 803793 43178 803799
rect 43030 796303 43082 796309
rect 43030 796245 43082 796251
rect 43030 796155 43082 796161
rect 43030 796097 43082 796103
rect 42934 794823 42986 794829
rect 42934 794765 42986 794771
rect 42934 794675 42986 794681
rect 42934 794617 42986 794623
rect 42192 790232 42302 790260
rect 42754 791986 42878 792014
rect 42262 790161 42314 790167
rect 42262 790103 42314 790109
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42178 788957 42206 789437
rect 42274 788410 42302 790103
rect 42754 789945 42782 791986
rect 42836 791902 42892 791911
rect 42946 791888 42974 794617
rect 43042 792165 43070 796097
rect 43138 793867 43166 803793
rect 43126 793861 43178 793867
rect 43126 793803 43178 793809
rect 43126 793713 43178 793719
rect 43126 793655 43178 793661
rect 43030 792159 43082 792165
rect 43030 792101 43082 792107
rect 42946 791860 43070 791888
rect 42836 791837 42892 791846
rect 42742 789939 42794 789945
rect 42742 789881 42794 789887
rect 42742 789199 42794 789205
rect 42742 789141 42794 789147
rect 42192 788382 42302 788410
rect 42166 786905 42218 786911
rect 42166 786847 42218 786853
rect 42178 786546 42206 786847
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42178 785921 42206 786403
rect 42070 785647 42122 785653
rect 42070 785589 42122 785595
rect 42082 785288 42110 785589
rect 42754 785209 42782 789141
rect 42850 786467 42878 791837
rect 42932 791754 42988 791763
rect 42932 791689 42988 791698
rect 42838 786461 42890 786467
rect 42838 786403 42890 786409
rect 42946 785653 42974 791689
rect 43042 789501 43070 791860
rect 43138 790167 43166 793655
rect 43126 790161 43178 790167
rect 43126 790103 43178 790109
rect 43126 790013 43178 790019
rect 43126 789955 43178 789961
rect 43030 789495 43082 789501
rect 43030 789437 43082 789443
rect 43138 786911 43166 789955
rect 43126 786905 43178 786911
rect 43126 786847 43178 786853
rect 42934 785647 42986 785653
rect 42934 785589 42986 785595
rect 42166 785203 42218 785209
rect 42166 785145 42218 785151
rect 42742 785203 42794 785209
rect 42742 785145 42794 785151
rect 42178 784725 42206 785145
rect 41588 774586 41644 774595
rect 41588 774521 41644 774530
rect 41492 773994 41548 774003
rect 41492 773929 41548 773938
rect 41506 771963 41534 773929
rect 41602 772185 41630 774521
rect 41780 773550 41836 773559
rect 41780 773485 41782 773494
rect 41834 773485 41836 773494
rect 41782 773453 41834 773459
rect 41780 772958 41836 772967
rect 41780 772893 41782 772902
rect 41834 772893 41836 772902
rect 41782 772861 41834 772867
rect 41780 772366 41836 772375
rect 41780 772301 41782 772310
rect 41834 772301 41836 772310
rect 41782 772269 41834 772275
rect 41590 772179 41642 772185
rect 41590 772121 41642 772127
rect 41494 771957 41546 771963
rect 41494 771899 41546 771905
rect 41506 769711 41534 771899
rect 41602 770747 41630 772121
rect 43234 772037 43262 814597
rect 44662 813471 44714 813477
rect 44662 813413 44714 813419
rect 44566 803777 44618 803783
rect 44566 803719 44618 803725
rect 43510 800891 43562 800897
rect 43510 800833 43562 800839
rect 43414 800817 43466 800823
rect 43414 800759 43466 800765
rect 43318 800225 43370 800231
rect 43318 800167 43370 800173
rect 43330 796161 43358 800167
rect 43318 796155 43370 796161
rect 43318 796097 43370 796103
rect 43426 794681 43454 800759
rect 43414 794675 43466 794681
rect 43414 794617 43466 794623
rect 43522 793719 43550 800833
rect 43702 800521 43754 800527
rect 43702 800463 43754 800469
rect 43510 793713 43562 793719
rect 43510 793655 43562 793661
rect 43714 790019 43742 800463
rect 43702 790013 43754 790019
rect 43702 789955 43754 789961
rect 41782 772031 41834 772037
rect 41780 771996 41782 772005
rect 43222 772031 43274 772037
rect 41834 771996 41836 772005
rect 43222 771973 43274 771979
rect 41780 771931 41836 771940
rect 41780 771478 41836 771487
rect 41780 771413 41782 771422
rect 41834 771413 41836 771422
rect 43222 771439 43274 771445
rect 41782 771381 41834 771387
rect 43222 771381 43274 771387
rect 41588 770738 41644 770747
rect 41588 770673 41644 770682
rect 41492 769702 41548 769711
rect 41492 769637 41548 769646
rect 41588 768814 41644 768823
rect 41588 768749 41644 768758
rect 38804 768074 38860 768083
rect 38804 768009 38860 768018
rect 34484 765854 34540 765863
rect 34484 765789 34540 765798
rect 28820 761266 28876 761275
rect 28820 761201 28876 761210
rect 28834 760831 28862 761201
rect 28820 760822 28876 760831
rect 28820 760757 28876 760766
rect 34498 758907 34526 765789
rect 34484 758898 34540 758907
rect 34484 758833 34540 758842
rect 38818 757575 38846 768009
rect 41602 767449 41630 768749
rect 41684 768222 41740 768231
rect 41684 768157 41740 768166
rect 41590 767443 41642 767449
rect 41590 767385 41642 767391
rect 41588 767334 41644 767343
rect 41588 767269 41644 767278
rect 40340 766594 40396 766603
rect 40340 766529 40396 766538
rect 38804 757566 38860 757575
rect 38804 757501 38860 757510
rect 40354 757385 40382 766529
rect 41602 766339 41630 767269
rect 41590 766333 41642 766339
rect 41590 766275 41642 766281
rect 41300 765114 41356 765123
rect 41300 765049 41356 765058
rect 41314 757459 41342 765049
rect 41588 761710 41644 761719
rect 41588 761645 41644 761654
rect 41602 760831 41630 761645
rect 41588 760822 41644 760831
rect 41588 760757 41590 760766
rect 41642 760757 41644 760766
rect 41590 760725 41642 760731
rect 41302 757453 41354 757459
rect 41302 757395 41354 757401
rect 41698 757385 41726 768157
rect 43030 767443 43082 767449
rect 43030 767385 43082 767391
rect 41972 766964 42028 766973
rect 41972 766899 42028 766908
rect 41780 765484 41836 765493
rect 41780 765419 41782 765428
rect 41834 765419 41836 765428
rect 41782 765387 41834 765393
rect 41876 764522 41932 764531
rect 41876 764457 41932 764466
rect 41780 763486 41836 763495
rect 41780 763421 41782 763430
rect 41834 763421 41836 763430
rect 41782 763389 41834 763395
rect 41780 762450 41836 762459
rect 41780 762385 41836 762394
rect 40342 757379 40394 757385
rect 40342 757321 40394 757327
rect 41686 757379 41738 757385
rect 41686 757321 41738 757327
rect 41794 757089 41822 762385
rect 41782 757083 41834 757089
rect 41782 757025 41834 757031
rect 41890 757015 41918 764457
rect 41986 757131 42014 766899
rect 42934 766333 42986 766339
rect 42934 766275 42986 766281
rect 42068 763930 42124 763939
rect 42068 763865 42124 763874
rect 42082 757163 42110 763865
rect 42838 763447 42890 763453
rect 42838 763389 42890 763395
rect 42164 763042 42220 763051
rect 42164 762977 42220 762986
rect 42178 757237 42206 762977
rect 42850 757700 42878 763389
rect 42946 757848 42974 766275
rect 43042 758019 43070 767385
rect 43126 765445 43178 765451
rect 43126 765387 43178 765393
rect 43028 758010 43084 758019
rect 43028 757945 43084 757954
rect 42946 757820 43070 757848
rect 42850 757672 42974 757700
rect 42838 757527 42890 757533
rect 42838 757469 42890 757475
rect 42742 757379 42794 757385
rect 42742 757321 42794 757327
rect 42166 757231 42218 757237
rect 42166 757173 42218 757179
rect 42070 757157 42122 757163
rect 41972 757122 42028 757131
rect 42070 757099 42122 757105
rect 41972 757057 42028 757066
rect 41878 757009 41930 757015
rect 41878 756951 41930 756957
rect 41782 756787 41834 756793
rect 41782 756729 41834 756735
rect 41794 756245 41822 756729
rect 42754 754943 42782 757321
rect 42070 754937 42122 754943
rect 42070 754879 42122 754885
rect 42742 754937 42794 754943
rect 42742 754879 42794 754885
rect 42082 754430 42110 754879
rect 42740 754754 42796 754763
rect 42740 754689 42796 754698
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 42178 753764 42206 754065
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42082 752580 42110 753029
rect 42166 752051 42218 752057
rect 42166 751993 42218 751999
rect 42178 751914 42206 751993
rect 42070 751829 42122 751835
rect 42070 751771 42122 751777
rect 42082 751396 42110 751771
rect 42070 751163 42122 751169
rect 42070 751105 42122 751111
rect 42082 750730 42110 751105
rect 42166 750645 42218 750651
rect 42166 750587 42218 750593
rect 42178 750064 42206 750587
rect 42754 749837 42782 754689
rect 42850 754129 42878 757469
rect 42946 757311 42974 757672
rect 43042 757385 43070 757820
rect 43030 757379 43082 757385
rect 43030 757321 43082 757327
rect 42934 757305 42986 757311
rect 43138 757279 43166 765387
rect 42934 757247 42986 757253
rect 43124 757270 43180 757279
rect 43124 757205 43180 757214
rect 43126 757157 43178 757163
rect 43126 757099 43178 757105
rect 43030 757083 43082 757089
rect 43030 757025 43082 757031
rect 42934 757009 42986 757015
rect 42934 756951 42986 756957
rect 42838 754123 42890 754129
rect 42838 754065 42890 754071
rect 42838 753975 42890 753981
rect 42838 753917 42890 753923
rect 42850 750651 42878 753917
rect 42946 753093 42974 756951
rect 42934 753087 42986 753093
rect 42934 753029 42986 753035
rect 42934 752939 42986 752945
rect 42934 752881 42986 752887
rect 42838 750645 42890 750651
rect 42838 750587 42890 750593
rect 42836 750462 42892 750471
rect 42836 750397 42892 750406
rect 42070 749831 42122 749837
rect 42070 749773 42122 749779
rect 42742 749831 42794 749837
rect 42742 749773 42794 749779
rect 42082 749546 42110 749773
rect 42166 747463 42218 747469
rect 42166 747405 42218 747411
rect 42178 747030 42206 747405
rect 42850 747321 42878 750397
rect 42838 747315 42890 747321
rect 42838 747257 42890 747263
rect 42836 747206 42892 747215
rect 42836 747141 42892 747150
rect 42166 746945 42218 746951
rect 42166 746887 42218 746893
rect 42740 746910 42796 746919
rect 42178 746401 42206 746887
rect 42740 746845 42796 746854
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42082 745772 42110 746073
rect 42358 745983 42410 745989
rect 42358 745925 42410 745931
rect 42166 745539 42218 745545
rect 42166 745481 42218 745487
rect 42178 745180 42206 745481
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42178 743365 42206 743779
rect 42070 743245 42122 743251
rect 42070 743187 42122 743193
rect 42082 742738 42110 743187
rect 42166 742653 42218 742659
rect 42166 742595 42218 742601
rect 42178 742072 42206 742595
rect 42370 741993 42398 745925
rect 42754 742659 42782 746845
rect 42850 743251 42878 747141
rect 42946 746951 42974 752881
rect 43042 751835 43070 757025
rect 43030 751829 43082 751835
rect 43030 751771 43082 751777
rect 43028 751646 43084 751655
rect 43028 751581 43084 751590
rect 42934 746945 42986 746951
rect 42934 746887 42986 746893
rect 42934 746797 42986 746803
rect 42934 746739 42986 746745
rect 42946 745545 42974 746739
rect 43042 746137 43070 751581
rect 43138 751169 43166 757099
rect 43126 751163 43178 751169
rect 43126 751105 43178 751111
rect 43126 751015 43178 751021
rect 43126 750957 43178 750963
rect 43138 747469 43166 750957
rect 43126 747463 43178 747469
rect 43126 747405 43178 747411
rect 43126 747315 43178 747321
rect 43126 747257 43178 747263
rect 43030 746131 43082 746137
rect 43030 746073 43082 746079
rect 42934 745539 42986 745545
rect 42934 745481 42986 745487
rect 43138 743843 43166 747257
rect 43126 743837 43178 743843
rect 43126 743779 43178 743785
rect 42838 743245 42890 743251
rect 42838 743187 42890 743193
rect 42742 742653 42794 742659
rect 42742 742595 42794 742601
rect 42166 741987 42218 741993
rect 42166 741929 42218 741935
rect 42358 741987 42410 741993
rect 42358 741929 42410 741935
rect 42178 741525 42206 741929
rect 41588 731518 41644 731527
rect 41588 731453 41644 731462
rect 41602 728969 41630 731453
rect 41684 731370 41740 731379
rect 41684 731305 41740 731314
rect 41590 728963 41642 728969
rect 41590 728905 41642 728911
rect 41602 727679 41630 728905
rect 41698 728747 41726 731305
rect 41780 730482 41836 730491
rect 41780 730417 41782 730426
rect 41834 730417 41836 730426
rect 41782 730385 41834 730391
rect 41780 729964 41836 729973
rect 41780 729899 41782 729908
rect 41834 729899 41836 729908
rect 41782 729867 41834 729873
rect 41780 729446 41836 729455
rect 41780 729381 41782 729390
rect 41834 729381 41836 729390
rect 41782 729349 41834 729355
rect 43234 729043 43262 771381
rect 43414 757453 43466 757459
rect 43414 757395 43466 757401
rect 43318 757231 43370 757237
rect 43318 757173 43370 757179
rect 43330 753981 43358 757173
rect 43318 753975 43370 753981
rect 43318 753917 43370 753923
rect 43426 752945 43454 757395
rect 43606 757379 43658 757385
rect 43606 757321 43658 757327
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43414 752939 43466 752945
rect 43414 752881 43466 752887
rect 43318 752051 43370 752057
rect 43318 751993 43370 751999
rect 43330 745619 43358 751993
rect 43522 751021 43550 757247
rect 43510 751015 43562 751021
rect 43510 750957 43562 750963
rect 43618 746803 43646 757321
rect 43606 746797 43658 746803
rect 43606 746739 43658 746745
rect 43318 745613 43370 745619
rect 43318 745555 43370 745561
rect 41782 729037 41834 729043
rect 41780 729002 41782 729011
rect 43222 729037 43274 729043
rect 41834 729002 41836 729011
rect 43222 728979 43274 728985
rect 41780 728937 41836 728946
rect 41686 728741 41738 728747
rect 41686 728683 41738 728689
rect 41588 727670 41644 727679
rect 41588 727605 41644 727614
rect 41698 726791 41726 728683
rect 41780 728410 41836 728419
rect 41780 728345 41782 728354
rect 41834 728345 41836 728354
rect 43318 728371 43370 728377
rect 41782 728313 41834 728319
rect 43318 728313 43370 728319
rect 41780 727966 41836 727975
rect 41780 727901 41782 727910
rect 41834 727901 41836 727910
rect 41782 727869 41834 727875
rect 41780 726930 41836 726939
rect 41780 726865 41782 726874
rect 41834 726865 41836 726874
rect 43222 726891 43274 726897
rect 41782 726833 41834 726839
rect 43222 726833 43274 726839
rect 41684 726782 41740 726791
rect 41684 726717 41740 726726
rect 41780 726042 41836 726051
rect 41780 725977 41782 725986
rect 41834 725977 41836 725986
rect 42934 726003 42986 726009
rect 41782 725945 41834 725951
rect 42934 725945 42986 725951
rect 41876 725450 41932 725459
rect 41876 725385 41932 725394
rect 39764 724710 39820 724719
rect 39764 724645 39820 724654
rect 34484 722786 34540 722795
rect 34484 722721 34540 722730
rect 28820 718198 28876 718207
rect 28820 718133 28876 718142
rect 28834 717763 28862 718133
rect 28820 717754 28876 717763
rect 28820 717689 28876 717698
rect 34498 715691 34526 722721
rect 34484 715682 34540 715691
rect 34484 715617 34540 715626
rect 39778 714951 39806 724645
rect 41684 724118 41740 724127
rect 41684 724053 41740 724062
rect 41588 721306 41644 721315
rect 41588 721241 41644 721250
rect 41602 721051 41630 721241
rect 41590 721045 41642 721051
rect 41590 720987 41642 720993
rect 41588 720714 41644 720723
rect 41588 720649 41590 720658
rect 41642 720649 41644 720658
rect 41590 720617 41642 720623
rect 41588 719826 41644 719835
rect 41588 719761 41644 719770
rect 41602 719349 41630 719761
rect 41590 719343 41642 719349
rect 41590 719285 41642 719291
rect 41588 719234 41644 719243
rect 41588 719169 41644 719178
rect 41492 717754 41548 717763
rect 41492 717689 41494 717698
rect 41546 717689 41548 717698
rect 41494 717657 41546 717663
rect 41602 717573 41630 719169
rect 41590 717567 41642 717573
rect 41590 717509 41642 717515
rect 39764 714942 39820 714951
rect 39764 714877 39820 714886
rect 41698 714095 41726 724053
rect 41780 723378 41836 723387
rect 41780 723313 41836 723322
rect 41686 714089 41738 714095
rect 41686 714031 41738 714037
rect 41794 713873 41822 723313
rect 41890 715649 41918 725385
rect 41972 724562 42028 724571
rect 41972 724497 42028 724506
rect 41878 715643 41930 715649
rect 41878 715585 41930 715591
rect 41986 714063 42014 724497
rect 42164 722490 42220 722499
rect 42164 722425 42220 722434
rect 42068 720418 42124 720427
rect 42068 720353 42124 720362
rect 41972 714054 42028 714063
rect 41972 713989 42028 713998
rect 42082 713915 42110 720353
rect 42178 719664 42206 722425
rect 42260 721898 42316 721907
rect 42260 721833 42316 721842
rect 42274 719793 42302 721833
rect 42946 720014 42974 725945
rect 43030 721045 43082 721051
rect 43030 720987 43082 720993
rect 42754 719986 42974 720014
rect 42262 719787 42314 719793
rect 42262 719729 42314 719735
rect 42178 719636 42302 719664
rect 42166 719491 42218 719497
rect 42166 719433 42218 719439
rect 42178 714211 42206 719433
rect 42164 714202 42220 714211
rect 42164 714137 42220 714146
rect 42068 713906 42124 713915
rect 41782 713867 41834 713873
rect 42068 713841 42124 713850
rect 41782 713809 41834 713815
rect 42274 713799 42302 719636
rect 42754 715839 42782 719986
rect 42838 719787 42890 719793
rect 42838 719729 42890 719735
rect 42740 715830 42796 715839
rect 42740 715765 42796 715774
rect 42742 715643 42794 715649
rect 42742 715585 42794 715591
rect 42262 713793 42314 713799
rect 42262 713735 42314 713741
rect 41782 713571 41834 713577
rect 41782 713513 41834 713519
rect 41794 713064 41822 713513
rect 42754 711727 42782 715585
rect 42850 714507 42878 719729
rect 42934 717567 42986 717573
rect 42934 717509 42986 717515
rect 42836 714498 42892 714507
rect 42836 714433 42892 714442
rect 42838 714311 42890 714317
rect 42838 714253 42890 714259
rect 42070 711721 42122 711727
rect 42070 711663 42122 711669
rect 42742 711721 42794 711727
rect 42742 711663 42794 711669
rect 42082 711214 42110 711663
rect 42742 711573 42794 711579
rect 42742 711515 42794 711521
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42754 709951 42782 711515
rect 42850 710913 42878 714253
rect 42946 711228 42974 717509
rect 43042 714243 43070 720987
rect 43126 720675 43178 720681
rect 43126 720617 43178 720623
rect 43138 719497 43166 720617
rect 43126 719491 43178 719497
rect 43126 719433 43178 719439
rect 43126 719343 43178 719349
rect 43126 719285 43178 719291
rect 43030 714237 43082 714243
rect 43030 714179 43082 714185
rect 43030 714089 43082 714095
rect 43030 714031 43082 714037
rect 43042 711357 43070 714031
rect 43030 711351 43082 711357
rect 43030 711293 43082 711299
rect 42946 711200 43070 711228
rect 42932 711094 42988 711103
rect 42932 711029 42988 711038
rect 42838 710907 42890 710913
rect 42838 710849 42890 710855
rect 42836 710798 42892 710807
rect 42836 710733 42892 710742
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42742 709945 42794 709951
rect 42742 709887 42794 709893
rect 42178 709364 42206 709887
rect 42742 709797 42794 709803
rect 42742 709739 42794 709745
rect 42082 708545 42110 708698
rect 42070 708539 42122 708545
rect 42070 708481 42122 708487
rect 42070 708391 42122 708397
rect 42070 708333 42122 708339
rect 42082 708180 42110 708333
rect 42164 707986 42220 707995
rect 42164 707921 42220 707930
rect 42178 707514 42206 707921
rect 42166 707429 42218 707435
rect 42166 707371 42218 707377
rect 42178 706881 42206 707371
rect 42754 706621 42782 709739
rect 42166 706615 42218 706621
rect 42166 706557 42218 706563
rect 42742 706615 42794 706621
rect 42742 706557 42794 706563
rect 42178 706330 42206 706557
rect 42740 705174 42796 705183
rect 42740 705109 42796 705118
rect 42358 704839 42410 704845
rect 42358 704781 42410 704787
rect 42166 704321 42218 704327
rect 42166 704263 42218 704269
rect 42178 703845 42206 704263
rect 42070 703581 42122 703587
rect 42070 703523 42122 703529
rect 42082 703222 42110 703523
rect 42370 702921 42398 704781
rect 42166 702915 42218 702921
rect 42166 702857 42218 702863
rect 42358 702915 42410 702921
rect 42358 702857 42410 702863
rect 42178 702556 42206 702857
rect 42166 702471 42218 702477
rect 42166 702413 42218 702419
rect 42178 702005 42206 702413
rect 42070 700547 42122 700553
rect 42070 700489 42122 700495
rect 42082 700188 42110 700489
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42178 699522 42206 700045
rect 42754 699443 42782 705109
rect 42850 702477 42878 710733
rect 42946 704327 42974 711029
rect 43042 708397 43070 711200
rect 43030 708391 43082 708397
rect 43030 708333 43082 708339
rect 43028 708282 43084 708291
rect 43028 708217 43084 708226
rect 42934 704321 42986 704327
rect 42934 704263 42986 704269
rect 42932 704138 42988 704147
rect 42932 704073 42988 704082
rect 42838 702471 42890 702477
rect 42838 702413 42890 702419
rect 42946 700109 42974 704073
rect 43042 703587 43070 708217
rect 43138 707435 43166 719285
rect 43126 707429 43178 707435
rect 43126 707371 43178 707377
rect 43124 707246 43180 707255
rect 43124 707181 43180 707190
rect 43030 703581 43082 703587
rect 43030 703523 43082 703529
rect 43138 700553 43166 707181
rect 43126 700547 43178 700553
rect 43126 700489 43178 700495
rect 42934 700103 42986 700109
rect 42934 700045 42986 700051
rect 42166 699437 42218 699443
rect 42166 699379 42218 699385
rect 42742 699437 42794 699443
rect 42742 699379 42794 699385
rect 42178 698856 42206 699379
rect 42070 698475 42122 698481
rect 42070 698417 42122 698423
rect 42082 698338 42110 698417
rect 41780 686896 41836 686905
rect 41780 686831 41782 686840
rect 41834 686831 41836 686840
rect 41782 686799 41834 686805
rect 41780 686378 41836 686387
rect 41780 686313 41782 686322
rect 41834 686313 41836 686322
rect 41782 686281 41834 686287
rect 41588 685638 41644 685647
rect 41588 685573 41590 685582
rect 41642 685573 41644 685582
rect 41590 685541 41642 685547
rect 41782 685377 41834 685383
rect 41780 685342 41782 685351
rect 41834 685342 41836 685351
rect 41780 685277 41836 685286
rect 41780 684898 41836 684907
rect 41780 684833 41782 684842
rect 41834 684833 41836 684842
rect 41782 684801 41834 684807
rect 41782 683897 41834 683903
rect 41780 683862 41782 683871
rect 41834 683862 41836 683871
rect 41780 683797 41836 683806
rect 43234 683015 43262 726833
rect 43330 685383 43358 728313
rect 43414 727927 43466 727933
rect 43414 727869 43466 727875
rect 43318 685377 43370 685383
rect 43318 685319 43370 685325
rect 43426 683903 43454 727869
rect 43510 714237 43562 714243
rect 43510 714179 43562 714185
rect 43522 711579 43550 714179
rect 43606 713793 43658 713799
rect 43606 713735 43658 713741
rect 43510 711573 43562 711579
rect 43510 711515 43562 711521
rect 43510 708539 43562 708545
rect 43510 708481 43562 708487
rect 43522 702699 43550 708481
rect 43618 704845 43646 713735
rect 43606 704839 43658 704845
rect 43606 704781 43658 704787
rect 43510 702693 43562 702699
rect 43510 702635 43562 702641
rect 43796 702066 43852 702075
rect 43796 702001 43852 702010
rect 43810 698481 43838 702001
rect 43798 698475 43850 698481
rect 43798 698417 43850 698423
rect 43606 684859 43658 684865
rect 43606 684801 43658 684807
rect 43414 683897 43466 683903
rect 43414 683839 43466 683845
rect 41590 683009 41642 683015
rect 41588 682974 41590 682983
rect 43222 683009 43274 683015
rect 41642 682974 41644 682983
rect 43222 682951 43274 682957
rect 41588 682909 41644 682918
rect 39764 682234 39820 682243
rect 39764 682169 39820 682178
rect 37364 680754 37420 680763
rect 37364 680689 37420 680698
rect 34484 678682 34540 678691
rect 34484 678617 34540 678626
rect 23060 674538 23116 674547
rect 23060 674473 23116 674482
rect 23074 674103 23102 674473
rect 23060 674094 23116 674103
rect 23060 674029 23116 674038
rect 34498 672581 34526 678617
rect 34486 672575 34538 672581
rect 34486 672517 34538 672523
rect 37378 671323 37406 680689
rect 39778 673913 39806 682169
rect 41780 681864 41836 681873
rect 41780 681799 41836 681808
rect 39860 681494 39916 681503
rect 39860 681429 39916 681438
rect 39766 673907 39818 673913
rect 39766 673849 39818 673855
rect 37366 671317 37418 671323
rect 37366 671259 37418 671265
rect 39874 671143 39902 681429
rect 41794 680721 41822 681799
rect 41782 680715 41834 680721
rect 41782 680657 41834 680663
rect 43030 680715 43082 680721
rect 43030 680657 43082 680663
rect 41972 680310 42028 680319
rect 41972 680245 42028 680254
rect 41780 679866 41836 679875
rect 41780 679801 41836 679810
rect 40244 679126 40300 679135
rect 40244 679061 40300 679070
rect 40258 673659 40286 679061
rect 41684 676610 41740 676619
rect 41684 676545 41740 676554
rect 41588 676166 41644 676175
rect 41588 676101 41590 676110
rect 41642 676101 41644 676110
rect 41590 676069 41642 676075
rect 41588 675722 41644 675731
rect 41588 675657 41644 675666
rect 41602 674357 41630 675657
rect 41590 674351 41642 674357
rect 41590 674293 41642 674299
rect 41588 674094 41644 674103
rect 41588 674029 41590 674038
rect 41642 674029 41644 674038
rect 41590 673997 41642 674003
rect 41494 673907 41546 673913
rect 41494 673849 41546 673855
rect 40244 673650 40300 673659
rect 40244 673585 40300 673594
rect 41506 671249 41534 673849
rect 41494 671243 41546 671249
rect 41494 671185 41546 671191
rect 39860 671134 39916 671143
rect 39860 671069 39916 671078
rect 41698 670995 41726 676545
rect 41684 670986 41740 670995
rect 41684 670921 41740 670930
rect 41794 670657 41822 679801
rect 41876 677942 41932 677951
rect 41876 677877 41932 677886
rect 41890 670847 41918 677877
rect 41986 671397 42014 680245
rect 42260 678386 42316 678395
rect 42260 678321 42316 678330
rect 42068 677350 42124 677359
rect 42068 677285 42124 677294
rect 41974 671391 42026 671397
rect 41974 671333 42026 671339
rect 41876 670838 41932 670847
rect 41876 670773 41932 670782
rect 42082 670699 42110 677285
rect 42166 672575 42218 672581
rect 42166 672517 42218 672523
rect 42178 671175 42206 672517
rect 42166 671169 42218 671175
rect 42166 671111 42218 671117
rect 42068 670690 42124 670699
rect 41782 670651 41834 670657
rect 42274 670657 42302 678321
rect 42934 674351 42986 674357
rect 42934 674293 42986 674299
rect 42838 671095 42890 671101
rect 42838 671037 42890 671043
rect 42068 670625 42124 670634
rect 42262 670651 42314 670657
rect 41782 670593 41834 670599
rect 42262 670593 42314 670599
rect 41782 670355 41834 670361
rect 41782 670297 41834 670303
rect 41794 669848 41822 670297
rect 42166 668579 42218 668585
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42850 667919 42878 671037
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42838 667913 42890 667919
rect 42838 667855 42890 667861
rect 42178 667361 42206 667855
rect 42838 667765 42890 667771
rect 42838 667707 42890 667713
rect 41876 666694 41932 666703
rect 41876 666629 41932 666638
rect 41890 666148 41918 666629
rect 42082 665329 42110 665521
rect 42166 665397 42218 665403
rect 42166 665339 42218 665345
rect 42070 665323 42122 665329
rect 42070 665265 42122 665271
rect 42178 664964 42206 665339
rect 42164 664770 42220 664779
rect 42164 664705 42220 664714
rect 42178 664298 42206 664705
rect 42070 663991 42122 663997
rect 42070 663933 42122 663939
rect 42082 663706 42110 663933
rect 42166 663399 42218 663405
rect 42166 663341 42218 663347
rect 42178 663114 42206 663341
rect 41780 660922 41836 660931
rect 41780 660857 41836 660866
rect 41794 660672 41822 660857
rect 42070 660439 42122 660445
rect 42070 660381 42122 660387
rect 42082 660006 42110 660381
rect 42850 659927 42878 667707
rect 42946 665403 42974 674293
rect 43042 668585 43070 680657
rect 43126 676127 43178 676133
rect 43126 676069 43178 676075
rect 43138 671564 43166 676069
rect 43138 671536 43262 671564
rect 43126 671391 43178 671397
rect 43126 671333 43178 671339
rect 43030 668579 43082 668585
rect 43030 668521 43082 668527
rect 43138 668511 43166 671333
rect 43126 668505 43178 668511
rect 43126 668447 43178 668453
rect 43234 668308 43262 671536
rect 43510 671243 43562 671249
rect 43510 671185 43562 671191
rect 43318 671169 43370 671175
rect 43318 671111 43370 671117
rect 43042 668280 43262 668308
rect 42934 665397 42986 665403
rect 42934 665339 42986 665345
rect 42934 665249 42986 665255
rect 42934 665191 42986 665197
rect 42946 660445 42974 665191
rect 43042 663997 43070 668280
rect 43126 668209 43178 668215
rect 43126 668151 43178 668157
rect 43030 663991 43082 663997
rect 43030 663933 43082 663939
rect 43138 663553 43166 668151
rect 43330 667771 43358 671111
rect 43414 670651 43466 670657
rect 43414 670593 43466 670599
rect 43318 667765 43370 667771
rect 43318 667707 43370 667713
rect 43426 665255 43454 670593
rect 43414 665249 43466 665255
rect 43414 665191 43466 665197
rect 43126 663547 43178 663553
rect 43126 663489 43178 663495
rect 43522 663424 43550 671185
rect 43042 663396 43550 663424
rect 42934 660439 42986 660445
rect 42934 660381 42986 660387
rect 42932 660330 42988 660339
rect 42932 660265 42988 660274
rect 42166 659921 42218 659927
rect 42166 659863 42218 659869
rect 42838 659921 42890 659927
rect 42838 659863 42890 659869
rect 42178 659340 42206 659863
rect 42836 659738 42892 659747
rect 42836 659673 42892 659682
rect 42070 659107 42122 659113
rect 42070 659049 42122 659055
rect 42082 658822 42110 659049
rect 42070 657405 42122 657411
rect 42070 657347 42122 657353
rect 42082 656972 42110 657347
rect 42850 656893 42878 659673
rect 42166 656887 42218 656893
rect 42166 656829 42218 656835
rect 42838 656887 42890 656893
rect 42838 656829 42890 656835
rect 42178 656306 42206 656829
rect 42946 656227 42974 660265
rect 43042 657411 43070 663396
rect 43126 663325 43178 663331
rect 43126 663267 43178 663273
rect 43138 659113 43166 663267
rect 43618 659534 43646 684801
rect 43702 671317 43754 671323
rect 43702 671259 43754 671265
rect 43714 663331 43742 671259
rect 43702 663325 43754 663331
rect 43702 663267 43754 663273
rect 43522 659506 43646 659534
rect 43126 659107 43178 659113
rect 43126 659049 43178 659055
rect 43030 657405 43082 657411
rect 43030 657347 43082 657353
rect 42166 656221 42218 656227
rect 42166 656163 42218 656169
rect 42934 656221 42986 656227
rect 42934 656163 42986 656169
rect 42178 655677 42206 656163
rect 42166 655555 42218 655561
rect 42166 655497 42218 655503
rect 42178 655122 42206 655497
rect 41492 645086 41548 645095
rect 41492 645021 41548 645030
rect 41506 642611 41534 645021
rect 41684 644938 41740 644947
rect 41684 644873 41740 644882
rect 41494 642605 41546 642611
rect 41494 642547 41546 642553
rect 41506 640951 41534 642547
rect 41698 642537 41726 644873
rect 41780 643754 41836 643763
rect 41780 643689 41782 643698
rect 41834 643689 41836 643698
rect 41782 643657 41834 643663
rect 41780 643162 41836 643171
rect 41780 643097 41782 643106
rect 41834 643097 41836 643106
rect 41782 643065 41834 643071
rect 41686 642531 41738 642537
rect 41686 642473 41738 642479
rect 41588 642422 41644 642431
rect 41588 642357 41590 642366
rect 41642 642357 41644 642366
rect 41590 642325 41642 642331
rect 41492 640942 41548 640951
rect 41492 640877 41548 640886
rect 41698 639915 41726 642473
rect 43522 642241 43550 659506
rect 41782 642235 41834 642241
rect 41780 642200 41782 642209
rect 43510 642235 43562 642241
rect 41834 642200 41836 642209
rect 43510 642177 43562 642183
rect 41780 642135 41836 642144
rect 41780 641682 41836 641691
rect 41780 641617 41782 641626
rect 41834 641617 41836 641626
rect 43606 641643 43658 641649
rect 41782 641585 41834 641591
rect 43606 641585 43658 641591
rect 41780 640202 41836 640211
rect 41780 640137 41782 640146
rect 41834 640137 41836 640146
rect 43414 640163 43466 640169
rect 41782 640105 41834 640111
rect 43414 640105 43466 640111
rect 41684 639906 41740 639915
rect 41684 639841 41740 639850
rect 43426 639374 43454 640105
rect 43330 639346 43454 639374
rect 37364 639018 37420 639027
rect 37364 638953 37420 638962
rect 34388 636058 34444 636067
rect 34388 635993 34444 636002
rect 23060 631470 23116 631479
rect 23060 631405 23116 631414
rect 23074 631035 23102 631405
rect 23060 631026 23116 631035
rect 23060 630961 23116 630970
rect 34402 628075 34430 635993
rect 34484 635466 34540 635475
rect 34484 635401 34540 635410
rect 34388 628066 34444 628075
rect 34388 628001 34444 628010
rect 34498 627959 34526 635401
rect 37378 628033 37406 638953
rect 40244 638278 40300 638287
rect 40244 638213 40300 638222
rect 40148 637538 40204 637547
rect 40148 637473 40204 637482
rect 37366 628027 37418 628033
rect 37366 627969 37418 627975
rect 34486 627953 34538 627959
rect 34486 627895 34538 627901
rect 40162 627885 40190 637473
rect 40258 627927 40286 638213
rect 41492 636946 41548 636955
rect 41492 636881 41548 636890
rect 40244 627918 40300 627927
rect 40150 627879 40202 627885
rect 40244 627853 40300 627862
rect 40150 627821 40202 627827
rect 41506 627737 41534 636881
rect 41780 636650 41836 636659
rect 41780 636585 41836 636594
rect 41588 633986 41644 633995
rect 41588 633921 41590 633930
rect 41642 633921 41644 633930
rect 41590 633889 41642 633895
rect 41588 630878 41644 630887
rect 41588 630813 41590 630822
rect 41642 630813 41644 630822
rect 41590 630781 41642 630787
rect 41494 627731 41546 627737
rect 41494 627673 41546 627679
rect 41794 627441 41822 636585
rect 42068 635170 42124 635179
rect 42068 635105 42124 635114
rect 41876 633246 41932 633255
rect 41876 633181 41932 633190
rect 41890 631141 41918 633181
rect 41878 631135 41930 631141
rect 41878 631077 41930 631083
rect 42082 627483 42110 635105
rect 42836 634726 42892 634735
rect 42836 634661 42892 634670
rect 42164 633690 42220 633699
rect 42164 633625 42220 633634
rect 42178 627589 42206 633625
rect 42260 632654 42316 632663
rect 42260 632589 42316 632598
rect 42274 627663 42302 632589
rect 42850 627793 42878 634661
rect 43126 633947 43178 633953
rect 43126 633889 43178 633895
rect 43030 631135 43082 631141
rect 43030 631077 43082 631083
rect 43042 628052 43070 631077
rect 43138 628181 43166 633889
rect 43330 630734 43358 639346
rect 43330 630706 43454 630734
rect 43126 628175 43178 628181
rect 43126 628117 43178 628123
rect 43042 628024 43166 628052
rect 43138 627904 43166 628024
rect 43138 627876 43262 627904
rect 42850 627765 42974 627793
rect 42262 627657 42314 627663
rect 42262 627599 42314 627605
rect 42166 627583 42218 627589
rect 42166 627525 42218 627531
rect 42068 627474 42124 627483
rect 41782 627435 41834 627441
rect 42068 627409 42124 627418
rect 41782 627377 41834 627383
rect 41782 627213 41834 627219
rect 41782 627155 41834 627161
rect 41794 626632 41822 627155
rect 42164 625254 42220 625263
rect 42164 625189 42220 625198
rect 42838 625215 42890 625221
rect 42178 624782 42206 625189
rect 42838 625157 42890 625163
rect 42740 624810 42796 624819
rect 42740 624745 42796 624754
rect 42166 624327 42218 624333
rect 42166 624269 42218 624275
rect 42178 624161 42206 624269
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42178 622965 42206 623455
rect 42178 622113 42206 622340
rect 42166 622107 42218 622113
rect 42166 622049 42218 622055
rect 42166 621959 42218 621965
rect 42166 621901 42218 621907
rect 42178 621748 42206 621901
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42178 621125 42206 621605
rect 42070 620923 42122 620929
rect 42070 620865 42122 620871
rect 42082 620490 42110 620865
rect 42166 620405 42218 620411
rect 42166 620347 42218 620353
rect 42178 619929 42206 620347
rect 42070 617889 42122 617895
rect 42070 617831 42122 617837
rect 42082 617456 42110 617831
rect 42754 617377 42782 624745
rect 42850 617895 42878 625157
rect 42946 623519 42974 627765
rect 43234 627737 43262 627876
rect 43126 627731 43178 627737
rect 43126 627673 43178 627679
rect 43222 627731 43274 627737
rect 43222 627673 43274 627679
rect 43030 627657 43082 627663
rect 43030 627599 43082 627605
rect 42934 623513 42986 623519
rect 42934 623455 42986 623461
rect 42934 623365 42986 623371
rect 42934 623307 42986 623313
rect 42946 621003 42974 623307
rect 43042 621965 43070 627599
rect 43030 621959 43082 621965
rect 43030 621901 43082 621907
rect 43030 621811 43082 621817
rect 43030 621753 43082 621759
rect 42934 620997 42986 621003
rect 42934 620939 42986 620945
rect 42934 620849 42986 620855
rect 42934 620791 42986 620797
rect 42838 617889 42890 617895
rect 42838 617831 42890 617837
rect 42836 617706 42892 617715
rect 42836 617641 42892 617650
rect 42742 617371 42794 617377
rect 42742 617313 42794 617319
rect 42740 617262 42796 617271
rect 42166 617223 42218 617229
rect 42740 617197 42796 617206
rect 42166 617165 42218 617171
rect 42178 616790 42206 617165
rect 42166 616705 42218 616711
rect 42166 616647 42218 616653
rect 42178 616157 42206 616647
rect 42166 616039 42218 616045
rect 42166 615981 42218 615987
rect 42178 615606 42206 615981
rect 42166 614189 42218 614195
rect 42166 614131 42218 614137
rect 42178 613756 42206 614131
rect 42166 613671 42218 613677
rect 42166 613613 42218 613619
rect 42178 613121 42206 613613
rect 42754 613011 42782 617197
rect 42850 613677 42878 617641
rect 42946 616711 42974 620791
rect 42934 616705 42986 616711
rect 42934 616647 42986 616653
rect 43042 616045 43070 621753
rect 43138 620411 43166 627673
rect 43426 627608 43454 630706
rect 43510 628175 43562 628181
rect 43510 628117 43562 628123
rect 43222 627583 43274 627589
rect 43222 627525 43274 627531
rect 43330 627580 43454 627608
rect 43234 625221 43262 627525
rect 43222 625215 43274 625221
rect 43222 625157 43274 625163
rect 43222 620701 43274 620707
rect 43222 620643 43274 620649
rect 43126 620405 43178 620411
rect 43126 620347 43178 620353
rect 43126 620257 43178 620263
rect 43126 620199 43178 620205
rect 43030 616039 43082 616045
rect 43030 615981 43082 615987
rect 43138 614195 43166 620199
rect 43126 614189 43178 614195
rect 43126 614131 43178 614137
rect 42838 613671 42890 613677
rect 42838 613613 42890 613619
rect 42070 613005 42122 613011
rect 42070 612947 42122 612953
rect 42742 613005 42794 613011
rect 42742 612947 42794 612953
rect 42082 612498 42110 612947
rect 42166 612413 42218 612419
rect 42166 612355 42218 612361
rect 42178 611906 42206 612355
rect 40340 602166 40396 602175
rect 40340 602101 40396 602110
rect 40354 597735 40382 602101
rect 41780 600538 41836 600547
rect 41780 600473 41782 600482
rect 41834 600473 41836 600482
rect 41782 600441 41834 600447
rect 41588 599798 41644 599807
rect 41588 599733 41590 599742
rect 41642 599733 41644 599742
rect 41590 599701 41642 599707
rect 41780 599428 41836 599437
rect 41780 599363 41782 599372
rect 41834 599363 41836 599372
rect 41782 599331 41834 599337
rect 41780 599058 41836 599067
rect 43234 599025 43262 620643
rect 41780 598993 41782 599002
rect 41834 598993 41836 599002
rect 43222 599019 43274 599025
rect 41782 598961 41834 598967
rect 43222 598961 43274 598967
rect 41588 598318 41644 598327
rect 41588 598253 41590 598262
rect 41642 598253 41644 598262
rect 41590 598221 41642 598227
rect 40340 597726 40396 597735
rect 40340 597661 40396 597670
rect 41588 596246 41644 596255
rect 43330 596213 43358 627580
rect 43414 627509 43466 627515
rect 43414 627451 43466 627457
rect 43426 623371 43454 627451
rect 43414 623365 43466 623371
rect 43414 623307 43466 623313
rect 43522 621669 43550 628117
rect 43510 621663 43562 621669
rect 43510 621605 43562 621611
rect 43618 620707 43646 641585
rect 43894 628027 43946 628033
rect 43894 627969 43946 627975
rect 43798 627953 43850 627959
rect 43798 627895 43850 627901
rect 43702 627879 43754 627885
rect 43702 627821 43754 627827
rect 43714 621817 43742 627821
rect 43702 621811 43754 621817
rect 43702 621753 43754 621759
rect 43810 620855 43838 627895
rect 43798 620849 43850 620855
rect 43798 620791 43850 620797
rect 43606 620701 43658 620707
rect 43606 620643 43658 620649
rect 43906 620263 43934 627969
rect 43894 620257 43946 620263
rect 43894 620199 43946 620205
rect 43510 598279 43562 598285
rect 43510 598221 43562 598227
rect 41588 596181 41590 596190
rect 41642 596181 41644 596190
rect 43318 596207 43370 596213
rect 41590 596149 41642 596155
rect 43318 596149 43370 596155
rect 41492 595802 41548 595811
rect 41492 595737 41548 595746
rect 34388 594766 34444 594775
rect 34388 594701 34444 594710
rect 23060 588254 23116 588263
rect 23060 588189 23116 588198
rect 23074 587819 23102 588189
rect 23060 587810 23116 587819
rect 23060 587745 23116 587754
rect 34402 584859 34430 594701
rect 34484 592842 34540 592851
rect 34484 592777 34540 592786
rect 34388 584850 34444 584859
rect 34388 584785 34444 584794
rect 34498 584711 34526 592777
rect 34484 584702 34540 584711
rect 34484 584637 34540 584646
rect 41506 584563 41534 595737
rect 41780 595506 41836 595515
rect 41780 595441 41836 595450
rect 41684 594322 41740 594331
rect 41684 594257 41740 594266
rect 41588 591362 41644 591371
rect 41588 591297 41644 591306
rect 41602 590589 41630 591297
rect 41590 590583 41642 590589
rect 41590 590525 41642 590531
rect 41588 589882 41644 589891
rect 41588 589817 41644 589826
rect 41602 589405 41630 589817
rect 41590 589399 41642 589405
rect 41590 589341 41642 589347
rect 41588 589290 41644 589299
rect 41588 589225 41644 589234
rect 41602 587925 41630 589225
rect 41590 587919 41642 587925
rect 41590 587861 41642 587867
rect 41588 587810 41644 587819
rect 41588 587745 41644 587754
rect 41602 587629 41630 587745
rect 41590 587623 41642 587629
rect 41590 587565 41642 587571
rect 41698 584563 41726 594257
rect 41794 593549 41822 595441
rect 42164 594026 42220 594035
rect 42164 593961 42220 593970
rect 41782 593543 41834 593549
rect 41782 593485 41834 593491
rect 41780 593434 41836 593443
rect 41780 593369 41836 593378
rect 41492 584554 41548 584563
rect 41492 584489 41548 584498
rect 41684 584554 41740 584563
rect 41684 584489 41740 584498
rect 41794 584225 41822 593369
rect 41972 592546 42028 592555
rect 41972 592481 42028 592490
rect 41876 590992 41932 591001
rect 41876 590927 41878 590936
rect 41930 590927 41932 590936
rect 41878 590895 41930 590901
rect 41986 590756 42014 592481
rect 42068 591954 42124 591963
rect 42068 591889 42124 591898
rect 41890 590728 42014 590756
rect 41890 584267 41918 590728
rect 41974 589547 42026 589553
rect 41974 589489 42026 589495
rect 41986 584711 42014 589489
rect 41972 584702 42028 584711
rect 41972 584637 42028 584646
rect 42082 584595 42110 591889
rect 42070 584589 42122 584595
rect 42070 584531 42122 584537
rect 42178 584521 42206 593961
rect 43030 593543 43082 593549
rect 43030 593485 43082 593491
rect 42838 590583 42890 590589
rect 42838 590525 42890 590531
rect 42356 590474 42412 590483
rect 42356 590409 42412 590418
rect 42850 590414 42878 590525
rect 42370 584669 42398 590409
rect 42850 590386 42974 590414
rect 42838 587919 42890 587925
rect 42838 587861 42890 587867
rect 42358 584663 42410 584669
rect 42358 584605 42410 584611
rect 42166 584515 42218 584521
rect 42166 584457 42218 584463
rect 41876 584258 41932 584267
rect 41782 584219 41834 584225
rect 41876 584193 41932 584202
rect 41782 584161 41834 584167
rect 41782 583997 41834 584003
rect 41782 583939 41834 583945
rect 41794 583445 41822 583939
rect 42166 582147 42218 582153
rect 42166 582089 42218 582095
rect 42178 581605 42206 582089
rect 42178 580895 42206 580974
rect 42166 580889 42218 580895
rect 42166 580831 42218 580837
rect 42070 580297 42122 580303
rect 42070 580239 42122 580245
rect 42082 579790 42110 580239
rect 42178 578971 42206 579124
rect 42166 578965 42218 578971
rect 42166 578907 42218 578913
rect 42850 578823 42878 587861
rect 42946 580303 42974 590386
rect 43042 582153 43070 593485
rect 43126 590953 43178 590959
rect 43126 590895 43178 590901
rect 43138 589553 43166 590895
rect 43126 589547 43178 589553
rect 43126 589489 43178 589495
rect 43126 589399 43178 589405
rect 43126 589341 43178 589347
rect 43030 582147 43082 582153
rect 43030 582089 43082 582095
rect 43030 581999 43082 582005
rect 43030 581941 43082 581947
rect 42934 580297 42986 580303
rect 42934 580239 42986 580245
rect 42934 580149 42986 580155
rect 42934 580091 42986 580097
rect 42166 578817 42218 578823
rect 42166 578759 42218 578765
rect 42838 578817 42890 578823
rect 42838 578759 42890 578765
rect 42178 578569 42206 578759
rect 42836 578634 42892 578643
rect 42836 578569 42892 578578
rect 42068 578190 42124 578199
rect 42068 578125 42124 578134
rect 42082 577940 42110 578125
rect 42166 577855 42218 577861
rect 42166 577797 42218 577803
rect 42178 577274 42206 577797
rect 42070 576967 42122 576973
rect 42070 576909 42122 576915
rect 42082 576756 42110 576909
rect 42166 574599 42218 574605
rect 42166 574541 42218 574547
rect 42178 574240 42206 574541
rect 42166 574155 42218 574161
rect 42166 574097 42218 574103
rect 42178 573574 42206 574097
rect 41780 573454 41836 573463
rect 41780 573389 41836 573398
rect 41794 572982 41822 573389
rect 42850 572681 42878 578569
rect 42946 574161 42974 580091
rect 43042 576973 43070 581941
rect 43138 577861 43166 589341
rect 43414 584663 43466 584669
rect 43414 584605 43466 584611
rect 43318 584589 43370 584595
rect 43318 584531 43370 584537
rect 43222 584515 43274 584521
rect 43222 584457 43274 584463
rect 43234 582005 43262 584457
rect 43222 581999 43274 582005
rect 43222 581941 43274 581947
rect 43330 580155 43358 584531
rect 43318 580149 43370 580155
rect 43318 580091 43370 580097
rect 43126 577855 43178 577861
rect 43126 577797 43178 577803
rect 43426 577732 43454 584605
rect 43138 577704 43454 577732
rect 43030 576967 43082 576973
rect 43030 576909 43082 576915
rect 43028 576858 43084 576867
rect 43028 576793 43084 576802
rect 42934 574155 42986 574161
rect 42934 574097 42986 574103
rect 42932 574046 42988 574055
rect 42932 573981 42988 573990
rect 42166 572675 42218 572681
rect 42166 572617 42218 572623
rect 42838 572675 42890 572681
rect 42838 572617 42890 572623
rect 42178 572390 42206 572617
rect 42082 570461 42110 570540
rect 42070 570455 42122 570461
rect 42070 570397 42122 570403
rect 42946 570387 42974 573981
rect 43042 570461 43070 576793
rect 43138 574605 43166 577704
rect 43126 574599 43178 574605
rect 43126 574541 43178 574547
rect 43124 574490 43180 574499
rect 43124 574425 43180 574434
rect 43030 570455 43082 570461
rect 43030 570397 43082 570403
rect 42166 570381 42218 570387
rect 42166 570323 42218 570329
rect 42934 570381 42986 570387
rect 42934 570323 42986 570329
rect 42178 570254 42206 570323
rect 43138 570254 43166 574425
rect 43522 570254 43550 598221
rect 42082 570226 42206 570254
rect 42946 570226 43166 570254
rect 43234 570226 43550 570254
rect 42082 569948 42110 570226
rect 42946 569721 42974 570226
rect 42070 569715 42122 569721
rect 42070 569657 42122 569663
rect 42934 569715 42986 569721
rect 42934 569657 42986 569663
rect 42082 569282 42110 569657
rect 42166 569197 42218 569203
rect 42166 569139 42218 569145
rect 42178 568725 42206 569139
rect 43028 544446 43084 544455
rect 43028 544381 43084 544390
rect 41588 543114 41644 543123
rect 41588 543049 41590 543058
rect 41642 543049 41644 543058
rect 41590 543017 41642 543023
rect 41780 542744 41836 542753
rect 41780 542679 41782 542688
rect 41834 542679 41836 542688
rect 41782 542647 41834 542653
rect 41780 542226 41836 542235
rect 41780 542161 41782 542170
rect 41834 542161 41836 542170
rect 41782 542129 41834 542135
rect 41782 541817 41834 541823
rect 41780 541782 41782 541791
rect 41834 541782 41836 541791
rect 41780 541717 41836 541726
rect 42742 541595 42794 541601
rect 42742 541537 42794 541543
rect 42178 539751 42206 540245
rect 42166 539745 42218 539751
rect 42166 539687 42218 539693
rect 41794 538239 41822 538424
rect 41780 538230 41836 538239
rect 42754 538197 42782 541537
rect 42838 541521 42890 541527
rect 42838 541463 42890 541469
rect 41780 538165 41836 538174
rect 42166 538191 42218 538197
rect 42166 538133 42218 538139
rect 42742 538191 42794 538197
rect 42742 538133 42794 538139
rect 42178 537758 42206 538133
rect 42740 536750 42796 536759
rect 42740 536685 42796 536694
rect 41794 536315 41822 536574
rect 42166 536489 42218 536495
rect 42166 536431 42218 536437
rect 41780 536306 41836 536315
rect 41780 536241 41836 536250
rect 42178 535908 42206 536431
rect 41986 534983 42014 535390
rect 41972 534974 42028 534983
rect 41972 534909 42028 534918
rect 41794 534243 41822 534724
rect 41780 534234 41836 534243
rect 41780 534169 41836 534178
rect 41794 533947 41822 534058
rect 41780 533938 41836 533947
rect 41780 533873 41836 533882
rect 42754 533757 42782 536685
rect 42850 536495 42878 541463
rect 42934 539745 42986 539751
rect 42934 539687 42986 539693
rect 42946 536611 42974 539687
rect 43042 539275 43070 544381
rect 43234 541823 43262 570226
rect 43222 541817 43274 541823
rect 43222 541759 43274 541765
rect 43508 541190 43564 541199
rect 43508 541125 43564 541134
rect 43412 540746 43468 540755
rect 43412 540681 43468 540690
rect 43028 539266 43084 539275
rect 43028 539201 43084 539210
rect 43124 538822 43180 538831
rect 43124 538757 43180 538766
rect 43028 537342 43084 537351
rect 43028 537277 43084 537286
rect 42932 536602 42988 536611
rect 42932 536537 42988 536546
rect 42838 536489 42890 536495
rect 42838 536431 42890 536437
rect 42836 534678 42892 534687
rect 42836 534613 42892 534622
rect 42070 533751 42122 533757
rect 42070 533693 42122 533699
rect 42742 533751 42794 533757
rect 42742 533693 42794 533699
rect 42082 533540 42110 533693
rect 42740 533198 42796 533207
rect 42740 533133 42796 533142
rect 42754 531537 42782 533133
rect 42166 531531 42218 531537
rect 42166 531473 42218 531479
rect 42742 531531 42794 531537
rect 42742 531473 42794 531479
rect 42178 531024 42206 531473
rect 42850 530945 42878 534613
rect 42932 532754 42988 532763
rect 42932 532689 42988 532698
rect 42166 530939 42218 530945
rect 42166 530881 42218 530887
rect 42838 530939 42890 530945
rect 42838 530881 42890 530887
rect 42178 530401 42206 530881
rect 42836 530682 42892 530691
rect 42836 530617 42892 530626
rect 41794 529655 41822 529766
rect 41780 529646 41836 529655
rect 41780 529581 41836 529590
rect 42166 529459 42218 529465
rect 42166 529401 42218 529407
rect 42178 529205 42206 529401
rect 42166 527831 42218 527837
rect 42166 527773 42218 527779
rect 42178 527365 42206 527773
rect 42850 527245 42878 530617
rect 42070 527239 42122 527245
rect 42070 527181 42122 527187
rect 42838 527239 42890 527245
rect 42838 527181 42890 527187
rect 42082 526732 42110 527181
rect 42946 526505 42974 532689
rect 43042 529465 43070 537277
rect 43030 529459 43082 529465
rect 43030 529401 43082 529407
rect 43138 527837 43166 538757
rect 43126 527831 43178 527837
rect 43126 527773 43178 527779
rect 42166 526499 42218 526505
rect 42166 526441 42218 526447
rect 42934 526499 42986 526505
rect 42934 526441 42986 526447
rect 42178 526066 42206 526441
rect 42070 525981 42122 525987
rect 42070 525923 42122 525929
rect 42082 525548 42110 525923
rect 41684 525058 41740 525067
rect 41684 524993 41740 525002
rect 41588 429302 41644 429311
rect 41588 429237 41590 429246
rect 41642 429237 41644 429246
rect 41590 429205 41642 429211
rect 41698 427271 41726 524993
rect 42274 524285 42398 524304
rect 42274 524279 42410 524285
rect 42274 524276 42358 524279
rect 42358 524221 42410 524227
rect 43426 519993 43454 540681
rect 43414 519987 43466 519993
rect 43414 519929 43466 519935
rect 43414 519765 43466 519771
rect 43414 519707 43466 519713
rect 43318 514141 43370 514147
rect 43318 514083 43370 514089
rect 41780 429006 41836 429015
rect 41780 428941 41782 428950
rect 41834 428941 41836 428950
rect 41782 428909 41834 428915
rect 41780 428414 41836 428423
rect 41780 428349 41782 428358
rect 41834 428349 41836 428358
rect 41782 428317 41834 428323
rect 43330 428011 43358 514083
rect 43426 429134 43454 519707
rect 43522 514147 43550 541125
rect 43510 514141 43562 514147
rect 43510 514083 43562 514089
rect 43426 429106 43550 429134
rect 41782 428005 41834 428011
rect 41780 427970 41782 427979
rect 43318 428005 43370 428011
rect 41834 427970 41836 427979
rect 43318 427947 43370 427953
rect 41780 427905 41836 427914
rect 41780 427452 41836 427461
rect 41780 427387 41782 427396
rect 41834 427387 41836 427396
rect 43414 427413 43466 427419
rect 41782 427355 41834 427361
rect 43414 427355 43466 427361
rect 41686 427265 41738 427271
rect 41686 427207 41738 427213
rect 41780 426934 41836 426943
rect 41780 426869 41782 426878
rect 41834 426869 41836 426878
rect 43318 426895 43370 426901
rect 41782 426837 41834 426843
rect 43318 426837 43370 426843
rect 25844 425602 25900 425611
rect 25844 425537 25900 425546
rect 25858 418803 25886 425537
rect 41780 425454 41836 425463
rect 41780 425389 41836 425398
rect 41684 422198 41740 422207
rect 41684 422133 41740 422142
rect 41588 420274 41644 420283
rect 41588 420209 41644 420218
rect 25844 418794 25900 418803
rect 25844 418729 25900 418738
rect 41602 417873 41630 420209
rect 41590 417867 41642 417873
rect 41590 417809 41642 417815
rect 28820 417166 28876 417175
rect 28820 417101 28876 417110
rect 28834 416731 28862 417101
rect 41698 416856 41726 422133
rect 41794 420463 41822 425389
rect 41782 420457 41834 420463
rect 41782 420399 41834 420405
rect 41780 419978 41836 419987
rect 41780 419913 41836 419922
rect 41794 419131 41822 419913
rect 41782 419125 41834 419131
rect 41782 419067 41834 419073
rect 42838 419125 42890 419131
rect 42838 419067 42890 419073
rect 41780 419016 41836 419025
rect 41780 418951 41836 418960
rect 41794 418613 41822 418951
rect 41782 418607 41834 418613
rect 41782 418549 41834 418555
rect 41780 418498 41836 418507
rect 41780 418433 41836 418442
rect 41794 417799 41822 418433
rect 41782 417793 41834 417799
rect 41782 417735 41834 417741
rect 41780 417018 41836 417027
rect 41780 416953 41782 416962
rect 41834 416953 41836 416962
rect 41782 416921 41834 416927
rect 41698 416828 41822 416856
rect 28820 416722 28876 416731
rect 28820 416657 28876 416666
rect 41794 413433 41822 416828
rect 41782 413427 41834 413433
rect 41782 413369 41834 413375
rect 41782 413205 41834 413211
rect 41782 413147 41834 413153
rect 41794 412624 41822 413147
rect 41876 411246 41932 411255
rect 41876 411181 41932 411190
rect 41890 410805 41918 411181
rect 42178 409733 42206 410182
rect 42850 409881 42878 419067
rect 43126 418607 43178 418613
rect 43126 418549 43178 418555
rect 42934 417867 42986 417873
rect 42934 417809 42986 417815
rect 42838 409875 42890 409881
rect 42838 409817 42890 409823
rect 42166 409727 42218 409733
rect 42166 409669 42218 409675
rect 42838 409727 42890 409733
rect 42838 409669 42890 409675
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42178 408965 42206 409447
rect 42070 408099 42122 408105
rect 42070 408041 42122 408047
rect 42082 407769 42110 408041
rect 42178 408031 42206 408332
rect 42166 408025 42218 408031
rect 42166 407967 42218 407973
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42166 406915 42218 406921
rect 42166 406857 42218 406863
rect 42178 406482 42206 406857
rect 42850 406107 42878 409669
rect 42946 409511 42974 417809
rect 43030 417793 43082 417799
rect 43030 417735 43082 417741
rect 42934 409505 42986 409511
rect 42934 409447 42986 409453
rect 42934 409357 42986 409363
rect 42934 409299 42986 409305
rect 42946 407976 42974 409299
rect 43042 408105 43070 417735
rect 43138 409363 43166 418549
rect 43222 409875 43274 409881
rect 43222 409817 43274 409823
rect 43126 409357 43178 409363
rect 43126 409299 43178 409305
rect 43234 409160 43262 409817
rect 43138 409132 43262 409160
rect 43030 408099 43082 408105
rect 43030 408041 43082 408047
rect 42946 407948 43070 407976
rect 42934 407877 42986 407883
rect 42934 407819 42986 407825
rect 42838 406101 42890 406107
rect 41876 406066 41932 406075
rect 42838 406043 42890 406049
rect 41876 406001 41932 406010
rect 41890 405929 41918 406001
rect 42068 403846 42124 403855
rect 42068 403781 42124 403790
rect 42082 403448 42110 403781
rect 41780 403106 41836 403115
rect 41780 403041 41836 403050
rect 41794 402782 41822 403041
rect 41780 402662 41836 402671
rect 42946 402629 42974 407819
rect 43042 406921 43070 407948
rect 43138 407513 43166 409132
rect 43222 409061 43274 409067
rect 43222 409003 43274 409009
rect 43126 407507 43178 407513
rect 43126 407449 43178 407455
rect 43030 406915 43082 406921
rect 43030 406857 43082 406863
rect 41780 402597 41836 402606
rect 42934 402623 42986 402629
rect 41794 402157 41822 402597
rect 42934 402565 42986 402571
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42082 394563 42110 397898
rect 42070 394557 42122 394563
rect 42070 394499 42122 394505
rect 41780 386530 41836 386539
rect 41780 386465 41782 386474
rect 41834 386465 41836 386474
rect 41782 386433 41834 386439
rect 41588 385790 41644 385799
rect 41588 385725 41590 385734
rect 41642 385725 41644 385734
rect 41590 385693 41642 385699
rect 41780 385420 41836 385429
rect 41780 385355 41782 385364
rect 41834 385355 41836 385364
rect 41782 385323 41834 385329
rect 43234 385239 43262 409003
rect 41590 385233 41642 385239
rect 41588 385198 41590 385207
rect 43222 385233 43274 385239
rect 41642 385198 41644 385207
rect 43222 385175 43274 385181
rect 41588 385133 41644 385142
rect 41780 384458 41836 384467
rect 41780 384393 41782 384402
rect 41834 384393 41836 384402
rect 41782 384361 41834 384367
rect 34484 383718 34540 383727
rect 34484 383653 34540 383662
rect 28724 381646 28780 381655
rect 34498 381613 34526 383653
rect 43330 383537 43358 426837
rect 43426 409067 43454 427355
rect 43522 426499 43550 429106
rect 43508 426490 43564 426499
rect 43508 426425 43564 426434
rect 43414 409061 43466 409067
rect 43414 409003 43466 409009
rect 43510 384419 43562 384425
rect 43510 384361 43562 384367
rect 41782 383531 41834 383537
rect 41780 383496 41782 383505
rect 43318 383531 43370 383537
rect 41834 383496 41836 383505
rect 43318 383473 43370 383479
rect 41780 383431 41836 383440
rect 40244 382682 40300 382691
rect 40244 382617 40300 382626
rect 28724 381581 28780 381590
rect 34486 381607 34538 381613
rect 23060 374246 23116 374255
rect 23060 374181 23116 374190
rect 23074 373811 23102 374181
rect 23060 373802 23116 373811
rect 23060 373737 23116 373746
rect 28738 372479 28766 381581
rect 34486 381549 34538 381555
rect 39380 380758 39436 380767
rect 39380 380693 39436 380702
rect 39284 379722 39340 379731
rect 39284 379657 39340 379666
rect 39298 374361 39326 379657
rect 39286 374355 39338 374361
rect 39286 374297 39338 374303
rect 39394 372775 39422 380693
rect 39860 379722 39916 379731
rect 39860 379657 39916 379666
rect 39764 378834 39820 378843
rect 39764 378769 39820 378778
rect 39476 378242 39532 378251
rect 39476 378177 39532 378186
rect 39490 373219 39518 378177
rect 39668 377206 39724 377215
rect 39668 377141 39724 377150
rect 39682 374287 39710 377141
rect 39670 374281 39722 374287
rect 39778 374255 39806 378769
rect 39670 374223 39722 374229
rect 39764 374246 39820 374255
rect 39764 374181 39820 374190
rect 39874 373811 39902 379657
rect 40258 377247 40286 382617
rect 43318 381607 43370 381613
rect 43318 381549 43370 381555
rect 40246 377241 40298 377247
rect 40246 377183 40298 377189
rect 41780 376984 41836 376993
rect 41780 376919 41782 376928
rect 41834 376919 41836 376928
rect 42934 376945 42986 376951
rect 41782 376887 41834 376893
rect 42934 376887 42986 376893
rect 41780 376022 41836 376031
rect 41780 375957 41836 375966
rect 41588 375282 41644 375291
rect 41588 375217 41644 375226
rect 41602 374657 41630 375217
rect 41794 374805 41822 375957
rect 41782 374799 41834 374805
rect 41782 374741 41834 374747
rect 41590 374651 41642 374657
rect 41590 374593 41642 374599
rect 42838 374651 42890 374657
rect 42838 374593 42890 374599
rect 41782 374355 41834 374361
rect 41782 374297 41834 374303
rect 39860 373802 39916 373811
rect 39860 373737 39916 373746
rect 39476 373210 39532 373219
rect 39476 373145 39532 373154
rect 39380 372766 39436 372775
rect 39380 372701 39436 372710
rect 28724 372470 28780 372479
rect 28724 372405 28780 372414
rect 41794 370217 41822 374297
rect 41876 373950 41932 373959
rect 41876 373885 41878 373894
rect 41930 373885 41932 373894
rect 41878 373853 41930 373859
rect 41782 370211 41834 370217
rect 41782 370153 41834 370159
rect 41782 369989 41834 369995
rect 41782 369931 41834 369937
rect 41794 369445 41822 369931
rect 41780 368178 41836 368187
rect 41780 368113 41836 368122
rect 41794 367632 41822 368113
rect 42178 366591 42206 366966
rect 42166 366585 42218 366591
rect 42166 366527 42218 366533
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42082 365782 42110 366231
rect 42082 364741 42110 365116
rect 42850 365037 42878 374593
rect 42946 366739 42974 376887
rect 43030 374799 43082 374805
rect 43030 374741 43082 374747
rect 42934 366733 42986 366739
rect 42934 366675 42986 366681
rect 42934 366585 42986 366591
rect 42934 366527 42986 366533
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42838 365031 42890 365037
rect 42838 364973 42890 364979
rect 42070 364735 42122 364741
rect 42070 364677 42122 364683
rect 42178 364569 42206 364973
rect 42838 364735 42890 364741
rect 42838 364677 42890 364683
rect 42070 364291 42122 364297
rect 42070 364233 42122 364239
rect 42082 363932 42110 364233
rect 42166 363847 42218 363853
rect 42166 363789 42218 363795
rect 42178 363266 42206 363789
rect 41780 362850 41836 362859
rect 41780 362785 41836 362794
rect 41794 362748 41822 362785
rect 41972 360630 42028 360639
rect 41972 360565 42028 360574
rect 41986 360232 42014 360565
rect 42850 360005 42878 364677
rect 42946 361485 42974 366527
rect 43042 363853 43070 374741
rect 43126 374281 43178 374287
rect 43126 374223 43178 374229
rect 43138 366295 43166 374223
rect 43222 366733 43274 366739
rect 43222 366675 43274 366681
rect 43126 366289 43178 366295
rect 43126 366231 43178 366237
rect 43234 366092 43262 366675
rect 43138 366064 43262 366092
rect 43138 364297 43166 366064
rect 43126 364291 43178 364297
rect 43126 364233 43178 364239
rect 43030 363847 43082 363853
rect 43030 363789 43082 363795
rect 42934 361479 42986 361485
rect 42934 361421 42986 361427
rect 42838 359999 42890 360005
rect 42838 359941 42890 359947
rect 41780 359890 41836 359899
rect 41780 359825 41836 359834
rect 41794 359601 41822 359825
rect 42068 359298 42124 359307
rect 42068 359233 42124 359242
rect 42082 358974 42110 359233
rect 41780 358854 41836 358863
rect 41780 358789 41836 358798
rect 41794 358382 41822 358789
rect 41876 356930 41932 356939
rect 41876 356865 41932 356874
rect 41890 356565 41918 356865
rect 41780 356190 41836 356199
rect 41780 356125 41836 356134
rect 41794 355940 41822 356125
rect 42164 355746 42220 355755
rect 42164 355681 42220 355690
rect 42178 355274 42206 355681
rect 42178 351347 42206 354725
rect 42166 351341 42218 351347
rect 42166 351283 42218 351289
rect 41588 343314 41644 343323
rect 41588 343249 41590 343258
rect 41642 343249 41644 343258
rect 41590 343217 41642 343223
rect 41780 342944 41836 342953
rect 41780 342879 41782 342888
rect 41834 342879 41836 342888
rect 41782 342847 41834 342853
rect 41780 342426 41836 342435
rect 41780 342361 41782 342370
rect 41834 342361 41836 342370
rect 41782 342329 41834 342335
rect 41782 342017 41834 342023
rect 41780 341982 41782 341991
rect 41834 341982 41836 341991
rect 41780 341917 41836 341926
rect 41780 341464 41836 341473
rect 41780 341399 41782 341408
rect 41834 341399 41836 341408
rect 43222 341425 43274 341431
rect 41782 341367 41834 341373
rect 43222 341367 43274 341373
rect 41780 340946 41836 340955
rect 41780 340881 41782 340890
rect 41834 340881 41836 340890
rect 41782 340849 41834 340855
rect 41782 340537 41834 340543
rect 41780 340502 41782 340511
rect 41834 340502 41836 340511
rect 41780 340437 41836 340446
rect 41780 339910 41836 339919
rect 41780 339845 41782 339854
rect 41834 339845 41836 339854
rect 41782 339813 41834 339819
rect 41590 339797 41642 339803
rect 41588 339762 41590 339771
rect 41642 339762 41644 339771
rect 41588 339697 41644 339706
rect 28724 338726 28780 338735
rect 28724 338661 28780 338670
rect 23060 331178 23116 331187
rect 23060 331113 23116 331122
rect 23074 330743 23102 331113
rect 23060 330734 23116 330743
rect 23060 330669 23116 330678
rect 28738 329263 28766 338661
rect 39284 337690 39340 337699
rect 39284 337625 39340 337634
rect 39298 331187 39326 337625
rect 41684 336210 41740 336219
rect 41684 336145 41740 336154
rect 41588 334138 41644 334147
rect 41588 334073 41644 334082
rect 39284 331178 39340 331187
rect 39284 331113 39340 331122
rect 28724 329254 28780 329263
rect 28724 329189 28780 329198
rect 41602 328777 41630 334073
rect 41698 331164 41726 336145
rect 41780 333990 41836 333999
rect 41780 333925 41836 333934
rect 41794 333143 41822 333925
rect 41782 333137 41834 333143
rect 41782 333079 41834 333085
rect 42742 333137 42794 333143
rect 42742 333079 42794 333085
rect 41780 332510 41836 332519
rect 41780 332445 41836 332454
rect 41794 331589 41822 332445
rect 41782 331583 41834 331589
rect 41782 331525 41834 331531
rect 41698 331136 41822 331164
rect 41590 328771 41642 328777
rect 41590 328713 41642 328719
rect 41794 327075 41822 331136
rect 41876 331030 41932 331039
rect 41876 330965 41878 330974
rect 41930 330965 41932 330974
rect 41878 330933 41930 330939
rect 42754 328334 42782 333079
rect 42934 331583 42986 331589
rect 42934 331525 42986 331531
rect 42754 328306 42878 328334
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 41782 326625 41834 326631
rect 41782 326567 41834 326573
rect 41794 326266 41822 326567
rect 42850 325688 42878 328306
rect 42946 325817 42974 331525
rect 43030 328771 43082 328777
rect 43030 328713 43082 328719
rect 42934 325811 42986 325817
rect 42934 325753 42986 325759
rect 42850 325660 42974 325688
rect 41780 324962 41836 324971
rect 41780 324897 41836 324906
rect 41794 324416 41822 324897
rect 42082 323375 42110 323750
rect 42070 323369 42122 323375
rect 42070 323311 42122 323317
rect 42454 323369 42506 323375
rect 42454 323311 42506 323317
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42178 322566 42206 323089
rect 42082 321692 42110 321900
rect 41974 321667 42026 321673
rect 42082 321664 42206 321692
rect 41974 321609 42026 321615
rect 41986 321382 42014 321609
rect 42178 321525 42206 321664
rect 42166 321519 42218 321525
rect 42166 321461 42218 321467
rect 42166 321297 42218 321303
rect 42166 321239 42218 321245
rect 42178 320716 42206 321239
rect 42164 320522 42220 320531
rect 42164 320457 42220 320466
rect 42178 320081 42206 320457
rect 41780 319782 41836 319791
rect 41780 319717 41836 319726
rect 41794 319532 41822 319717
rect 42466 319675 42494 323311
rect 42946 321692 42974 325660
rect 43042 323153 43070 328713
rect 43126 325811 43178 325817
rect 43126 325753 43178 325759
rect 43030 323147 43082 323153
rect 43030 323089 43082 323095
rect 42946 321664 43070 321692
rect 43138 321673 43166 325753
rect 43042 321303 43070 321664
rect 43126 321667 43178 321673
rect 43126 321609 43178 321615
rect 43126 321519 43178 321525
rect 43126 321461 43178 321467
rect 43030 321297 43082 321303
rect 43030 321239 43082 321245
rect 42454 319669 42506 319675
rect 42454 319611 42506 319617
rect 42164 317414 42220 317423
rect 42164 317349 42220 317358
rect 42178 317045 42206 317349
rect 41876 316822 41932 316831
rect 43138 316789 43166 321461
rect 41876 316757 41932 316766
rect 43126 316783 43178 316789
rect 41890 316424 41918 316757
rect 43126 316725 43178 316731
rect 41780 316082 41836 316091
rect 41780 316017 41836 316026
rect 41794 315758 41822 316017
rect 41780 315638 41836 315647
rect 41780 315573 41836 315582
rect 41794 315205 41822 315573
rect 42068 313714 42124 313723
rect 42068 313649 42124 313658
rect 42082 313390 42110 313649
rect 41780 313122 41836 313131
rect 41780 313057 41836 313066
rect 41794 312724 41822 313057
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42178 308131 42206 311540
rect 42166 308125 42218 308131
rect 42166 308067 42218 308073
rect 41588 299950 41644 299959
rect 41588 299885 41644 299894
rect 41602 299621 41630 299885
rect 41780 299802 41836 299811
rect 41780 299737 41782 299746
rect 41834 299737 41836 299746
rect 41782 299705 41834 299711
rect 41878 299689 41930 299695
rect 41878 299631 41930 299637
rect 41590 299615 41642 299621
rect 41590 299557 41642 299563
rect 39668 299506 39724 299515
rect 39668 299441 39724 299450
rect 28724 295510 28780 295519
rect 28724 295445 28780 295454
rect 23060 287962 23116 287971
rect 23060 287897 23116 287906
rect 23074 287527 23102 287897
rect 23060 287518 23116 287527
rect 23060 287453 23116 287462
rect 28738 285159 28766 295445
rect 39682 293775 39710 299441
rect 41782 298801 41834 298807
rect 41780 298766 41782 298775
rect 41834 298766 41836 298775
rect 41780 298701 41836 298710
rect 41780 298248 41836 298257
rect 41780 298183 41782 298192
rect 41834 298183 41836 298192
rect 41782 298151 41834 298157
rect 41780 297730 41836 297739
rect 41780 297665 41782 297674
rect 41834 297665 41836 297674
rect 41782 297633 41834 297639
rect 41890 297295 41918 299631
rect 43234 298807 43262 341367
rect 43330 340543 43358 381549
rect 43522 342023 43550 384361
rect 43510 342017 43562 342023
rect 43510 341959 43562 341965
rect 43414 340907 43466 340913
rect 43414 340849 43466 340855
rect 43318 340537 43370 340543
rect 43318 340479 43370 340485
rect 43426 300953 43454 340849
rect 43606 339871 43658 339877
rect 43606 339813 43658 339819
rect 43414 300947 43466 300953
rect 43414 300889 43466 300895
rect 43222 298801 43274 298807
rect 43222 298743 43274 298749
rect 43414 298209 43466 298215
rect 43414 298151 43466 298157
rect 43222 297691 43274 297697
rect 43222 297633 43274 297639
rect 41876 297286 41932 297295
rect 41876 297221 41932 297230
rect 39862 296803 39914 296809
rect 39862 296745 39914 296751
rect 41780 296768 41836 296777
rect 39874 296555 39902 296745
rect 41780 296703 41782 296712
rect 41834 296703 41836 296712
rect 41782 296671 41834 296677
rect 39860 296546 39916 296555
rect 39860 296481 39916 296490
rect 39670 293769 39722 293775
rect 39670 293711 39722 293717
rect 41684 292994 41740 293003
rect 41684 292929 41740 292938
rect 41588 291070 41644 291079
rect 41588 291005 41644 291014
rect 41602 285191 41630 291005
rect 41698 288014 41726 292929
rect 42452 290774 42508 290783
rect 42452 290709 42508 290718
rect 42466 290612 42494 290709
rect 42466 290584 42590 290612
rect 41780 289812 41836 289821
rect 41780 289747 41836 289756
rect 41794 289409 41822 289747
rect 41782 289403 41834 289409
rect 41782 289345 41834 289351
rect 41780 289294 41836 289303
rect 41780 289229 41836 289238
rect 41794 288225 41822 289229
rect 41782 288219 41834 288225
rect 41782 288161 41834 288167
rect 41698 287986 41822 288014
rect 41590 285185 41642 285191
rect 28724 285150 28780 285159
rect 41590 285127 41642 285133
rect 28724 285085 28780 285094
rect 41794 283859 41822 287986
rect 41876 287814 41932 287823
rect 41876 287749 41878 287758
rect 41930 287749 41932 287758
rect 41878 287717 41930 287723
rect 41782 283853 41834 283859
rect 41782 283795 41834 283801
rect 41782 283557 41834 283563
rect 41782 283499 41834 283505
rect 41794 283050 41822 283499
rect 42562 282254 42590 290584
rect 43126 289403 43178 289409
rect 43126 289345 43178 289351
rect 42934 288219 42986 288225
rect 42934 288161 42986 288167
rect 42946 288014 42974 288161
rect 42946 287986 43070 288014
rect 42934 285185 42986 285191
rect 42934 285127 42986 285133
rect 42466 282226 42590 282254
rect 41876 281746 41932 281755
rect 41876 281681 41932 281690
rect 41890 281200 41918 281681
rect 42466 281607 42494 282226
rect 42452 281598 42508 281607
rect 42452 281533 42508 281542
rect 42082 280159 42110 280534
rect 42070 280153 42122 280159
rect 42070 280095 42122 280101
rect 42838 280153 42890 280159
rect 42838 280095 42890 280101
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42082 278531 42110 278721
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42070 278525 42122 278531
rect 42070 278467 42122 278473
rect 42178 278166 42206 278541
rect 41972 278046 42028 278055
rect 41972 277981 42028 277990
rect 41986 277500 42014 277981
rect 42070 277267 42122 277273
rect 42070 277209 42122 277215
rect 42082 276908 42110 277209
rect 42164 276566 42220 276575
rect 42164 276501 42220 276510
rect 42178 276316 42206 276501
rect 42850 276459 42878 280095
rect 42946 279937 42974 285127
rect 42934 279931 42986 279937
rect 42934 279873 42986 279879
rect 43042 278605 43070 287986
rect 43030 278599 43082 278605
rect 43030 278541 43082 278547
rect 42934 278525 42986 278531
rect 42934 278467 42986 278473
rect 42838 276453 42890 276459
rect 42838 276395 42890 276401
rect 41780 274198 41836 274207
rect 41780 274133 41836 274142
rect 41794 273845 41822 274133
rect 41780 273606 41836 273615
rect 42946 273573 42974 278467
rect 43138 277273 43166 289345
rect 43126 277267 43178 277273
rect 43126 277209 43178 277215
rect 41780 273541 41836 273550
rect 42934 273567 42986 273573
rect 41794 273208 41822 273541
rect 42934 273509 42986 273515
rect 41780 272866 41836 272875
rect 41780 272801 41836 272810
rect 41794 272542 41822 272801
rect 41780 272274 41836 272283
rect 41780 272209 41836 272218
rect 41794 272024 41822 272209
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 41794 270174 41822 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 42164 269314 42220 269323
rect 42164 269249 42220 269258
rect 42178 268877 42206 269249
rect 42166 268609 42218 268615
rect 42166 268551 42218 268557
rect 42178 268324 42206 268551
rect 23158 265057 23210 265063
rect 23158 264999 23210 265005
rect 23062 263577 23114 263583
rect 23062 263519 23114 263525
rect 23074 253339 23102 263519
rect 23170 253931 23198 264999
rect 43234 264915 43262 297633
rect 43318 296729 43370 296735
rect 43318 296671 43370 296677
rect 43330 264989 43358 296671
rect 43318 264983 43370 264989
rect 43318 264925 43370 264931
rect 43222 264909 43274 264915
rect 43222 264851 43274 264857
rect 23542 263651 23594 263657
rect 23542 263593 23594 263599
rect 23350 262171 23402 262177
rect 23350 262113 23402 262119
rect 23362 254819 23390 262113
rect 23348 254810 23404 254819
rect 23348 254745 23404 254754
rect 23554 253931 23582 263593
rect 43316 263394 43372 263403
rect 43316 263329 43372 263338
rect 43330 262177 43358 263329
rect 43318 262171 43370 262177
rect 43318 262113 43370 262119
rect 41588 256882 41644 256891
rect 41588 256817 41644 256826
rect 41602 256405 41630 256817
rect 41780 256586 41836 256595
rect 41780 256521 41836 256530
rect 41794 256479 41822 256521
rect 41782 256473 41834 256479
rect 41782 256415 41834 256421
rect 41590 256399 41642 256405
rect 41590 256341 41642 256347
rect 41782 256029 41834 256035
rect 41780 255994 41782 256003
rect 41834 255994 41836 256003
rect 41780 255929 41836 255938
rect 41782 255585 41834 255591
rect 41780 255550 41782 255559
rect 41834 255550 41836 255559
rect 41780 255485 41836 255494
rect 41780 255106 41836 255115
rect 41780 255041 41782 255050
rect 41834 255041 41836 255050
rect 41782 255009 41834 255015
rect 23156 253922 23212 253931
rect 23156 253857 23212 253866
rect 23540 253922 23596 253931
rect 23540 253857 23596 253866
rect 23060 253330 23116 253339
rect 23060 253265 23116 253274
rect 41780 250074 41836 250083
rect 41780 250009 41836 250018
rect 41492 247854 41548 247863
rect 41492 247789 41548 247798
rect 41506 244713 41534 247789
rect 41588 247410 41644 247419
rect 41588 247345 41644 247354
rect 41602 245527 41630 247345
rect 41684 245930 41740 245939
rect 41684 245865 41740 245874
rect 41590 245521 41642 245527
rect 41590 245463 41642 245469
rect 41698 245453 41726 245865
rect 41686 245447 41738 245453
rect 41686 245389 41738 245395
rect 41684 245338 41740 245347
rect 41684 245273 41740 245282
rect 41590 244929 41642 244935
rect 41588 244894 41590 244903
rect 41642 244894 41644 244903
rect 41698 244861 41726 245273
rect 41588 244829 41644 244838
rect 41686 244855 41738 244861
rect 41686 244797 41738 244803
rect 41494 244707 41546 244713
rect 41494 244649 41546 244655
rect 41588 244302 41644 244311
rect 41588 244237 41644 244246
rect 41602 242641 41630 244237
rect 41590 242635 41642 242641
rect 41590 242577 41642 242583
rect 41794 240643 41822 250009
rect 41876 246670 41932 246679
rect 41876 246605 41932 246614
rect 41890 245083 41918 246605
rect 43030 245521 43082 245527
rect 43030 245463 43082 245469
rect 42838 245447 42890 245453
rect 42838 245389 42890 245395
rect 41878 245077 41930 245083
rect 41878 245019 41930 245025
rect 42742 244707 42794 244713
rect 42742 244649 42794 244655
rect 41782 240637 41834 240643
rect 41782 240579 41834 240585
rect 41782 240415 41834 240421
rect 41782 240357 41834 240363
rect 41794 239834 41822 240357
rect 41794 237947 41822 237984
rect 41780 237938 41836 237947
rect 41780 237873 41836 237882
rect 42754 236721 42782 244649
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42742 236715 42794 236721
rect 42742 236657 42794 236663
rect 42178 236165 42206 236657
rect 42742 236567 42794 236573
rect 42742 236509 42794 236515
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42754 234649 42782 236509
rect 42850 235463 42878 245389
rect 42934 245077 42986 245083
rect 42934 245019 42986 245025
rect 42838 235457 42890 235463
rect 42838 235399 42890 235405
rect 42166 234643 42218 234649
rect 42166 234585 42218 234591
rect 42742 234643 42794 234649
rect 42742 234585 42794 234591
rect 42178 234325 42206 234585
rect 42946 234057 42974 245019
rect 43042 236573 43070 245463
rect 43030 236567 43082 236573
rect 43030 236509 43082 236515
rect 42070 234051 42122 234057
rect 42070 233993 42122 233999
rect 42934 234051 42986 234057
rect 42934 233993 42986 233999
rect 42082 233692 42110 233993
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 41780 231130 41836 231139
rect 41780 231065 41836 231074
rect 41794 230658 41822 231065
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 229992 41822 230325
rect 41780 229650 41836 229659
rect 41780 229585 41836 229594
rect 41794 229357 41822 229585
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41780 227430 41836 227439
rect 41780 227365 41836 227374
rect 41794 226958 41822 227365
rect 41876 226838 41932 226847
rect 41876 226773 41932 226782
rect 41890 226321 41918 226773
rect 41780 225950 41836 225959
rect 41780 225885 41836 225894
rect 41794 225700 41822 225885
rect 42082 221773 42110 225108
rect 42070 221767 42122 221773
rect 42070 221709 42122 221715
rect 41782 213701 41834 213707
rect 41780 213666 41782 213675
rect 41834 213666 41836 213675
rect 41780 213601 41836 213610
rect 41782 213183 41834 213189
rect 41780 213148 41782 213157
rect 41834 213148 41836 213157
rect 41780 213083 41836 213092
rect 41590 212813 41642 212819
rect 41588 212778 41590 212787
rect 41642 212778 41644 212787
rect 41588 212713 41644 212722
rect 41782 212221 41834 212227
rect 41780 212186 41782 212195
rect 41834 212186 41836 212195
rect 41780 212121 41836 212130
rect 41782 211703 41834 211709
rect 41780 211668 41782 211677
rect 41834 211668 41836 211677
rect 41780 211603 41836 211612
rect 41590 211333 41642 211339
rect 41588 211298 41590 211307
rect 41642 211298 41644 211307
rect 41588 211233 41644 211242
rect 43330 210747 43358 262113
rect 43426 255591 43454 298151
rect 43618 298141 43646 339813
rect 44278 300947 44330 300953
rect 44278 300889 44330 300895
rect 44290 299695 44318 300889
rect 44278 299689 44330 299695
rect 44278 299631 44330 299637
rect 43606 298135 43658 298141
rect 43606 298077 43658 298083
rect 43618 296809 43646 298077
rect 43606 296803 43658 296809
rect 43606 296745 43658 296751
rect 43508 267242 43564 267251
rect 43508 267177 43564 267186
rect 43522 265063 43550 267177
rect 43510 265057 43562 265063
rect 43510 264999 43562 265005
rect 43414 255585 43466 255591
rect 43414 255527 43466 255533
rect 43414 255067 43466 255073
rect 43414 255009 43466 255015
rect 43426 212227 43454 255009
rect 43414 212221 43466 212227
rect 43414 212163 43466 212169
rect 41782 210741 41834 210747
rect 41780 210706 41782 210715
rect 43318 210741 43370 210747
rect 41834 210706 41836 210715
rect 43318 210683 43370 210689
rect 41780 210641 41836 210650
rect 41782 210149 41834 210155
rect 41780 210114 41782 210123
rect 41834 210114 41836 210123
rect 41780 210049 41836 210058
rect 43522 209859 43550 264999
rect 44278 264983 44330 264989
rect 44278 264925 44330 264931
rect 44182 264909 44234 264915
rect 44182 264851 44234 264857
rect 44194 263657 44222 264851
rect 44182 263651 44234 263657
rect 44182 263593 44234 263599
rect 44290 263583 44318 264925
rect 44278 263577 44330 263583
rect 44278 263519 44330 263525
rect 44578 246267 44606 803719
rect 44674 267399 44702 813413
rect 44758 812583 44810 812589
rect 44758 812525 44810 812531
rect 44770 275391 44798 812525
rect 44866 785579 44894 816077
rect 44950 815395 45002 815401
rect 44950 815337 45002 815343
rect 44962 789131 44990 815337
rect 44950 789125 45002 789131
rect 44950 789067 45002 789073
rect 44854 785573 44906 785579
rect 44854 785515 44906 785521
rect 47458 785431 47486 816595
rect 57718 800743 57770 800749
rect 57718 800685 57770 800691
rect 57622 800669 57674 800675
rect 57622 800611 57674 800617
rect 57634 789691 57662 800611
rect 57730 790875 57758 800685
rect 57716 790866 57772 790875
rect 57716 790801 57772 790810
rect 57620 789682 57676 789691
rect 57620 789617 57676 789626
rect 58198 789199 58250 789205
rect 58198 789141 58250 789147
rect 58210 788507 58238 789141
rect 58390 789125 58442 789131
rect 58390 789067 58442 789073
rect 58196 788498 58252 788507
rect 58196 788433 58252 788442
rect 58402 787323 58430 789067
rect 58388 787314 58444 787323
rect 58388 787249 58444 787258
rect 59158 785573 59210 785579
rect 59158 785515 59210 785521
rect 59636 785538 59692 785547
rect 47446 785425 47498 785431
rect 47446 785367 47498 785373
rect 59170 784955 59198 785515
rect 59636 785473 59692 785482
rect 59650 785431 59678 785473
rect 59638 785425 59690 785431
rect 59638 785367 59690 785373
rect 59156 784946 59212 784955
rect 59156 784881 59212 784890
rect 47446 773511 47498 773517
rect 47446 773453 47498 773459
rect 44950 772919 45002 772925
rect 44950 772861 45002 772867
rect 44854 760783 44906 760789
rect 44854 760725 44906 760731
rect 44756 275382 44812 275391
rect 44756 275317 44812 275326
rect 44660 267390 44716 267399
rect 44660 267325 44716 267334
rect 44866 246341 44894 760725
rect 44962 742955 44990 772861
rect 45046 772327 45098 772333
rect 45046 772269 45098 772275
rect 45058 745397 45086 772269
rect 45046 745391 45098 745397
rect 45046 745333 45098 745339
rect 47458 743029 47486 773453
rect 61846 772179 61898 772185
rect 61846 772121 61898 772127
rect 58678 757527 58730 757533
rect 58678 757469 58730 757475
rect 58690 747659 58718 757469
rect 58676 747650 58732 747659
rect 58676 747585 58732 747594
rect 54740 746022 54796 746031
rect 54646 745983 54698 745989
rect 54740 745957 54742 745966
rect 54646 745925 54698 745931
rect 54794 745957 54796 745966
rect 57622 745983 57674 745989
rect 54742 745925 54794 745931
rect 57622 745925 57674 745931
rect 54658 745883 54686 745925
rect 54644 745874 54700 745883
rect 54644 745809 54700 745818
rect 57634 745291 57662 745925
rect 59636 745726 59692 745735
rect 59636 745661 59692 745670
rect 59650 745619 59678 745661
rect 59638 745613 59690 745619
rect 59638 745555 59690 745561
rect 58486 745391 58538 745397
rect 58486 745333 58538 745339
rect 57620 745282 57676 745291
rect 57620 745217 57676 745226
rect 58498 744107 58526 745333
rect 58484 744098 58540 744107
rect 58484 744033 58540 744042
rect 47446 743023 47498 743029
rect 47446 742965 47498 742971
rect 59638 743023 59690 743029
rect 59638 742965 59690 742971
rect 44950 742949 45002 742955
rect 59650 742923 59678 742965
rect 59734 742949 59786 742955
rect 44950 742891 45002 742897
rect 59636 742914 59692 742923
rect 59734 742891 59786 742897
rect 59636 742849 59692 742858
rect 59746 741739 59774 742891
rect 59732 741730 59788 741739
rect 59732 741665 59788 741674
rect 47542 730443 47594 730449
rect 47542 730385 47594 730391
rect 44950 729925 45002 729931
rect 44950 729867 45002 729873
rect 44962 699739 44990 729867
rect 45046 729407 45098 729413
rect 45046 729349 45098 729355
rect 45058 702625 45086 729349
rect 47446 717715 47498 717721
rect 47446 717657 47498 717663
rect 45046 702619 45098 702625
rect 45046 702561 45098 702567
rect 44950 699733 45002 699739
rect 44950 699675 45002 699681
rect 44950 683897 45002 683903
rect 44950 683839 45002 683845
rect 44962 266511 44990 683839
rect 45142 683009 45194 683015
rect 45142 682951 45194 682957
rect 45046 665323 45098 665329
rect 45046 665265 45098 665271
rect 45058 659409 45086 665265
rect 45046 659403 45098 659409
rect 45046 659345 45098 659351
rect 45046 596207 45098 596213
rect 45046 596149 45098 596155
rect 45058 278647 45086 596149
rect 45044 278638 45100 278647
rect 45044 278573 45100 278582
rect 44948 266502 45004 266511
rect 44948 266437 45004 266446
rect 45154 266363 45182 682951
rect 45908 658850 45964 658859
rect 45908 658785 45964 658794
rect 45922 655561 45950 658785
rect 45910 655555 45962 655561
rect 45910 655497 45962 655503
rect 45908 615634 45964 615643
rect 45908 615569 45964 615578
rect 45922 612419 45950 615569
rect 45910 612413 45962 612419
rect 45910 612355 45962 612361
rect 46196 572418 46252 572427
rect 46196 572353 46252 572362
rect 46210 569203 46238 572353
rect 46198 569197 46250 569203
rect 46198 569139 46250 569145
rect 46676 529350 46732 529359
rect 46676 529285 46732 529294
rect 46690 525987 46718 529285
rect 46678 525981 46730 525987
rect 46678 525923 46730 525929
rect 45334 427265 45386 427271
rect 45334 427207 45386 427213
rect 45236 426490 45292 426499
rect 45236 426425 45292 426434
rect 45250 273319 45278 426425
rect 45346 282453 45374 427207
rect 45526 420457 45578 420463
rect 45526 420399 45578 420405
rect 45430 383531 45482 383537
rect 45430 383473 45482 383479
rect 45334 282447 45386 282453
rect 45334 282389 45386 282395
rect 45334 279487 45386 279493
rect 45334 279429 45386 279435
rect 45236 273310 45292 273319
rect 45236 273245 45292 273254
rect 45140 266354 45196 266363
rect 45140 266289 45196 266298
rect 44854 246335 44906 246341
rect 44854 246277 44906 246283
rect 44566 246261 44618 246267
rect 44566 246203 44618 246209
rect 44662 245003 44714 245009
rect 44662 244945 44714 244951
rect 44566 242709 44618 242715
rect 44566 242651 44618 242657
rect 41590 209853 41642 209859
rect 41588 209818 41590 209827
rect 43510 209853 43562 209859
rect 41642 209818 41644 209827
rect 43510 209795 43562 209801
rect 41588 209753 41644 209762
rect 25652 208930 25708 208939
rect 25652 208865 25708 208874
rect 25556 207894 25612 207903
rect 25556 207829 25612 207838
rect 25570 200059 25598 207829
rect 25666 200947 25694 208865
rect 25844 208338 25900 208347
rect 25844 208273 25900 208282
rect 25748 206858 25804 206867
rect 25748 206793 25804 206802
rect 25652 200938 25708 200947
rect 25652 200873 25708 200882
rect 25556 200050 25612 200059
rect 25556 199985 25612 199994
rect 25762 199763 25790 206793
rect 25858 200947 25886 208273
rect 34292 207450 34348 207459
rect 34292 207385 34348 207394
rect 34306 201539 34334 207385
rect 41876 206636 41932 206645
rect 41876 206571 41932 206580
rect 41588 204342 41644 204351
rect 41588 204277 41644 204286
rect 34292 201530 34348 201539
rect 34292 201465 34348 201474
rect 25844 200938 25900 200947
rect 25844 200873 25900 200882
rect 25748 199754 25804 199763
rect 25748 199689 25804 199698
rect 41602 198907 41630 204277
rect 41780 204194 41836 204203
rect 41780 204129 41836 204138
rect 41794 203347 41822 204129
rect 41782 203341 41834 203347
rect 41782 203283 41834 203289
rect 41780 203232 41836 203241
rect 41780 203167 41836 203176
rect 41794 202829 41822 203167
rect 41782 202823 41834 202829
rect 41782 202765 41834 202771
rect 41780 202714 41836 202723
rect 41780 202649 41836 202658
rect 41794 201645 41822 202649
rect 41782 201639 41834 201645
rect 41782 201581 41834 201587
rect 41782 201269 41834 201275
rect 41780 201234 41782 201243
rect 41834 201234 41836 201243
rect 41780 201169 41836 201178
rect 41590 198901 41642 198907
rect 41590 198843 41642 198849
rect 41890 197427 41918 206571
rect 43030 203341 43082 203347
rect 43030 203283 43082 203289
rect 42934 202823 42986 202829
rect 42934 202765 42986 202771
rect 41974 202157 42026 202163
rect 41972 202122 41974 202131
rect 42026 202122 42028 202131
rect 41972 202057 42028 202066
rect 41974 201713 42026 201719
rect 41972 201678 41974 201687
rect 42026 201678 42028 201687
rect 41972 201613 42028 201622
rect 42742 201639 42794 201645
rect 42742 201581 42794 201587
rect 41878 197421 41930 197427
rect 41878 197363 41930 197369
rect 41878 197199 41930 197205
rect 41878 197141 41930 197147
rect 41890 196618 41918 197141
rect 41780 195314 41836 195323
rect 41780 195249 41836 195258
rect 41794 194805 41822 195249
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42754 192247 42782 201581
rect 42838 198901 42890 198907
rect 42838 198843 42890 198849
rect 42850 193505 42878 198843
rect 42838 193499 42890 193505
rect 42838 193441 42890 193447
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42742 192241 42794 192247
rect 42742 192183 42794 192189
rect 42178 191769 42206 192183
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42082 191142 42110 191443
rect 42946 191063 42974 202765
rect 43042 191507 43070 203283
rect 44578 201275 44606 242651
rect 44674 202163 44702 244945
rect 44758 242857 44810 242863
rect 44758 242799 44810 242805
rect 44662 202157 44714 202163
rect 44662 202099 44714 202105
rect 44770 201719 44798 242799
rect 44854 242783 44906 242789
rect 44854 242725 44906 242731
rect 44866 211709 44894 242725
rect 45346 213707 45374 279429
rect 45442 270655 45470 383473
rect 45538 307835 45566 420399
rect 45622 377241 45674 377247
rect 45622 377183 45674 377189
rect 45634 339951 45662 377183
rect 45718 340537 45770 340543
rect 45718 340479 45770 340485
rect 45622 339945 45674 339951
rect 45622 339887 45674 339893
rect 45526 307829 45578 307835
rect 45526 307771 45578 307777
rect 45526 282373 45578 282379
rect 45526 282315 45578 282321
rect 45428 270646 45484 270655
rect 45428 270581 45484 270590
rect 45334 213701 45386 213707
rect 45334 213643 45386 213649
rect 45538 212819 45566 282315
rect 45622 279413 45674 279419
rect 45622 279355 45674 279361
rect 45634 213189 45662 279355
rect 45730 276279 45758 340479
rect 46102 307829 46154 307835
rect 46102 307771 46154 307777
rect 46114 302359 46142 307771
rect 46102 302353 46154 302359
rect 46102 302295 46154 302301
rect 45814 287775 45866 287781
rect 45814 287717 45866 287723
rect 45716 276270 45772 276279
rect 45716 276205 45772 276214
rect 45826 246415 45854 287717
rect 47458 246489 47486 717657
rect 47554 699813 47582 730385
rect 59638 714311 59690 714317
rect 59638 714253 59690 714259
rect 59650 704443 59678 714253
rect 59636 704434 59692 704443
rect 59636 704369 59692 704378
rect 58774 702693 58826 702699
rect 58772 702658 58774 702667
rect 58826 702658 58828 702667
rect 58678 702619 58730 702625
rect 58772 702593 58828 702602
rect 58678 702561 58730 702567
rect 58690 700891 58718 702561
rect 58676 700882 58732 700891
rect 58676 700817 58732 700826
rect 47542 699807 47594 699813
rect 47542 699749 47594 699755
rect 59254 699807 59306 699813
rect 59254 699749 59306 699755
rect 58870 699733 58922 699739
rect 59266 699707 59294 699749
rect 58870 699675 58922 699681
rect 59252 699698 59308 699707
rect 58882 698523 58910 699675
rect 59252 699633 59308 699642
rect 58868 698514 58924 698523
rect 58868 698449 58924 698458
rect 50326 686857 50378 686863
rect 50326 686799 50378 686805
rect 47638 686339 47690 686345
rect 47638 686281 47690 686287
rect 47542 674055 47594 674061
rect 47542 673997 47594 674003
rect 47554 246637 47582 673997
rect 47650 656597 47678 686281
rect 47734 685599 47786 685605
rect 47734 685541 47786 685547
rect 47746 659483 47774 685541
rect 47734 659477 47786 659483
rect 47734 659419 47786 659425
rect 50338 656671 50366 686799
rect 59638 671095 59690 671101
rect 59638 671037 59690 671043
rect 59650 661227 59678 671037
rect 59636 661218 59692 661227
rect 59636 661153 59692 661162
rect 59158 659477 59210 659483
rect 58772 659442 58828 659451
rect 59158 659419 59210 659425
rect 58772 659377 58774 659386
rect 58826 659377 58828 659386
rect 58774 659345 58826 659351
rect 59170 657675 59198 659419
rect 59156 657666 59212 657675
rect 59156 657601 59212 657610
rect 50326 656665 50378 656671
rect 50326 656607 50378 656613
rect 58198 656665 58250 656671
rect 58198 656607 58250 656613
rect 47638 656591 47690 656597
rect 47638 656533 47690 656539
rect 58210 656491 58238 656607
rect 58390 656591 58442 656597
rect 58390 656533 58442 656539
rect 58196 656482 58252 656491
rect 58196 656417 58252 656426
rect 58402 655307 58430 656533
rect 58388 655298 58444 655307
rect 58388 655233 58444 655242
rect 50326 643715 50378 643721
rect 50326 643657 50378 643663
rect 47734 643123 47786 643129
rect 47734 643065 47786 643071
rect 47638 630839 47690 630845
rect 47638 630781 47690 630787
rect 47542 246631 47594 246637
rect 47542 246573 47594 246579
rect 47650 246563 47678 630781
rect 47746 613381 47774 643065
rect 47830 642383 47882 642389
rect 47830 642325 47882 642331
rect 47842 616341 47870 642325
rect 47926 622107 47978 622113
rect 47926 622049 47978 622055
rect 47830 616335 47882 616341
rect 47830 616277 47882 616283
rect 47938 616267 47966 622049
rect 47926 616261 47978 616267
rect 47926 616203 47978 616209
rect 50338 613455 50366 643657
rect 58966 624327 59018 624333
rect 58966 624269 59018 624275
rect 58978 618011 59006 624269
rect 58964 618002 59020 618011
rect 58964 617937 59020 617946
rect 58966 616335 59018 616341
rect 58966 616277 59018 616283
rect 58978 614459 59006 616277
rect 59638 616261 59690 616267
rect 59636 616226 59638 616235
rect 59690 616226 59692 616235
rect 59636 616161 59692 616170
rect 58964 614450 59020 614459
rect 58964 614385 59020 614394
rect 50326 613449 50378 613455
rect 50326 613391 50378 613397
rect 59638 613449 59690 613455
rect 59638 613391 59690 613397
rect 47734 613375 47786 613381
rect 47734 613317 47786 613323
rect 59542 613375 59594 613381
rect 59542 613317 59594 613323
rect 59554 612091 59582 613317
rect 59650 613275 59678 613391
rect 59636 613266 59692 613275
rect 59636 613201 59692 613210
rect 59540 612082 59596 612091
rect 59540 612017 59596 612026
rect 50326 600499 50378 600505
rect 50326 600441 50378 600447
rect 47830 599759 47882 599765
rect 47830 599701 47882 599707
rect 47734 587623 47786 587629
rect 47734 587565 47786 587571
rect 47746 249153 47774 587565
rect 47842 570165 47870 599701
rect 47926 599389 47978 599395
rect 47926 599331 47978 599337
rect 47938 573125 47966 599331
rect 48022 578965 48074 578971
rect 48022 578907 48074 578913
rect 47926 573119 47978 573125
rect 47926 573061 47978 573067
rect 48034 573051 48062 578907
rect 48022 573045 48074 573051
rect 48022 572987 48074 572993
rect 50338 570239 50366 600441
rect 58966 580889 59018 580895
rect 58966 580831 59018 580837
rect 58978 574795 59006 580831
rect 58964 574786 59020 574795
rect 58964 574721 59020 574730
rect 58966 573119 59018 573125
rect 58966 573061 59018 573067
rect 58978 571243 59006 573061
rect 59638 573045 59690 573051
rect 59636 573010 59638 573019
rect 59690 573010 59692 573019
rect 59636 572945 59692 572954
rect 58964 571234 59020 571243
rect 58964 571169 59020 571178
rect 50326 570233 50378 570239
rect 50326 570175 50378 570181
rect 59350 570233 59402 570239
rect 59350 570175 59402 570181
rect 47830 570159 47882 570165
rect 47830 570101 47882 570107
rect 59362 570059 59390 570175
rect 59542 570159 59594 570165
rect 59542 570101 59594 570107
rect 59348 570050 59404 570059
rect 59348 569985 59404 569994
rect 59554 568875 59582 570101
rect 59540 568866 59596 568875
rect 59540 568801 59596 568810
rect 50518 543075 50570 543081
rect 50518 543017 50570 543023
rect 48790 542705 48842 542711
rect 48790 542647 48842 542653
rect 48802 525025 48830 542647
rect 48886 542187 48938 542193
rect 48886 542129 48938 542135
rect 48898 527541 48926 542129
rect 48886 527535 48938 527541
rect 48886 527477 48938 527483
rect 48790 525019 48842 525025
rect 48790 524961 48842 524967
rect 50530 524729 50558 543017
rect 57718 541595 57770 541601
rect 57718 541537 57770 541543
rect 57622 541521 57674 541527
rect 57622 541463 57674 541469
rect 57634 530543 57662 541463
rect 57730 531727 57758 541537
rect 57716 531718 57772 531727
rect 57716 531653 57772 531662
rect 57620 530534 57676 530543
rect 57620 530469 57676 530478
rect 59636 527574 59692 527583
rect 59636 527509 59638 527518
rect 59690 527509 59692 527518
rect 59638 527477 59690 527483
rect 59348 525946 59404 525955
rect 59348 525881 59404 525890
rect 59362 524729 59390 525881
rect 59636 525058 59692 525067
rect 59636 524993 59638 525002
rect 59690 524993 59692 525002
rect 59638 524961 59690 524967
rect 50518 524723 50570 524729
rect 50518 524665 50570 524671
rect 59350 524723 59402 524729
rect 59350 524665 59402 524671
rect 47830 524279 47882 524285
rect 47830 524221 47882 524227
rect 47842 263551 47870 524221
rect 53206 429263 53258 429269
rect 53206 429205 53258 429211
rect 50326 428967 50378 428973
rect 50326 428909 50378 428915
rect 48022 428375 48074 428381
rect 48022 428317 48074 428323
rect 47926 416979 47978 416985
rect 47926 416921 47978 416927
rect 47828 263542 47884 263551
rect 47828 263477 47884 263486
rect 47938 254999 47966 416921
rect 48034 400187 48062 428317
rect 50338 400261 50366 428909
rect 53218 400335 53246 429205
rect 58486 406101 58538 406107
rect 58486 406043 58538 406049
rect 58498 404151 58526 406043
rect 58484 404142 58540 404151
rect 58484 404077 58540 404086
rect 59350 402623 59402 402629
rect 59350 402565 59402 402571
rect 59362 402375 59390 402565
rect 59348 402366 59404 402375
rect 59348 402301 59404 402310
rect 57716 400590 57772 400599
rect 57716 400525 57772 400534
rect 53206 400329 53258 400335
rect 53206 400271 53258 400277
rect 50326 400255 50378 400261
rect 50326 400197 50378 400203
rect 48022 400181 48074 400187
rect 48022 400123 48074 400129
rect 57730 394563 57758 400525
rect 59734 400329 59786 400335
rect 59734 400271 59786 400277
rect 59542 400255 59594 400261
rect 59542 400197 59594 400203
rect 59554 398231 59582 400197
rect 59638 400181 59690 400187
rect 59638 400123 59690 400129
rect 59650 400007 59678 400123
rect 59636 399998 59692 400007
rect 59636 399933 59692 399942
rect 59746 399415 59774 400271
rect 59732 399406 59788 399415
rect 59732 399341 59788 399350
rect 59540 398222 59596 398231
rect 59540 398157 59596 398166
rect 57718 394557 57770 394563
rect 57718 394499 57770 394505
rect 53206 386491 53258 386497
rect 53206 386433 53258 386439
rect 50326 385751 50378 385757
rect 50326 385693 50378 385699
rect 48118 385381 48170 385387
rect 48118 385323 48170 385329
rect 48022 373911 48074 373917
rect 48022 373853 48074 373859
rect 47926 254993 47978 254999
rect 47926 254935 47978 254941
rect 48034 254925 48062 373853
rect 48130 356971 48158 385323
rect 50338 357045 50366 385693
rect 53218 357119 53246 386433
rect 58486 361479 58538 361485
rect 58486 361421 58538 361427
rect 58498 360935 58526 361421
rect 58484 360926 58540 360935
rect 58484 360861 58540 360870
rect 59158 359999 59210 360005
rect 59158 359941 59210 359947
rect 59170 359751 59198 359941
rect 59156 359742 59212 359751
rect 59156 359677 59212 359686
rect 57716 357522 57772 357531
rect 57716 357457 57772 357466
rect 53206 357113 53258 357119
rect 53206 357055 53258 357061
rect 50326 357039 50378 357045
rect 50326 356981 50378 356987
rect 48118 356965 48170 356971
rect 48118 356907 48170 356913
rect 57730 351347 57758 357457
rect 58390 357113 58442 357119
rect 58390 357055 58442 357061
rect 58402 356199 58430 357055
rect 58486 357039 58538 357045
rect 58486 356981 58538 356987
rect 58388 356190 58444 356199
rect 58388 356125 58444 356134
rect 58498 355015 58526 356981
rect 59638 356965 59690 356971
rect 59638 356907 59690 356913
rect 59650 356791 59678 356907
rect 59636 356782 59692 356791
rect 59636 356717 59692 356726
rect 58484 355006 58540 355015
rect 58484 354941 58540 354950
rect 57718 351341 57770 351347
rect 57718 351283 57770 351289
rect 53206 343275 53258 343281
rect 53206 343217 53258 343223
rect 50326 342905 50378 342911
rect 50326 342847 50378 342853
rect 48118 342387 48170 342393
rect 48118 342329 48170 342335
rect 48130 313755 48158 342329
rect 48214 330991 48266 330997
rect 48214 330933 48266 330939
rect 48118 313749 48170 313755
rect 48118 313691 48170 313697
rect 48118 282299 48170 282305
rect 48118 282241 48170 282247
rect 48022 254919 48074 254925
rect 48022 254861 48074 254867
rect 47734 249147 47786 249153
rect 47734 249089 47786 249095
rect 47638 246557 47690 246563
rect 47638 246499 47690 246505
rect 47446 246483 47498 246489
rect 47446 246425 47498 246431
rect 45814 246409 45866 246415
rect 45814 246351 45866 246357
rect 45622 213183 45674 213189
rect 45622 213125 45674 213131
rect 45526 212813 45578 212819
rect 45526 212755 45578 212761
rect 44854 211703 44906 211709
rect 44854 211645 44906 211651
rect 44758 201713 44810 201719
rect 44758 201655 44810 201661
rect 44566 201269 44618 201275
rect 44566 201211 44618 201217
rect 43030 191501 43082 191507
rect 43030 191443 43082 191449
rect 42166 191057 42218 191063
rect 42166 190999 42218 191005
rect 42934 191057 42986 191063
rect 42934 190999 42986 191005
rect 42178 190476 42206 190999
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 41876 187914 41932 187923
rect 41876 187849 41932 187858
rect 41890 187442 41918 187849
rect 41780 187174 41836 187183
rect 41780 187109 41836 187118
rect 41794 186776 41822 187109
rect 41780 186730 41836 186739
rect 41780 186665 41836 186674
rect 41794 186184 41822 186665
rect 41780 185842 41836 185851
rect 41780 185777 41836 185786
rect 41794 185592 41822 185777
rect 42164 184214 42220 184223
rect 42164 184149 42220 184158
rect 42178 183742 42206 184149
rect 41876 183622 41932 183631
rect 41876 183557 41932 183566
rect 41890 183121 41918 183557
rect 42068 182882 42124 182891
rect 42068 182817 42124 182826
rect 42082 182484 42110 182817
rect 48130 182257 48158 282241
rect 48226 249227 48254 330933
rect 50338 313829 50366 342847
rect 53218 313903 53246 343217
rect 58486 319669 58538 319675
rect 58486 319611 58538 319617
rect 58498 317719 58526 319611
rect 58484 317710 58540 317719
rect 58484 317645 58540 317654
rect 59158 316783 59210 316789
rect 59158 316725 59210 316731
rect 59170 316535 59198 316725
rect 59156 316526 59212 316535
rect 59156 316461 59212 316470
rect 59060 314158 59116 314167
rect 59060 314093 59116 314102
rect 53206 313897 53258 313903
rect 53206 313839 53258 313845
rect 50326 313823 50378 313829
rect 50326 313765 50378 313771
rect 59074 308131 59102 314093
rect 59734 313897 59786 313903
rect 59734 313839 59786 313845
rect 59542 313823 59594 313829
rect 59542 313765 59594 313771
rect 59554 311799 59582 313765
rect 59638 313749 59690 313755
rect 59638 313691 59690 313697
rect 59650 313575 59678 313691
rect 59636 313566 59692 313575
rect 59636 313501 59692 313510
rect 59746 312983 59774 313839
rect 59732 312974 59788 312983
rect 59732 312909 59788 312918
rect 59540 311790 59596 311799
rect 59540 311725 59596 311734
rect 59062 308125 59114 308131
rect 59062 308067 59114 308073
rect 54646 302353 54698 302359
rect 54646 302295 54698 302301
rect 50710 299763 50762 299769
rect 50710 299705 50762 299711
rect 48310 291031 48362 291037
rect 48310 290973 48362 290979
rect 48322 268615 48350 290973
rect 50722 288965 50750 299705
rect 53302 293917 53354 293923
rect 53302 293859 53354 293865
rect 50710 288959 50762 288965
rect 50710 288901 50762 288907
rect 50326 288071 50378 288077
rect 50326 288013 50378 288019
rect 48310 268609 48362 268615
rect 48310 268551 48362 268557
rect 48214 249221 48266 249227
rect 48214 249163 48266 249169
rect 50338 221773 50366 288013
rect 53206 285185 53258 285191
rect 53206 285127 53258 285133
rect 53014 282447 53066 282453
rect 53014 282389 53066 282395
rect 53026 278013 53054 282389
rect 53014 278007 53066 278013
rect 53014 277949 53066 277955
rect 50612 275234 50668 275243
rect 50612 275169 50668 275178
rect 50420 275086 50476 275095
rect 50420 275021 50476 275030
rect 50326 221767 50378 221773
rect 50326 221709 50378 221715
rect 50434 210155 50462 275021
rect 50626 211339 50654 275169
rect 53218 256035 53246 285127
rect 53314 276459 53342 293859
rect 54658 290963 54686 302295
rect 60214 299615 60266 299621
rect 60214 299557 60266 299563
rect 59252 295214 59308 295223
rect 59252 295149 59308 295158
rect 59266 293923 59294 295149
rect 59254 293917 59306 293923
rect 59254 293859 59306 293865
rect 56182 293843 56234 293849
rect 56182 293785 56234 293791
rect 54646 290957 54698 290963
rect 54646 290899 54698 290905
rect 56086 282447 56138 282453
rect 56086 282389 56138 282395
rect 53302 276453 53354 276459
rect 53302 276395 53354 276401
rect 56098 256479 56126 282389
rect 56194 273573 56222 293785
rect 58198 293769 58250 293775
rect 58198 293711 58250 293717
rect 58210 292707 58238 293711
rect 59636 292846 59692 292855
rect 59636 292781 59692 292790
rect 58196 292698 58252 292707
rect 58196 292633 58252 292642
rect 59650 291037 59678 292781
rect 60226 291523 60254 299557
rect 60308 294030 60364 294039
rect 60308 293965 60364 293974
rect 60322 293849 60350 293965
rect 60310 293843 60362 293849
rect 60310 293785 60362 293791
rect 60212 291514 60268 291523
rect 60212 291449 60268 291458
rect 59638 291031 59690 291037
rect 59638 290973 59690 290979
rect 58774 290883 58826 290889
rect 58774 290825 58826 290831
rect 57620 284558 57676 284567
rect 57620 284493 57676 284502
rect 57634 282453 57662 284493
rect 58580 283374 58636 283383
rect 58580 283309 58636 283318
rect 57622 282447 57674 282453
rect 57622 282389 57674 282395
rect 58594 282305 58622 283309
rect 58786 282305 58814 290825
rect 59540 289294 59596 289303
rect 59540 289229 59596 289238
rect 59554 288965 59582 289229
rect 59542 288959 59594 288965
rect 59542 288901 59594 288907
rect 59156 288110 59212 288119
rect 59156 288045 59158 288054
rect 59210 288045 59212 288054
rect 59158 288013 59210 288019
rect 59252 286926 59308 286935
rect 59252 286861 59308 286870
rect 58964 285742 59020 285751
rect 58964 285677 59020 285686
rect 58582 282299 58634 282305
rect 58582 282241 58634 282247
rect 58774 282299 58826 282305
rect 58774 282241 58826 282247
rect 58388 281006 58444 281015
rect 58388 280941 58444 280950
rect 58402 279493 58430 280941
rect 58580 279822 58636 279831
rect 58580 279757 58636 279766
rect 58390 279487 58442 279493
rect 58390 279429 58442 279435
rect 58594 279419 58622 279757
rect 58582 279413 58634 279419
rect 58582 279355 58634 279361
rect 56182 273567 56234 273573
rect 56182 273509 56234 273515
rect 56086 256473 56138 256479
rect 56086 256415 56138 256421
rect 58978 256405 59006 285677
rect 59266 285191 59294 286861
rect 59254 285185 59306 285191
rect 59254 285127 59306 285133
rect 59636 282486 59692 282495
rect 59636 282421 59692 282430
rect 59650 282379 59678 282421
rect 59638 282373 59690 282379
rect 59638 282315 59690 282321
rect 61858 266807 61886 772121
rect 62038 771957 62090 771963
rect 62038 771899 62090 771905
rect 61942 642605 61994 642611
rect 61942 642547 61994 642553
rect 61954 278499 61982 642547
rect 61940 278490 61996 278499
rect 61940 278425 61996 278434
rect 62050 266955 62078 771899
rect 62230 728963 62282 728969
rect 62230 728905 62282 728911
rect 62134 642531 62186 642537
rect 62134 642473 62186 642479
rect 62146 278351 62174 642473
rect 62132 278342 62188 278351
rect 62132 278277 62188 278286
rect 62036 266946 62092 266955
rect 62036 266881 62092 266890
rect 61844 266798 61900 266807
rect 61844 266733 61900 266742
rect 62242 266659 62270 728905
rect 62422 728741 62474 728747
rect 62422 728683 62474 728689
rect 62324 602166 62380 602175
rect 62324 602101 62380 602110
rect 62338 278203 62366 602101
rect 62324 278194 62380 278203
rect 62324 278129 62380 278138
rect 62434 267103 62462 728683
rect 62516 547258 62572 547267
rect 62516 547193 62572 547202
rect 62530 273467 62558 547193
rect 62708 544446 62764 544455
rect 62708 544381 62764 544390
rect 62614 339945 62666 339951
rect 62614 339887 62666 339893
rect 62626 278055 62654 339887
rect 62612 278046 62668 278055
rect 62612 277981 62668 277990
rect 62722 273615 62750 544381
rect 62902 300947 62954 300953
rect 62902 300889 62954 300895
rect 62914 277907 62942 300889
rect 62998 298135 63050 298141
rect 62998 298077 63050 298083
rect 62900 277898 62956 277907
rect 62900 277833 62956 277842
rect 63010 277759 63038 298077
rect 63382 282225 63434 282231
rect 63382 282167 63434 282173
rect 63394 277939 63422 282167
rect 314902 278377 314954 278383
rect 314902 278319 314954 278325
rect 408310 278377 408362 278383
rect 408362 278325 408624 278328
rect 408310 278319 408624 278325
rect 63382 277933 63434 277939
rect 63382 277875 63434 277881
rect 62996 277750 63052 277759
rect 62996 277685 63052 277694
rect 62708 273606 62764 273615
rect 62708 273541 62764 273550
rect 62516 273458 62572 273467
rect 62516 273393 62572 273402
rect 65890 272167 65918 278018
rect 65878 272161 65930 272167
rect 65878 272103 65930 272109
rect 67042 269471 67070 278018
rect 68290 273277 68318 278018
rect 68278 273271 68330 273277
rect 68278 273213 68330 273219
rect 69442 269619 69470 278018
rect 70594 272135 70622 278018
rect 70580 272126 70636 272135
rect 70580 272061 70636 272070
rect 69428 269610 69484 269619
rect 69428 269545 69484 269554
rect 67028 269462 67084 269471
rect 67028 269397 67084 269406
rect 71746 269323 71774 278018
rect 72994 272283 73022 278018
rect 72980 272274 73036 272283
rect 72980 272209 73036 272218
rect 71732 269314 71788 269323
rect 74146 269281 74174 278018
rect 75298 271649 75326 278018
rect 75286 271643 75338 271649
rect 75286 271585 75338 271591
rect 76546 271205 76574 278018
rect 77698 276494 77726 278018
rect 77602 276466 77726 276494
rect 76534 271199 76586 271205
rect 76534 271141 76586 271147
rect 77602 269767 77630 276466
rect 78850 272431 78878 278018
rect 80112 278004 80606 278032
rect 78836 272422 78892 272431
rect 78836 272357 78892 272366
rect 77686 271643 77738 271649
rect 77686 271585 77738 271591
rect 77588 269758 77644 269767
rect 77588 269693 77644 269702
rect 71732 269249 71788 269258
rect 74134 269275 74186 269281
rect 74134 269217 74186 269223
rect 62420 267094 62476 267103
rect 62420 267029 62476 267038
rect 62228 266650 62284 266659
rect 62228 266585 62284 266594
rect 58966 256399 59018 256405
rect 58966 256341 59018 256347
rect 53206 256029 53258 256035
rect 53206 255971 53258 255977
rect 77698 249301 77726 271585
rect 80578 249375 80606 278004
rect 81250 269355 81278 278018
rect 82402 269429 82430 278018
rect 83650 269577 83678 278018
rect 84802 272315 84830 278018
rect 84790 272309 84842 272315
rect 84790 272251 84842 272257
rect 85954 271057 85982 278018
rect 86326 272309 86378 272315
rect 86326 272251 86378 272257
rect 85942 271051 85994 271057
rect 85942 270993 85994 270999
rect 83638 269571 83690 269577
rect 83638 269513 83690 269519
rect 82390 269423 82442 269429
rect 82390 269365 82442 269371
rect 81238 269349 81290 269355
rect 81238 269291 81290 269297
rect 86338 252187 86366 272251
rect 87202 269503 87230 278018
rect 88354 272579 88382 278018
rect 88340 272570 88396 272579
rect 88340 272505 88396 272514
rect 89506 271575 89534 278018
rect 89494 271569 89546 271575
rect 89494 271511 89546 271517
rect 90658 269651 90686 278018
rect 91906 272727 91934 278018
rect 91892 272718 91948 272727
rect 91892 272653 91948 272662
rect 92086 271569 92138 271575
rect 92086 271511 92138 271517
rect 90646 269645 90698 269651
rect 90646 269587 90698 269593
rect 87190 269497 87242 269503
rect 87190 269439 87242 269445
rect 86326 252181 86378 252187
rect 86326 252123 86378 252129
rect 92098 252039 92126 271511
rect 93058 269725 93086 278018
rect 94210 270761 94238 278018
rect 94198 270755 94250 270761
rect 94198 270697 94250 270703
rect 94966 270755 95018 270761
rect 94966 270697 95018 270703
rect 93046 269719 93098 269725
rect 93046 269661 93098 269667
rect 94978 252113 95006 270697
rect 95458 269799 95486 278018
rect 96610 272389 96638 278018
rect 97776 278004 97886 278032
rect 96598 272383 96650 272389
rect 96598 272325 96650 272331
rect 95446 269793 95498 269799
rect 95446 269735 95498 269741
rect 97858 252409 97886 278004
rect 99010 272463 99038 278018
rect 98998 272457 99050 272463
rect 98998 272399 99050 272405
rect 100162 269873 100190 278018
rect 101314 271797 101342 278018
rect 101302 271791 101354 271797
rect 101302 271733 101354 271739
rect 102562 269947 102590 278018
rect 103714 272537 103742 278018
rect 103702 272531 103754 272537
rect 103702 272473 103754 272479
rect 104866 272315 104894 278018
rect 106114 272611 106142 278018
rect 106102 272605 106154 272611
rect 106102 272547 106154 272553
rect 104854 272309 104906 272315
rect 104854 272251 104906 272257
rect 106486 272309 106538 272315
rect 106486 272251 106538 272257
rect 103606 271791 103658 271797
rect 103606 271733 103658 271739
rect 102550 269941 102602 269947
rect 102550 269883 102602 269889
rect 100150 269867 100202 269873
rect 100150 269809 100202 269815
rect 97846 252403 97898 252409
rect 97846 252345 97898 252351
rect 103618 252335 103646 271733
rect 106498 252483 106526 272251
rect 107266 270021 107294 278018
rect 108418 270761 108446 278018
rect 108406 270755 108458 270761
rect 108406 270697 108458 270703
rect 109366 270755 109418 270761
rect 109366 270697 109418 270703
rect 107254 270015 107306 270021
rect 107254 269957 107306 269963
rect 106486 252477 106538 252483
rect 106486 252419 106538 252425
rect 103606 252329 103658 252335
rect 103606 252271 103658 252277
rect 109378 252261 109406 270697
rect 109570 270095 109598 278018
rect 110818 272685 110846 278018
rect 111984 278004 112286 278032
rect 110806 272679 110858 272685
rect 110806 272621 110858 272627
rect 109558 270089 109610 270095
rect 109558 270031 109610 270037
rect 109366 252255 109418 252261
rect 109366 252197 109418 252203
rect 94966 252107 95018 252113
rect 94966 252049 95018 252055
rect 92086 252033 92138 252039
rect 92086 251975 92138 251981
rect 80566 249369 80618 249375
rect 80566 249311 80618 249317
rect 77686 249295 77738 249301
rect 77686 249237 77738 249243
rect 112258 246711 112286 278004
rect 113122 272759 113150 278018
rect 113110 272753 113162 272759
rect 113110 272695 113162 272701
rect 114370 270243 114398 278018
rect 115522 271723 115550 278018
rect 116674 272907 116702 278018
rect 116662 272901 116714 272907
rect 116662 272843 116714 272849
rect 115510 271717 115562 271723
rect 115510 271659 115562 271665
rect 114358 270237 114410 270243
rect 114358 270179 114410 270185
rect 117922 270169 117950 278018
rect 118006 271717 118058 271723
rect 118006 271659 118058 271665
rect 117910 270163 117962 270169
rect 117910 270105 117962 270111
rect 118018 249671 118046 271659
rect 119074 270761 119102 278018
rect 120226 272833 120254 278018
rect 120214 272827 120266 272833
rect 120214 272769 120266 272775
rect 119062 270755 119114 270761
rect 119062 270697 119114 270703
rect 120886 270755 120938 270761
rect 120886 270697 120938 270703
rect 120898 249893 120926 270697
rect 121474 270317 121502 278018
rect 122626 270761 122654 278018
rect 123778 272981 123806 278018
rect 123766 272975 123818 272981
rect 123766 272917 123818 272923
rect 122614 270755 122666 270761
rect 122614 270697 122666 270703
rect 123766 270755 123818 270761
rect 123766 270697 123818 270703
rect 121462 270311 121514 270317
rect 121462 270253 121514 270259
rect 120886 249887 120938 249893
rect 120886 249829 120938 249835
rect 118006 249665 118058 249671
rect 118006 249607 118058 249613
rect 123778 249449 123806 270697
rect 125026 270391 125054 278018
rect 126192 278004 126686 278032
rect 125014 270385 125066 270391
rect 125014 270327 125066 270333
rect 126658 249523 126686 278004
rect 127330 273129 127358 278018
rect 127318 273123 127370 273129
rect 127318 273065 127370 273071
rect 128482 273055 128510 278018
rect 128470 273049 128522 273055
rect 128470 272991 128522 272997
rect 129730 271649 129758 278018
rect 130882 273499 130910 278018
rect 130870 273493 130922 273499
rect 130870 273435 130922 273441
rect 132034 273203 132062 278018
rect 133282 273351 133310 278018
rect 133270 273345 133322 273351
rect 133270 273287 133322 273293
rect 132022 273197 132074 273203
rect 132022 273139 132074 273145
rect 129718 271643 129770 271649
rect 129718 271585 129770 271591
rect 132406 271643 132458 271649
rect 132406 271585 132458 271591
rect 132418 249819 132446 271585
rect 134434 270465 134462 278018
rect 135586 273351 135614 278018
rect 135286 273345 135338 273351
rect 135286 273287 135338 273293
rect 135574 273345 135626 273351
rect 135574 273287 135626 273293
rect 134422 270459 134474 270465
rect 134422 270401 134474 270407
rect 132406 249813 132458 249819
rect 132406 249755 132458 249761
rect 135298 249745 135326 273287
rect 136834 270761 136862 278018
rect 136822 270755 136874 270761
rect 136822 270697 136874 270703
rect 137986 270539 138014 278018
rect 138262 278007 138314 278013
rect 138262 277949 138314 277955
rect 138274 270761 138302 277949
rect 138166 270755 138218 270761
rect 138166 270697 138218 270703
rect 138262 270755 138314 270761
rect 138262 270697 138314 270703
rect 137974 270533 138026 270539
rect 137974 270475 138026 270481
rect 135286 249739 135338 249745
rect 135286 249681 135338 249687
rect 138178 249597 138206 270697
rect 139138 269915 139166 278018
rect 140400 278004 141086 278032
rect 139124 269906 139180 269915
rect 139124 269841 139180 269850
rect 141058 252557 141086 278004
rect 141538 270613 141566 278018
rect 142690 273425 142718 278018
rect 142678 273419 142730 273425
rect 142678 273361 142730 273367
rect 142582 273271 142634 273277
rect 142582 273213 142634 273219
rect 141526 270607 141578 270613
rect 141526 270549 141578 270555
rect 141046 252551 141098 252557
rect 141046 252493 141098 252499
rect 138166 249591 138218 249597
rect 138166 249533 138218 249539
rect 126646 249517 126698 249523
rect 126646 249459 126698 249465
rect 123766 249443 123818 249449
rect 123766 249385 123818 249391
rect 112246 246705 112298 246711
rect 112246 246647 112298 246653
rect 142486 244929 142538 244935
rect 142486 244871 142538 244877
rect 50614 211333 50666 211339
rect 50614 211275 50666 211281
rect 50422 210149 50474 210155
rect 50422 210091 50474 210097
rect 142498 195854 142526 244871
rect 142594 216014 142622 273213
rect 142678 242635 142730 242641
rect 142678 242577 142730 242583
rect 142690 236174 142718 242577
rect 142690 236146 143102 236174
rect 143074 218887 143102 236146
rect 143062 218881 143114 218887
rect 143062 218823 143114 218829
rect 142594 215986 143102 216014
rect 143074 201571 143102 215986
rect 143062 201565 143114 201571
rect 143062 201507 143114 201513
rect 142498 195826 143102 195854
rect 42166 182251 42218 182257
rect 42166 182193 42218 182199
rect 48118 182251 48170 182257
rect 48118 182193 48170 182199
rect 42178 181925 42206 182193
rect 143074 175671 143102 195826
rect 143938 190101 143966 278018
rect 145090 270687 145118 278018
rect 145078 270681 145130 270687
rect 145078 270623 145130 270629
rect 146242 269207 146270 278018
rect 147394 271871 147422 278018
rect 147382 271865 147434 271871
rect 147382 271807 147434 271813
rect 146230 269201 146282 269207
rect 146230 269143 146282 269149
rect 148642 269133 148670 278018
rect 149686 271865 149738 271871
rect 149686 271807 149738 271813
rect 148630 269127 148682 269133
rect 148630 269069 148682 269075
rect 145558 249887 145610 249893
rect 145558 249829 145610 249835
rect 145462 249369 145514 249375
rect 145462 249311 145514 249317
rect 145366 249295 145418 249301
rect 145366 249237 145418 249243
rect 143926 190095 143978 190101
rect 143926 190037 143978 190043
rect 143062 175665 143114 175671
rect 143062 175607 143114 175613
rect 145378 175597 145406 249237
rect 145474 178557 145502 249311
rect 145570 184329 145598 249829
rect 148340 244598 148396 244607
rect 148340 244533 148396 244542
rect 148244 239714 148300 239723
rect 148244 239649 148300 239658
rect 147668 232314 147724 232323
rect 147668 232249 147724 232258
rect 147682 232059 147710 232249
rect 147670 232053 147722 232059
rect 147670 231995 147722 232001
rect 146900 229946 146956 229955
rect 146900 229881 146956 229890
rect 146914 229839 146942 229881
rect 146902 229833 146954 229839
rect 146902 229775 146954 229781
rect 147670 219103 147722 219109
rect 147670 219045 147722 219051
rect 147682 219003 147710 219045
rect 147668 218994 147724 219003
rect 147668 218929 147724 218938
rect 147284 217810 147340 217819
rect 147284 217745 147286 217754
rect 147338 217745 147340 217754
rect 147286 217713 147338 217719
rect 147380 214850 147436 214859
rect 147380 214785 147436 214794
rect 147394 213189 147422 214785
rect 147572 214110 147628 214119
rect 147572 214045 147628 214054
rect 147586 213337 147614 214045
rect 147574 213331 147626 213337
rect 147574 213273 147626 213279
rect 147382 213183 147434 213189
rect 147382 213125 147434 213131
rect 146900 212926 146956 212935
rect 146900 212861 146902 212870
rect 146954 212861 146956 212870
rect 146902 212829 146954 212835
rect 147380 211742 147436 211751
rect 147380 211677 147436 211686
rect 147394 210525 147422 211677
rect 147382 210519 147434 210525
rect 147382 210461 147434 210467
rect 147380 210410 147436 210419
rect 147380 210345 147382 210354
rect 147434 210345 147436 210354
rect 147382 210313 147434 210319
rect 146900 209226 146956 209235
rect 146900 209161 146956 209170
rect 146914 208379 146942 209161
rect 146902 208373 146954 208379
rect 146902 208315 146954 208321
rect 146996 208042 147052 208051
rect 146996 207977 147052 207986
rect 147010 207417 147038 207977
rect 146998 207411 147050 207417
rect 146998 207353 147050 207359
rect 147092 206414 147148 206423
rect 147092 206349 147148 206358
rect 147106 206307 147134 206349
rect 147094 206301 147146 206307
rect 147094 206243 147146 206249
rect 147668 204490 147724 204499
rect 147668 204425 147724 204434
rect 147682 204087 147710 204425
rect 147670 204081 147722 204087
rect 147670 204023 147722 204029
rect 147476 199606 147532 199615
rect 147476 199541 147532 199550
rect 147490 198833 147518 199541
rect 147478 198827 147530 198833
rect 147478 198769 147530 198775
rect 147286 196015 147338 196021
rect 147286 195957 147338 195963
rect 147298 195915 147326 195957
rect 147284 195906 147340 195915
rect 147284 195841 147340 195850
rect 147284 191022 147340 191031
rect 147284 190957 147340 190966
rect 147298 190175 147326 190957
rect 147286 190169 147338 190175
rect 147286 190111 147338 190117
rect 145558 184323 145610 184329
rect 145558 184265 145610 184271
rect 145462 178551 145514 178557
rect 145462 178493 145514 178499
rect 145366 175591 145418 175597
rect 145366 175533 145418 175539
rect 147668 175186 147724 175195
rect 147668 175121 147724 175130
rect 147682 175079 147710 175121
rect 147670 175073 147722 175079
rect 147670 175015 147722 175021
rect 148258 169751 148286 239649
rect 148354 172637 148382 244533
rect 148532 243414 148588 243423
rect 148532 243349 148588 243358
rect 148436 234830 148492 234839
rect 148436 234765 148492 234774
rect 148342 172631 148394 172637
rect 148342 172573 148394 172579
rect 148246 169745 148298 169751
rect 148246 169687 148298 169693
rect 148450 167013 148478 234765
rect 148546 172785 148574 243349
rect 148724 242082 148780 242091
rect 148724 242017 148780 242026
rect 148628 236754 148684 236763
rect 148628 236689 148684 236698
rect 148534 172779 148586 172785
rect 148534 172721 148586 172727
rect 148642 169899 148670 236689
rect 148738 172711 148766 242017
rect 149012 240898 149068 240907
rect 149012 240833 149068 240842
rect 148820 238530 148876 238539
rect 148820 238465 148876 238474
rect 148726 172705 148778 172711
rect 148726 172647 148778 172653
rect 148724 170302 148780 170311
rect 148724 170237 148780 170246
rect 148630 169893 148682 169899
rect 148630 169835 148682 169841
rect 148438 167007 148490 167013
rect 148438 166949 148490 166955
rect 148738 166717 148766 170237
rect 148834 169825 148862 238465
rect 148916 233646 148972 233655
rect 148916 233581 148972 233590
rect 148930 174117 148958 233581
rect 148918 174111 148970 174117
rect 148918 174053 148970 174059
rect 148916 174002 148972 174011
rect 148916 173937 148972 173946
rect 148822 169819 148874 169825
rect 148822 169761 148874 169767
rect 148726 166711 148778 166717
rect 148726 166653 148778 166659
rect 148724 166306 148780 166315
rect 148724 166241 148780 166250
rect 148532 165566 148588 165575
rect 148532 165501 148588 165510
rect 148340 164382 148396 164391
rect 148340 164317 148396 164326
rect 148244 161866 148300 161875
rect 148244 161801 148300 161810
rect 146900 159498 146956 159507
rect 146900 159433 146956 159442
rect 146914 159169 146942 159433
rect 146902 159163 146954 159169
rect 146902 159105 146954 159111
rect 147862 145473 147914 145479
rect 147862 145415 147914 145421
rect 147094 140219 147146 140225
rect 147094 140161 147146 140167
rect 147106 139971 147134 140161
rect 147092 139962 147148 139971
rect 147092 139897 147148 139906
rect 147188 130342 147244 130351
rect 147188 130277 147190 130286
rect 147242 130277 147244 130286
rect 147190 130245 147242 130251
rect 147874 123723 147902 145415
rect 148258 135374 148286 161801
rect 148354 145479 148382 164317
rect 148436 160682 148492 160691
rect 148436 160617 148492 160626
rect 148342 145473 148394 145479
rect 148342 145415 148394 145421
rect 148342 145325 148394 145331
rect 148342 145267 148394 145273
rect 148162 135346 148286 135374
rect 148162 125740 148190 135346
rect 148246 129415 148298 129421
rect 148246 129357 148298 129363
rect 147970 125712 148190 125740
rect 147862 123717 147914 123723
rect 147862 123659 147914 123665
rect 147970 120985 147998 125712
rect 148148 125458 148204 125467
rect 148148 125393 148204 125402
rect 147958 120979 148010 120985
rect 147958 120921 148010 120927
rect 147668 108438 147724 108447
rect 147668 108373 147670 108382
rect 147722 108373 147724 108382
rect 147670 108341 147722 108347
rect 146996 107254 147052 107263
rect 146996 107189 147052 107198
rect 147010 106629 147038 107189
rect 146998 106623 147050 106629
rect 146998 106565 147050 106571
rect 148162 100783 148190 125393
rect 148258 120911 148286 129357
rect 148354 123649 148382 145267
rect 148450 129421 148478 160617
rect 148438 129415 148490 129421
rect 148438 129357 148490 129363
rect 148546 129292 148574 165501
rect 148628 163198 148684 163207
rect 148628 163133 148684 163142
rect 148642 145553 148670 163133
rect 148630 145547 148682 145553
rect 148630 145489 148682 145495
rect 148738 145424 148766 166241
rect 148820 155798 148876 155807
rect 148820 155733 148876 155742
rect 148834 155691 148862 155733
rect 148822 155685 148874 155691
rect 148822 155627 148874 155633
rect 148930 155617 148958 173937
rect 149026 172563 149054 240833
rect 149108 236014 149164 236023
rect 149108 235949 149164 235958
rect 149014 172557 149066 172563
rect 149014 172499 149066 172505
rect 149122 171176 149150 235949
rect 149396 231130 149452 231139
rect 149396 231065 149398 231074
rect 149450 231065 149452 231074
rect 149398 231033 149450 231039
rect 149396 228170 149452 228179
rect 149396 228105 149452 228114
rect 149410 227619 149438 228105
rect 149398 227613 149450 227619
rect 149398 227555 149450 227561
rect 149300 227430 149356 227439
rect 149300 227365 149356 227374
rect 149314 224881 149342 227365
rect 149396 226394 149452 226403
rect 149396 226329 149452 226338
rect 149302 224875 149354 224881
rect 149302 224817 149354 224823
rect 149410 224807 149438 226329
rect 149492 225210 149548 225219
rect 149492 225145 149548 225154
rect 149398 224801 149450 224807
rect 149398 224743 149450 224749
rect 149506 224733 149534 225145
rect 149494 224727 149546 224733
rect 149494 224669 149546 224675
rect 149492 223878 149548 223887
rect 149492 223813 149548 223822
rect 149396 222694 149452 222703
rect 149396 222629 149452 222638
rect 149410 221847 149438 222629
rect 149506 221921 149534 223813
rect 149494 221915 149546 221921
rect 149494 221857 149546 221863
rect 149398 221841 149450 221847
rect 149398 221783 149450 221789
rect 149492 221510 149548 221519
rect 149492 221445 149548 221454
rect 149396 219734 149452 219743
rect 149396 219669 149452 219678
rect 149410 219035 149438 219669
rect 149398 219029 149450 219035
rect 149398 218971 149450 218977
rect 149506 218961 149534 221445
rect 149494 218955 149546 218961
rect 149494 218897 149546 218903
rect 149396 216626 149452 216635
rect 149396 216561 149452 216570
rect 149410 216445 149438 216561
rect 149398 216439 149450 216445
rect 149398 216381 149450 216387
rect 149396 205674 149452 205683
rect 149396 205609 149452 205618
rect 149410 204605 149438 205609
rect 149398 204599 149450 204605
rect 149398 204541 149450 204547
rect 149492 203306 149548 203315
rect 149492 203241 149548 203250
rect 149506 201719 149534 203241
rect 149494 201713 149546 201719
rect 149396 201678 149452 201687
rect 149494 201655 149546 201661
rect 149396 201613 149398 201622
rect 149450 201613 149452 201622
rect 149398 201581 149450 201587
rect 149396 200790 149452 200799
rect 149396 200725 149452 200734
rect 149410 198759 149438 200725
rect 149398 198753 149450 198759
rect 149398 198695 149450 198701
rect 149300 198422 149356 198431
rect 149300 198357 149356 198366
rect 149314 195873 149342 198357
rect 149396 197090 149452 197099
rect 149396 197025 149452 197034
rect 149410 195947 149438 197025
rect 149398 195941 149450 195947
rect 149398 195883 149450 195889
rect 149302 195867 149354 195873
rect 149302 195809 149354 195815
rect 149492 194722 149548 194731
rect 149492 194657 149548 194666
rect 149396 193390 149452 193399
rect 149396 193325 149452 193334
rect 149410 193209 149438 193325
rect 149398 193203 149450 193209
rect 149398 193145 149450 193151
rect 149506 193061 149534 194657
rect 149494 193055 149546 193061
rect 149494 192997 149546 193003
rect 149396 192206 149452 192215
rect 149396 192141 149452 192150
rect 149410 191137 149438 192141
rect 149398 191131 149450 191137
rect 149398 191073 149450 191079
rect 149698 190027 149726 271807
rect 149794 269059 149822 278018
rect 150946 271649 150974 278018
rect 150934 271643 150986 271649
rect 150934 271585 150986 271591
rect 151606 270755 151658 270761
rect 151606 270697 151658 270703
rect 149782 269053 149834 269059
rect 149782 268995 149834 269001
rect 151618 257811 151646 270697
rect 152194 268985 152222 278018
rect 153346 273277 153374 278018
rect 153334 273271 153386 273277
rect 153334 273213 153386 273219
rect 152374 271643 152426 271649
rect 152374 271585 152426 271591
rect 152182 268979 152234 268985
rect 152182 268921 152234 268927
rect 151606 257805 151658 257811
rect 151606 257747 151658 257753
rect 151222 229833 151274 229839
rect 151222 229775 151274 229781
rect 151126 226133 151178 226139
rect 151126 226075 151178 226081
rect 149686 190021 149738 190027
rect 149686 189963 149738 189969
rect 149396 189838 149452 189847
rect 149396 189773 149452 189782
rect 149300 187470 149356 187479
rect 149300 187405 149356 187414
rect 149204 186286 149260 186295
rect 149204 186221 149260 186230
rect 149218 180037 149246 186221
rect 149314 182997 149342 187405
rect 149410 185809 149438 189773
rect 149588 188062 149644 188071
rect 149588 187997 149644 188006
rect 149398 185803 149450 185809
rect 149398 185745 149450 185751
rect 149396 184510 149452 184519
rect 149396 184445 149452 184454
rect 149302 182991 149354 182997
rect 149302 182933 149354 182939
rect 149410 182868 149438 184445
rect 149492 183770 149548 183779
rect 149492 183705 149548 183714
rect 149314 182840 149438 182868
rect 149206 180031 149258 180037
rect 149206 179973 149258 179979
rect 149314 179908 149342 182840
rect 149396 182586 149452 182595
rect 149396 182521 149452 182530
rect 149410 181591 149438 182521
rect 149398 181585 149450 181591
rect 149398 181527 149450 181533
rect 149506 181517 149534 183705
rect 149602 182923 149630 187997
rect 149590 182917 149642 182923
rect 149590 182859 149642 182865
rect 149494 181511 149546 181517
rect 149494 181453 149546 181459
rect 149492 181402 149548 181411
rect 149492 181337 149548 181346
rect 149218 179880 149342 179908
rect 149218 174265 149246 179880
rect 149300 179626 149356 179635
rect 149300 179561 149356 179570
rect 149314 178631 149342 179561
rect 149396 178886 149452 178895
rect 149396 178821 149452 178830
rect 149410 178705 149438 178821
rect 149506 178779 149534 181337
rect 149494 178773 149546 178779
rect 149494 178715 149546 178721
rect 149398 178699 149450 178705
rect 149398 178641 149450 178647
rect 149302 178625 149354 178631
rect 149302 178567 149354 178573
rect 149492 177702 149548 177711
rect 149492 177637 149548 177646
rect 149396 176518 149452 176527
rect 149396 176453 149452 176462
rect 149410 175819 149438 176453
rect 149398 175813 149450 175819
rect 149398 175755 149450 175761
rect 149506 175745 149534 177637
rect 149494 175739 149546 175745
rect 149494 175681 149546 175687
rect 149206 174259 149258 174265
rect 149206 174201 149258 174207
rect 149398 174111 149450 174117
rect 149398 174053 149450 174059
rect 149122 171148 149342 171176
rect 149204 171042 149260 171051
rect 149204 170977 149260 170986
rect 149218 169548 149246 170977
rect 149314 169677 149342 171148
rect 149302 169671 149354 169677
rect 149302 169613 149354 169619
rect 149218 169520 149342 169548
rect 149012 168082 149068 168091
rect 149012 168017 149068 168026
rect 148918 155611 148970 155617
rect 148918 155553 148970 155559
rect 148450 129264 148574 129292
rect 148642 145396 148766 145424
rect 148450 123797 148478 129264
rect 148532 129158 148588 129167
rect 148532 129093 148588 129102
rect 148438 123791 148490 123797
rect 148438 123733 148490 123739
rect 148342 123643 148394 123649
rect 148342 123585 148394 123591
rect 148246 120905 148298 120911
rect 148246 120847 148298 120853
rect 148546 115255 148574 129093
rect 148642 123871 148670 145396
rect 149026 145276 149054 168017
rect 149314 166810 149342 169520
rect 149410 166939 149438 174053
rect 149588 172818 149644 172827
rect 149588 172753 149644 172762
rect 149492 169118 149548 169127
rect 149492 169053 149548 169062
rect 149398 166933 149450 166939
rect 149398 166875 149450 166881
rect 149314 166782 149438 166810
rect 149110 166711 149162 166717
rect 149110 166653 149162 166659
rect 148738 145248 149054 145276
rect 148738 126609 148766 145248
rect 148820 141294 148876 141303
rect 148820 141229 148822 141238
rect 148874 141229 148876 141238
rect 148822 141197 148874 141203
rect 149122 135374 149150 166653
rect 149300 157722 149356 157731
rect 149300 157657 149356 157666
rect 149314 155765 149342 157657
rect 149302 155759 149354 155765
rect 149302 155701 149354 155707
rect 149302 155611 149354 155617
rect 149302 155553 149354 155559
rect 149204 153134 149260 153143
rect 149204 153069 149260 153078
rect 149218 152805 149246 153069
rect 149206 152799 149258 152805
rect 149206 152741 149258 152747
rect 149204 152098 149260 152107
rect 149204 152033 149260 152042
rect 149218 151843 149246 152033
rect 149206 151837 149258 151843
rect 149206 151779 149258 151785
rect 149206 149913 149258 149919
rect 149204 149878 149206 149887
rect 149258 149878 149260 149887
rect 149204 149813 149260 149822
rect 149204 147362 149260 147371
rect 149204 147297 149260 147306
rect 149218 147033 149246 147297
rect 149206 147027 149258 147033
rect 149206 146969 149258 146975
rect 149204 144550 149260 144559
rect 149204 144485 149260 144494
rect 149218 144147 149246 144485
rect 149206 144141 149258 144147
rect 149206 144083 149258 144089
rect 149204 142478 149260 142487
rect 149204 142413 149260 142422
rect 149218 142297 149246 142413
rect 149206 142291 149258 142297
rect 149206 142233 149258 142239
rect 149204 138778 149260 138787
rect 149204 138713 149260 138722
rect 149218 138301 149246 138713
rect 149206 138295 149258 138301
rect 149206 138237 149258 138243
rect 149204 135966 149260 135975
rect 149204 135901 149260 135910
rect 149218 135489 149246 135901
rect 149206 135483 149258 135489
rect 149206 135425 149258 135431
rect 149314 135374 149342 155553
rect 149026 135346 149150 135374
rect 149218 135346 149342 135374
rect 148820 132710 148876 132719
rect 148820 132645 148876 132654
rect 148726 126603 148778 126609
rect 148726 126545 148778 126551
rect 148630 123865 148682 123871
rect 148630 123807 148682 123813
rect 148532 115246 148588 115255
rect 148532 115181 148588 115190
rect 148726 113727 148778 113733
rect 148726 113669 148778 113675
rect 148244 111990 148300 111999
rect 148244 111925 148300 111934
rect 148150 100777 148202 100783
rect 148150 100719 148202 100725
rect 148258 92051 148286 111925
rect 148436 110954 148492 110963
rect 148436 110889 148492 110898
rect 148340 104738 148396 104747
rect 148340 104673 148396 104682
rect 148246 92045 148298 92051
rect 148246 91987 148298 91993
rect 148354 86427 148382 104673
rect 148450 92125 148478 110889
rect 148532 106070 148588 106079
rect 148532 106005 148588 106014
rect 148438 92119 148490 92125
rect 148438 92061 148490 92067
rect 148546 89239 148574 106005
rect 148628 102370 148684 102379
rect 148628 102305 148684 102314
rect 148534 89233 148586 89239
rect 148534 89175 148586 89181
rect 148342 86421 148394 86427
rect 148342 86363 148394 86369
rect 148642 86353 148670 102305
rect 148738 97897 148766 113669
rect 148834 103595 148862 132645
rect 148916 130934 148972 130943
rect 148916 130869 148972 130878
rect 148930 103669 148958 130869
rect 149026 126683 149054 135346
rect 149218 129495 149246 135346
rect 149410 134028 149438 166782
rect 149506 135193 149534 169053
rect 149494 135187 149546 135193
rect 149494 135129 149546 135135
rect 149492 135078 149548 135087
rect 149492 135013 149548 135022
rect 149314 134000 149438 134028
rect 149314 129569 149342 134000
rect 149396 133894 149452 133903
rect 149396 133829 149452 133838
rect 149410 132603 149438 133829
rect 149398 132597 149450 132603
rect 149398 132539 149450 132545
rect 149506 132529 149534 135013
rect 149494 132523 149546 132529
rect 149494 132465 149546 132471
rect 149302 129563 149354 129569
rect 149302 129505 149354 129511
rect 149206 129489 149258 129495
rect 149206 129431 149258 129437
rect 149602 129421 149630 172753
rect 149684 156982 149740 156991
rect 149684 156917 149740 156926
rect 149698 155617 149726 156917
rect 149686 155611 149738 155617
rect 149686 155553 149738 155559
rect 149684 154614 149740 154623
rect 149684 154549 149740 154558
rect 149698 152731 149726 154549
rect 149686 152725 149738 152731
rect 149686 152667 149738 152673
rect 149684 150914 149740 150923
rect 149684 150849 149740 150858
rect 149698 149845 149726 150849
rect 149686 149839 149738 149845
rect 149686 149781 149738 149787
rect 149684 148546 149740 148555
rect 149684 148481 149740 148490
rect 149698 146959 149726 148481
rect 149686 146953 149738 146959
rect 149686 146895 149738 146901
rect 149684 146178 149740 146187
rect 149684 146113 149740 146122
rect 149698 144073 149726 146113
rect 149686 144067 149738 144073
rect 149686 144009 149738 144015
rect 149684 143662 149740 143671
rect 149684 143597 149740 143606
rect 149698 142371 149726 143597
rect 149686 142365 149738 142371
rect 149686 142307 149738 142313
rect 151138 140225 151166 226075
rect 151234 163905 151262 229775
rect 151798 217771 151850 217777
rect 151798 217713 151850 217719
rect 151702 213331 151754 213337
rect 151702 213273 151754 213279
rect 151510 213183 151562 213189
rect 151510 213125 151562 213131
rect 151414 210371 151466 210377
rect 151414 210313 151466 210319
rect 151318 207411 151370 207417
rect 151318 207353 151370 207359
rect 151222 163899 151274 163905
rect 151222 163841 151274 163847
rect 151222 159163 151274 159169
rect 151222 159105 151274 159111
rect 151126 140219 151178 140225
rect 151126 140161 151178 140167
rect 149684 137594 149740 137603
rect 149684 137529 149740 137538
rect 149698 135415 149726 137529
rect 149686 135409 149738 135415
rect 149686 135351 149738 135357
rect 149686 135187 149738 135193
rect 149686 135129 149738 135135
rect 149590 129415 149642 129421
rect 149590 129357 149642 129363
rect 149108 127974 149164 127983
rect 149108 127909 149164 127918
rect 149014 126677 149066 126683
rect 149014 126619 149066 126625
rect 149012 122498 149068 122507
rect 149012 122433 149068 122442
rect 149026 113733 149054 122433
rect 149014 113727 149066 113733
rect 149014 113669 149066 113675
rect 149014 113579 149066 113585
rect 149014 113521 149066 113527
rect 148918 103663 148970 103669
rect 148918 103605 148970 103611
rect 148822 103589 148874 103595
rect 148822 103531 148874 103537
rect 148726 97891 148778 97897
rect 148726 97833 148778 97839
rect 149026 97823 149054 113521
rect 149122 100635 149150 127909
rect 149588 126642 149644 126651
rect 149588 126577 149644 126586
rect 149300 124274 149356 124283
rect 149300 124209 149356 124218
rect 149204 121758 149260 121767
rect 149204 121693 149260 121702
rect 149218 113585 149246 121693
rect 149206 113579 149258 113585
rect 149206 113521 149258 113527
rect 149314 113456 149342 124209
rect 149396 120574 149452 120583
rect 149396 120509 149452 120518
rect 149410 118321 149438 120509
rect 149492 119390 149548 119399
rect 149492 119325 149548 119334
rect 149398 118315 149450 118321
rect 149398 118257 149450 118263
rect 149506 118247 149534 119325
rect 149494 118241 149546 118247
rect 149396 118206 149452 118215
rect 149494 118183 149546 118189
rect 149396 118141 149398 118150
rect 149450 118141 149452 118150
rect 149398 118109 149450 118115
rect 149396 116874 149452 116883
rect 149396 116809 149452 116818
rect 149410 115361 149438 116809
rect 149492 115690 149548 115699
rect 149492 115625 149548 115634
rect 149398 115355 149450 115361
rect 149398 115297 149450 115303
rect 149506 115287 149534 115625
rect 149494 115281 149546 115287
rect 149396 115246 149452 115255
rect 149494 115223 149546 115229
rect 149396 115181 149452 115190
rect 149602 115214 149630 126577
rect 149698 126535 149726 135129
rect 151126 130303 151178 130309
rect 151126 130245 151178 130251
rect 149686 126529 149738 126535
rect 149686 126471 149738 126477
rect 149602 115186 149726 115214
rect 149218 113428 149342 113456
rect 149218 100709 149246 113428
rect 149410 113308 149438 115181
rect 149492 114506 149548 114515
rect 149492 114441 149548 114450
rect 149314 113280 149438 113308
rect 149314 103521 149342 113280
rect 149396 113174 149452 113183
rect 149396 113109 149452 113118
rect 149410 112919 149438 113109
rect 149398 112913 149450 112919
rect 149398 112855 149450 112861
rect 149506 112401 149534 114441
rect 149494 112395 149546 112401
rect 149494 112337 149546 112343
rect 149396 109622 149452 109631
rect 149396 109557 149398 109566
rect 149450 109557 149452 109566
rect 149398 109525 149450 109531
rect 149588 103554 149644 103563
rect 149302 103515 149354 103521
rect 149588 103489 149644 103498
rect 149302 103457 149354 103463
rect 149396 100890 149452 100899
rect 149396 100825 149398 100834
rect 149450 100825 149452 100834
rect 149398 100793 149450 100799
rect 149206 100703 149258 100709
rect 149206 100645 149258 100651
rect 149110 100629 149162 100635
rect 149110 100571 149162 100577
rect 149492 99854 149548 99863
rect 149492 99789 149548 99798
rect 149396 98670 149452 98679
rect 149396 98605 149452 98614
rect 149410 98045 149438 98605
rect 149398 98039 149450 98045
rect 149398 97981 149450 97987
rect 149506 97971 149534 99789
rect 149494 97965 149546 97971
rect 149494 97907 149546 97913
rect 149014 97817 149066 97823
rect 149014 97759 149066 97765
rect 149492 97486 149548 97495
rect 149492 97421 149548 97430
rect 149396 95710 149452 95719
rect 149396 95645 149452 95654
rect 149410 95085 149438 95645
rect 149506 95159 149534 97421
rect 149494 95153 149546 95159
rect 149494 95095 149546 95101
rect 149398 95079 149450 95085
rect 149398 95021 149450 95027
rect 149492 93786 149548 93795
rect 149492 93721 149548 93730
rect 149396 92602 149452 92611
rect 149396 92537 149452 92546
rect 149410 92421 149438 92537
rect 149398 92415 149450 92421
rect 149398 92357 149450 92363
rect 149506 92199 149534 93721
rect 149494 92193 149546 92199
rect 149494 92135 149546 92141
rect 149204 91418 149260 91427
rect 149204 91353 149260 91362
rect 148724 86534 148780 86543
rect 148724 86469 148726 86478
rect 148778 86469 148780 86478
rect 148726 86437 148778 86443
rect 148630 86347 148682 86353
rect 148630 86289 148682 86295
rect 148436 85350 148492 85359
rect 148436 85285 148492 85294
rect 147092 84166 147148 84175
rect 147092 84101 147148 84110
rect 147106 83615 147134 84101
rect 147094 83609 147146 83615
rect 147094 83551 147146 83557
rect 148244 81650 148300 81659
rect 148244 81585 148300 81594
rect 148258 71997 148286 81585
rect 148450 74883 148478 85285
rect 149108 82390 149164 82399
rect 149108 82325 149164 82334
rect 148820 77950 148876 77959
rect 148820 77885 148876 77894
rect 148438 74877 148490 74883
rect 148438 74819 148490 74825
rect 148246 71991 148298 71997
rect 148246 71933 148298 71939
rect 148834 69111 148862 77885
rect 149122 74809 149150 82325
rect 149218 77769 149246 91353
rect 149300 90234 149356 90243
rect 149300 90169 149356 90178
rect 149206 77763 149258 77769
rect 149206 77705 149258 77711
rect 149314 77695 149342 90169
rect 149396 89050 149452 89059
rect 149396 88985 149452 88994
rect 149302 77689 149354 77695
rect 149302 77631 149354 77637
rect 149410 77621 149438 88985
rect 149492 87422 149548 87431
rect 149492 87357 149548 87366
rect 149506 87093 149534 87357
rect 149494 87087 149546 87093
rect 149494 87029 149546 87035
rect 149602 86279 149630 103489
rect 149698 100561 149726 115186
rect 151138 105149 151166 130245
rect 151234 115213 151262 159105
rect 151330 149771 151358 207353
rect 151426 152657 151454 210313
rect 151522 155469 151550 213125
rect 151606 210519 151658 210525
rect 151606 210461 151658 210467
rect 151510 155463 151562 155469
rect 151510 155405 151562 155411
rect 151414 152651 151466 152657
rect 151414 152593 151466 152599
rect 151618 152583 151646 210461
rect 151714 155543 151742 213273
rect 151810 158429 151838 217713
rect 152086 212887 152138 212893
rect 152086 212829 152138 212835
rect 151990 208373 152042 208379
rect 151990 208315 152042 208321
rect 151894 206301 151946 206307
rect 151894 206243 151946 206249
rect 151798 158423 151850 158429
rect 151798 158365 151850 158371
rect 151702 155537 151754 155543
rect 151702 155479 151754 155485
rect 151606 152577 151658 152583
rect 151606 152519 151658 152525
rect 151318 149765 151370 149771
rect 151318 149707 151370 149713
rect 151906 149697 151934 206243
rect 152002 152509 152030 208315
rect 152098 155395 152126 212829
rect 152182 198827 152234 198833
rect 152182 198769 152234 198775
rect 152086 155389 152138 155395
rect 152086 155331 152138 155337
rect 151990 152503 152042 152509
rect 151990 152445 152042 152451
rect 151894 149691 151946 149697
rect 151894 149633 151946 149639
rect 152194 146663 152222 198769
rect 152386 192987 152414 271585
rect 154498 270761 154526 278018
rect 154486 270755 154538 270761
rect 154486 270697 154538 270703
rect 155446 270755 155498 270761
rect 155446 270697 155498 270703
rect 154006 252403 154058 252409
rect 154006 252345 154058 252351
rect 152374 192981 152426 192987
rect 152374 192923 152426 192929
rect 154018 181443 154046 252345
rect 154102 232053 154154 232059
rect 154102 231995 154154 232001
rect 154006 181437 154058 181443
rect 154006 181379 154058 181385
rect 154006 175073 154058 175079
rect 154006 175015 154058 175021
rect 152182 146657 152234 146663
rect 152182 146599 152234 146605
rect 154018 129347 154046 175015
rect 154114 166865 154142 231995
rect 154198 204081 154250 204087
rect 154198 204023 154250 204029
rect 154102 166859 154154 166865
rect 154102 166801 154154 166807
rect 154210 149623 154238 204023
rect 155458 192913 155486 270697
rect 155746 268911 155774 278018
rect 155734 268905 155786 268911
rect 155734 268847 155786 268853
rect 156898 268837 156926 278018
rect 158050 276494 158078 278018
rect 158050 276466 158174 276494
rect 156886 268831 156938 268837
rect 156886 268773 156938 268779
rect 156886 252477 156938 252483
rect 156886 252419 156938 252425
rect 155446 192907 155498 192913
rect 155446 192849 155498 192855
rect 154294 190169 154346 190175
rect 154294 190111 154346 190117
rect 154198 149617 154250 149623
rect 154198 149559 154250 149565
rect 154102 141255 154154 141261
rect 154102 141197 154154 141203
rect 154006 129341 154058 129347
rect 154006 129283 154058 129289
rect 151222 115207 151274 115213
rect 151222 115149 151274 115155
rect 154114 115139 154142 141197
rect 154306 141113 154334 190111
rect 156898 181369 156926 252419
rect 156982 249665 157034 249671
rect 156982 249607 157034 249613
rect 156994 184255 157022 249607
rect 157078 204599 157130 204605
rect 157078 204541 157130 204547
rect 156982 184249 157034 184255
rect 156982 184191 157034 184197
rect 156886 181363 156938 181369
rect 156886 181305 156938 181311
rect 156886 175813 156938 175819
rect 156886 175755 156938 175761
rect 154294 141107 154346 141113
rect 154294 141049 154346 141055
rect 156898 132233 156926 175755
rect 157090 149549 157118 204541
rect 158146 192839 158174 276466
rect 159298 271945 159326 278018
rect 160450 273573 160478 278018
rect 160438 273567 160490 273573
rect 160438 273509 160490 273515
rect 159286 271939 159338 271945
rect 159286 271881 159338 271887
rect 161602 271353 161630 278018
rect 161590 271347 161642 271353
rect 161590 271289 161642 271295
rect 162850 268763 162878 278018
rect 163894 271347 163946 271353
rect 163894 271289 163946 271295
rect 162838 268757 162890 268763
rect 162838 268699 162890 268705
rect 159766 252329 159818 252335
rect 159766 252271 159818 252277
rect 158134 192833 158186 192839
rect 158134 192775 158186 192781
rect 157174 191131 157226 191137
rect 157174 191073 157226 191079
rect 157078 149543 157130 149549
rect 157078 149485 157130 149491
rect 156982 142291 157034 142297
rect 156982 142233 157034 142239
rect 156886 132227 156938 132233
rect 156886 132169 156938 132175
rect 154102 115133 154154 115139
rect 154102 115075 154154 115081
rect 156994 115065 157022 142233
rect 157186 141039 157214 191073
rect 159778 181295 159806 252271
rect 162742 249813 162794 249819
rect 162742 249755 162794 249761
rect 159958 244855 160010 244861
rect 159958 244797 160010 244803
rect 159862 231091 159914 231097
rect 159862 231033 159914 231039
rect 159766 181289 159818 181295
rect 159766 181231 159818 181237
rect 159874 164053 159902 231033
rect 159970 221773 159998 244797
rect 162646 221915 162698 221921
rect 162646 221857 162698 221863
rect 159958 221767 160010 221773
rect 159958 221709 160010 221715
rect 159958 216439 160010 216445
rect 159958 216381 160010 216387
rect 159862 164047 159914 164053
rect 159862 163989 159914 163995
rect 159970 155321 159998 216381
rect 160054 193203 160106 193209
rect 160054 193145 160106 193151
rect 159958 155315 160010 155321
rect 159958 155257 160010 155263
rect 159958 151837 160010 151843
rect 159958 151779 160010 151785
rect 159862 142365 159914 142371
rect 159862 142307 159914 142313
rect 157174 141033 157226 141039
rect 157174 140975 157226 140981
rect 159766 135483 159818 135489
rect 159766 135425 159818 135431
rect 156982 115059 157034 115065
rect 156982 115001 157034 115007
rect 156886 109583 156938 109589
rect 156886 109525 156938 109531
rect 154006 108399 154058 108405
rect 154006 108341 154058 108347
rect 151222 106623 151274 106629
rect 151222 106565 151274 106571
rect 151126 105143 151178 105149
rect 151126 105085 151178 105091
rect 149686 100555 149738 100561
rect 149686 100497 149738 100503
rect 149684 94970 149740 94979
rect 149684 94905 149740 94914
rect 149590 86273 149642 86279
rect 149590 86215 149642 86221
rect 149698 80655 149726 94905
rect 151234 89165 151262 106565
rect 151222 89159 151274 89165
rect 151222 89101 151274 89107
rect 154018 89091 154046 108341
rect 154006 89085 154058 89091
rect 154006 89027 154058 89033
rect 156898 89017 156926 109525
rect 159778 106555 159806 135425
rect 159874 118099 159902 142307
rect 159970 133935 159998 151779
rect 160066 140965 160094 193145
rect 162658 161241 162686 221857
rect 162754 187215 162782 249755
rect 162838 193055 162890 193061
rect 162838 192997 162890 193003
rect 162742 187209 162794 187215
rect 162742 187151 162794 187157
rect 162742 178773 162794 178779
rect 162742 178715 162794 178721
rect 162646 161235 162698 161241
rect 162646 161177 162698 161183
rect 160054 140959 160106 140965
rect 160054 140901 160106 140907
rect 162646 135409 162698 135415
rect 162646 135351 162698 135357
rect 159958 133929 160010 133935
rect 159958 133871 160010 133877
rect 159862 118093 159914 118099
rect 159862 118035 159914 118041
rect 159862 112913 159914 112919
rect 159862 112855 159914 112861
rect 159766 106549 159818 106555
rect 159766 106491 159818 106497
rect 159574 92415 159626 92421
rect 159574 92357 159626 92363
rect 156886 89011 156938 89017
rect 156886 88953 156938 88959
rect 156406 87087 156458 87093
rect 156406 87029 156458 87035
rect 154102 86495 154154 86501
rect 154102 86437 154154 86443
rect 151126 83609 151178 83615
rect 151126 83551 151178 83557
rect 149686 80649 149738 80655
rect 149686 80591 149738 80597
rect 149588 80466 149644 80475
rect 149588 80401 149644 80410
rect 149398 77615 149450 77621
rect 149398 77557 149450 77563
rect 149204 76766 149260 76775
rect 149204 76701 149260 76710
rect 149110 74803 149162 74809
rect 149110 74745 149162 74751
rect 149012 73066 149068 73075
rect 149012 73001 149068 73010
rect 148822 69105 148874 69111
rect 148822 69047 148874 69053
rect 149026 66003 149054 73001
rect 149108 72030 149164 72039
rect 149108 71965 149164 71974
rect 149122 66225 149150 71965
rect 149218 69037 149246 76701
rect 149396 75582 149452 75591
rect 149396 75517 149452 75526
rect 149410 74894 149438 75517
rect 149410 74866 149534 74894
rect 149300 73806 149356 73815
rect 149300 73741 149356 73750
rect 149206 69031 149258 69037
rect 149206 68973 149258 68979
rect 149314 68889 149342 73741
rect 149506 70980 149534 74866
rect 149602 71849 149630 80401
rect 149684 79282 149740 79291
rect 149684 79217 149740 79226
rect 149698 71923 149726 79217
rect 151138 74735 151166 83551
rect 151126 74729 151178 74735
rect 151126 74671 151178 74677
rect 154114 74661 154142 86437
rect 156418 77547 156446 87029
rect 159586 80581 159614 92357
rect 159874 91977 159902 112855
rect 162658 106481 162686 135351
rect 162754 135341 162782 178715
rect 162850 143999 162878 192997
rect 163906 192765 163934 271289
rect 164002 268689 164030 278018
rect 165154 272241 165182 278018
rect 165142 272235 165194 272241
rect 165142 272177 165194 272183
rect 166306 271871 166334 278018
rect 166966 272235 167018 272241
rect 166966 272177 167018 272183
rect 166294 271865 166346 271871
rect 166294 271807 166346 271813
rect 163990 268683 164042 268689
rect 163990 268625 164042 268631
rect 165526 252181 165578 252187
rect 165526 252123 165578 252129
rect 163894 192759 163946 192765
rect 163894 192701 163946 192707
rect 165538 178483 165566 252123
rect 165622 224875 165674 224881
rect 165622 224817 165674 224823
rect 165526 178477 165578 178483
rect 165526 178419 165578 178425
rect 165634 163979 165662 224817
rect 165718 198753 165770 198759
rect 165718 198695 165770 198701
rect 165622 163973 165674 163979
rect 165622 163915 165674 163921
rect 165730 146811 165758 198695
rect 166978 195799 167006 272177
rect 167554 272093 167582 278018
rect 167542 272087 167594 272093
rect 167542 272029 167594 272035
rect 168706 270761 168734 278018
rect 169762 278004 169872 278032
rect 168694 270755 168746 270761
rect 168694 270697 168746 270703
rect 169762 268615 169790 278004
rect 169846 270755 169898 270761
rect 169846 270697 169898 270703
rect 169750 268609 169802 268615
rect 169750 268551 169802 268557
rect 169750 257805 169802 257811
rect 169750 257747 169802 257753
rect 168502 249739 168554 249745
rect 168502 249681 168554 249687
rect 168406 221841 168458 221847
rect 168406 221783 168458 221789
rect 166966 195793 167018 195799
rect 166966 195735 167018 195741
rect 165814 181585 165866 181591
rect 165814 181527 165866 181533
rect 165718 146805 165770 146811
rect 165718 146747 165770 146753
rect 162934 144141 162986 144147
rect 162934 144083 162986 144089
rect 162838 143993 162890 143999
rect 162838 143935 162890 143941
rect 162742 135335 162794 135341
rect 162742 135277 162794 135283
rect 162946 118025 162974 144083
rect 165622 144067 165674 144073
rect 165622 144009 165674 144015
rect 165526 138295 165578 138301
rect 165526 138237 165578 138243
rect 162934 118019 162986 118025
rect 162934 117961 162986 117967
rect 162742 112395 162794 112401
rect 162742 112337 162794 112343
rect 162646 106475 162698 106481
rect 162646 106417 162698 106423
rect 162358 92193 162410 92199
rect 162358 92135 162410 92141
rect 159862 91971 159914 91977
rect 159862 91913 159914 91919
rect 159574 80575 159626 80581
rect 159574 80517 159626 80523
rect 162370 80507 162398 92135
rect 162754 91903 162782 112337
rect 165538 109441 165566 138237
rect 165634 117951 165662 144009
rect 165826 135267 165854 181527
rect 168418 161167 168446 221783
rect 168514 187141 168542 249681
rect 169762 243085 169790 257747
rect 169750 243079 169802 243085
rect 169750 243021 169802 243027
rect 168598 196015 168650 196021
rect 168598 195957 168650 195963
rect 168502 187135 168554 187141
rect 168502 187077 168554 187083
rect 168502 175739 168554 175745
rect 168502 175681 168554 175687
rect 168406 161161 168458 161167
rect 168406 161103 168458 161109
rect 168406 147027 168458 147033
rect 168406 146969 168458 146975
rect 165814 135261 165866 135267
rect 165814 135203 165866 135209
rect 165622 117945 165674 117951
rect 165622 117887 165674 117893
rect 168418 117877 168446 146969
rect 168514 132381 168542 175681
rect 168610 143925 168638 195957
rect 169858 195725 169886 270697
rect 171106 268541 171134 278018
rect 172272 278004 172766 278032
rect 171094 268535 171146 268541
rect 171094 268477 171146 268483
rect 171382 252551 171434 252557
rect 171382 252493 171434 252499
rect 171286 224801 171338 224807
rect 171286 224743 171338 224749
rect 169846 195719 169898 195725
rect 169846 195661 169898 195667
rect 171298 161093 171326 224743
rect 171394 189953 171422 252493
rect 171478 195941 171530 195947
rect 171478 195883 171530 195889
rect 171382 189947 171434 189953
rect 171382 189889 171434 189895
rect 171382 178699 171434 178705
rect 171382 178641 171434 178647
rect 171286 161087 171338 161093
rect 171286 161029 171338 161035
rect 168598 143919 168650 143925
rect 168598 143861 168650 143867
rect 171286 132597 171338 132603
rect 171286 132539 171338 132545
rect 168502 132375 168554 132381
rect 168502 132317 168554 132323
rect 168502 118315 168554 118321
rect 168502 118257 168554 118263
rect 168406 117871 168458 117877
rect 168406 117813 168458 117819
rect 165718 115355 165770 115361
rect 165718 115297 165770 115303
rect 165526 109435 165578 109441
rect 165526 109377 165578 109383
rect 165526 95153 165578 95159
rect 165526 95095 165578 95101
rect 162742 91897 162794 91903
rect 162742 91839 162794 91845
rect 165538 83541 165566 95095
rect 165730 94789 165758 115297
rect 168406 100851 168458 100857
rect 168406 100793 168458 100799
rect 165718 94783 165770 94789
rect 165718 94725 165770 94731
rect 165526 83535 165578 83541
rect 165526 83477 165578 83483
rect 168418 83467 168446 100793
rect 168514 97749 168542 118257
rect 171298 106407 171326 132539
rect 171394 132307 171422 178641
rect 171490 143851 171518 195883
rect 172738 195651 172766 278004
rect 173410 271797 173438 278018
rect 174658 272019 174686 278018
rect 174646 272013 174698 272019
rect 174646 271955 174698 271961
rect 173398 271791 173450 271797
rect 173398 271733 173450 271739
rect 175810 271205 175838 278018
rect 175798 271199 175850 271205
rect 175798 271141 175850 271147
rect 176962 268467 176990 278018
rect 176950 268461 177002 268467
rect 176950 268403 177002 268409
rect 178210 268393 178238 278018
rect 178294 271199 178346 271205
rect 178294 271141 178346 271147
rect 178198 268387 178250 268393
rect 178198 268329 178250 268335
rect 177046 252255 177098 252261
rect 177046 252197 177098 252203
rect 174166 252107 174218 252113
rect 174166 252049 174218 252055
rect 172726 195645 172778 195651
rect 172726 195587 172778 195593
rect 174178 181221 174206 252049
rect 174454 249443 174506 249449
rect 174454 249385 174506 249391
rect 174262 224727 174314 224733
rect 174262 224669 174314 224675
rect 174166 181215 174218 181221
rect 174166 181157 174218 181163
rect 174274 161019 174302 224669
rect 174358 219103 174410 219109
rect 174358 219045 174410 219051
rect 174262 161013 174314 161019
rect 174262 160955 174314 160961
rect 174370 158355 174398 219045
rect 174466 187067 174494 249385
rect 174454 187061 174506 187067
rect 174454 187003 174506 187009
rect 177058 184181 177086 252197
rect 177238 249517 177290 249523
rect 177238 249459 177290 249465
rect 177142 219029 177194 219035
rect 177142 218971 177194 218977
rect 177046 184175 177098 184181
rect 177046 184117 177098 184123
rect 174454 181511 174506 181517
rect 174454 181453 174506 181459
rect 174358 158349 174410 158355
rect 174358 158291 174410 158297
rect 174166 149913 174218 149919
rect 174166 149855 174218 149861
rect 171574 146953 171626 146959
rect 171574 146895 171626 146901
rect 171478 143845 171530 143851
rect 171478 143787 171530 143793
rect 171382 132301 171434 132307
rect 171382 132243 171434 132249
rect 171586 120837 171614 146895
rect 171574 120831 171626 120837
rect 171574 120773 171626 120779
rect 174178 120763 174206 149855
rect 174466 135193 174494 181453
rect 177154 158207 177182 218971
rect 177250 186993 177278 249459
rect 178306 198611 178334 271141
rect 179362 270761 179390 278018
rect 180514 271575 180542 278018
rect 181762 271649 181790 278018
rect 181750 271643 181802 271649
rect 181750 271585 181802 271591
rect 180502 271569 180554 271575
rect 180502 271511 180554 271517
rect 182914 270761 182942 278018
rect 184066 271279 184094 278018
rect 185218 271501 185246 278018
rect 185206 271495 185258 271501
rect 185206 271437 185258 271443
rect 184054 271273 184106 271279
rect 184054 271215 184106 271221
rect 186466 270761 186494 278018
rect 187618 271131 187646 278018
rect 188770 271353 188798 278018
rect 189730 278004 190032 278032
rect 188758 271347 188810 271353
rect 188758 271289 188810 271295
rect 187606 271125 187658 271131
rect 187606 271067 187658 271073
rect 179350 270755 179402 270761
rect 179350 270697 179402 270703
rect 181366 270755 181418 270761
rect 181366 270697 181418 270703
rect 182902 270755 182954 270761
rect 182902 270697 182954 270703
rect 184246 270755 184298 270761
rect 184246 270697 184298 270703
rect 185494 270755 185546 270761
rect 185494 270697 185546 270703
rect 186454 270755 186506 270761
rect 186454 270697 186506 270703
rect 180022 249591 180074 249597
rect 180022 249533 180074 249539
rect 179926 218955 179978 218961
rect 179926 218897 179978 218903
rect 178294 198605 178346 198611
rect 178294 198547 178346 198553
rect 177334 195867 177386 195873
rect 177334 195809 177386 195815
rect 177238 186987 177290 186993
rect 177238 186929 177290 186935
rect 177142 158201 177194 158207
rect 177142 158143 177194 158149
rect 174550 155759 174602 155765
rect 174550 155701 174602 155707
rect 174454 135187 174506 135193
rect 174454 135129 174506 135135
rect 174562 134009 174590 155701
rect 177046 152799 177098 152805
rect 177046 152741 177098 152747
rect 174550 134003 174602 134009
rect 174550 133945 174602 133951
rect 174262 132523 174314 132529
rect 174262 132465 174314 132471
rect 174166 120757 174218 120763
rect 174166 120699 174218 120705
rect 171286 106401 171338 106407
rect 171286 106343 171338 106349
rect 174274 106333 174302 132465
rect 174358 118241 174410 118247
rect 174358 118183 174410 118189
rect 174262 106327 174314 106333
rect 174262 106269 174314 106275
rect 168502 97743 168554 97749
rect 168502 97685 168554 97691
rect 174370 94937 174398 118183
rect 177058 109367 177086 152741
rect 177142 152725 177194 152731
rect 177142 152667 177194 152673
rect 177154 112179 177182 152667
rect 177346 143777 177374 195809
rect 179938 158281 179966 218897
rect 180034 189879 180062 249533
rect 180118 243079 180170 243085
rect 180118 243021 180170 243027
rect 180130 212893 180158 243021
rect 180118 212887 180170 212893
rect 180118 212829 180170 212835
rect 180118 201713 180170 201719
rect 180118 201655 180170 201661
rect 180022 189873 180074 189879
rect 180022 189815 180074 189821
rect 179926 158275 179978 158281
rect 179926 158217 179978 158223
rect 180022 155685 180074 155691
rect 180022 155627 180074 155633
rect 179926 149839 179978 149845
rect 179926 149781 179978 149787
rect 177334 143771 177386 143777
rect 177334 143713 177386 143719
rect 179938 123575 179966 149781
rect 179926 123569 179978 123575
rect 179926 123511 179978 123517
rect 179926 115281 179978 115287
rect 179926 115223 179978 115229
rect 177142 112173 177194 112179
rect 177142 112115 177194 112121
rect 177046 109361 177098 109367
rect 177046 109303 177098 109309
rect 174358 94931 174410 94937
rect 174358 94873 174410 94879
rect 179938 94641 179966 115223
rect 180034 112253 180062 155627
rect 180130 146737 180158 201655
rect 181378 198685 181406 270697
rect 182806 252033 182858 252039
rect 182806 251975 182858 251981
rect 181366 198679 181418 198685
rect 181366 198621 181418 198627
rect 182818 178409 182846 251975
rect 182902 227613 182954 227619
rect 182902 227555 182954 227561
rect 182806 178403 182858 178409
rect 182806 178345 182858 178351
rect 182914 164127 182942 227555
rect 182998 201639 183050 201645
rect 182998 201581 183050 201587
rect 182902 164121 182954 164127
rect 182902 164063 182954 164069
rect 182806 155611 182858 155617
rect 182806 155553 182858 155559
rect 180118 146731 180170 146737
rect 180118 146673 180170 146679
rect 182818 112327 182846 155553
rect 183010 146885 183038 201581
rect 184258 197691 184286 270697
rect 184342 221767 184394 221773
rect 184342 221709 184394 221715
rect 184354 219595 184382 221709
rect 184340 219586 184396 219595
rect 184340 219521 184396 219530
rect 184342 218881 184394 218887
rect 184340 218846 184342 218855
rect 184394 218846 184396 218855
rect 184340 218781 184396 218790
rect 184342 201565 184394 201571
rect 184342 201507 184394 201513
rect 184354 199763 184382 201507
rect 184340 199754 184396 199763
rect 184340 199689 184396 199698
rect 184438 198679 184490 198685
rect 184438 198621 184490 198627
rect 184342 198605 184394 198611
rect 184342 198547 184394 198553
rect 184244 197682 184300 197691
rect 184244 197617 184300 197626
rect 184354 196063 184382 198547
rect 184450 196803 184478 198621
rect 185506 198283 185534 270697
rect 189730 257811 189758 278004
rect 191170 272167 191198 278018
rect 191158 272161 191210 272167
rect 191158 272103 191210 272109
rect 192322 271723 192350 278018
rect 192982 273493 193034 273499
rect 192982 273435 193034 273441
rect 192406 272235 192458 272241
rect 192406 272177 192458 272183
rect 192310 271717 192362 271723
rect 192310 271659 192362 271665
rect 192418 263810 192446 272177
rect 192596 269462 192652 269471
rect 192596 269397 192652 269406
rect 192610 263824 192638 269397
rect 192994 268245 193022 273435
rect 193570 271427 193598 278018
rect 194420 272274 194476 272283
rect 194722 272241 194750 278018
rect 195874 273499 195902 278018
rect 195862 273493 195914 273499
rect 195862 273435 195914 273441
rect 196628 272422 196684 272431
rect 196628 272357 196684 272366
rect 194420 272209 194476 272218
rect 194710 272235 194762 272241
rect 193748 272126 193804 272135
rect 193748 272061 193804 272070
rect 193558 271421 193610 271427
rect 193558 271363 193610 271369
rect 193076 269610 193132 269619
rect 193076 269545 193132 269554
rect 192982 268239 193034 268245
rect 192982 268181 193034 268187
rect 193090 263824 193118 269545
rect 192610 263796 192864 263824
rect 193090 263796 193344 263824
rect 193762 263810 193790 272061
rect 194228 269314 194284 269323
rect 194228 269249 194284 269258
rect 194242 263810 194270 269249
rect 194434 263824 194462 272209
rect 194710 272177 194762 272183
rect 195670 271199 195722 271205
rect 195670 271141 195722 271147
rect 194998 269275 195050 269281
rect 194998 269217 195050 269223
rect 195010 263824 195038 269217
rect 194434 263796 194736 263824
rect 195010 263796 195264 263824
rect 195682 263810 195710 271141
rect 196148 269758 196204 269767
rect 196148 269693 196204 269702
rect 196162 263810 196190 269693
rect 196642 263810 196670 272357
rect 196822 269349 196874 269355
rect 196822 269291 196874 269297
rect 196834 263824 196862 269291
rect 197122 269281 197150 278018
rect 198274 272315 198302 278018
rect 199220 272570 199276 272579
rect 199220 272505 199276 272514
rect 199126 272457 199178 272463
rect 199126 272399 199178 272405
rect 198262 272309 198314 272315
rect 198262 272251 198314 272257
rect 198646 271939 198698 271945
rect 198646 271881 198698 271887
rect 198550 271051 198602 271057
rect 198550 270993 198602 270999
rect 198070 269571 198122 269577
rect 198070 269513 198122 269519
rect 197398 269423 197450 269429
rect 197398 269365 197450 269371
rect 197110 269275 197162 269281
rect 197110 269217 197162 269223
rect 197410 263824 197438 269365
rect 196834 263796 197088 263824
rect 197410 263796 197664 263824
rect 198082 263810 198110 269513
rect 198562 263810 198590 270993
rect 198658 268319 198686 271881
rect 199030 269497 199082 269503
rect 199030 269439 199082 269445
rect 198646 268313 198698 268319
rect 198646 268255 198698 268261
rect 199042 263810 199070 269439
rect 199138 267875 199166 272399
rect 199126 267869 199178 267875
rect 199126 267811 199178 267817
rect 199234 263824 199262 272505
rect 199426 271205 199454 278018
rect 200468 272718 200524 272727
rect 200468 272653 200524 272662
rect 199414 271199 199466 271205
rect 199414 271141 199466 271147
rect 199702 269645 199754 269651
rect 199702 269587 199754 269593
rect 199714 263824 199742 269587
rect 199234 263796 199488 263824
rect 199714 263796 199968 263824
rect 200482 263810 200510 272653
rect 200674 269355 200702 278018
rect 201622 272383 201674 272389
rect 201622 272325 201674 272331
rect 201526 271865 201578 271871
rect 201526 271807 201578 271813
rect 201538 269799 201566 271807
rect 201142 269793 201194 269799
rect 201142 269735 201194 269741
rect 201526 269793 201578 269799
rect 201526 269735 201578 269741
rect 200950 269719 201002 269725
rect 200950 269661 201002 269667
rect 200662 269349 200714 269355
rect 200662 269291 200714 269297
rect 200962 263810 200990 269661
rect 201154 263824 201182 269735
rect 201634 263824 201662 272325
rect 201826 271945 201854 278018
rect 201814 271939 201866 271945
rect 201814 271881 201866 271887
rect 202870 269867 202922 269873
rect 202870 269809 202922 269815
rect 202294 267869 202346 267875
rect 202294 267811 202346 267817
rect 201154 263796 201408 263824
rect 201634 263796 201888 263824
rect 202306 263810 202334 267811
rect 202882 263810 202910 269809
rect 202978 269503 203006 278018
rect 204022 272605 204074 272611
rect 204022 272547 204074 272553
rect 203542 272531 203594 272537
rect 203542 272473 203594 272479
rect 203350 269941 203402 269947
rect 203350 269883 203402 269889
rect 202966 269497 203018 269503
rect 202966 269439 203018 269445
rect 203362 263810 203390 269883
rect 203554 263824 203582 272473
rect 204034 263824 204062 272547
rect 204130 269429 204158 278018
rect 205378 271871 205406 278018
rect 206230 272753 206282 272759
rect 206230 272695 206282 272701
rect 205462 272679 205514 272685
rect 205462 272621 205514 272627
rect 205366 271865 205418 271871
rect 205366 271807 205418 271813
rect 205270 270089 205322 270095
rect 205270 270031 205322 270037
rect 204694 270015 204746 270021
rect 204694 269957 204746 269963
rect 204118 269423 204170 269429
rect 204118 269365 204170 269371
rect 203554 263796 203808 263824
rect 204034 263796 204288 263824
rect 204706 263810 204734 269957
rect 205282 263810 205310 270031
rect 205474 263824 205502 272621
rect 206038 271791 206090 271797
rect 206038 271733 206090 271739
rect 205846 271569 205898 271575
rect 205846 271511 205898 271517
rect 205750 271273 205802 271279
rect 205750 271215 205802 271221
rect 205762 269651 205790 271215
rect 205858 269947 205886 271511
rect 205942 271125 205994 271131
rect 205942 271067 205994 271073
rect 205846 269941 205898 269947
rect 205846 269883 205898 269889
rect 205954 269725 205982 271067
rect 206050 269873 206078 271733
rect 206038 269867 206090 269873
rect 206038 269809 206090 269815
rect 205942 269719 205994 269725
rect 205942 269661 205994 269667
rect 205750 269645 205802 269651
rect 205750 269587 205802 269593
rect 206242 264120 206270 272695
rect 206422 270237 206474 270243
rect 206422 270179 206474 270185
rect 206194 264092 206270 264120
rect 205474 263796 205776 263824
rect 206194 263810 206222 264092
rect 206434 263824 206462 270179
rect 206530 269577 206558 278018
rect 207478 273567 207530 273573
rect 207478 273509 207530 273515
rect 207382 273271 207434 273277
rect 207382 273213 207434 273219
rect 207094 272901 207146 272907
rect 207094 272843 207146 272849
rect 206518 269571 206570 269577
rect 206518 269513 206570 269519
rect 206434 263796 206688 263824
rect 207106 263810 207134 272843
rect 207394 268097 207422 273213
rect 207382 268091 207434 268097
rect 207382 268033 207434 268039
rect 207490 267875 207518 273509
rect 207682 272389 207710 278018
rect 208150 273419 208202 273425
rect 208150 273361 208202 273367
rect 207862 272827 207914 272833
rect 207862 272769 207914 272775
rect 207670 272383 207722 272389
rect 207670 272325 207722 272331
rect 207574 270163 207626 270169
rect 207574 270105 207626 270111
rect 207478 267869 207530 267875
rect 207478 267811 207530 267817
rect 207586 263810 207614 270105
rect 207874 263824 207902 272769
rect 208162 268139 208190 273361
rect 208930 272611 208958 278018
rect 209782 273345 209834 273351
rect 209782 273287 209834 273293
rect 209014 272975 209066 272981
rect 209014 272917 209066 272923
rect 208918 272605 208970 272611
rect 208918 272547 208970 272553
rect 208342 270311 208394 270317
rect 208342 270253 208394 270259
rect 208148 268130 208204 268139
rect 208148 268065 208204 268074
rect 208354 263824 208382 270253
rect 207874 263796 208128 263824
rect 208354 263796 208608 263824
rect 209026 263810 209054 272917
rect 209494 270385 209546 270391
rect 209494 270327 209546 270333
rect 209506 263810 209534 270327
rect 209794 268171 209822 273287
rect 209878 273197 209930 273203
rect 209878 273139 209930 273145
rect 209782 268165 209834 268171
rect 209782 268107 209834 268113
rect 209890 268023 209918 273139
rect 209974 273123 210026 273129
rect 209974 273065 210026 273071
rect 209878 268017 209930 268023
rect 209878 267959 209930 267965
rect 209986 263810 210014 273065
rect 210082 272537 210110 278018
rect 210166 273049 210218 273055
rect 210166 272991 210218 272997
rect 210070 272531 210122 272537
rect 210070 272473 210122 272479
rect 210178 267968 210206 272991
rect 211234 272759 211262 278018
rect 212482 272833 212510 278018
rect 213634 272907 213662 278018
rect 213622 272901 213674 272907
rect 213622 272843 213674 272849
rect 212470 272827 212522 272833
rect 212470 272769 212522 272775
rect 211222 272753 211274 272759
rect 211222 272695 211274 272701
rect 214786 272685 214814 278018
rect 216034 273129 216062 278018
rect 216022 273123 216074 273129
rect 216022 273065 216074 273071
rect 217186 272981 217214 278018
rect 218338 273203 218366 278018
rect 219586 273425 219614 278018
rect 219574 273419 219626 273425
rect 219574 273361 219626 273367
rect 218326 273197 218378 273203
rect 218326 273139 218378 273145
rect 220738 273055 220766 278018
rect 221494 273493 221546 273499
rect 221494 273435 221546 273441
rect 220726 273049 220778 273055
rect 220726 272991 220778 272997
rect 217174 272975 217226 272981
rect 217174 272917 217226 272923
rect 214774 272679 214826 272685
rect 214774 272621 214826 272627
rect 210646 272087 210698 272093
rect 210646 272029 210698 272035
rect 210550 272013 210602 272019
rect 210550 271955 210602 271961
rect 210454 271643 210506 271649
rect 210454 271585 210506 271591
rect 210358 271495 210410 271501
rect 210358 271437 210410 271443
rect 210262 271347 210314 271353
rect 210262 271289 210314 271295
rect 210274 270021 210302 271289
rect 210370 270095 210398 271437
rect 210466 270169 210494 271585
rect 210562 270317 210590 271955
rect 210550 270311 210602 270317
rect 210550 270253 210602 270259
rect 210454 270163 210506 270169
rect 210454 270105 210506 270111
rect 210358 270089 210410 270095
rect 210358 270031 210410 270037
rect 210262 270015 210314 270021
rect 210262 269957 210314 269963
rect 210178 267940 210302 267968
rect 210658 267949 210686 272029
rect 214486 270681 214538 270687
rect 214486 270623 214538 270629
rect 213814 270607 213866 270613
rect 213814 270549 213866 270555
rect 212662 270533 212714 270539
rect 212662 270475 212714 270481
rect 211894 270459 211946 270465
rect 211894 270401 211946 270407
rect 210742 268239 210794 268245
rect 210742 268181 210794 268187
rect 210274 263824 210302 267940
rect 210646 267943 210698 267949
rect 210646 267885 210698 267891
rect 210754 263824 210782 268181
rect 211414 268017 211466 268023
rect 211414 267959 211466 267965
rect 210274 263796 210528 263824
rect 210754 263796 211008 263824
rect 211426 263810 211454 267959
rect 211906 263810 211934 270401
rect 212374 268165 212426 268171
rect 212374 268107 212426 268113
rect 212470 268165 212522 268171
rect 212470 268107 212522 268113
rect 212386 263810 212414 268107
rect 212482 267875 212510 268107
rect 212470 267869 212522 267875
rect 212470 267811 212522 267817
rect 212674 263824 212702 270475
rect 213332 269906 213388 269915
rect 213332 269841 213388 269850
rect 212674 263796 212928 263824
rect 213346 263810 213374 269841
rect 213826 263810 213854 270549
rect 214292 268130 214348 268139
rect 214292 268065 214348 268074
rect 214306 263810 214334 268065
rect 214498 263824 214526 270623
rect 220534 269793 220586 269799
rect 220534 269735 220586 269741
rect 214966 269201 215018 269207
rect 214966 269143 215018 269149
rect 214978 263824 215006 269143
rect 215734 269127 215786 269133
rect 215734 269069 215786 269075
rect 214498 263796 214752 263824
rect 214978 263796 215232 263824
rect 215746 263810 215774 269069
rect 216214 269053 216266 269059
rect 216214 268995 216266 269001
rect 216226 263810 216254 268995
rect 216694 268979 216746 268985
rect 216694 268921 216746 268927
rect 216706 263810 216734 268921
rect 217366 268905 217418 268911
rect 217366 268847 217418 268853
rect 216886 268091 216938 268097
rect 216886 268033 216938 268039
rect 216898 263824 216926 268033
rect 217378 263824 217406 268847
rect 218134 268831 218186 268837
rect 218134 268773 218186 268779
rect 216898 263796 217152 263824
rect 217378 263796 217632 263824
rect 218146 263810 218174 268773
rect 219286 268757 219338 268763
rect 219286 268699 219338 268705
rect 218614 268313 218666 268319
rect 218614 268255 218666 268261
rect 218626 263810 218654 268255
rect 218902 268165 218954 268171
rect 218902 268107 218954 268113
rect 218914 263824 218942 268107
rect 219298 263824 219326 268699
rect 219958 268683 220010 268689
rect 219958 268625 220010 268631
rect 218914 263796 219072 263824
rect 219298 263796 219552 263824
rect 219970 263810 219998 268625
rect 220546 263810 220574 269735
rect 221206 268609 221258 268615
rect 221206 268551 221258 268557
rect 221014 267943 221066 267949
rect 221014 267885 221066 267891
rect 221026 263810 221054 267885
rect 221218 263824 221246 268551
rect 221506 268319 221534 273435
rect 221686 271421 221738 271427
rect 221686 271363 221738 271369
rect 221590 271199 221642 271205
rect 221590 271141 221642 271147
rect 221494 268313 221546 268319
rect 221494 268255 221546 268261
rect 221602 268023 221630 271141
rect 221590 268017 221642 268023
rect 221590 267959 221642 267965
rect 221698 267949 221726 271363
rect 221890 271057 221918 278018
rect 221878 271051 221930 271057
rect 221878 270993 221930 270999
rect 223042 270983 223070 278018
rect 223702 271939 223754 271945
rect 223702 271881 223754 271887
rect 223030 270977 223082 270983
rect 223030 270919 223082 270925
rect 222838 270311 222890 270317
rect 222838 270253 222890 270259
rect 222358 269867 222410 269873
rect 222358 269809 222410 269815
rect 221782 268535 221834 268541
rect 221782 268477 221834 268483
rect 221686 267943 221738 267949
rect 221686 267885 221738 267891
rect 221794 263824 221822 268477
rect 221218 263796 221472 263824
rect 221794 263796 221952 263824
rect 222370 263810 222398 269809
rect 222850 263810 222878 270253
rect 223414 268461 223466 268467
rect 223414 268403 223466 268409
rect 223426 263810 223454 268403
rect 223606 268387 223658 268393
rect 223606 268329 223658 268335
rect 223618 263824 223646 268329
rect 223714 268245 223742 271881
rect 224290 270909 224318 278018
rect 224374 272309 224426 272315
rect 224374 272251 224426 272257
rect 224278 270903 224330 270909
rect 224278 270845 224330 270851
rect 224086 269941 224138 269947
rect 224086 269883 224138 269889
rect 223702 268239 223754 268245
rect 223702 268181 223754 268187
rect 224098 263824 224126 269883
rect 224386 268171 224414 272251
rect 224470 272235 224522 272241
rect 224470 272177 224522 272183
rect 224374 268165 224426 268171
rect 224374 268107 224426 268113
rect 224482 268097 224510 272177
rect 224566 271717 224618 271723
rect 224566 271659 224618 271665
rect 224470 268091 224522 268097
rect 224470 268033 224522 268039
rect 224578 267875 224606 271659
rect 225442 270835 225470 278018
rect 225430 270829 225482 270835
rect 225430 270771 225482 270777
rect 226594 270761 226622 278018
rect 227842 272315 227870 278018
rect 227830 272309 227882 272315
rect 227830 272251 227882 272257
rect 228994 272167 229022 278018
rect 230146 273573 230174 278018
rect 230134 273567 230186 273573
rect 230134 273509 230186 273515
rect 227158 272161 227210 272167
rect 227158 272103 227210 272109
rect 228982 272161 229034 272167
rect 228982 272103 229034 272109
rect 226582 270755 226634 270761
rect 226582 270697 226634 270703
rect 224758 270163 224810 270169
rect 224758 270105 224810 270111
rect 224566 267869 224618 267875
rect 224566 267811 224618 267817
rect 223618 263796 223872 263824
rect 224098 263796 224352 263824
rect 224770 263810 224798 270105
rect 225526 270089 225578 270095
rect 225526 270031 225578 270037
rect 225238 269645 225290 269651
rect 225238 269587 225290 269593
rect 225250 263810 225278 269587
rect 225538 263824 225566 270031
rect 226678 270015 226730 270021
rect 226678 269957 226730 269963
rect 226006 269719 226058 269725
rect 226006 269661 226058 269667
rect 226018 263824 226046 269661
rect 225538 263796 225792 263824
rect 226018 263796 226272 263824
rect 226690 263810 226718 269957
rect 227170 263810 227198 272103
rect 231394 272019 231422 278018
rect 232546 272463 232574 278018
rect 232534 272457 232586 272463
rect 232534 272399 232586 272405
rect 231382 272013 231434 272019
rect 231382 271955 231434 271961
rect 233698 271945 233726 278018
rect 234358 272605 234410 272611
rect 234358 272547 234410 272553
rect 233878 272383 233930 272389
rect 233878 272325 233930 272331
rect 233686 271939 233738 271945
rect 233686 271881 233738 271887
rect 232630 271865 232682 271871
rect 232630 271807 232682 271813
rect 231958 269497 232010 269503
rect 231958 269439 232010 269445
rect 230998 269349 231050 269355
rect 230998 269291 231050 269297
rect 229558 269275 229610 269281
rect 229558 269217 229610 269223
rect 229078 268313 229130 268319
rect 229078 268255 229130 268261
rect 228406 268091 228458 268097
rect 228406 268033 228458 268039
rect 227830 267943 227882 267949
rect 227830 267885 227882 267891
rect 227638 267869 227690 267875
rect 227638 267811 227690 267817
rect 227650 263810 227678 267811
rect 227842 263824 227870 267885
rect 228418 263824 228446 268033
rect 227842 263796 228096 263824
rect 228418 263796 228672 263824
rect 229090 263810 229118 268255
rect 229570 263810 229598 269217
rect 230038 268165 230090 268171
rect 230038 268107 230090 268113
rect 230050 263810 230078 268107
rect 230518 268017 230570 268023
rect 230518 267959 230570 267965
rect 230530 264120 230558 267959
rect 230482 264092 230558 264120
rect 230482 263810 230510 264092
rect 231010 263810 231038 269291
rect 231478 268239 231530 268245
rect 231478 268181 231530 268187
rect 231490 263810 231518 268181
rect 231970 263810 231998 269439
rect 232150 269423 232202 269429
rect 232150 269365 232202 269371
rect 232162 263824 232190 269365
rect 232642 263824 232670 271807
rect 233398 269571 233450 269577
rect 233398 269513 233450 269519
rect 232162 263796 232416 263824
rect 232642 263796 232896 263824
rect 233410 263810 233438 269513
rect 233890 263810 233918 272325
rect 234370 263810 234398 272547
rect 234946 272537 234974 278018
rect 235702 272827 235754 272833
rect 235702 272769 235754 272775
rect 235030 272753 235082 272759
rect 235030 272695 235082 272701
rect 234550 272531 234602 272537
rect 234550 272473 234602 272479
rect 234934 272531 234986 272537
rect 234934 272473 234986 272479
rect 234562 263824 234590 272473
rect 235042 263824 235070 272695
rect 234562 263796 234816 263824
rect 235042 263796 235296 263824
rect 235714 263810 235742 272769
rect 236098 272389 236126 278018
rect 236950 273123 237002 273129
rect 236950 273065 237002 273071
rect 236278 272901 236330 272907
rect 236278 272843 236330 272849
rect 236086 272383 236138 272389
rect 236086 272325 236138 272331
rect 236290 263810 236318 272843
rect 236470 272679 236522 272685
rect 236470 272621 236522 272627
rect 236482 263824 236510 272621
rect 236962 263824 236990 273065
rect 237250 271279 237278 278018
rect 238102 273197 238154 273203
rect 238102 273139 238154 273145
rect 237622 272975 237674 272981
rect 237622 272917 237674 272923
rect 237238 271273 237290 271279
rect 237238 271215 237290 271221
rect 236482 263796 236736 263824
rect 236962 263796 237216 263824
rect 237634 263810 237662 272917
rect 238114 263810 238142 273139
rect 238498 271205 238526 278018
rect 238678 273419 238730 273425
rect 238678 273361 238730 273367
rect 238486 271199 238538 271205
rect 238486 271141 238538 271147
rect 238690 263810 238718 273361
rect 239158 273049 239210 273055
rect 239158 272991 239210 272997
rect 239170 263824 239198 272991
rect 239350 271051 239402 271057
rect 239350 270993 239402 270999
rect 239542 271051 239594 271057
rect 239542 270993 239594 270999
rect 239136 263796 239198 263824
rect 239362 263824 239390 270993
rect 239554 270761 239582 270993
rect 239650 270761 239678 278018
rect 240802 271131 240830 278018
rect 240790 271125 240842 271131
rect 240790 271067 240842 271073
rect 241954 271057 241982 278018
rect 242902 273567 242954 273573
rect 242902 273509 242954 273515
rect 242134 272309 242186 272315
rect 242134 272251 242186 272257
rect 241270 271051 241322 271057
rect 241270 270993 241322 270999
rect 241942 271051 241994 271057
rect 241942 270993 241994 270999
rect 240022 270977 240074 270983
rect 240022 270919 240074 270925
rect 239542 270755 239594 270761
rect 239542 270697 239594 270703
rect 239638 270755 239690 270761
rect 239638 270697 239690 270703
rect 239362 263796 239616 263824
rect 240034 263810 240062 270919
rect 240502 270903 240554 270909
rect 240502 270845 240554 270851
rect 240514 263810 240542 270845
rect 241078 270829 241130 270835
rect 241078 270771 241130 270777
rect 241090 263810 241118 270771
rect 241282 263824 241310 270993
rect 242146 263824 242174 272251
rect 242422 272161 242474 272167
rect 242422 272103 242474 272109
rect 241282 263796 241536 263824
rect 242016 263796 242174 263824
rect 242434 263810 242462 272103
rect 242914 263810 242942 273509
rect 243094 272013 243146 272019
rect 243094 271955 243146 271961
rect 243106 263824 243134 271955
rect 243202 270983 243230 278018
rect 243670 272457 243722 272463
rect 243670 272399 243722 272405
rect 243190 270977 243242 270983
rect 243190 270919 243242 270925
rect 243682 263824 243710 272399
rect 244054 271939 244106 271945
rect 244054 271881 244106 271887
rect 244066 263824 244094 271881
rect 244354 270909 244382 278018
rect 244822 272531 244874 272537
rect 244822 272473 244874 272479
rect 244342 270903 244394 270909
rect 244342 270845 244394 270851
rect 243106 263796 243360 263824
rect 243682 263796 243936 263824
rect 244066 263796 244368 263824
rect 244834 263810 244862 272473
rect 245302 272383 245354 272389
rect 245302 272325 245354 272331
rect 245314 263810 245342 272325
rect 245506 270835 245534 278018
rect 245590 271273 245642 271279
rect 245590 271215 245642 271221
rect 245494 270829 245546 270835
rect 245494 270771 245546 270777
rect 245602 263824 245630 271215
rect 246070 271199 246122 271205
rect 246070 271141 246122 271147
rect 246082 263824 246110 271141
rect 246754 270761 246782 278018
rect 247222 271125 247274 271131
rect 247222 271067 247274 271073
rect 246454 270755 246506 270761
rect 246454 270697 246506 270703
rect 246742 270755 246794 270761
rect 246742 270697 246794 270703
rect 246466 263824 246494 270697
rect 245602 263796 245760 263824
rect 246082 263796 246336 263824
rect 246466 263796 246768 263824
rect 247234 263810 247262 271067
rect 247702 271051 247754 271057
rect 247702 270993 247754 270999
rect 247714 263810 247742 270993
rect 247906 268393 247934 278018
rect 247990 270977 248042 270983
rect 247990 270919 248042 270925
rect 247894 268387 247946 268393
rect 247894 268329 247946 268335
rect 248002 263824 248030 270919
rect 248662 270903 248714 270909
rect 248662 270845 248714 270851
rect 248002 263796 248160 263824
rect 248674 263810 248702 270845
rect 249058 269651 249086 278018
rect 250320 278004 250526 278032
rect 249142 270829 249194 270835
rect 249142 270771 249194 270777
rect 250498 270780 250526 278004
rect 249046 269645 249098 269651
rect 249046 269587 249098 269593
rect 249154 263810 249182 270771
rect 249622 270755 249674 270761
rect 250498 270752 250718 270780
rect 249622 270697 249674 270703
rect 249634 263810 249662 270697
rect 250294 269645 250346 269651
rect 250294 269587 250346 269593
rect 249814 268387 249866 268393
rect 249814 268329 249866 268335
rect 249826 263824 249854 268329
rect 250306 263824 250334 269587
rect 250690 263824 250718 270752
rect 251458 263824 251486 278018
rect 252322 278004 252624 278032
rect 252322 263824 252350 278004
rect 253366 269127 253418 269133
rect 253366 269069 253418 269075
rect 253174 268535 253226 268541
rect 253174 268477 253226 268483
rect 252694 268091 252746 268097
rect 252694 268033 252746 268039
rect 252706 263824 252734 268033
rect 253186 263824 253214 268477
rect 249826 263796 250080 263824
rect 250306 263796 250560 263824
rect 250690 263796 250992 263824
rect 251458 263796 251568 263824
rect 252048 263796 252350 263824
rect 252480 263796 252734 263824
rect 252960 263796 253214 263824
rect 253378 263810 253406 269069
rect 253762 268097 253790 278018
rect 253942 270459 253994 270465
rect 253942 270401 253994 270407
rect 253750 268091 253802 268097
rect 253750 268033 253802 268039
rect 253954 263810 253982 270401
rect 254614 268683 254666 268689
rect 254614 268625 254666 268631
rect 254626 263824 254654 268625
rect 255010 268541 255038 278018
rect 255286 270311 255338 270317
rect 255286 270253 255338 270259
rect 254998 268535 255050 268541
rect 254998 268477 255050 268483
rect 255094 268387 255146 268393
rect 255094 268329 255146 268335
rect 255106 263824 255134 268329
rect 254400 263796 254654 263824
rect 254880 263796 255134 263824
rect 255298 263810 255326 270253
rect 255766 269645 255818 269651
rect 255766 269587 255818 269593
rect 255778 263810 255806 269587
rect 256162 269133 256190 278018
rect 257314 270465 257342 278018
rect 257302 270459 257354 270465
rect 257302 270401 257354 270407
rect 256246 269793 256298 269799
rect 256246 269735 256298 269741
rect 256150 269127 256202 269133
rect 256150 269069 256202 269075
rect 256258 263810 256286 269735
rect 257014 269127 257066 269133
rect 257014 269069 257066 269075
rect 257026 263824 257054 269069
rect 258166 268831 258218 268837
rect 258166 268773 258218 268779
rect 257686 268757 257738 268763
rect 257686 268699 257738 268705
rect 257494 268239 257546 268245
rect 257494 268181 257546 268187
rect 257506 263824 257534 268181
rect 256800 263796 257054 263824
rect 257280 263796 257534 263824
rect 257698 263810 257726 268699
rect 258178 263810 258206 268773
rect 258562 268689 258590 278018
rect 258646 269423 258698 269429
rect 258646 269365 258698 269371
rect 258550 268683 258602 268689
rect 258550 268625 258602 268631
rect 258658 263810 258686 269365
rect 259414 268683 259466 268689
rect 259414 268625 259466 268631
rect 259426 263824 259454 268625
rect 259714 268393 259742 278018
rect 260866 270317 260894 278018
rect 262006 270459 262058 270465
rect 262006 270401 262058 270407
rect 260854 270311 260906 270317
rect 260854 270253 260906 270259
rect 261814 269941 261866 269947
rect 261814 269883 261866 269889
rect 261238 269867 261290 269873
rect 261238 269809 261290 269815
rect 259894 269719 259946 269725
rect 259894 269661 259946 269667
rect 259702 268387 259754 268393
rect 259702 268329 259754 268335
rect 259906 263824 259934 269661
rect 260566 269275 260618 269281
rect 260566 269217 260618 269223
rect 260086 268979 260138 268985
rect 260086 268921 260138 268927
rect 259200 263796 259454 263824
rect 259680 263796 259934 263824
rect 260098 263810 260126 268921
rect 260578 263810 260606 269217
rect 261250 263824 261278 269809
rect 261826 263824 261854 269883
rect 261024 263796 261278 263824
rect 261600 263796 261854 263824
rect 262018 263810 262046 270401
rect 262114 269651 262142 278018
rect 262486 270385 262538 270391
rect 262486 270327 262538 270333
rect 262102 269645 262154 269651
rect 262102 269587 262154 269593
rect 262498 263810 262526 270327
rect 262966 270311 263018 270317
rect 262966 270253 263018 270259
rect 262978 263810 263006 270253
rect 263266 269799 263294 278018
rect 263254 269793 263306 269799
rect 263254 269735 263306 269741
rect 264418 269133 264446 278018
rect 264694 270533 264746 270539
rect 264694 270475 264746 270481
rect 264406 269127 264458 269133
rect 264406 269069 264458 269075
rect 264118 268387 264170 268393
rect 264118 268329 264170 268335
rect 263638 268165 263690 268171
rect 263638 268107 263690 268113
rect 263650 263824 263678 268107
rect 264130 263824 264158 268329
rect 264706 263824 264734 270475
rect 264886 270237 264938 270243
rect 264886 270179 264938 270185
rect 263424 263796 263678 263824
rect 263904 263796 264158 263824
rect 264432 263796 264734 263824
rect 264898 263810 264926 270179
rect 265366 270163 265418 270169
rect 265366 270105 265418 270111
rect 265378 263810 265406 270105
rect 265666 268245 265694 278018
rect 266518 270089 266570 270095
rect 266518 270031 266570 270037
rect 266038 269053 266090 269059
rect 266038 268995 266090 269001
rect 265654 268239 265706 268245
rect 265654 268181 265706 268187
rect 266050 263824 266078 268995
rect 266530 263824 266558 270031
rect 266818 268763 266846 278018
rect 267766 269793 267818 269799
rect 267766 269735 267818 269741
rect 267094 269201 267146 269207
rect 267094 269143 267146 269149
rect 266806 268757 266858 268763
rect 266806 268699 266858 268705
rect 267106 263824 267134 269143
rect 267286 268535 267338 268541
rect 267286 268477 267338 268483
rect 265824 263796 266078 263824
rect 266304 263796 266558 263824
rect 266832 263796 267134 263824
rect 267298 263810 267326 268477
rect 267778 263824 267806 269735
rect 267970 268837 267998 278018
rect 269122 269429 269150 278018
rect 270262 273567 270314 273573
rect 270262 273509 270314 273515
rect 269686 269645 269738 269651
rect 269686 269587 269738 269593
rect 269206 269571 269258 269577
rect 269206 269513 269258 269519
rect 269110 269423 269162 269429
rect 269110 269365 269162 269371
rect 268630 269349 268682 269355
rect 268630 269291 268682 269297
rect 268438 269127 268490 269133
rect 268438 269069 268490 269075
rect 267958 268831 268010 268837
rect 267958 268773 268010 268779
rect 268450 263824 268478 269069
rect 267744 263796 267806 263824
rect 268224 263796 268478 263824
rect 268642 263810 268670 269291
rect 269218 263810 269246 269513
rect 269698 263810 269726 269587
rect 270274 263824 270302 273509
rect 270370 268689 270398 278018
rect 270550 272605 270602 272611
rect 270550 272547 270602 272553
rect 270358 268683 270410 268689
rect 270358 268625 270410 268631
rect 270144 263796 270302 263824
rect 270562 263824 270590 272547
rect 271030 272087 271082 272093
rect 271030 272029 271082 272035
rect 270562 263796 270624 263824
rect 271042 263810 271070 272029
rect 271522 269725 271550 278018
rect 272278 272531 272330 272537
rect 272278 272473 272330 272479
rect 271510 269719 271562 269725
rect 271510 269661 271562 269667
rect 271702 269645 271754 269651
rect 271702 269587 271754 269593
rect 271510 269497 271562 269503
rect 271510 269439 271562 269445
rect 271522 263810 271550 269439
rect 271714 269355 271742 269587
rect 271702 269349 271754 269355
rect 271702 269291 271754 269297
rect 272290 263824 272318 272473
rect 272674 268985 272702 278018
rect 272758 272457 272810 272463
rect 272758 272399 272810 272405
rect 272662 268979 272714 268985
rect 272662 268921 272714 268927
rect 272770 263824 272798 272399
rect 273430 272383 273482 272389
rect 273430 272325 273482 272331
rect 272950 269423 273002 269429
rect 272950 269365 273002 269371
rect 272064 263796 272318 263824
rect 272544 263796 272798 263824
rect 272962 263810 272990 269365
rect 273442 263810 273470 272325
rect 273922 269281 273950 278018
rect 274198 272975 274250 272981
rect 274198 272917 274250 272923
rect 273910 269275 273962 269281
rect 273910 269217 273962 269223
rect 274210 263824 274238 272917
rect 275074 269873 275102 278018
rect 275350 273493 275402 273499
rect 275350 273435 275402 273441
rect 275158 272309 275210 272315
rect 275158 272251 275210 272257
rect 275062 269867 275114 269873
rect 275062 269809 275114 269815
rect 274678 268609 274730 268615
rect 274678 268551 274730 268557
rect 274690 263824 274718 268551
rect 275170 263824 275198 272251
rect 275254 269867 275306 269873
rect 275254 269809 275306 269815
rect 275266 269207 275294 269809
rect 275254 269201 275306 269207
rect 275254 269143 275306 269149
rect 273936 263796 274238 263824
rect 274464 263796 274718 263824
rect 274944 263796 275198 263824
rect 275362 263810 275390 273435
rect 276226 269947 276254 278018
rect 277078 273419 277130 273425
rect 277078 273361 277130 273367
rect 276310 272235 276362 272241
rect 276310 272177 276362 272183
rect 276214 269941 276266 269947
rect 276214 269883 276266 269889
rect 275830 268683 275882 268689
rect 275830 268625 275882 268631
rect 275842 263810 275870 268625
rect 276322 263810 276350 272177
rect 276406 269941 276458 269947
rect 276406 269883 276458 269889
rect 276418 269133 276446 269883
rect 276406 269127 276458 269133
rect 276406 269069 276458 269075
rect 277090 263824 277118 273361
rect 277474 270465 277502 278018
rect 278230 273271 278282 273277
rect 278230 273213 278282 273219
rect 277750 272161 277802 272167
rect 277750 272103 277802 272109
rect 277462 270459 277514 270465
rect 277462 270401 277514 270407
rect 277558 269201 277610 269207
rect 277558 269143 277610 269149
rect 277570 263824 277598 269143
rect 276864 263796 277118 263824
rect 277344 263796 277598 263824
rect 277762 263810 277790 272103
rect 278242 263810 278270 273213
rect 278626 270391 278654 278018
rect 279670 273345 279722 273351
rect 279670 273287 279722 273293
rect 279286 270681 279338 270687
rect 279286 270623 279338 270629
rect 278614 270385 278666 270391
rect 278614 270327 278666 270333
rect 278902 269349 278954 269355
rect 278902 269291 278954 269297
rect 278914 263824 278942 269291
rect 279298 263824 279326 270623
rect 278688 263796 278942 263824
rect 279168 263796 279326 263824
rect 279682 263810 279710 273287
rect 279778 270317 279806 278018
rect 280150 270607 280202 270613
rect 280150 270549 280202 270555
rect 279766 270311 279818 270317
rect 279766 270253 279818 270259
rect 280162 263810 280190 270549
rect 280630 270459 280682 270465
rect 280630 270401 280682 270407
rect 280642 263810 280670 270401
rect 281026 268245 281054 278018
rect 281782 274899 281834 274905
rect 281782 274841 281834 274847
rect 281302 269127 281354 269133
rect 281302 269069 281354 269075
rect 281014 268239 281066 268245
rect 281014 268181 281066 268187
rect 281314 263824 281342 269069
rect 281794 263824 281822 274841
rect 282070 268979 282122 268985
rect 282070 268921 282122 268927
rect 281088 263796 281342 263824
rect 281568 263796 281822 263824
rect 282082 263810 282110 268921
rect 282178 268393 282206 278018
rect 283030 274973 283082 274979
rect 283030 274915 283082 274921
rect 282166 268387 282218 268393
rect 282166 268329 282218 268335
rect 282550 267869 282602 267875
rect 282550 267811 282602 267817
rect 282562 263810 282590 267811
rect 283042 263810 283070 274915
rect 283330 270539 283358 278018
rect 284470 276379 284522 276385
rect 284470 276321 284522 276327
rect 283318 270533 283370 270539
rect 283318 270475 283370 270481
rect 283702 270459 283754 270465
rect 283702 270401 283754 270407
rect 283714 263824 283742 270401
rect 284182 270385 284234 270391
rect 284182 270327 284234 270333
rect 284194 263824 284222 270327
rect 283488 263796 283742 263824
rect 283968 263796 284222 263824
rect 284482 263810 284510 276321
rect 284578 270243 284606 278018
rect 285622 273197 285674 273203
rect 285622 273139 285674 273145
rect 284950 271865 285002 271871
rect 284950 271807 285002 271813
rect 284566 270237 284618 270243
rect 284566 270179 284618 270185
rect 284962 263810 284990 271807
rect 285634 263824 285662 273139
rect 285730 270095 285758 278018
rect 286102 276453 286154 276459
rect 286102 276395 286154 276401
rect 285718 270089 285770 270095
rect 285718 270031 285770 270037
rect 286114 263824 286142 276395
rect 286774 273123 286826 273129
rect 286774 273065 286826 273071
rect 286294 270311 286346 270317
rect 286294 270253 286346 270259
rect 285408 263796 285662 263824
rect 285888 263796 286142 263824
rect 286306 263810 286334 270253
rect 286786 263810 286814 273065
rect 286882 269059 286910 278018
rect 287350 276305 287402 276311
rect 287350 276247 287402 276253
rect 286870 269053 286922 269059
rect 286870 268995 286922 269001
rect 287362 263810 287390 276247
rect 287926 270237 287978 270243
rect 287926 270179 287978 270185
rect 287938 263824 287966 270179
rect 288034 270021 288062 278018
rect 288694 276231 288746 276237
rect 288694 276173 288746 276179
rect 288502 270163 288554 270169
rect 288502 270105 288554 270111
rect 288022 270015 288074 270021
rect 288022 269957 288074 269963
rect 288514 263824 288542 270105
rect 287808 263796 287966 263824
rect 288288 263796 288542 263824
rect 288706 263810 288734 276173
rect 289282 269873 289310 278018
rect 290326 276083 290378 276089
rect 290326 276025 290378 276031
rect 289942 273049 289994 273055
rect 289942 272991 289994 272997
rect 289270 269867 289322 269873
rect 289270 269809 289322 269815
rect 289174 268831 289226 268837
rect 289174 268773 289226 268779
rect 289186 263810 289214 268773
rect 289954 263824 289982 272991
rect 290338 263824 290366 276025
rect 290434 268541 290462 278018
rect 290614 270015 290666 270021
rect 290614 269957 290666 269963
rect 290422 268535 290474 268541
rect 290422 268477 290474 268483
rect 289728 263796 289982 263824
rect 290208 263796 290366 263824
rect 290626 263810 290654 269957
rect 291094 269941 291146 269947
rect 291094 269883 291146 269889
rect 291106 263810 291134 269883
rect 291586 269799 291614 278018
rect 291862 276157 291914 276163
rect 291862 276099 291914 276105
rect 291574 269793 291626 269799
rect 291574 269735 291626 269741
rect 291874 263824 291902 276099
rect 292246 272901 292298 272907
rect 292246 272843 292298 272849
rect 292258 263824 292286 272843
rect 292726 272827 292778 272833
rect 292726 272769 292778 272775
rect 292738 263824 292766 272769
rect 292834 270095 292862 278018
rect 293794 278004 294000 278032
rect 293014 276009 293066 276015
rect 293014 275951 293066 275957
rect 292918 270237 292970 270243
rect 292918 270179 292970 270185
rect 292930 270095 292958 270179
rect 292822 270089 292874 270095
rect 292822 270031 292874 270037
rect 292918 270089 292970 270095
rect 292918 270031 292970 270037
rect 291600 263796 291902 263824
rect 292032 263796 292286 263824
rect 292608 263796 292766 263824
rect 293026 263810 293054 275951
rect 293302 270681 293354 270687
rect 293302 270623 293354 270629
rect 293398 270681 293450 270687
rect 293398 270623 293450 270629
rect 293314 270465 293342 270623
rect 293302 270459 293354 270465
rect 293302 270401 293354 270407
rect 293410 269355 293438 270623
rect 293494 269793 293546 269799
rect 293494 269735 293546 269741
rect 293398 269349 293450 269355
rect 293398 269291 293450 269297
rect 293506 263810 293534 269735
rect 293794 269651 293822 278004
rect 294646 275935 294698 275941
rect 294646 275877 294698 275883
rect 293974 269867 294026 269873
rect 293974 269809 294026 269815
rect 293782 269645 293834 269651
rect 293782 269587 293834 269593
rect 293986 263810 294014 269809
rect 294658 263824 294686 275877
rect 295138 269577 295166 278018
rect 295894 275713 295946 275719
rect 295894 275655 295946 275661
rect 295414 272753 295466 272759
rect 295414 272695 295466 272701
rect 295126 269571 295178 269577
rect 295126 269513 295178 269519
rect 295222 268757 295274 268763
rect 295222 268699 295274 268705
rect 295234 263824 295262 268699
rect 294432 263796 294686 263824
rect 295008 263796 295262 263824
rect 295426 263810 295454 272695
rect 295906 263810 295934 275655
rect 296386 269725 296414 278018
rect 296470 275861 296522 275867
rect 296470 275803 296522 275809
rect 296374 269719 296426 269725
rect 296374 269661 296426 269667
rect 296482 263824 296510 275803
rect 297334 275787 297386 275793
rect 297334 275729 297386 275735
rect 297046 269719 297098 269725
rect 297046 269661 297098 269667
rect 297058 263824 297086 269661
rect 296352 263796 296510 263824
rect 296832 263796 297086 263824
rect 297346 263810 297374 275729
rect 297538 273573 297566 278018
rect 297814 275565 297866 275571
rect 297814 275507 297866 275513
rect 297526 273567 297578 273573
rect 297526 273509 297578 273515
rect 297826 263810 297854 275507
rect 298294 272753 298346 272759
rect 298294 272695 298346 272701
rect 298306 263810 298334 272695
rect 298690 272611 298718 278018
rect 298966 275639 299018 275645
rect 298966 275581 299018 275587
rect 298678 272605 298730 272611
rect 298678 272547 298730 272553
rect 298978 263824 299006 275581
rect 299158 275417 299210 275423
rect 299158 275359 299210 275365
rect 298752 263796 299006 263824
rect 299170 263676 299198 275359
rect 299350 273567 299402 273573
rect 299350 273509 299402 273515
rect 299362 268985 299390 273509
rect 299938 272093 299966 278018
rect 300214 275491 300266 275497
rect 300214 275433 300266 275439
rect 299926 272087 299978 272093
rect 299926 272029 299978 272035
rect 299446 272013 299498 272019
rect 299446 271955 299498 271961
rect 299350 268979 299402 268985
rect 299350 268921 299402 268927
rect 299458 267875 299486 271955
rect 299638 269645 299690 269651
rect 299638 269587 299690 269593
rect 299446 267869 299498 267875
rect 299446 267811 299498 267817
rect 299650 263810 299678 269587
rect 300226 263810 300254 275433
rect 301090 269503 301118 278018
rect 301954 278004 302256 278032
rect 301366 272605 301418 272611
rect 301366 272547 301418 272553
rect 301078 269497 301130 269503
rect 301078 269439 301130 269445
rect 300694 268905 300746 268911
rect 300694 268847 300746 268853
rect 300706 263810 300734 268847
rect 301378 263824 301406 272547
rect 301954 272537 301982 278004
rect 303286 275343 303338 275349
rect 303286 275285 303338 275291
rect 302050 272685 302366 272704
rect 302038 272679 302378 272685
rect 302090 272676 302326 272679
rect 302038 272621 302090 272627
rect 302326 272621 302378 272627
rect 301942 272531 301994 272537
rect 301942 272473 301994 272479
rect 302326 272013 302378 272019
rect 302326 271955 302378 271961
rect 302338 269133 302366 271955
rect 302614 269571 302666 269577
rect 302614 269513 302666 269519
rect 302326 269127 302378 269133
rect 302326 269069 302378 269075
rect 302038 268979 302090 268985
rect 302038 268921 302090 268927
rect 301846 266907 301898 266913
rect 301846 266849 301898 266855
rect 301858 263824 301886 266849
rect 301152 263796 301406 263824
rect 301632 263796 301886 263824
rect 302050 263810 302078 268921
rect 302626 263810 302654 269513
rect 303298 263824 303326 275285
rect 303490 272463 303518 278018
rect 304438 275269 304490 275275
rect 304438 275211 304490 275217
rect 303478 272457 303530 272463
rect 303478 272399 303530 272405
rect 303958 271939 304010 271945
rect 303958 271881 304010 271887
rect 303766 269053 303818 269059
rect 303766 268995 303818 269001
rect 303778 263824 303806 268995
rect 303072 263796 303326 263824
rect 303552 263796 303806 263824
rect 303970 263810 303998 271881
rect 304450 263810 304478 275211
rect 304642 269429 304670 278018
rect 305302 273567 305354 273573
rect 305302 273509 305354 273515
rect 305314 272981 305342 273509
rect 305302 272975 305354 272981
rect 305302 272917 305354 272923
rect 305794 272389 305822 278018
rect 306946 273573 306974 278018
rect 307318 275195 307370 275201
rect 307318 275137 307370 275143
rect 306934 273567 306986 273573
rect 306934 273509 306986 273515
rect 306646 273123 306698 273129
rect 306646 273065 306698 273071
rect 305782 272383 305834 272389
rect 305782 272325 305834 272331
rect 306658 271871 306686 273065
rect 306838 272975 306890 272981
rect 306838 272917 306890 272923
rect 306646 271865 306698 271871
rect 306646 271807 306698 271813
rect 305686 269497 305738 269503
rect 305686 269439 305738 269445
rect 304630 269423 304682 269429
rect 304630 269365 304682 269371
rect 305014 266833 305066 266839
rect 305014 266775 305066 266781
rect 305026 263810 305054 266775
rect 305698 263824 305726 269439
rect 306358 269127 306410 269133
rect 306358 269069 306410 269075
rect 306166 266759 306218 266765
rect 306166 266701 306218 266707
rect 306178 263824 306206 266701
rect 305472 263796 305726 263824
rect 305952 263796 306206 263824
rect 306370 263810 306398 269069
rect 306850 268763 306878 272917
rect 307126 272457 307178 272463
rect 307126 272399 307178 272405
rect 306838 268757 306890 268763
rect 306838 268699 306890 268705
rect 307138 263824 307166 272399
rect 306864 263796 307166 263824
rect 307330 263810 307358 275137
rect 308194 268615 308222 278018
rect 309346 272315 309374 278018
rect 310390 275121 310442 275127
rect 310390 275063 310442 275069
rect 309910 272383 309962 272389
rect 309910 272325 309962 272331
rect 309334 272309 309386 272315
rect 309334 272251 309386 272257
rect 308278 269423 308330 269429
rect 308278 269365 308330 269371
rect 308182 268609 308234 268615
rect 308182 268551 308234 268557
rect 308086 266685 308138 266691
rect 308086 266627 308138 266633
rect 308098 263824 308126 266627
rect 307872 263796 308126 263824
rect 308290 263810 308318 269365
rect 309238 268313 309290 268319
rect 309238 268255 309290 268261
rect 308758 266611 308810 266617
rect 308758 266553 308810 266559
rect 308770 263810 308798 266553
rect 309250 263810 309278 268255
rect 309922 263824 309950 272325
rect 310402 263824 310430 275063
rect 310498 273499 310526 278018
rect 311638 275047 311690 275053
rect 311638 274989 311690 274995
rect 310486 273493 310538 273499
rect 310486 273435 310538 273441
rect 310582 273493 310634 273499
rect 310582 273435 310634 273441
rect 310594 268837 310622 273435
rect 311158 269349 311210 269355
rect 311158 269291 311210 269297
rect 310582 268831 310634 268837
rect 310582 268773 310634 268779
rect 310678 266537 310730 266543
rect 310678 266479 310730 266485
rect 309696 263796 309950 263824
rect 310272 263796 310430 263824
rect 310690 263810 310718 266479
rect 311170 263810 311198 269291
rect 311650 263810 311678 274989
rect 311746 268689 311774 278018
rect 312790 272309 312842 272315
rect 312790 272251 312842 272257
rect 311734 268683 311786 268689
rect 311734 268625 311786 268631
rect 312310 268239 312362 268245
rect 312310 268181 312362 268187
rect 312322 263824 312350 268181
rect 312802 263824 312830 272251
rect 312898 272241 312926 278018
rect 314050 273425 314078 278018
rect 314710 274159 314762 274165
rect 314710 274101 314762 274107
rect 314038 273419 314090 273425
rect 314038 273361 314090 273367
rect 312886 272235 312938 272241
rect 312886 272177 312938 272183
rect 314230 269275 314282 269281
rect 314230 269217 314282 269223
rect 313078 266463 313130 266469
rect 313078 266405 313130 266411
rect 312096 263796 312350 263824
rect 312672 263796 312830 263824
rect 313090 263810 313118 266405
rect 313558 266389 313610 266395
rect 313558 266331 313610 266337
rect 313570 263810 313598 266331
rect 314242 263824 314270 269217
rect 314722 263824 314750 274101
rect 314016 263796 314270 263824
rect 314496 263796 314750 263824
rect 314914 263810 314942 278319
rect 381046 278303 381098 278309
rect 408322 278300 408624 278319
rect 571426 278309 571728 278328
rect 571414 278303 571728 278309
rect 381046 278245 381098 278251
rect 571466 278300 571728 278303
rect 571414 278245 571466 278251
rect 319510 278229 319562 278235
rect 319510 278171 319562 278177
rect 315298 269207 315326 278018
rect 315958 274307 316010 274313
rect 315958 274249 316010 274255
rect 315478 272161 315530 272167
rect 315478 272103 315530 272109
rect 315286 269201 315338 269207
rect 315286 269143 315338 269149
rect 315490 263810 315518 272103
rect 315970 263810 315998 274249
rect 316450 272241 316478 278018
rect 316630 276897 316682 276903
rect 316630 276839 316682 276845
rect 316438 272235 316490 272241
rect 316438 272177 316490 272183
rect 316642 263824 316670 276839
rect 317302 274233 317354 274239
rect 317302 274175 317354 274181
rect 317110 268387 317162 268393
rect 317110 268329 317162 268335
rect 317122 263824 317150 268329
rect 316416 263796 316670 263824
rect 316896 263796 317150 263824
rect 317314 263810 317342 274175
rect 317602 273277 317630 278018
rect 317878 277785 317930 277791
rect 317878 277727 317930 277733
rect 317590 273271 317642 273277
rect 317590 273213 317642 273219
rect 317890 263810 317918 277727
rect 318358 271273 318410 271279
rect 318358 271215 318410 271221
rect 318370 263810 318398 271215
rect 318850 270687 318878 278018
rect 318838 270681 318890 270687
rect 318838 270623 318890 270629
rect 319030 265501 319082 265507
rect 319030 265443 319082 265449
rect 319042 263824 319070 265443
rect 319522 263824 319550 278171
rect 320950 278155 321002 278161
rect 320950 278097 321002 278103
rect 320002 270465 320030 278018
rect 320182 274381 320234 274387
rect 320182 274323 320234 274329
rect 319990 270459 320042 270465
rect 319990 270401 320042 270407
rect 319702 268461 319754 268467
rect 319702 268403 319754 268409
rect 318816 263796 319070 263824
rect 319296 263796 319550 263824
rect 319714 263810 319742 268403
rect 320194 263810 320222 274323
rect 320962 263824 320990 278097
rect 321154 273351 321182 278018
rect 322102 276601 322154 276607
rect 322102 276543 322154 276549
rect 321142 273345 321194 273351
rect 321142 273287 321194 273293
rect 321430 271347 321482 271353
rect 321430 271289 321482 271295
rect 321442 263824 321470 271289
rect 321622 265575 321674 265581
rect 321622 265517 321674 265523
rect 320736 263796 320990 263824
rect 321216 263796 321470 263824
rect 321634 263810 321662 265517
rect 322114 263810 322142 276543
rect 322402 270613 322430 278018
rect 323350 274455 323402 274461
rect 323350 274397 323402 274403
rect 322390 270607 322442 270613
rect 322390 270549 322442 270555
rect 322582 268535 322634 268541
rect 322582 268477 322634 268483
rect 322594 263810 322622 268477
rect 323362 263824 323390 274397
rect 323554 270539 323582 278018
rect 323830 278007 323882 278013
rect 323830 277949 323882 277955
rect 323542 270533 323594 270539
rect 323542 270475 323594 270481
rect 323842 263824 323870 277949
rect 324706 272019 324734 278018
rect 325858 274905 325886 278018
rect 326422 277859 326474 277865
rect 326422 277801 326474 277807
rect 325846 274899 325898 274905
rect 325846 274841 325898 274847
rect 325942 274529 325994 274535
rect 325942 274471 325994 274477
rect 324694 272013 324746 272019
rect 324694 271955 324746 271961
rect 324022 271421 324074 271427
rect 324022 271363 324074 271369
rect 323136 263796 323390 263824
rect 323616 263796 323870 263824
rect 324034 263810 324062 271363
rect 325750 268609 325802 268615
rect 325750 268551 325802 268557
rect 324502 265649 324554 265655
rect 324502 265591 324554 265597
rect 324514 263810 324542 265591
rect 325366 264761 325418 264767
rect 325366 264703 325418 264709
rect 325378 263824 325406 264703
rect 325762 263824 325790 268551
rect 325008 263796 325406 263824
rect 325536 263796 325790 263824
rect 325954 263810 325982 274471
rect 326434 263810 326462 277801
rect 326806 273937 326858 273943
rect 326806 273879 326858 273885
rect 326818 268911 326846 273879
rect 327106 273573 327134 278018
rect 327094 273567 327146 273573
rect 327094 273509 327146 273515
rect 326902 272457 326954 272463
rect 326902 272399 326954 272405
rect 326914 271945 326942 272399
rect 328258 272093 328286 278018
rect 329302 277711 329354 277717
rect 329302 277653 329354 277659
rect 328822 274603 328874 274609
rect 328822 274545 328874 274551
rect 328246 272087 328298 272093
rect 328246 272029 328298 272035
rect 326902 271939 326954 271945
rect 326902 271881 326954 271887
rect 326902 271495 326954 271501
rect 326902 271437 326954 271443
rect 326806 268905 326858 268911
rect 326806 268847 326858 268853
rect 326914 263810 326942 271437
rect 328342 268683 328394 268689
rect 328342 268625 328394 268631
rect 327574 265723 327626 265729
rect 327574 265665 327626 265671
rect 327586 263824 327614 265665
rect 328054 264539 328106 264545
rect 328054 264481 328106 264487
rect 328066 263824 328094 264481
rect 327360 263796 327614 263824
rect 327840 263796 328094 263824
rect 328354 263810 328382 268625
rect 328834 263810 328862 274545
rect 329314 263810 329342 277653
rect 329410 274979 329438 278018
rect 329398 274973 329450 274979
rect 329398 274915 329450 274921
rect 330454 274677 330506 274683
rect 330454 274619 330506 274625
rect 329974 271569 330026 271575
rect 329974 271511 330026 271517
rect 329986 263824 330014 271511
rect 330466 263824 330494 274619
rect 330658 270391 330686 278018
rect 331222 273715 331274 273721
rect 331222 273657 331274 273663
rect 330646 270385 330698 270391
rect 330646 270327 330698 270333
rect 331234 268985 331262 273657
rect 331810 270317 331838 278018
rect 332374 277637 332426 277643
rect 332374 277579 332426 277585
rect 331798 270311 331850 270317
rect 331798 270253 331850 270259
rect 331222 268979 331274 268985
rect 331222 268921 331274 268927
rect 331222 268757 331274 268763
rect 331222 268699 331274 268705
rect 330742 268165 330794 268171
rect 330742 268107 330794 268113
rect 329760 263796 330014 263824
rect 330240 263796 330494 263824
rect 330754 263810 330782 268107
rect 331234 263810 331262 268699
rect 331894 265871 331946 265877
rect 331894 265813 331946 265819
rect 331906 263824 331934 265813
rect 332386 263824 332414 277579
rect 332962 276385 332990 278018
rect 332950 276379 333002 276385
rect 332950 276321 333002 276327
rect 333142 274751 333194 274757
rect 333142 274693 333194 274699
rect 332566 271643 332618 271649
rect 332566 271585 332618 271591
rect 331680 263796 331934 263824
rect 332160 263796 332414 263824
rect 332578 263810 332606 271585
rect 333154 263810 333182 274693
rect 334210 273129 334238 278018
rect 334966 277563 335018 277569
rect 334966 277505 335018 277511
rect 334294 273863 334346 273869
rect 334294 273805 334346 273811
rect 334198 273123 334250 273129
rect 334198 273065 334250 273071
rect 334102 271051 334154 271057
rect 334102 270993 334154 270999
rect 334114 270243 334142 270993
rect 334102 270237 334154 270243
rect 334102 270179 334154 270185
rect 334306 269059 334334 273805
rect 334294 269053 334346 269059
rect 334294 268995 334346 269001
rect 334294 268831 334346 268837
rect 334294 268773 334346 268779
rect 333622 268091 333674 268097
rect 333622 268033 333674 268039
rect 333634 263810 333662 268033
rect 334306 263824 334334 268773
rect 334774 265945 334826 265951
rect 334774 265887 334826 265893
rect 334786 263824 334814 265887
rect 334080 263796 334334 263824
rect 334560 263796 334814 263824
rect 334978 263810 335006 277505
rect 335362 273203 335390 278018
rect 336514 276459 336542 278018
rect 336502 276453 336554 276459
rect 336502 276395 336554 276401
rect 336022 274825 336074 274831
rect 336022 274767 336074 274773
rect 335350 273197 335402 273203
rect 335350 273139 335402 273145
rect 335446 271717 335498 271723
rect 335446 271659 335498 271665
rect 335458 263810 335486 271659
rect 336034 263810 336062 274767
rect 337762 271057 337790 278018
rect 337846 277489 337898 277495
rect 337846 277431 337898 277437
rect 337750 271051 337802 271057
rect 337750 270993 337802 270999
rect 336886 268905 336938 268911
rect 336886 268847 336938 268853
rect 336694 268017 336746 268023
rect 336694 267959 336746 267965
rect 336706 263824 336734 267959
rect 336480 263796 336734 263824
rect 336898 263824 336926 268847
rect 337366 266019 337418 266025
rect 337366 265961 337418 265967
rect 336898 263796 336960 263824
rect 337378 263810 337406 265961
rect 337858 263810 337886 277431
rect 338914 273055 338942 278018
rect 340066 276311 340094 278018
rect 341014 277415 341066 277421
rect 341014 277357 341066 277363
rect 340054 276305 340106 276311
rect 340054 276247 340106 276253
rect 339094 274899 339146 274905
rect 339094 274841 339146 274847
rect 338902 273049 338954 273055
rect 338902 272991 338954 272997
rect 338614 271199 338666 271205
rect 338614 271141 338666 271147
rect 338626 263824 338654 271141
rect 338710 270903 338762 270909
rect 338710 270845 338762 270851
rect 338722 270095 338750 270845
rect 338710 270089 338762 270095
rect 338710 270031 338762 270037
rect 339106 263824 339134 274841
rect 339766 268979 339818 268985
rect 339766 268921 339818 268927
rect 339286 267943 339338 267949
rect 339286 267885 339338 267891
rect 338400 263796 338654 263824
rect 338880 263796 339134 263824
rect 339298 263810 339326 267885
rect 339778 263810 339806 268921
rect 340246 266093 340298 266099
rect 340246 266035 340298 266041
rect 340258 263810 340286 266035
rect 341026 263824 341054 277357
rect 341206 274011 341258 274017
rect 341206 273953 341258 273959
rect 341218 269133 341246 273953
rect 341314 270909 341342 278018
rect 341684 274494 341740 274503
rect 341684 274429 341740 274438
rect 341494 271791 341546 271797
rect 341494 271733 341546 271739
rect 341302 270903 341354 270909
rect 341302 270845 341354 270851
rect 341206 269127 341258 269133
rect 341206 269069 341258 269075
rect 341506 263824 341534 271733
rect 340800 263796 341054 263824
rect 341280 263796 341534 263824
rect 341698 263810 341726 274429
rect 342466 270169 342494 278018
rect 343618 276237 343646 278018
rect 343894 277341 343946 277347
rect 343894 277283 343946 277289
rect 343606 276231 343658 276237
rect 343606 276173 343658 276179
rect 342742 270829 342794 270835
rect 342742 270771 342794 270777
rect 342454 270163 342506 270169
rect 342454 270105 342506 270111
rect 342754 270021 342782 270771
rect 342742 270015 342794 270021
rect 342742 269957 342794 269963
rect 342646 269053 342698 269059
rect 342646 268995 342698 269001
rect 342166 267869 342218 267875
rect 342166 267811 342218 267817
rect 342178 263810 342206 267811
rect 342658 263810 342686 268995
rect 343798 268165 343850 268171
rect 343798 268107 343850 268113
rect 343318 266167 343370 266173
rect 343318 266109 343370 266115
rect 343330 263824 343358 266109
rect 343810 264471 343838 268107
rect 343798 264465 343850 264471
rect 343798 264407 343850 264413
rect 343906 263824 343934 277283
rect 344566 274973 344618 274979
rect 344566 274915 344618 274921
rect 344086 271939 344138 271945
rect 344086 271881 344138 271887
rect 343104 263796 343358 263824
rect 343632 263796 343934 263824
rect 344098 263810 344126 271881
rect 344578 263810 344606 274915
rect 344770 273499 344798 278018
rect 344758 273493 344810 273499
rect 344758 273435 344810 273441
rect 346018 272907 346046 278018
rect 347170 276089 347198 278018
rect 347158 276083 347210 276089
rect 347158 276025 347210 276031
rect 347636 274642 347692 274651
rect 347636 274577 347692 274586
rect 347062 273789 347114 273795
rect 347062 273731 347114 273737
rect 346006 272901 346058 272907
rect 346006 272843 346058 272849
rect 346966 272087 347018 272093
rect 346966 272029 347018 272035
rect 346486 272013 346538 272019
rect 346486 271955 346538 271961
rect 345430 269201 345482 269207
rect 345430 269143 345482 269149
rect 345238 269127 345290 269133
rect 345238 269069 345290 269075
rect 345250 263824 345278 269069
rect 345024 263796 345278 263824
rect 345442 263676 345470 269143
rect 346006 266241 346058 266247
rect 346006 266183 346058 266189
rect 346018 263810 346046 266183
rect 346498 263810 346526 271955
rect 346978 263810 347006 272029
rect 347074 268319 347102 273731
rect 347062 268313 347114 268319
rect 347062 268255 347114 268261
rect 347650 263824 347678 274577
rect 348322 270835 348350 278018
rect 348502 274085 348554 274091
rect 348502 274027 348554 274033
rect 348310 270829 348362 270835
rect 348310 270771 348362 270777
rect 348118 270681 348170 270687
rect 348118 270623 348170 270629
rect 348130 263824 348158 270623
rect 348406 270607 348458 270613
rect 348406 270549 348458 270555
rect 347424 263796 347678 263824
rect 347904 263796 348158 263824
rect 348418 263810 348446 270549
rect 348514 268245 348542 274027
rect 349462 273567 349514 273573
rect 349462 273509 349514 273515
rect 348502 268239 348554 268245
rect 348502 268181 348554 268187
rect 348886 266315 348938 266321
rect 348886 266257 348938 266263
rect 348898 263810 348926 266257
rect 349474 263824 349502 273509
rect 349570 269947 349598 278018
rect 350722 276163 350750 278018
rect 350710 276157 350762 276163
rect 350710 276099 350762 276105
rect 350228 274790 350284 274799
rect 350228 274725 350284 274734
rect 350038 273493 350090 273499
rect 350038 273435 350090 273441
rect 349558 269941 349610 269947
rect 349558 269883 349610 269889
rect 350050 263824 350078 273435
rect 349344 263796 349502 263824
rect 349824 263796 350078 263824
rect 350242 263810 350270 274725
rect 351874 272833 351902 278018
rect 352438 273419 352490 273425
rect 352438 273361 352490 273367
rect 351862 272827 351914 272833
rect 351862 272769 351914 272775
rect 351382 271865 351434 271871
rect 351382 271807 351434 271813
rect 350710 270533 350762 270539
rect 350710 270475 350762 270481
rect 350722 263810 350750 270475
rect 351286 270459 351338 270465
rect 351286 270401 351338 270407
rect 351298 263810 351326 270401
rect 351394 269799 351422 271807
rect 351382 269793 351434 269799
rect 351382 269735 351434 269741
rect 351382 268091 351434 268097
rect 351382 268033 351434 268039
rect 351394 264397 351422 268033
rect 351958 267721 352010 267727
rect 351958 267663 352010 267669
rect 351382 264391 351434 264397
rect 351382 264333 351434 264339
rect 351970 263824 351998 267663
rect 352450 263824 352478 273361
rect 352630 273345 352682 273351
rect 352630 273287 352682 273293
rect 351744 263796 351998 263824
rect 352224 263796 352478 263824
rect 352642 263810 352670 273287
rect 353122 272759 353150 278018
rect 354274 276015 354302 278018
rect 354262 276009 354314 276015
rect 354262 275951 354314 275957
rect 353396 274938 353452 274947
rect 353396 274873 353452 274882
rect 353110 272753 353162 272759
rect 353110 272695 353162 272701
rect 353410 263824 353438 274873
rect 355030 273197 355082 273203
rect 355030 273139 355082 273145
rect 354070 270385 354122 270391
rect 354070 270327 354122 270333
rect 353686 270311 353738 270317
rect 353686 270253 353738 270259
rect 353136 263796 353438 263824
rect 353698 263810 353726 270253
rect 354082 264120 354110 270327
rect 354838 267647 354890 267653
rect 354838 267589 354890 267595
rect 354082 264092 354158 264120
rect 354130 263810 354158 264092
rect 354850 263824 354878 267589
rect 354624 263796 354878 263824
rect 355042 263810 355070 273139
rect 355426 271871 355454 278018
rect 356182 276453 356234 276459
rect 356182 276395 356234 276401
rect 355510 273271 355562 273277
rect 355510 273213 355562 273219
rect 355414 271865 355466 271871
rect 355414 271807 355466 271813
rect 355522 263810 355550 273213
rect 355606 271791 355658 271797
rect 355606 271733 355658 271739
rect 355618 271205 355646 271733
rect 355606 271199 355658 271205
rect 355606 271141 355658 271147
rect 356194 263824 356222 276395
rect 356674 269873 356702 278018
rect 357826 275941 357854 278018
rect 357814 275935 357866 275941
rect 357814 275877 357866 275883
rect 358582 273123 358634 273129
rect 358582 273065 358634 273071
rect 357910 271199 357962 271205
rect 357910 271141 357962 271147
rect 356758 270237 356810 270243
rect 356758 270179 356810 270185
rect 356662 269867 356714 269873
rect 356662 269809 356714 269815
rect 356770 263824 356798 270179
rect 356950 270163 357002 270169
rect 356950 270105 357002 270111
rect 355968 263796 356222 263824
rect 356544 263796 356798 263824
rect 356962 263810 356990 270105
rect 357622 268017 357674 268023
rect 357622 267959 357674 267965
rect 357430 267573 357482 267579
rect 357430 267515 357482 267521
rect 357442 263810 357470 267515
rect 357634 264619 357662 267959
rect 357622 264613 357674 264619
rect 357622 264555 357674 264561
rect 357922 263810 357950 271141
rect 358594 263824 358622 273065
rect 358978 272981 359006 278018
rect 359158 276379 359210 276385
rect 359158 276321 359210 276327
rect 358966 272975 359018 272981
rect 358966 272917 359018 272923
rect 359170 263824 359198 276321
rect 360226 272685 360254 278018
rect 361378 275719 361406 278018
rect 361750 276305 361802 276311
rect 361750 276247 361802 276253
rect 361366 275713 361418 275719
rect 361366 275655 361418 275661
rect 360982 273049 361034 273055
rect 360982 272991 361034 272997
rect 360214 272679 360266 272685
rect 360214 272621 360266 272627
rect 359830 270089 359882 270095
rect 359830 270031 359882 270037
rect 359350 270015 359402 270021
rect 359350 269957 359402 269963
rect 358368 263796 358622 263824
rect 358944 263796 359198 263824
rect 359362 263810 359390 269957
rect 359842 263810 359870 270031
rect 360310 267499 360362 267505
rect 360310 267441 360362 267447
rect 360322 263810 360350 267441
rect 360994 263824 361022 272991
rect 361270 272975 361322 272981
rect 361270 272917 361322 272923
rect 360768 263796 361022 263824
rect 361282 263810 361310 272917
rect 361762 263810 361790 276247
rect 362530 275867 362558 278018
rect 362518 275861 362570 275867
rect 362518 275803 362570 275809
rect 363574 272901 363626 272907
rect 363574 272843 363626 272849
rect 362710 269941 362762 269947
rect 362710 269883 362762 269889
rect 362230 269867 362282 269873
rect 362230 269809 362282 269815
rect 362242 263810 362270 269809
rect 362722 263824 362750 269883
rect 362806 267943 362858 267949
rect 362806 267885 362858 267891
rect 362818 264693 362846 267885
rect 363382 267425 363434 267431
rect 363382 267367 363434 267373
rect 362806 264687 362858 264693
rect 362806 264629 362858 264635
rect 363394 263824 363422 267367
rect 362688 263796 362750 263824
rect 363168 263796 363422 263824
rect 363586 263810 363614 272843
rect 363682 269725 363710 278018
rect 364630 276231 364682 276237
rect 364630 276173 364682 276179
rect 364150 272827 364202 272833
rect 364150 272769 364202 272775
rect 363670 269719 363722 269725
rect 363670 269661 363722 269667
rect 364162 263810 364190 272769
rect 364642 263810 364670 276173
rect 364930 275793 364958 278018
rect 364918 275787 364970 275793
rect 364918 275729 364970 275735
rect 366082 275571 366110 278018
rect 366070 275565 366122 275571
rect 366070 275507 366122 275513
rect 366550 272753 366602 272759
rect 366550 272695 366602 272701
rect 365302 269793 365354 269799
rect 365302 269735 365354 269741
rect 365314 263824 365342 269735
rect 365494 269719 365546 269725
rect 365494 269661 365546 269667
rect 365088 263796 365342 263824
rect 365506 263824 365534 269661
rect 365686 267869 365738 267875
rect 365686 267811 365738 267817
rect 365698 264841 365726 267811
rect 365974 267351 366026 267357
rect 365974 267293 366026 267299
rect 365686 264835 365738 264841
rect 365686 264777 365738 264783
rect 365506 263796 365568 263824
rect 365986 263810 366014 267293
rect 366562 263810 366590 272695
rect 367126 272679 367178 272685
rect 367126 272621 367178 272627
rect 367138 263824 367166 272621
rect 367234 272611 367262 278018
rect 367702 276157 367754 276163
rect 367702 276099 367754 276105
rect 367222 272605 367274 272611
rect 367222 272547 367274 272553
rect 367714 263824 367742 276099
rect 368482 275645 368510 278018
rect 368470 275639 368522 275645
rect 368470 275581 368522 275587
rect 369634 275423 369662 278018
rect 370294 275935 370346 275941
rect 370294 275877 370346 275883
rect 369622 275417 369674 275423
rect 369622 275359 369674 275365
rect 370100 271682 370156 271691
rect 370100 271617 370156 271626
rect 369620 271534 369676 271543
rect 369620 271469 369676 271478
rect 367892 270498 367948 270507
rect 367892 270433 367948 270442
rect 367008 263796 367166 263824
rect 367488 263796 367742 263824
rect 367906 263810 367934 270433
rect 368372 269166 368428 269175
rect 368372 269101 368428 269110
rect 368386 263810 368414 269101
rect 368950 267277 369002 267283
rect 368950 267219 369002 267225
rect 368962 263810 368990 267219
rect 369634 263824 369662 271469
rect 370114 263824 370142 271617
rect 369408 263796 369662 263824
rect 369888 263796 370142 263824
rect 370306 263810 370334 275877
rect 370786 269651 370814 278018
rect 371926 276083 371978 276089
rect 371926 276025 371978 276031
rect 371062 276009 371114 276015
rect 371062 275951 371114 275957
rect 370774 269645 370826 269651
rect 370774 269587 370826 269593
rect 371074 263824 371102 275951
rect 371254 268165 371306 268171
rect 371254 268107 371306 268113
rect 370800 263796 371102 263824
rect 371266 263810 371294 268107
rect 371938 263824 371966 276025
rect 372034 275497 372062 278018
rect 372022 275491 372074 275497
rect 372022 275433 372074 275439
rect 373186 273943 373214 278018
rect 373846 277267 373898 277273
rect 373846 277209 373898 277215
rect 373462 275861 373514 275867
rect 373462 275803 373514 275809
rect 373174 273937 373226 273943
rect 373174 273879 373226 273885
rect 372694 272605 372746 272611
rect 372694 272547 372746 272553
rect 372502 267203 372554 267209
rect 372502 267145 372554 267151
rect 372514 263824 372542 267145
rect 371808 263796 371966 263824
rect 372288 263796 372542 263824
rect 372706 263810 372734 272547
rect 373474 263824 373502 275803
rect 373858 263824 373886 277209
rect 374338 272537 374366 278018
rect 375298 278004 375600 278032
rect 375094 277193 375146 277199
rect 375094 277135 375146 277141
rect 374614 275787 374666 275793
rect 374614 275729 374666 275735
rect 374518 272753 374570 272759
rect 374518 272695 374570 272701
rect 374530 272611 374558 272695
rect 374518 272605 374570 272611
rect 374518 272547 374570 272553
rect 374326 272531 374378 272537
rect 374326 272473 374378 272479
rect 374324 268870 374380 268879
rect 374324 268805 374380 268814
rect 374338 263824 374366 268805
rect 373200 263796 373502 263824
rect 373632 263796 373886 263824
rect 374208 263796 374366 263824
rect 374626 263810 374654 275729
rect 375106 263810 375134 277135
rect 375190 273123 375242 273129
rect 375190 273065 375242 273071
rect 375202 271205 375230 273065
rect 375190 271199 375242 271205
rect 375190 271141 375242 271147
rect 375298 266913 375326 278004
rect 376246 275639 376298 275645
rect 376246 275581 376298 275587
rect 375572 271830 375628 271839
rect 375572 271765 375628 271774
rect 375286 266907 375338 266913
rect 375286 266849 375338 266855
rect 375586 263810 375614 271765
rect 376258 263824 376286 275581
rect 376738 273721 376766 278018
rect 376822 277119 376874 277125
rect 376822 277061 376874 277067
rect 376726 273715 376778 273721
rect 376726 273657 376778 273663
rect 376834 263824 376862 277061
rect 377494 275713 377546 275719
rect 377494 275655 377546 275661
rect 377012 270350 377068 270359
rect 377012 270285 377068 270294
rect 376032 263796 376286 263824
rect 376608 263796 376862 263824
rect 377026 263810 377054 270285
rect 377506 263810 377534 275655
rect 377890 269577 377918 278018
rect 377974 277045 378026 277051
rect 377974 276987 378026 276993
rect 377878 269571 377930 269577
rect 377878 269513 377930 269519
rect 377986 263810 378014 276987
rect 379028 276122 379084 276131
rect 379028 276057 379084 276066
rect 378644 271978 378700 271987
rect 378644 271913 378700 271922
rect 378658 263824 378686 271913
rect 379042 263824 379070 276057
rect 379138 275349 379166 278018
rect 379414 276971 379466 276977
rect 379414 276913 379466 276919
rect 379126 275343 379178 275349
rect 379126 275285 379178 275291
rect 378432 263796 378686 263824
rect 378912 263796 379070 263824
rect 379426 263810 379454 276913
rect 380290 273869 380318 278018
rect 380566 275565 380618 275571
rect 380566 275507 380618 275513
rect 380278 273863 380330 273869
rect 380278 273805 380330 273811
rect 379894 269571 379946 269577
rect 379894 269513 379946 269519
rect 379606 269497 379658 269503
rect 379658 269445 379838 269448
rect 379606 269439 379838 269445
rect 379618 269429 379838 269439
rect 379618 269423 379850 269429
rect 379618 269420 379798 269423
rect 379798 269365 379850 269371
rect 379906 263810 379934 269513
rect 380578 263824 380606 275507
rect 381058 263824 381086 278245
rect 418966 278229 419018 278235
rect 419018 278177 419280 278180
rect 418966 278171 419280 278177
rect 418978 278152 419280 278171
rect 422530 278161 422832 278180
rect 422518 278155 422832 278161
rect 422570 278152 422832 278155
rect 422518 278097 422570 278103
rect 386518 278081 386570 278087
rect 381442 272463 381470 278018
rect 382390 277933 382442 277939
rect 382390 277875 382442 277881
rect 382294 276823 382346 276829
rect 382294 276765 382346 276771
rect 381814 275491 381866 275497
rect 381814 275433 381866 275439
rect 381430 272457 381482 272463
rect 381430 272399 381482 272405
rect 381526 272457 381578 272463
rect 381526 272399 381578 272405
rect 381538 263824 381566 272399
rect 380352 263796 380606 263824
rect 380832 263796 381086 263824
rect 381264 263796 381566 263824
rect 381826 263810 381854 275433
rect 382306 263810 382334 276765
rect 382402 270803 382430 277875
rect 382594 275275 382622 278018
rect 383554 278004 383856 278032
rect 585622 278081 585674 278087
rect 386518 278023 386570 278029
rect 383444 275974 383500 275983
rect 383444 275909 383500 275918
rect 382582 275269 382634 275275
rect 382582 275211 382634 275217
rect 382964 273162 383020 273171
rect 382964 273097 383020 273106
rect 382388 270794 382444 270803
rect 382388 270729 382444 270738
rect 382978 263824 383006 273097
rect 383458 263824 383486 275909
rect 383554 266839 383582 278004
rect 383638 276749 383690 276755
rect 383638 276691 383690 276697
rect 383542 266833 383594 266839
rect 383542 266775 383594 266781
rect 382752 263796 383006 263824
rect 383232 263796 383486 263824
rect 383650 263810 383678 276691
rect 384118 269497 384170 269503
rect 384118 269439 384170 269445
rect 384130 263810 384158 269439
rect 384994 269429 385022 278018
rect 385366 276675 385418 276681
rect 385366 276617 385418 276623
rect 385078 269645 385130 269651
rect 385078 269587 385130 269593
rect 385090 269429 385118 269587
rect 384982 269423 385034 269429
rect 384982 269365 385034 269371
rect 385078 269423 385130 269429
rect 385078 269365 385130 269371
rect 384886 267129 384938 267135
rect 384886 267071 384938 267077
rect 384898 263824 384926 267071
rect 385378 263824 385406 276617
rect 385556 270202 385612 270211
rect 385556 270137 385612 270146
rect 384672 263796 384926 263824
rect 385152 263796 385406 263824
rect 385570 263810 385598 270137
rect 386038 267055 386090 267061
rect 386038 266997 386090 267003
rect 386050 263810 386078 266997
rect 386146 266765 386174 278018
rect 386134 266759 386186 266765
rect 386134 266701 386186 266707
rect 386530 263810 386558 278023
rect 387394 274017 387422 278018
rect 387958 276527 388010 276533
rect 387958 276469 388010 276475
rect 387382 274011 387434 274017
rect 387382 273953 387434 273959
rect 387286 271199 387338 271205
rect 387286 271141 387338 271147
rect 387298 263824 387326 271141
rect 387382 269645 387434 269651
rect 387382 269587 387434 269593
rect 387394 269355 387422 269587
rect 387382 269349 387434 269355
rect 387382 269291 387434 269297
rect 387766 266981 387818 266987
rect 387766 266923 387818 266929
rect 387778 263824 387806 266923
rect 387072 263796 387326 263824
rect 387552 263796 387806 263824
rect 387970 263810 387998 276469
rect 388546 272389 388574 278018
rect 388918 275417 388970 275423
rect 388918 275359 388970 275365
rect 388534 272383 388586 272389
rect 388534 272325 388586 272331
rect 388724 270794 388780 270803
rect 388724 270729 388780 270738
rect 388436 270054 388492 270063
rect 388436 269989 388492 269998
rect 388450 263810 388478 269989
rect 388738 267801 388766 270729
rect 388726 267795 388778 267801
rect 388726 267737 388778 267743
rect 388930 263810 388958 275359
rect 389590 275343 389642 275349
rect 389590 275285 389642 275291
rect 389602 263824 389630 275285
rect 389698 275201 389726 278018
rect 390356 275826 390412 275835
rect 390356 275761 390412 275770
rect 389686 275195 389738 275201
rect 389686 275137 389738 275143
rect 390164 273014 390220 273023
rect 390164 272949 390220 272958
rect 390178 263824 390206 272949
rect 389472 263796 389630 263824
rect 389952 263796 390206 263824
rect 390370 263810 390398 275761
rect 390946 266691 390974 278018
rect 391990 275269 392042 275275
rect 391990 275211 392042 275217
rect 391508 269906 391564 269915
rect 391508 269841 391564 269850
rect 390934 266685 390986 266691
rect 390934 266627 390986 266633
rect 390838 264021 390890 264027
rect 390838 263963 390890 263969
rect 390850 263810 390878 263963
rect 391522 263824 391550 269841
rect 392002 263824 392030 275211
rect 392098 269429 392126 278018
rect 392962 278004 393264 278032
rect 392756 272866 392812 272875
rect 392756 272801 392812 272810
rect 392086 269423 392138 269429
rect 392086 269365 392138 269371
rect 392278 263947 392330 263953
rect 392278 263889 392330 263895
rect 391296 263796 391550 263824
rect 391776 263796 392030 263824
rect 392290 263810 392318 263889
rect 392770 263810 392798 272801
rect 392962 266617 392990 278004
rect 393908 276714 393964 276723
rect 393908 276649 393964 276658
rect 393238 266907 393290 266913
rect 393238 266849 393290 266855
rect 392950 266611 393002 266617
rect 392950 266553 393002 266559
rect 393250 263810 393278 266849
rect 393922 263824 393950 276649
rect 394498 273795 394526 278018
rect 394486 273789 394538 273795
rect 394486 273731 394538 273737
rect 395650 272315 395678 278018
rect 396692 276566 396748 276575
rect 396692 276501 396748 276510
rect 396310 275195 396362 275201
rect 396310 275137 396362 275143
rect 395638 272309 395690 272315
rect 395638 272251 395690 272257
rect 395926 272309 395978 272315
rect 395926 272251 395978 272257
rect 394390 269423 394442 269429
rect 394390 269365 394442 269371
rect 394402 263824 394430 269365
rect 394678 266833 394730 266839
rect 394678 266775 394730 266781
rect 393696 263796 393950 263824
rect 394176 263796 394430 263824
rect 394690 263810 394718 266775
rect 395446 263873 395498 263879
rect 395184 263821 395446 263824
rect 395938 263824 395966 272251
rect 396322 263824 396350 275137
rect 396706 263824 396734 276501
rect 396802 275127 396830 278018
rect 396790 275121 396842 275127
rect 396790 275063 396842 275069
rect 397076 269018 397132 269027
rect 397076 268953 397132 268962
rect 395184 263815 395498 263821
rect 395184 263796 395486 263815
rect 395664 263796 395966 263824
rect 396096 263796 396350 263824
rect 396576 263796 396734 263824
rect 397090 263810 397118 268953
rect 397558 266759 397610 266765
rect 397558 266701 397610 266707
rect 397570 263810 397598 266701
rect 398050 266543 398078 278018
rect 398900 275678 398956 275687
rect 398900 275613 398956 275622
rect 398708 272718 398764 272727
rect 398708 272653 398764 272662
rect 398230 266685 398282 266691
rect 398230 266627 398282 266633
rect 398038 266537 398090 266543
rect 398038 266479 398090 266485
rect 398242 263824 398270 266627
rect 398722 263824 398750 272653
rect 398016 263796 398270 263824
rect 398496 263796 398750 263824
rect 398914 263810 398942 275613
rect 399202 269651 399230 278018
rect 400354 275053 400382 278018
rect 400342 275047 400394 275053
rect 400342 274989 400394 274995
rect 401506 274091 401534 278018
rect 402548 276862 402604 276871
rect 402548 276797 402604 276806
rect 401782 275121 401834 275127
rect 401782 275063 401834 275069
rect 401494 274085 401546 274091
rect 401494 274027 401546 274033
rect 399190 269645 399242 269651
rect 399190 269587 399242 269593
rect 399958 269349 400010 269355
rect 399958 269291 400010 269297
rect 399382 264095 399434 264101
rect 399382 264037 399434 264043
rect 399394 263810 399422 264037
rect 399970 263810 399998 269291
rect 401302 267869 401354 267875
rect 401302 267811 401354 267817
rect 400630 266611 400682 266617
rect 400630 266553 400682 266559
rect 400642 263824 400670 266553
rect 400416 263796 400670 263824
rect 400896 263805 401150 263824
rect 401314 263810 401342 267811
rect 401794 263810 401822 275063
rect 402562 263824 402590 276797
rect 402754 272241 402782 278018
rect 402742 272235 402794 272241
rect 402742 272177 402794 272183
rect 402934 272235 402986 272241
rect 402934 272177 402986 272183
rect 402946 267875 402974 272177
rect 403028 269758 403084 269767
rect 403028 269693 403084 269702
rect 402934 267869 402986 267875
rect 402934 267811 402986 267817
rect 403042 263824 403070 269693
rect 403222 266537 403274 266543
rect 403222 266479 403274 266485
rect 400896 263799 401162 263805
rect 400896 263796 401110 263799
rect 402336 263796 402590 263824
rect 402816 263796 403070 263824
rect 403234 263810 403262 266479
rect 403906 266469 403934 278018
rect 404950 275047 405002 275053
rect 404950 274989 405002 274995
rect 404180 272570 404236 272579
rect 404180 272505 404236 272514
rect 403894 266463 403946 266469
rect 403894 266405 403946 266411
rect 404194 263810 404222 272505
rect 404962 263824 404990 274989
rect 405058 266395 405086 278018
rect 405620 269610 405676 269619
rect 405620 269545 405676 269554
rect 405046 266389 405098 266395
rect 405046 266331 405098 266337
rect 404736 263796 404990 263824
rect 405634 263810 405662 269545
rect 406306 269281 406334 278018
rect 407458 274165 407486 278018
rect 408886 277933 408938 277939
rect 408886 277875 408938 277881
rect 407828 275530 407884 275539
rect 407828 275465 407884 275474
rect 407446 274159 407498 274165
rect 407446 274101 407498 274107
rect 406582 273641 406634 273647
rect 406582 273583 406634 273589
rect 406294 269275 406346 269281
rect 406294 269217 406346 269223
rect 406102 266463 406154 266469
rect 406102 266405 406154 266411
rect 406114 263810 406142 266405
rect 406594 263810 406622 273583
rect 407252 272422 407308 272431
rect 407252 272357 407308 272366
rect 407446 272383 407498 272389
rect 407266 263824 407294 272357
rect 407446 272325 407498 272331
rect 407458 271205 407486 272325
rect 407446 271199 407498 271205
rect 407446 271141 407498 271147
rect 407842 263824 407870 275465
rect 408898 273319 408926 277875
rect 408884 273310 408940 273319
rect 408884 273245 408940 273254
rect 409858 272167 409886 278018
rect 411010 274313 411038 278018
rect 412162 276903 412190 278018
rect 412150 276897 412202 276903
rect 412150 276839 412202 276845
rect 410998 274307 411050 274313
rect 410998 274249 411050 274255
rect 410900 272274 410956 272283
rect 410900 272209 410956 272218
rect 409846 272161 409898 272167
rect 409846 272103 409898 272109
rect 408982 270755 409034 270761
rect 408982 270697 409034 270703
rect 408994 268393 409022 270697
rect 410420 269462 410476 269471
rect 410420 269397 410476 269406
rect 408982 268387 409034 268393
rect 408982 268329 409034 268335
rect 408502 268239 408554 268245
rect 408502 268181 408554 268187
rect 408022 265797 408074 265803
rect 408022 265739 408074 265745
rect 407040 263796 407294 263824
rect 407616 263796 407870 263824
rect 408034 263810 408062 265739
rect 408514 263810 408542 268181
rect 409942 267869 409994 267875
rect 409942 267811 409994 267817
rect 409174 266389 409226 266395
rect 409174 266331 409226 266337
rect 409186 263824 409214 266331
rect 408960 263796 409214 263824
rect 409954 263810 409982 267811
rect 410434 263810 410462 269397
rect 410914 263810 410942 272209
rect 411764 272126 411820 272135
rect 411764 272061 411820 272070
rect 411572 269314 411628 269323
rect 411572 269249 411628 269258
rect 411586 263824 411614 269249
rect 411670 264095 411722 264101
rect 411670 264037 411722 264043
rect 411360 263796 411614 263824
rect 411682 263805 411710 264037
rect 411778 263824 411806 272061
rect 413410 270761 413438 278018
rect 414562 274239 414590 278018
rect 415714 277791 415742 278018
rect 415702 277785 415754 277791
rect 415702 277727 415754 277733
rect 414550 274233 414602 274239
rect 414550 274175 414602 274181
rect 413686 272161 413738 272167
rect 413686 272103 413738 272109
rect 413398 270755 413450 270761
rect 413398 270697 413450 270703
rect 413698 267875 413726 272103
rect 416962 271279 416990 278018
rect 416950 271273 417002 271279
rect 416950 271215 417002 271221
rect 413686 267869 413738 267875
rect 413686 267811 413738 267817
rect 418114 265507 418142 278018
rect 420514 268467 420542 278018
rect 421666 274387 421694 278018
rect 421654 274381 421706 274387
rect 421654 274323 421706 274329
rect 423970 271353 423998 278018
rect 423958 271347 424010 271353
rect 423958 271289 424010 271295
rect 420502 268461 420554 268467
rect 420502 268403 420554 268409
rect 425218 265581 425246 278018
rect 426370 276607 426398 278018
rect 426358 276601 426410 276607
rect 426358 276543 426410 276549
rect 427522 268541 427550 278018
rect 428770 274461 428798 278018
rect 429634 278013 429936 278032
rect 585674 278029 585936 278032
rect 585622 278023 585936 278029
rect 429622 278007 429936 278013
rect 429674 278004 429936 278007
rect 429622 277949 429674 277955
rect 428758 274455 428810 274461
rect 428758 274397 428810 274403
rect 431074 271427 431102 278018
rect 431062 271421 431114 271427
rect 431062 271363 431114 271369
rect 427510 268535 427562 268541
rect 427510 268477 427562 268483
rect 432322 265655 432350 278018
rect 432310 265649 432362 265655
rect 432310 265591 432362 265597
rect 425206 265575 425258 265581
rect 425206 265517 425258 265523
rect 418102 265501 418154 265507
rect 418102 265443 418154 265449
rect 433474 264767 433502 278018
rect 434626 268615 434654 278018
rect 435874 274535 435902 278018
rect 437026 277865 437054 278018
rect 437014 277859 437066 277865
rect 437014 277801 437066 277807
rect 435862 274529 435914 274535
rect 435862 274471 435914 274477
rect 438178 271501 438206 278018
rect 438166 271495 438218 271501
rect 438166 271437 438218 271443
rect 434614 268609 434666 268615
rect 434614 268551 434666 268557
rect 439330 265729 439358 278018
rect 439318 265723 439370 265729
rect 439318 265665 439370 265671
rect 433462 264761 433514 264767
rect 433462 264703 433514 264709
rect 440578 264545 440606 278018
rect 441730 268689 441758 278018
rect 442882 274609 442910 278018
rect 444130 277717 444158 278018
rect 444118 277711 444170 277717
rect 444118 277653 444170 277659
rect 442870 274603 442922 274609
rect 442870 274545 442922 274551
rect 445282 271575 445310 278018
rect 446434 274683 446462 278018
rect 446422 274677 446474 274683
rect 446422 274619 446474 274625
rect 445270 271569 445322 271575
rect 445270 271511 445322 271517
rect 441718 268683 441770 268689
rect 441718 268625 441770 268631
rect 440566 264539 440618 264545
rect 440566 264481 440618 264487
rect 447682 264471 447710 278018
rect 448834 268763 448862 278018
rect 448822 268757 448874 268763
rect 448822 268699 448874 268705
rect 449986 265877 450014 278018
rect 451234 277643 451262 278018
rect 451222 277637 451274 277643
rect 451222 277579 451274 277585
rect 452386 271649 452414 278018
rect 453538 274757 453566 278018
rect 453526 274751 453578 274757
rect 453526 274693 453578 274699
rect 452374 271643 452426 271649
rect 452374 271585 452426 271591
rect 449974 265871 450026 265877
rect 449974 265813 450026 265819
rect 447670 264465 447722 264471
rect 447670 264407 447722 264413
rect 454786 264397 454814 278018
rect 455938 268837 455966 278018
rect 455926 268831 455978 268837
rect 455926 268773 455978 268779
rect 457090 265951 457118 278018
rect 458242 277569 458270 278018
rect 458230 277563 458282 277569
rect 458230 277505 458282 277511
rect 459490 271723 459518 278018
rect 460642 274831 460670 278018
rect 460630 274825 460682 274831
rect 460630 274767 460682 274773
rect 459478 271717 459530 271723
rect 459478 271659 459530 271665
rect 457078 265945 457130 265951
rect 457078 265887 457130 265893
rect 461794 264619 461822 278018
rect 463042 268911 463070 278018
rect 463030 268905 463082 268911
rect 463030 268847 463082 268853
rect 464194 266025 464222 278018
rect 465346 277495 465374 278018
rect 465334 277489 465386 277495
rect 465334 277431 465386 277437
rect 466594 271797 466622 278018
rect 467746 274905 467774 278018
rect 467734 274899 467786 274905
rect 467734 274841 467786 274847
rect 466582 271791 466634 271797
rect 466582 271733 466634 271739
rect 464182 266019 464234 266025
rect 464182 265961 464234 265967
rect 468898 264693 468926 278018
rect 470146 268985 470174 278018
rect 470134 268979 470186 268985
rect 470134 268921 470186 268927
rect 471298 266099 471326 278018
rect 472450 277421 472478 278018
rect 472438 277415 472490 277421
rect 472438 277357 472490 277363
rect 473698 271871 473726 278018
rect 474850 274503 474878 278018
rect 474836 274494 474892 274503
rect 474836 274429 474892 274438
rect 473686 271865 473738 271871
rect 473686 271807 473738 271813
rect 471286 266093 471338 266099
rect 471286 266035 471338 266041
rect 476002 264841 476030 278018
rect 477154 269059 477182 278018
rect 477142 269053 477194 269059
rect 477142 268995 477194 269001
rect 478402 266173 478430 278018
rect 479554 277347 479582 278018
rect 479542 277341 479594 277347
rect 479542 277283 479594 277289
rect 480706 271945 480734 278018
rect 481954 274979 481982 278018
rect 481942 274973 481994 274979
rect 481942 274915 481994 274921
rect 480694 271939 480746 271945
rect 480694 271881 480746 271887
rect 483106 269133 483134 278018
rect 484258 269207 484286 278018
rect 484246 269201 484298 269207
rect 484246 269143 484298 269149
rect 483094 269127 483146 269133
rect 483094 269069 483146 269075
rect 485506 266247 485534 278018
rect 486658 272019 486686 278018
rect 487810 272093 487838 278018
rect 489058 274651 489086 278018
rect 489044 274642 489100 274651
rect 489044 274577 489100 274586
rect 487798 272087 487850 272093
rect 487798 272029 487850 272035
rect 486646 272013 486698 272019
rect 486646 271955 486698 271961
rect 490210 270687 490238 278018
rect 490198 270681 490250 270687
rect 490198 270623 490250 270629
rect 491362 270613 491390 278018
rect 491350 270607 491402 270613
rect 491350 270549 491402 270555
rect 492610 266321 492638 278018
rect 493762 273573 493790 278018
rect 493750 273567 493802 273573
rect 493750 273509 493802 273515
rect 494914 273499 494942 278018
rect 496066 274799 496094 278018
rect 496052 274790 496108 274799
rect 496052 274725 496108 274734
rect 494902 273493 494954 273499
rect 494902 273435 494954 273441
rect 497314 270539 497342 278018
rect 497302 270533 497354 270539
rect 497302 270475 497354 270481
rect 498466 270465 498494 278018
rect 498454 270459 498506 270465
rect 498454 270401 498506 270407
rect 499618 267727 499646 278018
rect 500866 273425 500894 278018
rect 500854 273419 500906 273425
rect 500854 273361 500906 273367
rect 502018 273351 502046 278018
rect 503170 274947 503198 278018
rect 503156 274938 503212 274947
rect 503156 274873 503212 274882
rect 502006 273345 502058 273351
rect 502006 273287 502058 273293
rect 504418 270317 504446 278018
rect 505570 270391 505598 278018
rect 505558 270385 505610 270391
rect 505558 270327 505610 270333
rect 504406 270311 504458 270317
rect 504406 270253 504458 270259
rect 499606 267721 499658 267727
rect 499606 267663 499658 267669
rect 506722 267653 506750 278018
rect 507970 273203 507998 278018
rect 509122 273277 509150 278018
rect 510274 276459 510302 278018
rect 510262 276453 510314 276459
rect 510262 276395 510314 276401
rect 509110 273271 509162 273277
rect 509110 273213 509162 273219
rect 507958 273197 508010 273203
rect 507958 273139 508010 273145
rect 508246 273197 508298 273203
rect 508246 273139 508298 273145
rect 508258 268879 508286 273139
rect 511522 270243 511550 278018
rect 511510 270237 511562 270243
rect 511510 270179 511562 270185
rect 512674 270169 512702 278018
rect 512662 270163 512714 270169
rect 512662 270105 512714 270111
rect 508244 268870 508300 268879
rect 508244 268805 508300 268814
rect 506710 267647 506762 267653
rect 506710 267589 506762 267595
rect 513826 267579 513854 278018
rect 514978 273129 515006 278018
rect 514966 273123 515018 273129
rect 514966 273065 515018 273071
rect 516226 273055 516254 278018
rect 517378 276385 517406 278018
rect 517366 276379 517418 276385
rect 517366 276321 517418 276327
rect 516214 273049 516266 273055
rect 516214 272991 516266 272997
rect 518530 270021 518558 278018
rect 519778 270095 519806 278018
rect 519766 270089 519818 270095
rect 519766 270031 519818 270037
rect 518518 270015 518570 270021
rect 518518 269957 518570 269963
rect 513814 267573 513866 267579
rect 513814 267515 513866 267521
rect 520930 267505 520958 278018
rect 522082 272981 522110 278018
rect 522070 272975 522122 272981
rect 522070 272917 522122 272923
rect 523330 272907 523358 278018
rect 524482 276311 524510 278018
rect 524470 276305 524522 276311
rect 524470 276247 524522 276253
rect 523318 272901 523370 272907
rect 523318 272843 523370 272849
rect 523990 272901 524042 272907
rect 523990 272843 524042 272849
rect 520918 267499 520970 267505
rect 520918 267441 520970 267447
rect 492598 266315 492650 266321
rect 492598 266257 492650 266263
rect 485494 266241 485546 266247
rect 485494 266183 485546 266189
rect 478390 266167 478442 266173
rect 478390 266109 478442 266115
rect 524002 265803 524030 272843
rect 525634 269873 525662 278018
rect 526882 269947 526910 278018
rect 526964 276862 527020 276871
rect 526964 276797 527020 276806
rect 526978 273499 527006 276797
rect 526966 273493 527018 273499
rect 526966 273435 527018 273441
rect 526870 269941 526922 269947
rect 526870 269883 526922 269889
rect 525622 269867 525674 269873
rect 525622 269809 525674 269815
rect 528034 267431 528062 278018
rect 529186 272833 529214 278018
rect 529174 272827 529226 272833
rect 529174 272769 529226 272775
rect 530434 272759 530462 278018
rect 531586 276237 531614 278018
rect 531574 276231 531626 276237
rect 531574 276173 531626 276179
rect 530422 272753 530474 272759
rect 530422 272695 530474 272701
rect 532738 269799 532766 278018
rect 532822 272753 532874 272759
rect 532822 272695 532874 272701
rect 532726 269793 532778 269799
rect 532726 269735 532778 269741
rect 532834 269027 532862 272695
rect 533890 269725 533918 278018
rect 533878 269719 533930 269725
rect 533878 269661 533930 269667
rect 532820 269018 532876 269027
rect 532820 268953 532876 268962
rect 528022 267425 528074 267431
rect 528022 267367 528074 267373
rect 535138 267357 535166 278018
rect 536290 272611 536318 278018
rect 537442 272685 537470 278018
rect 538690 276163 538718 278018
rect 538678 276157 538730 276163
rect 538678 276099 538730 276105
rect 537430 272679 537482 272685
rect 537430 272621 537482 272627
rect 536278 272605 536330 272611
rect 536278 272547 536330 272553
rect 539842 270507 539870 278018
rect 539828 270498 539884 270507
rect 539828 270433 539884 270442
rect 540994 269175 541022 278018
rect 540980 269166 541036 269175
rect 540980 269101 541036 269110
rect 535126 267351 535178 267357
rect 535126 267293 535178 267299
rect 542242 267283 542270 278018
rect 543394 271543 543422 278018
rect 544546 271691 544574 278018
rect 545794 275941 545822 278018
rect 546946 276015 546974 278018
rect 546934 276009 546986 276015
rect 546934 275951 546986 275957
rect 545782 275935 545834 275941
rect 545782 275877 545834 275883
rect 544532 271682 544588 271691
rect 544532 271617 544588 271626
rect 543380 271534 543436 271543
rect 543380 271469 543436 271478
rect 548098 268171 548126 278018
rect 549346 276089 549374 278018
rect 549334 276083 549386 276089
rect 549334 276025 549386 276031
rect 548086 268165 548138 268171
rect 548086 268107 548138 268113
rect 542230 267277 542282 267283
rect 542230 267219 542282 267225
rect 550498 267209 550526 278018
rect 551650 272537 551678 278018
rect 552802 275867 552830 278018
rect 554050 277273 554078 278018
rect 554038 277267 554090 277273
rect 554038 277209 554090 277215
rect 552790 275861 552842 275867
rect 552790 275803 552842 275809
rect 555202 273203 555230 278018
rect 556354 275793 556382 278018
rect 557602 277199 557630 278018
rect 557590 277193 557642 277199
rect 557590 277135 557642 277141
rect 556342 275787 556394 275793
rect 556342 275729 556394 275735
rect 555190 273197 555242 273203
rect 555190 273139 555242 273145
rect 551638 272531 551690 272537
rect 551638 272473 551690 272479
rect 558754 271839 558782 278018
rect 559906 275645 559934 278018
rect 561154 277125 561182 278018
rect 561142 277119 561194 277125
rect 561142 277061 561194 277067
rect 559894 275639 559946 275645
rect 559894 275581 559946 275587
rect 558740 271830 558796 271839
rect 558740 271765 558796 271774
rect 562306 270359 562334 278018
rect 563458 275719 563486 278018
rect 564706 277051 564734 278018
rect 564694 277045 564746 277051
rect 564694 276987 564746 276993
rect 563446 275713 563498 275719
rect 563446 275655 563498 275661
rect 565858 271987 565886 278018
rect 567010 276131 567038 278018
rect 568258 276977 568286 278018
rect 568246 276971 568298 276977
rect 568246 276913 568298 276919
rect 566996 276122 567052 276131
rect 566996 276057 567052 276066
rect 565844 271978 565900 271987
rect 565844 271913 565900 271922
rect 562292 270350 562348 270359
rect 562292 270285 562348 270294
rect 569410 269577 569438 278018
rect 570562 275571 570590 278018
rect 570550 275565 570602 275571
rect 570550 275507 570602 275513
rect 572962 272463 572990 278018
rect 574114 275497 574142 278018
rect 575266 276829 575294 278018
rect 575254 276823 575306 276829
rect 575254 276765 575306 276771
rect 574102 275491 574154 275497
rect 574102 275433 574154 275439
rect 576514 273171 576542 278018
rect 577666 275983 577694 278018
rect 578818 276755 578846 278018
rect 578806 276749 578858 276755
rect 578806 276691 578858 276697
rect 577652 275974 577708 275983
rect 577652 275909 577708 275918
rect 576500 273162 576556 273171
rect 576500 273097 576556 273106
rect 572950 272457 573002 272463
rect 572950 272399 573002 272405
rect 569398 269571 569450 269577
rect 569398 269513 569450 269519
rect 580066 269503 580094 278018
rect 580054 269497 580106 269503
rect 580054 269439 580106 269445
rect 550486 267203 550538 267209
rect 550486 267145 550538 267151
rect 581218 267135 581246 278018
rect 582370 276681 582398 278018
rect 582358 276675 582410 276681
rect 582358 276617 582410 276623
rect 583618 270211 583646 278018
rect 583604 270202 583660 270211
rect 583604 270137 583660 270146
rect 581206 267129 581258 267135
rect 581206 267071 581258 267077
rect 584770 267061 584798 278018
rect 585634 278004 585936 278023
rect 587170 272389 587198 278018
rect 587158 272383 587210 272389
rect 587158 272325 587210 272331
rect 584758 267055 584810 267061
rect 584758 266997 584810 267003
rect 588322 266987 588350 278018
rect 589474 276533 589502 278018
rect 589462 276527 589514 276533
rect 589462 276469 589514 276475
rect 590626 270063 590654 278018
rect 591874 275423 591902 278018
rect 591862 275417 591914 275423
rect 591862 275359 591914 275365
rect 593026 275349 593054 278018
rect 593014 275343 593066 275349
rect 593014 275285 593066 275291
rect 594178 273023 594206 278018
rect 595426 275835 595454 278018
rect 595412 275826 595468 275835
rect 595412 275761 595468 275770
rect 594164 273014 594220 273023
rect 594164 272949 594220 272958
rect 590612 270054 590668 270063
rect 590612 269989 590668 269998
rect 588310 266981 588362 266987
rect 588310 266923 588362 266929
rect 523990 265797 524042 265803
rect 523990 265739 524042 265745
rect 475990 264835 476042 264841
rect 475990 264777 476042 264783
rect 468886 264687 468938 264693
rect 468886 264629 468938 264635
rect 461782 264613 461834 264619
rect 461782 264555 461834 264561
rect 454774 264391 454826 264397
rect 454774 264333 454826 264339
rect 596578 264027 596606 278018
rect 597730 269915 597758 278018
rect 598978 275275 599006 278018
rect 598966 275269 599018 275275
rect 598966 275211 599018 275217
rect 597716 269906 597772 269915
rect 597716 269841 597772 269850
rect 596566 264021 596618 264027
rect 596566 263963 596618 263969
rect 600130 263953 600158 278018
rect 601282 272875 601310 278018
rect 601268 272866 601324 272875
rect 601268 272801 601324 272810
rect 602530 266913 602558 278018
rect 603682 276723 603710 278018
rect 603668 276714 603724 276723
rect 603668 276649 603724 276658
rect 604834 269429 604862 278018
rect 604822 269423 604874 269429
rect 604822 269365 604874 269371
rect 602518 266907 602570 266913
rect 602518 266849 602570 266855
rect 606082 266839 606110 278018
rect 606070 266833 606122 266839
rect 606070 266775 606122 266781
rect 600118 263947 600170 263953
rect 600118 263889 600170 263895
rect 607234 263879 607262 278018
rect 608386 272315 608414 278018
rect 609538 275201 609566 278018
rect 610786 276575 610814 278018
rect 610772 276566 610828 276575
rect 610772 276501 610828 276510
rect 609526 275195 609578 275201
rect 609526 275137 609578 275143
rect 611938 272759 611966 278018
rect 611926 272753 611978 272759
rect 611926 272695 611978 272701
rect 608374 272309 608426 272315
rect 608374 272251 608426 272257
rect 613090 266765 613118 278018
rect 613078 266759 613130 266765
rect 613078 266701 613130 266707
rect 614338 266691 614366 278018
rect 615490 272727 615518 278018
rect 616642 275687 616670 278018
rect 616628 275678 616684 275687
rect 616628 275613 616684 275622
rect 615476 272718 615532 272727
rect 615476 272653 615532 272662
rect 614326 266685 614378 266691
rect 614326 266627 614378 266633
rect 607222 263873 607274 263879
rect 411670 263799 411722 263805
rect 401110 263741 401162 263747
rect 411778 263796 411840 263824
rect 607222 263815 607274 263821
rect 617890 263805 617918 278018
rect 619042 269355 619070 278018
rect 619030 269349 619082 269355
rect 619030 269291 619082 269297
rect 620194 266617 620222 278018
rect 620182 266611 620234 266617
rect 620182 266553 620234 266559
rect 617878 263799 617930 263805
rect 411670 263741 411722 263747
rect 617878 263741 617930 263747
rect 621442 263731 621470 278018
rect 622594 272241 622622 278018
rect 623746 275127 623774 278018
rect 623734 275121 623786 275127
rect 623734 275063 623786 275069
rect 624994 273499 625022 278018
rect 624982 273493 625034 273499
rect 624982 273435 625034 273441
rect 622582 272235 622634 272241
rect 622582 272177 622634 272183
rect 626146 269767 626174 278018
rect 626132 269758 626188 269767
rect 626132 269693 626188 269702
rect 627298 266543 627326 278018
rect 627286 266537 627338 266543
rect 627286 266479 627338 266485
rect 403990 263725 404042 263731
rect 299170 263648 299232 263676
rect 345442 263648 345504 263676
rect 403728 263673 403990 263676
rect 621430 263725 621482 263731
rect 403728 263667 404042 263673
rect 403728 263648 404030 263667
rect 405216 263657 405470 263676
rect 621430 263667 621482 263673
rect 628450 263657 628478 278018
rect 629698 272579 629726 278018
rect 630850 275053 630878 278018
rect 630838 275047 630890 275053
rect 630838 274989 630890 274995
rect 629684 272570 629740 272579
rect 629684 272505 629740 272514
rect 405216 263651 405482 263657
rect 405216 263648 405430 263651
rect 405430 263593 405482 263599
rect 628438 263651 628490 263657
rect 628438 263593 628490 263599
rect 632002 263583 632030 278018
rect 633250 269619 633278 278018
rect 633236 269610 633292 269619
rect 633236 269545 633292 269554
rect 634402 266469 634430 278018
rect 635554 273573 635582 278018
rect 635542 273567 635594 273573
rect 635542 273509 635594 273515
rect 636802 272431 636830 278018
rect 637954 275539 637982 278018
rect 637940 275530 637996 275539
rect 637940 275465 637996 275474
rect 639106 272907 639134 278018
rect 639094 272901 639146 272907
rect 639094 272843 639146 272849
rect 636788 272422 636844 272431
rect 636788 272357 636844 272366
rect 640354 268245 640382 278018
rect 640342 268239 640394 268245
rect 640342 268181 640394 268187
rect 634390 266463 634442 266469
rect 634390 266405 634442 266411
rect 641506 266395 641534 278018
rect 641494 266389 641546 266395
rect 641494 266331 641546 266337
rect 409654 263577 409706 263583
rect 409440 263525 409654 263528
rect 409440 263519 409706 263525
rect 631990 263577 632042 263583
rect 631990 263519 632042 263525
rect 409440 263500 409694 263519
rect 642658 263509 642686 278018
rect 643906 272167 643934 278018
rect 643894 272161 643946 272167
rect 643894 272103 643946 272109
rect 645058 269471 645086 278018
rect 646210 272283 646238 278018
rect 646484 275382 646540 275391
rect 646484 275317 646540 275326
rect 646196 272274 646252 272283
rect 646196 272209 646252 272218
rect 645238 270903 645290 270909
rect 645238 270845 645290 270851
rect 645044 269462 645100 269471
rect 645044 269397 645100 269406
rect 645250 267801 645278 270845
rect 645238 267795 645290 267801
rect 645238 267737 645290 267743
rect 642646 263503 642698 263509
rect 642646 263445 642698 263451
rect 420404 262210 420460 262219
rect 420404 262145 420406 262154
rect 420458 262145 420460 262154
rect 606166 262171 606218 262177
rect 420406 262113 420458 262119
rect 606166 262113 606218 262119
rect 420404 259842 420460 259851
rect 420404 259777 420460 259786
rect 191540 259398 191596 259407
rect 191540 259333 191596 259342
rect 187222 257805 187274 257811
rect 187222 257747 187274 257753
rect 189718 257805 189770 257811
rect 189718 257747 189770 257753
rect 186070 254993 186122 254999
rect 186070 254935 186122 254941
rect 185782 246705 185834 246711
rect 185782 246647 185834 246653
rect 185686 242857 185738 242863
rect 185686 242799 185738 242805
rect 185492 198274 185548 198283
rect 185492 198209 185548 198218
rect 184436 196794 184492 196803
rect 184436 196729 184492 196738
rect 184340 196054 184396 196063
rect 184340 195989 184396 195998
rect 184534 195793 184586 195799
rect 184534 195735 184586 195741
rect 184438 195719 184490 195725
rect 184438 195661 184490 195667
rect 184342 195645 184394 195651
rect 184342 195587 184394 195593
rect 184354 195323 184382 195587
rect 184340 195314 184396 195323
rect 184340 195249 184396 195258
rect 184450 194435 184478 195661
rect 184436 194426 184492 194435
rect 184436 194361 184492 194370
rect 184546 193843 184574 195735
rect 184532 193834 184588 193843
rect 184532 193769 184588 193778
rect 184630 192981 184682 192987
rect 184436 192946 184492 192955
rect 184630 192923 184682 192929
rect 184436 192881 184492 192890
rect 184534 192907 184586 192913
rect 184342 192833 184394 192839
rect 184342 192775 184394 192781
rect 184354 192363 184382 192775
rect 184450 192765 184478 192881
rect 184534 192849 184586 192855
rect 184438 192759 184490 192765
rect 184438 192701 184490 192707
rect 184340 192354 184396 192363
rect 184340 192289 184396 192298
rect 184546 191475 184574 192849
rect 184532 191466 184588 191475
rect 184532 191401 184588 191410
rect 184642 190735 184670 192923
rect 184628 190726 184684 190735
rect 184628 190661 184684 190670
rect 184534 190095 184586 190101
rect 184534 190037 184586 190043
rect 184342 190021 184394 190027
rect 184340 189986 184342 189995
rect 184394 189986 184396 189995
rect 184340 189921 184396 189930
rect 184438 189947 184490 189953
rect 184438 189889 184490 189895
rect 184342 189873 184394 189879
rect 184342 189815 184394 189821
rect 184354 187627 184382 189815
rect 184450 188515 184478 189889
rect 184546 189255 184574 190037
rect 184532 189246 184588 189255
rect 184532 189181 184588 189190
rect 184436 188506 184492 188515
rect 184436 188441 184492 188450
rect 184340 187618 184396 187627
rect 184340 187553 184396 187562
rect 184438 187209 184490 187215
rect 184438 187151 184490 187157
rect 184342 187135 184394 187141
rect 184342 187077 184394 187083
rect 184354 186887 184382 187077
rect 184340 186878 184396 186887
rect 184340 186813 184396 186822
rect 184450 186147 184478 187151
rect 184534 187061 184586 187067
rect 184534 187003 184586 187009
rect 184436 186138 184492 186147
rect 184436 186073 184492 186082
rect 184546 184667 184574 187003
rect 184630 186987 184682 186993
rect 184630 186929 184682 186935
rect 184642 185407 184670 186929
rect 184628 185398 184684 185407
rect 184628 185333 184684 185342
rect 184532 184658 184588 184667
rect 184532 184593 184588 184602
rect 184342 184323 184394 184329
rect 184342 184265 184394 184271
rect 184354 183927 184382 184265
rect 184438 184249 184490 184255
rect 184438 184191 184490 184197
rect 184340 183918 184396 183927
rect 184340 183853 184396 183862
rect 184450 183187 184478 184191
rect 184534 184175 184586 184181
rect 184534 184117 184586 184123
rect 184436 183178 184492 183187
rect 184436 183113 184492 183122
rect 184546 181559 184574 184117
rect 184532 181550 184588 181559
rect 184532 181485 184588 181494
rect 184630 181437 184682 181443
rect 184630 181379 184682 181385
rect 184342 181363 184394 181369
rect 184342 181305 184394 181311
rect 184354 180819 184382 181305
rect 184438 181289 184490 181295
rect 184438 181231 184490 181237
rect 184340 180810 184396 180819
rect 184340 180745 184396 180754
rect 184450 180079 184478 181231
rect 184534 181215 184586 181221
rect 184534 181157 184586 181163
rect 184436 180070 184492 180079
rect 184436 180005 184492 180014
rect 183094 178625 183146 178631
rect 184546 178599 184574 181157
rect 184642 179339 184670 181379
rect 185494 180031 185546 180037
rect 185494 179973 185546 179979
rect 184628 179330 184684 179339
rect 184628 179265 184684 179274
rect 183094 178567 183146 178573
rect 184532 178590 184588 178599
rect 182998 146879 183050 146885
rect 182998 146821 183050 146827
rect 183106 132455 183134 178567
rect 184438 178551 184490 178557
rect 184532 178525 184588 178534
rect 184438 178493 184490 178499
rect 184342 178477 184394 178483
rect 184342 178419 184394 178425
rect 184354 177119 184382 178419
rect 184340 177110 184396 177119
rect 184340 177045 184396 177054
rect 184450 176231 184478 178493
rect 184436 176222 184492 176231
rect 184436 176157 184492 176166
rect 184438 175665 184490 175671
rect 184340 175630 184396 175639
rect 184438 175607 184490 175613
rect 184340 175565 184342 175574
rect 184394 175565 184396 175574
rect 184342 175533 184394 175539
rect 184450 174011 184478 175607
rect 184436 174002 184492 174011
rect 184436 173937 184492 173946
rect 184534 172779 184586 172785
rect 184534 172721 184586 172727
rect 184342 172631 184394 172637
rect 184342 172573 184394 172579
rect 184354 172531 184382 172573
rect 184438 172557 184490 172563
rect 184340 172522 184396 172531
rect 184438 172499 184490 172505
rect 184340 172457 184396 172466
rect 184450 170311 184478 172499
rect 184546 171791 184574 172721
rect 184630 172705 184682 172711
rect 184630 172647 184682 172653
rect 184532 171782 184588 171791
rect 184532 171717 184588 171726
rect 184642 170903 184670 172647
rect 184628 170894 184684 170903
rect 184628 170829 184684 170838
rect 184436 170302 184492 170311
rect 184436 170237 184492 170246
rect 184630 169893 184682 169899
rect 184630 169835 184682 169841
rect 184438 169819 184490 169825
rect 184438 169761 184490 169767
rect 184342 169745 184394 169751
rect 184342 169687 184394 169693
rect 184354 169423 184382 169687
rect 184340 169414 184396 169423
rect 184340 169349 184396 169358
rect 184450 168683 184478 169761
rect 184534 169671 184586 169677
rect 184534 169613 184586 169619
rect 184436 168674 184492 168683
rect 184436 168609 184492 168618
rect 184546 167203 184574 169613
rect 184642 167943 184670 169835
rect 184628 167934 184684 167943
rect 184628 167869 184684 167878
rect 184532 167194 184588 167203
rect 184532 167129 184588 167138
rect 184342 167007 184394 167013
rect 184342 166949 184394 166955
rect 184354 166463 184382 166949
rect 184438 166933 184490 166939
rect 184438 166875 184490 166881
rect 184340 166454 184396 166463
rect 184340 166389 184396 166398
rect 184450 165723 184478 166875
rect 184534 166859 184586 166865
rect 184534 166801 184586 166807
rect 184436 165714 184492 165723
rect 184436 165649 184492 165658
rect 184546 164835 184574 166801
rect 184532 164826 184588 164835
rect 184532 164761 184588 164770
rect 185302 164121 185354 164127
rect 184340 164086 184396 164095
rect 185302 164063 185354 164069
rect 184340 164021 184342 164030
rect 184394 164021 184396 164030
rect 184342 163989 184394 163995
rect 184438 163973 184490 163979
rect 184438 163915 184490 163921
rect 184342 163899 184394 163905
rect 184342 163841 184394 163847
rect 184354 163355 184382 163841
rect 184340 163346 184396 163355
rect 184340 163281 184396 163290
rect 184450 161875 184478 163915
rect 185314 162615 185342 164063
rect 185300 162606 185356 162615
rect 185300 162541 185356 162550
rect 184436 161866 184492 161875
rect 184436 161801 184492 161810
rect 184534 161235 184586 161241
rect 184534 161177 184586 161183
rect 184342 161087 184394 161093
rect 184342 161029 184394 161035
rect 184354 160987 184382 161029
rect 184438 161013 184490 161019
rect 184340 160978 184396 160987
rect 184438 160955 184490 160961
rect 184340 160913 184396 160922
rect 184450 160395 184478 160955
rect 184436 160386 184492 160395
rect 184436 160321 184492 160330
rect 184546 159507 184574 161177
rect 184630 161161 184682 161167
rect 184630 161103 184682 161109
rect 184532 159498 184588 159507
rect 184532 159433 184588 159442
rect 184642 158915 184670 161103
rect 184628 158906 184684 158915
rect 184628 158841 184684 158850
rect 184438 158423 184490 158429
rect 184438 158365 184490 158371
rect 184342 158349 184394 158355
rect 184342 158291 184394 158297
rect 184354 156547 184382 158291
rect 184340 156538 184396 156547
rect 184340 156473 184396 156482
rect 184450 155659 184478 158365
rect 184534 158275 184586 158281
rect 184534 158217 184586 158223
rect 184546 158027 184574 158217
rect 184630 158201 184682 158207
rect 184630 158143 184682 158149
rect 184532 158018 184588 158027
rect 184532 157953 184588 157962
rect 184642 157435 184670 158143
rect 184628 157426 184684 157435
rect 184628 157361 184684 157370
rect 184436 155650 184492 155659
rect 184436 155585 184492 155594
rect 184534 155537 184586 155543
rect 184534 155479 184586 155485
rect 184438 155463 184490 155469
rect 184438 155405 184490 155411
rect 184342 155315 184394 155321
rect 184342 155257 184394 155263
rect 184354 155067 184382 155257
rect 184340 155058 184396 155067
rect 184340 154993 184396 155002
rect 184450 154179 184478 155405
rect 184436 154170 184492 154179
rect 184436 154105 184492 154114
rect 184546 153587 184574 155479
rect 184630 155389 184682 155395
rect 184630 155331 184682 155337
rect 184532 153578 184588 153587
rect 184532 153513 184588 153522
rect 184642 152699 184670 155331
rect 184628 152690 184684 152699
rect 184534 152651 184586 152657
rect 184628 152625 184684 152634
rect 184534 152593 184586 152599
rect 184342 152577 184394 152583
rect 184342 152519 184394 152525
rect 184354 151959 184382 152519
rect 184438 152503 184490 152509
rect 184438 152445 184490 152451
rect 184340 151950 184396 151959
rect 184340 151885 184396 151894
rect 184450 150479 184478 152445
rect 184546 151219 184574 152593
rect 184532 151210 184588 151219
rect 184532 151145 184588 151154
rect 184436 150470 184492 150479
rect 184436 150405 184492 150414
rect 184342 149765 184394 149771
rect 184340 149730 184342 149739
rect 184394 149730 184396 149739
rect 184340 149665 184396 149674
rect 184438 149691 184490 149697
rect 184438 149633 184490 149639
rect 184342 149543 184394 149549
rect 184342 149485 184394 149491
rect 184354 148111 184382 149485
rect 184450 148999 184478 149633
rect 184534 149617 184586 149623
rect 184534 149559 184586 149565
rect 184436 148990 184492 148999
rect 184436 148925 184492 148934
rect 184340 148102 184396 148111
rect 184340 148037 184396 148046
rect 184546 147371 184574 149559
rect 184532 147362 184588 147371
rect 184532 147297 184588 147306
rect 184342 146805 184394 146811
rect 184342 146747 184394 146753
rect 184354 145151 184382 146747
rect 185398 146731 185450 146737
rect 185398 146673 185450 146679
rect 184438 146657 184490 146663
rect 185410 146631 185438 146673
rect 184438 146599 184490 146605
rect 185396 146622 185452 146631
rect 184340 145142 184396 145151
rect 184340 145077 184396 145086
rect 184450 144411 184478 146599
rect 185396 146557 185452 146566
rect 184436 144402 184492 144411
rect 184436 144337 184492 144346
rect 184534 143993 184586 143999
rect 184534 143935 184586 143941
rect 184438 143919 184490 143925
rect 184438 143861 184490 143867
rect 184342 143845 184394 143851
rect 184342 143787 184394 143793
rect 184354 142783 184382 143787
rect 184340 142774 184396 142783
rect 184340 142709 184396 142718
rect 184450 142191 184478 143861
rect 184436 142182 184492 142191
rect 184436 142117 184492 142126
rect 184546 141303 184574 143935
rect 184630 143771 184682 143777
rect 184630 143713 184682 143719
rect 184642 143671 184670 143713
rect 184628 143662 184684 143671
rect 184628 143597 184684 143606
rect 184532 141294 184588 141303
rect 184532 141229 184588 141238
rect 184534 141107 184586 141113
rect 184534 141049 184586 141055
rect 184438 141033 184490 141039
rect 184438 140975 184490 140981
rect 184342 140959 184394 140965
rect 184342 140901 184394 140907
rect 184354 140563 184382 140901
rect 184340 140554 184396 140563
rect 184340 140489 184396 140498
rect 184450 139823 184478 140975
rect 184436 139814 184492 139823
rect 184436 139749 184492 139758
rect 184546 138935 184574 141049
rect 184532 138926 184588 138935
rect 184532 138861 184588 138870
rect 185506 135975 185534 179973
rect 185698 175694 185726 242799
rect 185794 182447 185822 246647
rect 185974 246261 186026 246267
rect 185974 246203 186026 246209
rect 185878 242783 185930 242789
rect 185878 242725 185930 242731
rect 185890 195854 185918 242725
rect 185986 202871 186014 246203
rect 186082 213527 186110 254935
rect 186262 254919 186314 254925
rect 186262 254861 186314 254867
rect 186166 246335 186218 246341
rect 186166 246277 186218 246283
rect 186068 213518 186124 213527
rect 186068 213453 186124 213462
rect 186178 204351 186206 246277
rect 186274 215007 186302 254861
rect 186742 249221 186794 249227
rect 186742 249163 186794 249169
rect 186454 249147 186506 249153
rect 186454 249089 186506 249095
rect 186358 246631 186410 246637
rect 186358 246573 186410 246579
rect 186260 214998 186316 215007
rect 186260 214933 186316 214942
rect 186370 207311 186398 246573
rect 186466 210567 186494 249089
rect 186646 246557 186698 246563
rect 186646 246499 186698 246505
rect 186550 246483 186602 246489
rect 186550 246425 186602 246431
rect 186452 210558 186508 210567
rect 186452 210493 186508 210502
rect 186356 207302 186412 207311
rect 186356 207237 186412 207246
rect 186562 205239 186590 246425
rect 186658 209087 186686 246499
rect 186754 216487 186782 249163
rect 186934 246409 186986 246415
rect 186934 246351 186986 246357
rect 186838 245003 186890 245009
rect 186838 244945 186890 244951
rect 186850 221075 186878 244945
rect 186836 221066 186892 221075
rect 186836 221001 186892 221010
rect 186946 218115 186974 246351
rect 187124 243414 187180 243423
rect 187124 243349 187180 243358
rect 187030 242709 187082 242715
rect 187030 242651 187082 242657
rect 187042 220335 187070 242651
rect 187138 227545 187166 243349
rect 187126 227539 187178 227545
rect 187126 227481 187178 227487
rect 187138 226139 187166 227481
rect 187126 226133 187178 226139
rect 187126 226075 187178 226081
rect 187028 220326 187084 220335
rect 187028 220261 187084 220270
rect 186932 218106 186988 218115
rect 186932 218041 186988 218050
rect 186740 216478 186796 216487
rect 186740 216413 186796 216422
rect 187030 212887 187082 212893
rect 187030 212829 187082 212835
rect 187042 212047 187070 212829
rect 187028 212038 187084 212047
rect 187028 211973 187084 211982
rect 186644 209078 186700 209087
rect 186644 209013 186700 209022
rect 186548 205230 186604 205239
rect 186548 205165 186604 205174
rect 186164 204342 186220 204351
rect 186164 204277 186220 204286
rect 185972 202862 186028 202871
rect 185972 202797 186028 202806
rect 187234 199171 187262 257747
rect 190196 251702 190252 251711
rect 190196 251637 190252 251646
rect 190210 228581 190238 251637
rect 190198 228575 190250 228581
rect 190198 228517 190250 228523
rect 190774 227539 190826 227545
rect 190774 227481 190826 227487
rect 190786 221792 190814 227481
rect 190786 221764 190862 221792
rect 190834 221482 190862 221764
rect 191554 221482 191582 259333
rect 420418 259291 420446 259777
rect 420406 259285 420458 259291
rect 420406 259227 420458 259233
rect 420404 257030 420460 257039
rect 420404 256965 420460 256974
rect 420418 256405 420446 256965
rect 420406 256399 420458 256405
rect 420406 256341 420458 256347
rect 420404 255254 420460 255263
rect 420404 255189 420460 255198
rect 420418 253519 420446 255189
rect 420406 253513 420458 253519
rect 420406 253455 420458 253461
rect 603286 253513 603338 253519
rect 603286 253455 603338 253461
rect 420404 252886 420460 252895
rect 420404 252821 420460 252830
rect 420418 250633 420446 252821
rect 420406 250627 420458 250633
rect 420406 250569 420458 250575
rect 420308 250518 420364 250527
rect 420308 250453 420364 250462
rect 420322 247821 420350 250453
rect 420404 248150 420460 248159
rect 420404 248085 420460 248094
rect 420310 247815 420362 247821
rect 420310 247757 420362 247763
rect 420418 247747 420446 248085
rect 420406 247741 420458 247747
rect 420406 247683 420458 247689
rect 420404 245338 420460 245347
rect 420404 245273 420460 245282
rect 420418 244861 420446 245273
rect 420406 244855 420458 244861
rect 420406 244797 420458 244803
rect 420308 243562 420364 243571
rect 420308 243497 420364 243506
rect 420322 241975 420350 243497
rect 420310 241969 420362 241975
rect 420310 241911 420362 241917
rect 600406 241969 600458 241975
rect 600406 241911 600458 241917
rect 412436 241490 412492 241499
rect 412436 241425 412492 241434
rect 567380 241490 567436 241499
rect 567380 241425 567436 241434
rect 412244 240750 412300 240759
rect 412244 240685 412300 240694
rect 412148 240454 412204 240463
rect 412148 240389 412204 240398
rect 412052 240306 412108 240315
rect 412052 240241 412108 240250
rect 368592 239977 368702 239996
rect 412066 239977 412094 240241
rect 368592 239971 368714 239977
rect 368592 239968 368662 239971
rect 368662 239913 368714 239919
rect 412054 239971 412106 239977
rect 412054 239913 412106 239919
rect 412162 239903 412190 240389
rect 409558 239897 409610 239903
rect 350448 239829 350750 239848
rect 409344 239845 409558 239848
rect 409344 239839 409610 239845
rect 412150 239897 412202 239903
rect 412150 239839 412202 239845
rect 350448 239823 350762 239829
rect 350448 239820 350710 239823
rect 409344 239820 409598 239839
rect 350710 239765 350762 239771
rect 360022 239749 360074 239755
rect 192418 233391 192446 239686
rect 192768 239672 192926 239700
rect 192898 233613 192926 239672
rect 192994 239672 193152 239700
rect 192886 233607 192938 233613
rect 192886 233549 192938 233555
rect 192406 233385 192458 233391
rect 192406 233327 192458 233333
rect 192310 228575 192362 228581
rect 192310 228517 192362 228523
rect 192322 221482 192350 228517
rect 192994 221792 193022 239672
rect 193474 233317 193502 239686
rect 193858 233391 193886 239686
rect 194242 233539 194270 239686
rect 194230 233533 194282 233539
rect 194230 233475 194282 233481
rect 194626 233465 194654 239686
rect 194976 239672 195230 239700
rect 195360 239672 195614 239700
rect 194614 233459 194666 233465
rect 194614 233401 194666 233407
rect 193750 233385 193802 233391
rect 193750 233327 193802 233333
rect 193846 233385 193898 233391
rect 193846 233327 193898 233333
rect 193462 233311 193514 233317
rect 193462 233253 193514 233259
rect 192994 221764 193070 221792
rect 193042 221482 193070 221764
rect 193762 221482 193790 233327
rect 195202 233317 195230 239672
rect 195586 233613 195614 239672
rect 195682 233687 195710 239686
rect 195670 233681 195722 233687
rect 195670 233623 195722 233629
rect 195286 233607 195338 233613
rect 195286 233549 195338 233555
rect 195574 233607 195626 233613
rect 195574 233549 195626 233555
rect 194614 233311 194666 233317
rect 194614 233253 194666 233259
rect 195190 233311 195242 233317
rect 195190 233253 195242 233259
rect 194626 221482 194654 233253
rect 195298 221792 195326 233549
rect 196054 233459 196106 233465
rect 196054 233401 196106 233407
rect 195862 233311 195914 233317
rect 195862 233253 195914 233259
rect 195298 221764 195374 221792
rect 195346 221482 195374 221764
rect 195766 221767 195818 221773
rect 195874 221755 195902 233253
rect 195818 221727 195902 221755
rect 195766 221709 195818 221715
rect 196066 221482 196094 233401
rect 196162 233317 196190 239686
rect 196546 233465 196574 239686
rect 196930 233835 196958 239686
rect 197280 239672 197534 239700
rect 197664 239672 197918 239700
rect 197506 233909 197534 239672
rect 197494 233903 197546 233909
rect 197494 233845 197546 233851
rect 196918 233829 196970 233835
rect 196918 233771 196970 233777
rect 196534 233459 196586 233465
rect 196534 233401 196586 233407
rect 197890 233391 197918 239672
rect 197986 233761 198014 239686
rect 198370 233983 198398 239686
rect 198754 234057 198782 239686
rect 198742 234051 198794 234057
rect 198742 233993 198794 233999
rect 198358 233977 198410 233983
rect 198358 233919 198410 233925
rect 197974 233755 198026 233761
rect 197974 233697 198026 233703
rect 199138 233539 199166 239686
rect 199488 239672 199742 239700
rect 199968 239672 200222 239700
rect 198358 233533 198410 233539
rect 198358 233475 198410 233481
rect 199126 233533 199178 233539
rect 199126 233475 199178 233481
rect 196822 233385 196874 233391
rect 196822 233327 196874 233333
rect 197878 233385 197930 233391
rect 197878 233327 197930 233333
rect 196150 233311 196202 233317
rect 196150 233253 196202 233259
rect 196834 221482 196862 233327
rect 197542 221767 197594 221773
rect 197542 221709 197594 221715
rect 197554 221482 197582 221709
rect 198370 221482 198398 233475
rect 199714 233317 199742 239672
rect 200194 234131 200222 239672
rect 200290 234205 200318 239686
rect 200278 234199 200330 234205
rect 200278 234141 200330 234147
rect 200182 234125 200234 234131
rect 200182 234067 200234 234073
rect 199798 233607 199850 233613
rect 199798 233549 199850 233555
rect 199126 233311 199178 233317
rect 199126 233253 199178 233259
rect 199702 233311 199754 233317
rect 199702 233253 199754 233259
rect 199138 221482 199166 233253
rect 199810 221792 199838 233549
rect 200674 233465 200702 239686
rect 201058 233613 201086 239686
rect 201408 239672 201566 239700
rect 201792 239672 202046 239700
rect 202176 239672 202430 239700
rect 201538 234353 201566 239672
rect 202018 234649 202046 239672
rect 202006 234643 202058 234649
rect 202006 234585 202058 234591
rect 201526 234347 201578 234353
rect 201526 234289 201578 234295
rect 201334 233681 201386 233687
rect 201334 233623 201386 233629
rect 201046 233607 201098 233613
rect 201046 233549 201098 233555
rect 200566 233459 200618 233465
rect 200566 233401 200618 233407
rect 200662 233459 200714 233465
rect 200662 233401 200714 233407
rect 199810 221764 199886 221792
rect 199858 221482 199886 221764
rect 200578 221482 200606 233401
rect 201346 221482 201374 233623
rect 202402 233391 202430 239672
rect 202498 233687 202526 239686
rect 202882 234797 202910 239686
rect 203266 235093 203294 239686
rect 203712 239672 203966 239700
rect 204096 239672 204254 239700
rect 203254 235087 203306 235093
rect 203254 235029 203306 235035
rect 202870 234791 202922 234797
rect 202870 234733 202922 234739
rect 202870 233829 202922 233835
rect 202870 233771 202922 233777
rect 202486 233681 202538 233687
rect 202486 233623 202538 233629
rect 202102 233385 202154 233391
rect 202102 233327 202154 233333
rect 202390 233385 202442 233391
rect 202390 233327 202442 233333
rect 202114 221792 202142 233327
rect 202114 221764 202190 221792
rect 202162 221482 202190 221764
rect 202882 221482 202910 233771
rect 203938 233761 203966 239672
rect 204226 234575 204254 239672
rect 204418 239672 204480 239700
rect 204214 234569 204266 234575
rect 204214 234511 204266 234517
rect 204418 234427 204446 239672
rect 204802 234723 204830 239686
rect 204790 234717 204842 234723
rect 204790 234659 204842 234665
rect 204406 234421 204458 234427
rect 204406 234363 204458 234369
rect 204310 233903 204362 233909
rect 204310 233845 204362 233851
rect 203638 233755 203690 233761
rect 203638 233697 203690 233703
rect 203926 233755 203978 233761
rect 203926 233697 203978 233703
rect 203650 221482 203678 233697
rect 204322 221755 204350 233845
rect 205186 233835 205214 239686
rect 205174 233829 205226 233835
rect 205174 233771 205226 233777
rect 205570 233539 205598 239686
rect 205920 239672 206174 239700
rect 206304 239672 206558 239700
rect 206688 239672 206942 239700
rect 206146 235167 206174 239672
rect 206134 235161 206186 235167
rect 206134 235103 206186 235109
rect 206530 234501 206558 239672
rect 206518 234495 206570 234501
rect 206518 234437 206570 234443
rect 206914 233983 206942 239672
rect 207010 235389 207038 239686
rect 207490 235981 207518 239686
rect 207478 235975 207530 235981
rect 207478 235917 207530 235923
rect 206998 235383 207050 235389
rect 206998 235325 207050 235331
rect 207874 234279 207902 239686
rect 208224 239672 208478 239700
rect 208608 239672 208862 239700
rect 208450 236055 208478 239672
rect 208438 236049 208490 236055
rect 208438 235991 208490 235997
rect 208834 235019 208862 239672
rect 208930 235833 208958 239686
rect 208918 235827 208970 235833
rect 208918 235769 208970 235775
rect 208822 235013 208874 235019
rect 208822 234955 208874 234961
rect 209314 234871 209342 239686
rect 209698 235907 209726 239686
rect 209686 235901 209738 235907
rect 209686 235843 209738 235849
rect 210082 235611 210110 239686
rect 210432 239672 210686 239700
rect 210816 239672 211070 239700
rect 210658 235685 210686 239672
rect 210646 235679 210698 235685
rect 210646 235621 210698 235627
rect 210070 235605 210122 235611
rect 210070 235547 210122 235553
rect 211042 234945 211070 239672
rect 211234 235759 211262 239686
rect 211222 235753 211274 235759
rect 211222 235695 211274 235701
rect 211510 235087 211562 235093
rect 211510 235029 211562 235035
rect 211030 234939 211082 234945
rect 211030 234881 211082 234887
rect 209302 234865 209354 234871
rect 209302 234807 209354 234813
rect 210166 234421 210218 234427
rect 210166 234363 210218 234369
rect 207862 234273 207914 234279
rect 207862 234215 207914 234221
rect 210178 234131 210206 234363
rect 210358 234199 210410 234205
rect 210358 234141 210410 234147
rect 208822 234125 208874 234131
rect 208822 234067 208874 234073
rect 210166 234125 210218 234131
rect 210166 234067 210218 234073
rect 207382 234051 207434 234057
rect 207382 233993 207434 233999
rect 205942 233977 205994 233983
rect 205942 233919 205994 233925
rect 206902 233977 206954 233983
rect 206902 233919 206954 233925
rect 205078 233533 205130 233539
rect 205078 233475 205130 233481
rect 205558 233533 205610 233539
rect 205558 233475 205610 233481
rect 204322 221727 204446 221755
rect 204418 221681 204446 221727
rect 204370 221653 204446 221681
rect 204370 221482 204398 221653
rect 205090 221482 205118 233475
rect 205954 221496 205982 233919
rect 206614 233311 206666 233317
rect 206614 233253 206666 233259
rect 205920 221468 205982 221496
rect 206626 221496 206654 233253
rect 206626 221468 206688 221496
rect 207394 221482 207422 233993
rect 208150 233459 208202 233465
rect 208150 233401 208202 233407
rect 208162 221496 208190 233401
rect 208128 221468 208190 221496
rect 208834 221496 208862 234067
rect 209686 233607 209738 233613
rect 209686 233549 209738 233555
rect 208834 221468 208896 221496
rect 209698 221482 209726 233549
rect 210370 221681 210398 234141
rect 211522 233983 211550 235029
rect 211510 233977 211562 233983
rect 211510 233919 211562 233925
rect 211618 233835 211646 239686
rect 212002 235463 212030 239686
rect 211990 235457 212042 235463
rect 211990 235399 212042 235405
rect 211894 234347 211946 234353
rect 211894 234289 211946 234295
rect 211606 233829 211658 233835
rect 211606 233771 211658 233777
rect 211126 233385 211178 233391
rect 211126 233327 211178 233333
rect 210370 221653 210446 221681
rect 210418 221482 210446 221653
rect 211138 221482 211166 233327
rect 211906 221482 211934 234289
rect 212386 227027 212414 239686
rect 212736 239672 212990 239700
rect 212962 235537 212990 239672
rect 213058 239672 213120 239700
rect 212950 235531 213002 235537
rect 212950 235473 213002 235479
rect 212566 233681 212618 233687
rect 212566 233623 212618 233629
rect 212374 227021 212426 227027
rect 212374 226963 212426 226969
rect 212578 221681 212606 233623
rect 213058 226065 213086 239672
rect 213442 235093 213470 239686
rect 213430 235087 213482 235093
rect 213430 235029 213482 235035
rect 213430 234643 213482 234649
rect 213430 234585 213482 234591
rect 213046 226059 213098 226065
rect 213046 226001 213098 226007
rect 212578 221653 212654 221681
rect 212626 221482 212654 221653
rect 213442 221482 213470 234585
rect 213826 227545 213854 239686
rect 214210 235315 214238 239686
rect 214198 235309 214250 235315
rect 214198 235251 214250 235257
rect 214486 233903 214538 233909
rect 214486 233845 214538 233851
rect 214198 233755 214250 233761
rect 214198 233697 214250 233703
rect 213814 227539 213866 227545
rect 213814 227481 213866 227487
rect 214210 221482 214238 233697
rect 214498 233687 214526 233845
rect 214486 233681 214538 233687
rect 214486 233623 214538 233629
rect 214594 226361 214622 239686
rect 215040 239672 215294 239700
rect 215424 239672 215678 239700
rect 214774 234791 214826 234797
rect 214774 234733 214826 234739
rect 214582 226355 214634 226361
rect 214582 226297 214634 226303
rect 214786 221792 214814 234733
rect 214870 234717 214922 234723
rect 214870 234659 214922 234665
rect 214882 234279 214910 234659
rect 214870 234273 214922 234279
rect 214870 234215 214922 234221
rect 215266 229543 215294 239672
rect 215542 234569 215594 234575
rect 215542 234511 215594 234517
rect 215254 229537 215306 229543
rect 215254 229479 215306 229485
rect 215554 226084 215582 234511
rect 215650 226213 215678 239672
rect 215746 227397 215774 239686
rect 215926 235161 215978 235167
rect 215926 235103 215978 235109
rect 215938 234427 215966 235103
rect 215926 234421 215978 234427
rect 215926 234363 215978 234369
rect 216130 227471 216158 239686
rect 216514 236174 216542 239686
rect 216864 239672 217118 239700
rect 217248 239672 217502 239700
rect 217632 239672 217886 239700
rect 216514 236146 216638 236174
rect 216502 233977 216554 233983
rect 216502 233919 216554 233925
rect 216118 227465 216170 227471
rect 216118 227407 216170 227413
rect 215734 227391 215786 227397
rect 215734 227333 215786 227339
rect 215638 226207 215690 226213
rect 215638 226149 215690 226155
rect 215554 226056 215678 226084
rect 214786 221764 214958 221792
rect 214930 221482 214958 221764
rect 215650 221482 215678 226056
rect 216514 221482 216542 233919
rect 216610 232725 216638 236146
rect 216598 232719 216650 232725
rect 216598 232661 216650 232667
rect 217090 225843 217118 239672
rect 217174 233681 217226 233687
rect 217174 233623 217226 233629
rect 217078 225837 217130 225843
rect 217078 225779 217130 225785
rect 217186 221792 217214 233623
rect 217474 225991 217502 239672
rect 217858 226287 217886 239672
rect 217954 236174 217982 239686
rect 217954 236146 218078 236174
rect 217942 234125 217994 234131
rect 217942 234067 217994 234073
rect 217846 226281 217898 226287
rect 217846 226223 217898 226229
rect 217462 225985 217514 225991
rect 217462 225927 217514 225933
rect 217186 221764 217262 221792
rect 217234 221482 217262 221764
rect 217954 221482 217982 234067
rect 218050 232577 218078 236146
rect 218038 232571 218090 232577
rect 218038 232513 218090 232519
rect 218338 226139 218366 239686
rect 218710 233755 218762 233761
rect 218710 233697 218762 233703
rect 218326 226133 218378 226139
rect 218326 226075 218378 226081
rect 218722 221482 218750 233697
rect 218818 225917 218846 239686
rect 219168 239672 219422 239700
rect 219552 239672 219806 239700
rect 219936 239672 220190 239700
rect 219394 236174 219422 239672
rect 219394 236146 219518 236174
rect 219382 234273 219434 234279
rect 219382 234215 219434 234221
rect 218806 225911 218858 225917
rect 218806 225853 218858 225859
rect 219394 221792 219422 234215
rect 219490 227175 219518 236146
rect 219778 232651 219806 239672
rect 219766 232645 219818 232651
rect 219766 232587 219818 232593
rect 220162 229765 220190 239672
rect 220258 236174 220286 239686
rect 220258 236146 220382 236174
rect 220246 234051 220298 234057
rect 220246 233993 220298 233999
rect 220150 229759 220202 229765
rect 220150 229701 220202 229707
rect 219478 227169 219530 227175
rect 219478 227111 219530 227117
rect 219394 221764 219470 221792
rect 219442 221482 219470 221764
rect 220258 221482 220286 233993
rect 220354 227249 220382 236146
rect 220642 235241 220670 239686
rect 221026 236174 221054 239686
rect 221376 239672 221630 239700
rect 221026 236146 221150 236174
rect 220630 235235 220682 235241
rect 220630 235177 220682 235183
rect 221014 234421 221066 234427
rect 221014 234363 221066 234369
rect 220342 227243 220394 227249
rect 220342 227185 220394 227191
rect 221026 221482 221054 234363
rect 221122 232429 221150 236146
rect 221110 232423 221162 232429
rect 221110 232365 221162 232371
rect 221602 229691 221630 239672
rect 221746 239404 221774 239686
rect 222144 239672 222398 239700
rect 221698 239376 221774 239404
rect 221590 229685 221642 229691
rect 221590 229627 221642 229633
rect 221698 226953 221726 239376
rect 221782 235383 221834 235389
rect 221782 235325 221834 235331
rect 221686 226947 221738 226953
rect 221686 226889 221738 226895
rect 221794 221792 221822 235325
rect 222370 234723 222398 239672
rect 222358 234717 222410 234723
rect 222358 234659 222410 234665
rect 222454 234347 222506 234353
rect 222454 234289 222506 234295
rect 221746 221764 221822 221792
rect 221746 221482 221774 221764
rect 222466 221482 222494 234289
rect 222562 232503 222590 239686
rect 222550 232497 222602 232503
rect 222550 232439 222602 232445
rect 222946 232355 222974 239686
rect 223222 236049 223274 236055
rect 223222 235991 223274 235997
rect 222934 232349 222986 232355
rect 222934 232291 222986 232297
rect 223234 221482 223262 235991
rect 223330 226805 223358 239686
rect 223680 239672 223934 239700
rect 224064 239672 224318 239700
rect 223906 235389 223934 239672
rect 223990 235975 224042 235981
rect 223990 235917 224042 235923
rect 223894 235383 223946 235389
rect 223894 235325 223946 235331
rect 223318 226799 223370 226805
rect 223318 226741 223370 226747
rect 224002 221792 224030 235917
rect 224290 232207 224318 239672
rect 224278 232201 224330 232207
rect 224278 232143 224330 232149
rect 224386 228507 224414 239686
rect 224770 236174 224798 239686
rect 224770 236146 224894 236174
rect 224758 235013 224810 235019
rect 224758 234955 224810 234961
rect 224374 228501 224426 228507
rect 224374 228443 224426 228449
rect 224002 221764 224078 221792
rect 224050 221482 224078 221764
rect 224770 221482 224798 234955
rect 224866 226879 224894 236146
rect 225154 234797 225182 239686
rect 225538 235019 225566 239686
rect 225984 239672 226238 239700
rect 226368 239672 226622 239700
rect 226210 236174 226238 239672
rect 226210 236146 226334 236174
rect 226198 235901 226250 235907
rect 226198 235843 226250 235849
rect 225526 235013 225578 235019
rect 225526 234955 225578 234961
rect 225142 234791 225194 234797
rect 225142 234733 225194 234739
rect 225526 234199 225578 234205
rect 225526 234141 225578 234147
rect 224854 226873 224906 226879
rect 224854 226815 224906 226821
rect 225538 221482 225566 234141
rect 226210 221792 226238 235843
rect 226306 232281 226334 236146
rect 226294 232275 226346 232281
rect 226294 232217 226346 232223
rect 226594 226731 226622 239672
rect 226690 233317 226718 239686
rect 226966 235827 227018 235833
rect 226966 235769 227018 235775
rect 226678 233311 226730 233317
rect 226678 233253 226730 233259
rect 226582 226725 226634 226731
rect 226582 226667 226634 226673
rect 226210 221764 226286 221792
rect 226258 221482 226286 221764
rect 226978 221482 227006 235769
rect 227074 232133 227102 239686
rect 227062 232127 227114 232133
rect 227062 232069 227114 232075
rect 227458 229987 227486 239686
rect 227842 236174 227870 239686
rect 228192 239672 228446 239700
rect 228576 239672 228830 239700
rect 227842 236146 227966 236174
rect 227830 235605 227882 235611
rect 227830 235547 227882 235553
rect 227446 229981 227498 229987
rect 227446 229923 227498 229929
rect 227842 221482 227870 235547
rect 227938 226657 227966 236146
rect 228418 233391 228446 239672
rect 228502 234865 228554 234871
rect 228502 234807 228554 234813
rect 228406 233385 228458 233391
rect 228406 233327 228458 233333
rect 227926 226651 227978 226657
rect 227926 226593 227978 226599
rect 228514 221792 228542 234807
rect 228802 228581 228830 239672
rect 228898 230357 228926 239686
rect 229296 239672 229598 239700
rect 229270 235753 229322 235759
rect 229270 235695 229322 235701
rect 228886 230351 228938 230357
rect 228886 230293 228938 230299
rect 228790 228575 228842 228581
rect 228790 228517 228842 228523
rect 228514 221764 228590 221792
rect 228562 221482 228590 221764
rect 229282 221482 229310 235695
rect 229570 226509 229598 239672
rect 229762 234871 229790 239686
rect 230112 239672 230366 239700
rect 230496 239672 230750 239700
rect 230880 239672 231134 239700
rect 230038 235679 230090 235685
rect 230038 235621 230090 235627
rect 229750 234865 229802 234871
rect 229750 234807 229802 234813
rect 229558 226503 229610 226509
rect 229558 226445 229610 226451
rect 230050 221482 230078 235621
rect 230338 228655 230366 239672
rect 230722 236174 230750 239672
rect 230722 236146 230846 236174
rect 230710 233829 230762 233835
rect 230710 233771 230762 233777
rect 230326 228649 230378 228655
rect 230326 228591 230378 228597
rect 230722 221792 230750 233771
rect 230818 229321 230846 236146
rect 230806 229315 230858 229321
rect 230806 229257 230858 229263
rect 231106 226583 231134 239672
rect 231202 235759 231230 239686
rect 231600 239672 231902 239700
rect 231190 235753 231242 235759
rect 231190 235695 231242 235701
rect 231574 234939 231626 234945
rect 231574 234881 231626 234887
rect 231094 226577 231146 226583
rect 231094 226519 231146 226525
rect 230722 221764 230798 221792
rect 230770 221482 230798 221764
rect 231586 221482 231614 234881
rect 231874 229395 231902 239672
rect 231862 229389 231914 229395
rect 231862 229331 231914 229337
rect 231970 229173 231998 239686
rect 232320 239672 232574 239700
rect 232704 239672 232958 239700
rect 233088 239672 233246 239700
rect 232342 235531 232394 235537
rect 232342 235473 232394 235479
rect 231958 229167 232010 229173
rect 231958 229109 232010 229115
rect 232354 221482 232382 235473
rect 232546 226435 232574 239672
rect 232930 235167 232958 239672
rect 233014 235457 233066 235463
rect 233014 235399 233066 235405
rect 232918 235161 232970 235167
rect 232918 235103 232970 235109
rect 232534 226429 232586 226435
rect 232534 226371 232586 226377
rect 233026 221792 233054 235399
rect 233218 231911 233246 239672
rect 233398 235087 233450 235093
rect 233398 235029 233450 235035
rect 233410 233465 233438 235029
rect 233398 233459 233450 233465
rect 233398 233401 233450 233407
rect 233206 231905 233258 231911
rect 233206 231847 233258 231853
rect 233506 229247 233534 239686
rect 233890 232059 233918 239686
rect 234274 235907 234302 239686
rect 234624 239672 234878 239700
rect 235008 239672 235262 239700
rect 235392 239672 235646 239700
rect 234262 235901 234314 235907
rect 234262 235843 234314 235849
rect 233878 232053 233930 232059
rect 233878 231995 233930 232001
rect 234850 231985 234878 239672
rect 234838 231979 234890 231985
rect 234838 231921 234890 231927
rect 233494 229241 233546 229247
rect 233494 229183 233546 229189
rect 235234 229099 235262 239672
rect 235318 235309 235370 235315
rect 235318 235251 235370 235257
rect 235222 229093 235274 229099
rect 235222 229035 235274 229041
rect 234550 227021 234602 227027
rect 234550 226963 234602 226969
rect 233782 226059 233834 226065
rect 233782 226001 233834 226007
rect 233026 221764 233102 221792
rect 233074 221482 233102 221764
rect 233794 221482 233822 226001
rect 234562 221482 234590 226963
rect 235330 221496 235358 235251
rect 235618 234427 235646 239672
rect 235714 235093 235742 239686
rect 235702 235087 235754 235093
rect 235702 235029 235754 235035
rect 235606 234421 235658 234427
rect 235606 234363 235658 234369
rect 235990 233459 236042 233465
rect 235990 233401 236042 233407
rect 236002 228008 236030 233401
rect 236098 231837 236126 239686
rect 236482 235611 236510 239686
rect 236832 239672 237086 239700
rect 237312 239672 237566 239700
rect 236470 235605 236522 235611
rect 236470 235547 236522 235553
rect 237058 234575 237086 239672
rect 237538 235833 237566 239672
rect 237526 235827 237578 235833
rect 237526 235769 237578 235775
rect 237046 234569 237098 234575
rect 237046 234511 237098 234517
rect 236374 233385 236426 233391
rect 236374 233327 236426 233333
rect 236086 231831 236138 231837
rect 236086 231773 236138 231779
rect 236002 227980 236126 228008
rect 235330 221468 235392 221496
rect 236098 221482 236126 227980
rect 236386 227027 236414 233327
rect 237634 232873 237662 239686
rect 238018 235537 238046 239686
rect 238006 235531 238058 235537
rect 238006 235473 238058 235479
rect 237622 232867 237674 232873
rect 237622 232809 237674 232815
rect 238402 229025 238430 239686
rect 238390 229019 238442 229025
rect 238390 228961 238442 228967
rect 237526 227539 237578 227545
rect 237526 227481 237578 227487
rect 236374 227021 236426 227027
rect 236374 226963 236426 226969
rect 236854 226355 236906 226361
rect 236854 226297 236906 226303
rect 236866 221496 236894 226297
rect 236832 221468 236894 221496
rect 237538 221496 237566 227481
rect 238390 227391 238442 227397
rect 238390 227333 238442 227339
rect 237538 221468 237600 221496
rect 238402 221482 238430 227333
rect 238786 227101 238814 239686
rect 239136 239672 239390 239700
rect 239520 239672 239774 239700
rect 239362 235315 239390 239672
rect 239350 235309 239402 235315
rect 239350 235251 239402 235257
rect 238966 233311 239018 233317
rect 238966 233253 239018 233259
rect 238774 227095 238826 227101
rect 238774 227037 238826 227043
rect 238978 226065 239006 233253
rect 239746 229839 239774 239672
rect 239842 234353 239870 239686
rect 240226 236129 240254 239686
rect 240214 236123 240266 236129
rect 240214 236065 240266 236071
rect 239830 234347 239882 234353
rect 239830 234289 239882 234295
rect 240610 233539 240638 239686
rect 240598 233533 240650 233539
rect 240598 233475 240650 233481
rect 239734 229833 239786 229839
rect 239734 229775 239786 229781
rect 241090 229617 241118 239686
rect 241440 239672 241694 239700
rect 241078 229611 241130 229617
rect 241078 229553 241130 229559
rect 239062 229537 239114 229543
rect 239062 229479 239114 229485
rect 238966 226059 239018 226065
rect 238966 226001 239018 226007
rect 239074 221792 239102 229479
rect 241666 228729 241694 239672
rect 241810 239404 241838 239686
rect 241810 239376 241886 239404
rect 241858 236174 241886 239376
rect 241762 236146 241886 236174
rect 241654 228723 241706 228729
rect 241654 228665 241706 228671
rect 239830 227465 239882 227471
rect 239830 227407 239882 227413
rect 239074 221764 239150 221792
rect 239122 221482 239150 221764
rect 239842 221482 239870 227407
rect 241762 226361 241790 236146
rect 242146 235463 242174 239686
rect 242134 235457 242186 235463
rect 242134 235399 242186 235405
rect 241846 235235 241898 235241
rect 241846 235177 241898 235183
rect 241750 226355 241802 226361
rect 241750 226297 241802 226303
rect 240598 226207 240650 226213
rect 240598 226149 240650 226155
rect 240610 221482 240638 226149
rect 241270 225985 241322 225991
rect 241270 225927 241322 225933
rect 241282 221792 241310 225927
rect 241858 225399 241886 235177
rect 242134 232719 242186 232725
rect 242134 232661 242186 232667
rect 241846 225393 241898 225399
rect 241846 225335 241898 225341
rect 241282 221764 241358 221792
rect 241330 221482 241358 221764
rect 242146 221482 242174 232661
rect 242530 228803 242558 239686
rect 242914 233835 242942 239686
rect 243298 235981 243326 239686
rect 243648 239672 243902 239700
rect 244032 239672 244286 239700
rect 243286 235975 243338 235981
rect 243286 235917 243338 235923
rect 243874 234945 243902 239672
rect 243862 234939 243914 234945
rect 243862 234881 243914 234887
rect 243958 234717 244010 234723
rect 243958 234659 244010 234665
rect 242902 233829 242954 233835
rect 242902 233771 242954 233777
rect 242518 228797 242570 228803
rect 242518 228739 242570 228745
rect 242902 226281 242954 226287
rect 242902 226223 242954 226229
rect 242914 221482 242942 226223
rect 243574 225837 243626 225843
rect 243574 225779 243626 225785
rect 243586 221792 243614 225779
rect 243970 225473 243998 234659
rect 244258 229543 244286 239672
rect 244354 234279 244382 239686
rect 244726 235383 244778 235389
rect 244726 235325 244778 235331
rect 244342 234273 244394 234279
rect 244342 234215 244394 234221
rect 244246 229537 244298 229543
rect 244246 229479 244298 229485
rect 244738 225917 244766 235325
rect 244834 226065 244862 239686
rect 245110 232571 245162 232577
rect 245110 232513 245162 232519
rect 244822 226059 244874 226065
rect 244822 226001 244874 226007
rect 244342 225911 244394 225917
rect 244342 225853 244394 225859
rect 244726 225911 244778 225917
rect 244726 225853 244778 225859
rect 243958 225467 244010 225473
rect 243958 225409 244010 225415
rect 243586 221764 243662 221792
rect 243634 221482 243662 221764
rect 244354 221482 244382 225853
rect 245122 221482 245150 232513
rect 245218 231023 245246 239686
rect 245568 239672 245822 239700
rect 245952 239672 246206 239700
rect 246336 239672 246590 239700
rect 245206 231017 245258 231023
rect 245206 230959 245258 230965
rect 245794 228951 245822 239672
rect 245782 228945 245834 228951
rect 245782 228887 245834 228893
rect 246178 228877 246206 239672
rect 246166 228871 246218 228877
rect 246166 228813 246218 228819
rect 245878 227169 245930 227175
rect 245878 227111 245930 227117
rect 245890 221792 245918 227111
rect 246562 226213 246590 239672
rect 246658 234723 246686 239686
rect 246646 234717 246698 234723
rect 246646 234659 246698 234665
rect 247042 230283 247070 239686
rect 247426 234131 247454 239686
rect 247776 239672 248030 239700
rect 248160 239672 248414 239700
rect 248640 239672 248798 239700
rect 248002 236055 248030 239672
rect 247990 236049 248042 236055
rect 247990 235991 248042 235997
rect 247702 234791 247754 234797
rect 247702 234733 247754 234739
rect 247414 234125 247466 234131
rect 247414 234067 247466 234073
rect 247030 230277 247082 230283
rect 247030 230219 247082 230225
rect 247714 227249 247742 234733
rect 248086 232645 248138 232651
rect 248086 232587 248138 232593
rect 247414 227243 247466 227249
rect 247414 227185 247466 227191
rect 247702 227243 247754 227249
rect 247702 227185 247754 227191
rect 246550 226207 246602 226213
rect 246550 226149 246602 226155
rect 246646 226133 246698 226139
rect 246646 226075 246698 226081
rect 245890 221764 245966 221792
rect 245938 221482 245966 221764
rect 246658 221482 246686 226075
rect 247426 221482 247454 227185
rect 248098 221792 248126 232587
rect 248386 231541 248414 239672
rect 248374 231535 248426 231541
rect 248374 231477 248426 231483
rect 248770 230209 248798 239672
rect 248962 230431 248990 239686
rect 248950 230425 249002 230431
rect 248950 230367 249002 230373
rect 248758 230203 248810 230209
rect 248758 230145 248810 230151
rect 249346 227545 249374 239686
rect 249730 235241 249758 239686
rect 250080 239672 250238 239700
rect 249718 235235 249770 235241
rect 249718 235177 249770 235183
rect 249718 229759 249770 229765
rect 249718 229701 249770 229707
rect 249334 227539 249386 227545
rect 249334 227481 249386 227487
rect 248854 225393 248906 225399
rect 248854 225335 248906 225341
rect 248098 221764 248174 221792
rect 248146 221482 248174 221764
rect 248866 221482 248894 225335
rect 249730 221482 249758 229701
rect 250210 227915 250238 239672
rect 250450 239404 250478 239686
rect 250848 239672 251102 239700
rect 250450 239376 250526 239404
rect 250498 234501 250526 239376
rect 251074 234649 251102 239672
rect 251170 234797 251198 239686
rect 251158 234791 251210 234797
rect 251158 234733 251210 234739
rect 251062 234643 251114 234649
rect 251062 234585 251114 234591
rect 250486 234495 250538 234501
rect 250486 234437 250538 234443
rect 250582 234421 250634 234427
rect 250582 234363 250634 234369
rect 250594 228285 250622 234363
rect 251158 232423 251210 232429
rect 251158 232365 251210 232371
rect 250582 228279 250634 228285
rect 250582 228221 250634 228227
rect 250198 227909 250250 227915
rect 250198 227851 250250 227857
rect 250390 226947 250442 226953
rect 250390 226889 250442 226895
rect 250402 221792 250430 226889
rect 250402 221764 250478 221792
rect 250450 221482 250478 221764
rect 251170 221482 251198 232365
rect 251554 230061 251582 239686
rect 251938 230135 251966 239686
rect 252384 239672 252638 239700
rect 252768 239672 253022 239700
rect 252610 236174 252638 239672
rect 252610 236146 252734 236174
rect 251926 230129 251978 230135
rect 251926 230071 251978 230077
rect 251542 230055 251594 230061
rect 251542 229997 251594 230003
rect 252598 229685 252650 229691
rect 252598 229627 252650 229633
rect 251926 225467 251978 225473
rect 251926 225409 251978 225415
rect 251938 221482 251966 225409
rect 252610 221792 252638 229627
rect 252706 225103 252734 236146
rect 252994 231097 253022 239672
rect 252982 231091 253034 231097
rect 252982 231033 253034 231039
rect 253090 229913 253118 239686
rect 253474 233909 253502 239686
rect 253558 234865 253610 234871
rect 253558 234807 253610 234813
rect 253462 233903 253514 233909
rect 253462 233845 253514 233851
rect 253078 229907 253130 229913
rect 253078 229849 253130 229855
rect 253570 226953 253598 234807
rect 253858 227471 253886 239686
rect 254242 235389 254270 239686
rect 254592 239672 254846 239700
rect 254976 239672 255230 239700
rect 254230 235383 254282 235389
rect 254230 235325 254282 235331
rect 254230 232497 254282 232503
rect 254230 232439 254282 232445
rect 253846 227465 253898 227471
rect 253846 227407 253898 227413
rect 253558 226947 253610 226953
rect 253558 226889 253610 226895
rect 253462 226799 253514 226805
rect 253462 226741 253514 226747
rect 252694 225097 252746 225103
rect 252694 225039 252746 225045
rect 252610 221764 252686 221792
rect 252658 221482 252686 221764
rect 253474 221482 253502 226741
rect 254242 221482 254270 232439
rect 254818 229691 254846 239672
rect 255202 229765 255230 239672
rect 255298 234427 255326 239686
rect 255286 234421 255338 234427
rect 255286 234363 255338 234369
rect 255670 232349 255722 232355
rect 255670 232291 255722 232297
rect 255190 229759 255242 229765
rect 255190 229701 255242 229707
rect 254806 229685 254858 229691
rect 254806 229627 254858 229633
rect 254902 227095 254954 227101
rect 254902 227037 254954 227043
rect 254914 226361 254942 227037
rect 254902 226355 254954 226361
rect 254902 226297 254954 226303
rect 254998 226281 255050 226287
rect 254998 226223 255050 226229
rect 255010 226065 255038 226223
rect 254998 226059 255050 226065
rect 254998 226001 255050 226007
rect 254902 225911 254954 225917
rect 254902 225853 254954 225859
rect 254914 221792 254942 225853
rect 254914 221764 254990 221792
rect 254962 221482 254990 221764
rect 255682 221482 255710 232291
rect 255778 231615 255806 239686
rect 255766 231609 255818 231615
rect 255766 231551 255818 231557
rect 256162 231171 256190 239686
rect 256546 234205 256574 239686
rect 256896 239672 257150 239700
rect 257280 239672 257534 239700
rect 256534 234199 256586 234205
rect 256534 234141 256586 234147
rect 256150 231165 256202 231171
rect 256150 231107 256202 231113
rect 256438 226873 256490 226879
rect 256438 226815 256490 226821
rect 256450 221482 256478 226815
rect 257122 226065 257150 239672
rect 257506 234871 257534 239672
rect 257494 234865 257546 234871
rect 257494 234807 257546 234813
rect 257206 232201 257258 232207
rect 257206 232143 257258 232149
rect 257110 226059 257162 226065
rect 257110 226001 257162 226007
rect 257218 221792 257246 232143
rect 257602 231245 257630 239686
rect 257986 233317 258014 239686
rect 258070 234569 258122 234575
rect 258070 234511 258122 234517
rect 257974 233311 258026 233317
rect 257974 233253 258026 233259
rect 257590 231239 257642 231245
rect 257590 231181 257642 231187
rect 258082 228137 258110 234511
rect 258370 233761 258398 239686
rect 258358 233755 258410 233761
rect 258358 233697 258410 233703
rect 258754 231689 258782 239686
rect 259104 239672 259166 239700
rect 259584 239672 259838 239700
rect 259030 235753 259082 235759
rect 259030 235695 259082 235701
rect 258742 231683 258794 231689
rect 258742 231625 258794 231631
rect 258742 228501 258794 228507
rect 258742 228443 258794 228449
rect 258070 228131 258122 228137
rect 258070 228073 258122 228079
rect 257974 227243 258026 227249
rect 257974 227185 258026 227191
rect 257218 221764 257294 221792
rect 257266 221482 257294 221764
rect 257986 221482 258014 227185
rect 258754 221482 258782 228443
rect 259042 227101 259070 235695
rect 259138 231763 259166 239672
rect 259810 234057 259838 239672
rect 259798 234051 259850 234057
rect 259798 233993 259850 233999
rect 259906 233613 259934 239686
rect 260290 235019 260318 239686
rect 260182 235013 260234 235019
rect 260182 234955 260234 234961
rect 260278 235013 260330 235019
rect 260278 234955 260330 234961
rect 259894 233607 259946 233613
rect 259894 233549 259946 233555
rect 259126 231757 259178 231763
rect 259126 231699 259178 231705
rect 259030 227095 259082 227101
rect 259030 227037 259082 227043
rect 259414 226725 259466 226731
rect 259414 226667 259466 226673
rect 259426 221792 259454 226667
rect 259426 221764 259502 221792
rect 259474 221482 259502 221764
rect 260194 221482 260222 234955
rect 260470 234347 260522 234353
rect 260470 234289 260522 234295
rect 260482 228507 260510 234289
rect 260674 233169 260702 239686
rect 261024 239672 261278 239700
rect 261408 239672 261662 239700
rect 261792 239672 261950 239700
rect 261250 234353 261278 239672
rect 261238 234347 261290 234353
rect 261238 234289 261290 234295
rect 260854 233829 260906 233835
rect 260854 233771 260906 233777
rect 260662 233163 260714 233169
rect 260662 233105 260714 233111
rect 260470 228501 260522 228507
rect 260470 228443 260522 228449
rect 260866 228359 260894 233771
rect 261634 233391 261662 239672
rect 261622 233385 261674 233391
rect 261622 233327 261674 233333
rect 261718 232275 261770 232281
rect 261718 232217 261770 232223
rect 260854 228353 260906 228359
rect 260854 228295 260906 228301
rect 261046 225985 261098 225991
rect 261046 225927 261098 225933
rect 261058 221482 261086 225927
rect 261730 221792 261758 232217
rect 261922 223771 261950 239672
rect 262006 235161 262058 235167
rect 262006 235103 262058 235109
rect 262018 225473 262046 235103
rect 262114 233243 262142 239686
rect 262498 234575 262526 239686
rect 262882 235759 262910 239686
rect 263328 239672 263582 239700
rect 263712 239672 263966 239700
rect 264096 239672 264350 239700
rect 262870 235753 262922 235759
rect 262870 235695 262922 235701
rect 262486 234569 262538 234575
rect 262486 234511 262538 234517
rect 262102 233237 262154 233243
rect 262102 233179 262154 233185
rect 263254 232127 263306 232133
rect 263254 232069 263306 232075
rect 262486 226651 262538 226657
rect 262486 226593 262538 226599
rect 262006 225467 262058 225473
rect 262006 225409 262058 225415
rect 261910 223765 261962 223771
rect 261910 223707 261962 223713
rect 261730 221764 261806 221792
rect 261778 221482 261806 221764
rect 262498 221482 262526 226593
rect 263266 221482 263294 232069
rect 263554 223845 263582 239672
rect 263734 236123 263786 236129
rect 263734 236065 263786 236071
rect 263746 227175 263774 236065
rect 263938 232947 263966 239672
rect 263926 232941 263978 232947
rect 263926 232883 263978 232889
rect 264322 229469 264350 239672
rect 264418 233465 264446 239686
rect 264610 239672 264816 239700
rect 264406 233459 264458 233465
rect 264406 233401 264458 233407
rect 264310 229463 264362 229469
rect 264310 229405 264362 229411
rect 263734 227169 263786 227175
rect 263734 227111 263786 227117
rect 264022 227021 264074 227027
rect 264022 226963 264074 226969
rect 263542 223839 263594 223845
rect 263542 223781 263594 223787
rect 264034 221496 264062 226963
rect 264610 223549 264638 239672
rect 264694 235901 264746 235907
rect 264694 235843 264746 235849
rect 264706 226657 264734 235843
rect 264886 234273 264938 234279
rect 264886 234215 264938 234221
rect 264790 229981 264842 229987
rect 264790 229923 264842 229929
rect 264694 226651 264746 226657
rect 264694 226593 264746 226599
rect 264598 223543 264650 223549
rect 264598 223485 264650 223491
rect 264034 221468 264096 221496
rect 264802 221482 264830 229923
rect 264898 228433 264926 234215
rect 265186 232799 265214 239686
rect 265536 239672 265790 239700
rect 265920 239672 266174 239700
rect 266304 239672 266558 239700
rect 265270 235087 265322 235093
rect 265270 235029 265322 235035
rect 265174 232793 265226 232799
rect 265174 232735 265226 232741
rect 264886 228427 264938 228433
rect 264886 228369 264938 228375
rect 265282 225547 265310 235029
rect 265762 233095 265790 239672
rect 266146 235167 266174 239672
rect 266134 235161 266186 235167
rect 266134 235103 266186 235109
rect 266326 234125 266378 234131
rect 266326 234067 266378 234073
rect 265750 233089 265802 233095
rect 265750 233031 265802 233037
rect 266338 228581 266366 234067
rect 266230 228575 266282 228581
rect 266230 228517 266282 228523
rect 266326 228575 266378 228581
rect 266326 228517 266378 228523
rect 265558 226503 265610 226509
rect 265558 226445 265610 226451
rect 265270 225541 265322 225547
rect 265270 225483 265322 225489
rect 265570 221496 265598 226445
rect 265536 221468 265598 221496
rect 266242 221496 266270 228517
rect 266530 223697 266558 239672
rect 266626 232725 266654 239686
rect 267106 234131 267134 239686
rect 267094 234125 267146 234131
rect 267094 234067 267146 234073
rect 267490 233835 267518 239686
rect 267840 239672 268094 239700
rect 268224 239672 268478 239700
rect 267958 235827 268010 235833
rect 267958 235769 268010 235775
rect 267478 233829 267530 233835
rect 267478 233771 267530 233777
rect 267766 233607 267818 233613
rect 267766 233549 267818 233555
rect 266614 232719 266666 232725
rect 266614 232661 266666 232667
rect 266998 226947 267050 226953
rect 266998 226889 267050 226895
rect 266518 223691 266570 223697
rect 266518 223633 266570 223639
rect 266242 221468 266304 221496
rect 267010 221482 267038 226889
rect 267778 225843 267806 233549
rect 267862 230351 267914 230357
rect 267862 230293 267914 230299
rect 267766 225837 267818 225843
rect 267766 225779 267818 225785
rect 267874 221792 267902 230293
rect 267970 224733 267998 235769
rect 267958 224727 268010 224733
rect 267958 224669 268010 224675
rect 268066 223623 268094 239672
rect 268450 232651 268478 239672
rect 268546 234279 268574 239686
rect 268930 235093 268958 239686
rect 269314 236174 269342 239686
rect 269314 236146 269534 236174
rect 268918 235087 268970 235093
rect 268918 235029 268970 235035
rect 269398 234495 269450 234501
rect 269398 234437 269450 234443
rect 268534 234273 268586 234279
rect 268534 234215 268586 234221
rect 269014 233385 269066 233391
rect 269014 233327 269066 233333
rect 268438 232645 268490 232651
rect 268438 232587 268490 232593
rect 268534 226577 268586 226583
rect 268534 226519 268586 226525
rect 268054 223617 268106 223623
rect 268054 223559 268106 223565
rect 267826 221764 267902 221792
rect 267826 221482 267854 221764
rect 268546 221482 268574 226519
rect 269026 225917 269054 233327
rect 269110 233311 269162 233317
rect 269110 233253 269162 233259
rect 269122 230357 269150 233253
rect 269110 230351 269162 230357
rect 269110 230293 269162 230299
rect 269410 228655 269438 234437
rect 269302 228649 269354 228655
rect 269302 228591 269354 228597
rect 269398 228649 269450 228655
rect 269398 228591 269450 228597
rect 269014 225911 269066 225917
rect 269014 225853 269066 225859
rect 269314 221482 269342 228591
rect 269506 223475 269534 236146
rect 269698 232503 269726 239686
rect 270048 239672 270302 239700
rect 270432 239672 270590 239700
rect 270864 239672 271166 239700
rect 270274 233317 270302 239672
rect 270562 233391 270590 239672
rect 270934 235975 270986 235981
rect 270934 235917 270986 235923
rect 270838 233903 270890 233909
rect 270838 233845 270890 233851
rect 270550 233385 270602 233391
rect 270550 233327 270602 233333
rect 270262 233311 270314 233317
rect 270262 233253 270314 233259
rect 269686 232497 269738 232503
rect 269686 232439 269738 232445
rect 270742 229315 270794 229321
rect 270742 229257 270794 229263
rect 269974 227095 270026 227101
rect 269974 227037 270026 227043
rect 269494 223469 269546 223475
rect 269494 223411 269546 223417
rect 269986 221792 270014 227037
rect 269986 221764 270062 221792
rect 270034 221482 270062 221764
rect 270754 221482 270782 229257
rect 270850 228211 270878 233845
rect 270838 228205 270890 228211
rect 270838 228147 270890 228153
rect 270946 226583 270974 235917
rect 270934 226577 270986 226583
rect 270934 226519 270986 226525
rect 271138 223401 271166 239672
rect 271234 232429 271262 239686
rect 271618 234501 271646 239686
rect 271606 234495 271658 234501
rect 271606 234437 271658 234443
rect 271894 233459 271946 233465
rect 271894 233401 271946 233407
rect 271222 232423 271274 232429
rect 271222 232365 271274 232371
rect 271906 226731 271934 233401
rect 272002 227249 272030 239686
rect 272352 239672 272606 239700
rect 272736 239672 272990 239700
rect 272278 229389 272330 229395
rect 272278 229331 272330 229337
rect 271990 227243 272042 227249
rect 271990 227185 272042 227191
rect 271894 226725 271946 226731
rect 271894 226667 271946 226673
rect 271606 226429 271658 226435
rect 271606 226371 271658 226377
rect 271126 223395 271178 223401
rect 271126 223337 271178 223343
rect 271618 221482 271646 226371
rect 272290 221792 272318 229331
rect 272578 223253 272606 239672
rect 272962 232355 272990 239672
rect 273058 236129 273086 239686
rect 273046 236123 273098 236129
rect 273046 236065 273098 236071
rect 272950 232349 273002 232355
rect 272950 232291 273002 232297
rect 273442 226953 273470 239686
rect 273840 239672 274142 239700
rect 273718 236049 273770 236055
rect 273718 235991 273770 235997
rect 273622 234643 273674 234649
rect 273622 234585 273674 234591
rect 273526 233311 273578 233317
rect 273526 233253 273578 233259
rect 273538 229395 273566 233253
rect 273526 229389 273578 229395
rect 273526 229331 273578 229337
rect 273430 226947 273482 226953
rect 273430 226889 273482 226895
rect 273634 225621 273662 234585
rect 273622 225615 273674 225621
rect 273622 225557 273674 225563
rect 273730 225473 273758 235991
rect 273814 229167 273866 229173
rect 273814 229109 273866 229115
rect 273046 225467 273098 225473
rect 273046 225409 273098 225415
rect 273718 225467 273770 225473
rect 273718 225409 273770 225415
rect 272566 223247 272618 223253
rect 272566 223189 272618 223195
rect 272290 221764 272366 221792
rect 272338 221482 272366 221764
rect 273058 221482 273086 225409
rect 273826 221482 273854 229109
rect 274114 222291 274142 239672
rect 274210 232281 274238 239686
rect 274656 239672 274910 239700
rect 275040 239672 275294 239700
rect 274678 233385 274730 233391
rect 274678 233327 274730 233333
rect 274198 232275 274250 232281
rect 274198 232217 274250 232223
rect 274486 232053 274538 232059
rect 274486 231995 274538 232001
rect 274102 222285 274154 222291
rect 274102 222227 274154 222233
rect 274498 221792 274526 231995
rect 274690 227323 274718 233327
rect 274882 232577 274910 239672
rect 274870 232571 274922 232577
rect 274870 232513 274922 232519
rect 274678 227317 274730 227323
rect 274678 227259 274730 227265
rect 275266 227101 275294 239672
rect 275362 237683 275390 239686
rect 275350 237677 275402 237683
rect 275350 237619 275402 237625
rect 275746 232133 275774 239686
rect 276130 235907 276158 239686
rect 276480 239672 276734 239700
rect 276864 239672 277118 239700
rect 277248 239672 277502 239700
rect 276118 235901 276170 235907
rect 276118 235843 276170 235849
rect 275734 232127 275786 232133
rect 275734 232069 275786 232075
rect 275350 231905 275402 231911
rect 275350 231847 275402 231853
rect 275254 227095 275306 227101
rect 275254 227037 275306 227043
rect 274498 221764 274574 221792
rect 274546 221482 274574 221764
rect 275362 221482 275390 231847
rect 276502 228279 276554 228285
rect 276502 228221 276554 228227
rect 276118 226651 276170 226657
rect 276118 226593 276170 226599
rect 276130 221482 276158 226593
rect 276514 224215 276542 228221
rect 276706 227027 276734 239672
rect 277090 237609 277118 239672
rect 277078 237603 277130 237609
rect 277078 237545 277130 237551
rect 277078 234421 277130 234427
rect 277078 234363 277130 234369
rect 276790 229241 276842 229247
rect 276790 229183 276842 229189
rect 276694 227021 276746 227027
rect 276694 226963 276746 226969
rect 276502 224209 276554 224215
rect 276502 224151 276554 224157
rect 276802 221792 276830 229183
rect 277090 225251 277118 234363
rect 277474 232207 277502 239672
rect 277570 235981 277598 239686
rect 277558 235975 277610 235981
rect 277558 235917 277610 235923
rect 277462 232201 277514 232207
rect 277462 232143 277514 232149
rect 277954 226879 277982 239686
rect 278434 236795 278462 239686
rect 278784 239672 279038 239700
rect 279168 239672 279326 239700
rect 279552 239672 279806 239700
rect 278422 236789 278474 236795
rect 278422 236731 278474 236737
rect 278230 233755 278282 233761
rect 278230 233697 278282 233703
rect 277942 226873 277994 226879
rect 277942 226815 277994 226821
rect 278242 225695 278270 233697
rect 279010 231985 279038 239672
rect 279298 235833 279326 239672
rect 279286 235827 279338 235833
rect 279286 235769 279338 235775
rect 279286 234199 279338 234205
rect 279286 234141 279338 234147
rect 278326 231979 278378 231985
rect 278326 231921 278378 231927
rect 278998 231979 279050 231985
rect 278998 231921 279050 231927
rect 278230 225689 278282 225695
rect 278230 225631 278282 225637
rect 277078 225245 277130 225251
rect 277078 225187 277130 225193
rect 277558 224209 277610 224215
rect 277558 224151 277610 224157
rect 276802 221764 276878 221792
rect 276850 221482 276878 221764
rect 277570 221482 277598 224151
rect 278338 221482 278366 231921
rect 279298 227619 279326 234141
rect 279286 227613 279338 227619
rect 279286 227555 279338 227561
rect 279778 226805 279806 239672
rect 279874 236869 279902 239686
rect 279862 236863 279914 236869
rect 279862 236805 279914 236811
rect 280258 232059 280286 239686
rect 280642 234649 280670 239686
rect 280992 239672 281246 239700
rect 281376 239672 281630 239700
rect 281760 239672 282014 239700
rect 280630 234643 280682 234649
rect 280630 234585 280682 234591
rect 280246 232053 280298 232059
rect 280246 231995 280298 232001
rect 281218 231319 281246 239672
rect 281302 231831 281354 231837
rect 281302 231773 281354 231779
rect 281206 231313 281258 231319
rect 281206 231255 281258 231261
rect 279862 229093 279914 229099
rect 279862 229035 279914 229041
rect 279766 226799 279818 226805
rect 279766 226741 279818 226747
rect 279094 225541 279146 225547
rect 279094 225483 279146 225489
rect 279106 221792 279134 225483
rect 279106 221764 279182 221792
rect 279154 221482 279182 221764
rect 279874 221482 279902 229035
rect 280630 228131 280682 228137
rect 280630 228073 280682 228079
rect 280642 221482 280670 228073
rect 281314 221792 281342 231773
rect 281602 222365 281630 239672
rect 281878 234051 281930 234057
rect 281878 233993 281930 233999
rect 281890 227989 281918 233993
rect 281986 231911 282014 239672
rect 281974 231905 282026 231911
rect 281974 231847 282026 231853
rect 282178 229247 282206 239686
rect 282166 229241 282218 229247
rect 282166 229183 282218 229189
rect 281878 227983 281930 227989
rect 281878 227925 281930 227931
rect 282562 224733 282590 239686
rect 282960 239672 283166 239700
rect 283296 239672 283550 239700
rect 283680 239672 283934 239700
rect 282934 235605 282986 235611
rect 282934 235547 282986 235553
rect 282070 224727 282122 224733
rect 282070 224669 282122 224675
rect 282550 224727 282602 224733
rect 282550 224669 282602 224675
rect 281590 222359 281642 222365
rect 281590 222301 281642 222307
rect 281314 221764 281390 221792
rect 281362 221482 281390 221764
rect 282082 221482 282110 224669
rect 282946 221482 282974 235547
rect 283138 222439 283166 239672
rect 283522 229321 283550 239672
rect 283906 234205 283934 239672
rect 284002 234427 284030 239686
rect 284400 239672 284702 239700
rect 283990 234421 284042 234427
rect 283990 234363 284042 234369
rect 283894 234199 283946 234205
rect 283894 234141 283946 234147
rect 284374 232867 284426 232873
rect 284374 232809 284426 232815
rect 283510 229315 283562 229321
rect 283510 229257 283562 229263
rect 283606 229019 283658 229025
rect 283606 228961 283658 228967
rect 283126 222433 283178 222439
rect 283126 222375 283178 222381
rect 283618 221792 283646 228961
rect 283618 221764 283694 221792
rect 283666 221482 283694 221764
rect 284386 221482 284414 232809
rect 284674 227397 284702 239672
rect 284770 229173 284798 239686
rect 285154 235685 285182 239686
rect 285504 239672 285758 239700
rect 285984 239672 286238 239700
rect 285142 235679 285194 235685
rect 285142 235621 285194 235627
rect 285046 233829 285098 233835
rect 285046 233771 285098 233777
rect 284758 229167 284810 229173
rect 284758 229109 284810 229115
rect 284662 227391 284714 227397
rect 284662 227333 284714 227339
rect 285058 225769 285086 233771
rect 285730 226657 285758 239672
rect 285910 235531 285962 235537
rect 285910 235473 285962 235479
rect 285718 226651 285770 226657
rect 285718 226593 285770 226599
rect 285142 226355 285194 226361
rect 285142 226297 285194 226303
rect 285046 225763 285098 225769
rect 285046 225705 285098 225711
rect 285154 221482 285182 226297
rect 285922 221792 285950 235473
rect 286210 223179 286238 239672
rect 286306 229099 286334 239686
rect 286690 235611 286718 239686
rect 287074 236055 287102 239686
rect 287062 236049 287114 236055
rect 287062 235991 287114 235997
rect 286678 235605 286730 235611
rect 286678 235547 286730 235553
rect 287350 235309 287402 235315
rect 287350 235251 287402 235257
rect 286294 229093 286346 229099
rect 286294 229035 286346 229041
rect 286678 228501 286730 228507
rect 286678 228443 286730 228449
rect 286198 223173 286250 223179
rect 286198 223115 286250 223121
rect 285922 221764 285998 221792
rect 285970 221482 285998 221764
rect 286690 221482 286718 228443
rect 287362 228156 287390 235251
rect 287458 233687 287486 239686
rect 287808 239672 287966 239700
rect 288192 239672 288446 239700
rect 287446 233681 287498 233687
rect 287446 233623 287498 233629
rect 287938 229025 287966 239672
rect 288022 234347 288074 234353
rect 288022 234289 288074 234295
rect 287926 229019 287978 229025
rect 287926 228961 287978 228967
rect 288034 228285 288062 234289
rect 288418 233613 288446 239672
rect 288406 233607 288458 233613
rect 288406 233549 288458 233555
rect 288022 228279 288074 228285
rect 288022 228221 288074 228227
rect 287362 228128 287486 228156
rect 287458 221482 287486 228128
rect 288118 227169 288170 227175
rect 288118 227111 288170 227117
rect 288130 221792 288158 227111
rect 288514 226509 288542 239686
rect 288898 235315 288926 239686
rect 288886 235309 288938 235315
rect 288886 235251 288938 235257
rect 289270 231313 289322 231319
rect 289270 231255 289322 231261
rect 288886 229833 288938 229839
rect 288886 229775 288938 229781
rect 288502 226503 288554 226509
rect 288502 226445 288554 226451
rect 288130 221764 288206 221792
rect 288178 221482 288206 221764
rect 288898 221482 288926 229775
rect 289282 227175 289310 231255
rect 289378 228507 289406 239686
rect 289728 239672 289982 239700
rect 290112 239672 290366 239700
rect 290496 239672 290750 239700
rect 289954 232873 289982 239672
rect 290338 235537 290366 239672
rect 290326 235531 290378 235537
rect 290326 235473 290378 235479
rect 290422 233533 290474 233539
rect 290422 233475 290474 233481
rect 289942 232867 289994 232873
rect 289942 232809 289994 232815
rect 289750 228723 289802 228729
rect 289750 228665 289802 228671
rect 289366 228501 289418 228507
rect 289366 228443 289418 228449
rect 289270 227169 289322 227175
rect 289270 227111 289322 227117
rect 289762 221482 289790 228665
rect 290434 221792 290462 233475
rect 290722 230875 290750 239672
rect 290818 233021 290846 239686
rect 290902 234569 290954 234575
rect 290902 234511 290954 234517
rect 290806 233015 290858 233021
rect 290806 232957 290858 232963
rect 290710 230869 290762 230875
rect 290710 230811 290762 230817
rect 290914 229987 290942 234511
rect 290998 234125 291050 234131
rect 290998 234067 291050 234073
rect 290902 229981 290954 229987
rect 290902 229923 290954 229929
rect 291010 228063 291038 234067
rect 291202 229839 291230 239686
rect 291190 229833 291242 229839
rect 291190 229775 291242 229781
rect 290998 228057 291050 228063
rect 290998 227999 291050 228005
rect 291586 226435 291614 239686
rect 291936 239672 292190 239700
rect 292320 239672 292574 239700
rect 292704 239672 292958 239700
rect 291958 229611 292010 229617
rect 291958 229553 292010 229559
rect 291574 226429 291626 226435
rect 291574 226371 291626 226377
rect 291190 226207 291242 226213
rect 291190 226149 291242 226155
rect 290434 221764 290510 221792
rect 290482 221482 290510 221764
rect 291202 221482 291230 226149
rect 291970 221482 291998 229553
rect 292162 228919 292190 239672
rect 292546 231467 292574 239672
rect 292930 233465 292958 239672
rect 292918 233459 292970 233465
rect 292918 233401 292970 233407
rect 292534 231461 292586 231467
rect 292534 231403 292586 231409
rect 293122 231393 293150 239686
rect 293398 235457 293450 235463
rect 293398 235399 293450 235405
rect 293110 231387 293162 231393
rect 293110 231329 293162 231335
rect 292148 228910 292204 228919
rect 292148 228845 292204 228854
rect 292630 228353 292682 228359
rect 292630 228295 292682 228301
rect 292642 221792 292670 228295
rect 293410 228156 293438 235399
rect 293506 231319 293534 239686
rect 293782 234273 293834 234279
rect 293782 234215 293834 234221
rect 293494 231313 293546 231319
rect 293494 231255 293546 231261
rect 293410 228128 293534 228156
rect 292642 221764 292718 221792
rect 292690 221482 292718 221764
rect 293506 221482 293534 228128
rect 293794 227841 293822 234215
rect 293890 228359 293918 239686
rect 294240 239672 294494 239700
rect 294624 239672 294878 239700
rect 295008 239672 295262 239700
rect 294466 233909 294494 239672
rect 294850 234131 294878 239672
rect 295234 235463 295262 239672
rect 295222 235457 295274 235463
rect 295222 235399 295274 235405
rect 294838 234125 294890 234131
rect 294838 234067 294890 234073
rect 294454 233903 294506 233909
rect 294454 233845 294506 233851
rect 295330 231837 295358 239686
rect 295714 234575 295742 239686
rect 295702 234569 295754 234575
rect 295702 234511 295754 234517
rect 296098 233983 296126 239686
rect 296448 239672 296606 239700
rect 296928 239672 297182 239700
rect 296578 234945 296606 239672
rect 296470 234939 296522 234945
rect 296470 234881 296522 234887
rect 296566 234939 296618 234945
rect 296566 234881 296618 234887
rect 296086 233977 296138 233983
rect 296086 233919 296138 233925
rect 295318 231831 295370 231837
rect 295318 231773 295370 231779
rect 294934 228797 294986 228803
rect 294934 228739 294986 228745
rect 293878 228353 293930 228359
rect 293878 228295 293930 228301
rect 293782 227835 293834 227841
rect 293782 227777 293834 227783
rect 294262 226577 294314 226583
rect 294262 226519 294314 226525
rect 294274 221496 294302 226519
rect 294240 221468 294302 221496
rect 294946 221496 294974 228739
rect 295702 228427 295754 228433
rect 295702 228369 295754 228375
rect 294946 221468 295008 221496
rect 295714 221482 295742 228369
rect 296482 221496 296510 234881
rect 297154 233539 297182 239672
rect 297250 233835 297278 239686
rect 297238 233829 297290 233835
rect 297238 233771 297290 233777
rect 297142 233533 297194 233539
rect 297142 233475 297194 233481
rect 297430 230869 297482 230875
rect 297430 230811 297482 230817
rect 297442 226583 297470 230811
rect 297430 226577 297482 226583
rect 297430 226519 297482 226525
rect 297634 226287 297662 239686
rect 298018 236174 298046 239686
rect 298018 236146 298142 236174
rect 298114 229617 298142 236146
rect 298102 229611 298154 229617
rect 298102 229553 298154 229559
rect 298402 229543 298430 239686
rect 298752 239672 299006 239700
rect 299136 239672 299390 239700
rect 298978 234691 299006 239672
rect 299362 234987 299390 239672
rect 299348 234978 299404 234987
rect 299348 234913 299404 234922
rect 299458 234839 299486 239686
rect 299444 234830 299500 234839
rect 299444 234765 299500 234774
rect 299350 234717 299402 234723
rect 298964 234682 299020 234691
rect 299350 234659 299402 234665
rect 298964 234617 299020 234626
rect 299362 230505 299390 234659
rect 299842 234057 299870 239686
rect 300226 236943 300254 239686
rect 300214 236937 300266 236943
rect 300214 236879 300266 236885
rect 299830 234051 299882 234057
rect 299830 233993 299882 233999
rect 299446 231017 299498 231023
rect 299446 230959 299498 230965
rect 299350 230499 299402 230505
rect 299350 230441 299402 230447
rect 298006 229537 298058 229543
rect 298006 229479 298058 229485
rect 298390 229537 298442 229543
rect 298390 229479 298442 229485
rect 297238 226281 297290 226287
rect 297238 226223 297290 226229
rect 297622 226281 297674 226287
rect 297622 226223 297674 226229
rect 296448 221468 296510 221496
rect 297250 221482 297278 226223
rect 298018 221482 298046 229479
rect 298678 228871 298730 228877
rect 298678 228813 298730 228819
rect 298690 221792 298718 228813
rect 298690 221764 298766 221792
rect 298738 221482 298766 221764
rect 299458 221482 299486 230959
rect 300706 226213 300734 239686
rect 301056 239672 301310 239700
rect 301440 239672 301694 239700
rect 301282 236174 301310 239672
rect 301282 236146 301406 236174
rect 301270 234495 301322 234501
rect 301270 234437 301322 234443
rect 300982 228945 301034 228951
rect 300982 228887 301034 228893
rect 300694 226207 300746 226213
rect 300694 226149 300746 226155
rect 300214 226133 300266 226139
rect 300214 226075 300266 226081
rect 300226 221482 300254 226075
rect 300994 221792 301022 228887
rect 301282 227767 301310 234437
rect 301270 227761 301322 227767
rect 301270 227703 301322 227709
rect 301378 226139 301406 236146
rect 301666 235135 301694 239672
rect 301652 235126 301708 235135
rect 301652 235061 301708 235070
rect 301762 234723 301790 239686
rect 301750 234717 301802 234723
rect 301750 234659 301802 234665
rect 301750 228575 301802 228581
rect 301750 228517 301802 228523
rect 301366 226133 301418 226139
rect 301366 226075 301418 226081
rect 300994 221764 301070 221792
rect 301042 221482 301070 221764
rect 301762 221482 301790 228517
rect 302146 225325 302174 239686
rect 302544 239672 302846 239700
rect 302326 235235 302378 235241
rect 302326 235177 302378 235183
rect 302338 230653 302366 235177
rect 302326 230647 302378 230653
rect 302326 230589 302378 230595
rect 302518 230499 302570 230505
rect 302518 230441 302570 230447
rect 302134 225319 302186 225325
rect 302134 225261 302186 225267
rect 302530 221482 302558 230441
rect 302818 222513 302846 239672
rect 302914 231139 302942 239686
rect 303264 239672 303518 239700
rect 303648 239672 303902 239700
rect 303984 239672 304286 239700
rect 302900 231130 302956 231139
rect 302900 231065 302956 231074
rect 303490 228433 303518 239672
rect 303478 228427 303530 228433
rect 303478 228369 303530 228375
rect 303190 225541 303242 225547
rect 303190 225483 303242 225489
rect 302806 222507 302858 222513
rect 302806 222449 302858 222455
rect 303202 221792 303230 225483
rect 303874 225399 303902 239672
rect 304150 234791 304202 234797
rect 304150 234733 304202 234739
rect 304162 230505 304190 234733
rect 304150 230499 304202 230505
rect 304150 230441 304202 230447
rect 303958 230277 304010 230283
rect 303958 230219 304010 230225
rect 303862 225393 303914 225399
rect 303862 225335 303914 225341
rect 303202 221764 303278 221792
rect 303250 221482 303278 221764
rect 303970 221482 303998 230219
rect 304258 222587 304286 239672
rect 304450 228581 304478 239686
rect 304834 233761 304862 239686
rect 305184 239672 305246 239700
rect 305568 239672 305822 239700
rect 305952 239672 306206 239700
rect 305110 236123 305162 236129
rect 305110 236065 305162 236071
rect 305014 235753 305066 235759
rect 305014 235695 305066 235701
rect 304822 233755 304874 233761
rect 304822 233697 304874 233703
rect 304822 230425 304874 230431
rect 304822 230367 304874 230373
rect 304438 228575 304490 228581
rect 304438 228517 304490 228523
rect 304246 222581 304298 222587
rect 304246 222523 304298 222529
rect 304834 221482 304862 230367
rect 305026 225177 305054 235695
rect 305122 230283 305150 236065
rect 305218 235241 305246 239672
rect 305794 237017 305822 239672
rect 305782 237011 305834 237017
rect 305782 236953 305834 236959
rect 305206 235235 305258 235241
rect 305206 235177 305258 235183
rect 305494 231535 305546 231541
rect 305494 231477 305546 231483
rect 305110 230277 305162 230283
rect 305110 230219 305162 230225
rect 305014 225171 305066 225177
rect 305014 225113 305066 225119
rect 305506 221792 305534 231477
rect 306178 228729 306206 239672
rect 306274 234501 306302 239686
rect 306262 234495 306314 234501
rect 306262 234437 306314 234443
rect 306166 228723 306218 228729
rect 306166 228665 306218 228671
rect 306658 227564 306686 239686
rect 307056 239672 307262 239700
rect 307392 239672 307646 239700
rect 307776 239672 308030 239700
rect 308256 239672 308510 239700
rect 306742 235383 306794 235389
rect 306742 235325 306794 235331
rect 306754 230579 306782 235325
rect 306742 230573 306794 230579
rect 306742 230515 306794 230521
rect 307030 230203 307082 230209
rect 307030 230145 307082 230151
rect 306262 227539 306314 227545
rect 306658 227536 306782 227564
rect 306262 227481 306314 227487
rect 305506 221764 305582 221792
rect 305554 221482 305582 221764
rect 306274 221482 306302 227481
rect 306646 227391 306698 227397
rect 306646 227333 306698 227339
rect 306658 226435 306686 227333
rect 306646 226429 306698 226435
rect 306646 226371 306698 226377
rect 306754 225473 306782 227536
rect 306742 225467 306794 225473
rect 306742 225409 306794 225415
rect 307042 221482 307070 230145
rect 307234 222661 307262 239672
rect 307618 231287 307646 239672
rect 307604 231278 307660 231287
rect 307604 231213 307660 231222
rect 307702 228649 307754 228655
rect 307702 228591 307754 228597
rect 307222 222655 307274 222661
rect 307222 222597 307274 222603
rect 307714 221792 307742 228591
rect 308002 222809 308030 239672
rect 308182 234865 308234 234871
rect 308182 234807 308234 234813
rect 308194 231023 308222 234807
rect 308482 234353 308510 239672
rect 308578 237165 308606 239686
rect 308566 237159 308618 237165
rect 308566 237101 308618 237107
rect 308470 234347 308522 234353
rect 308470 234289 308522 234295
rect 308182 231017 308234 231023
rect 308182 230959 308234 230965
rect 308566 230647 308618 230653
rect 308566 230589 308618 230595
rect 307990 222803 308042 222809
rect 307990 222745 308042 222751
rect 307714 221764 307790 221792
rect 307762 221482 307790 221764
rect 308578 221482 308606 230589
rect 308962 228803 308990 239686
rect 308950 228797 309002 228803
rect 308950 228739 309002 228745
rect 309346 228729 309374 239686
rect 309696 239672 309950 239700
rect 310080 239672 310334 239700
rect 310464 239672 310718 239700
rect 309334 228723 309386 228729
rect 309334 228665 309386 228671
rect 309334 225615 309386 225621
rect 309334 225557 309386 225563
rect 309346 221482 309374 225557
rect 309922 225547 309950 239672
rect 310102 235901 310154 235907
rect 310102 235843 310154 235849
rect 310114 227915 310142 235843
rect 310006 227909 310058 227915
rect 310006 227851 310058 227857
rect 310102 227909 310154 227915
rect 310102 227851 310154 227857
rect 309910 225541 309962 225547
rect 309910 225483 309962 225489
rect 310018 221792 310046 227851
rect 310306 222883 310334 239672
rect 310690 228327 310718 239672
rect 310786 237091 310814 239686
rect 310774 237085 310826 237091
rect 310774 237027 310826 237033
rect 311062 233459 311114 233465
rect 311062 233401 311114 233407
rect 310774 230129 310826 230135
rect 310774 230071 310826 230077
rect 310676 228318 310732 228327
rect 310676 228253 310732 228262
rect 310294 222877 310346 222883
rect 310294 222819 310346 222825
rect 310018 221764 310094 221792
rect 310066 221482 310094 221764
rect 310786 221482 310814 230071
rect 311074 228137 311102 233401
rect 311170 233391 311198 239686
rect 311554 237239 311582 239686
rect 312000 239672 312254 239700
rect 312384 239672 312638 239700
rect 311542 237233 311594 237239
rect 311542 237175 311594 237181
rect 311350 234421 311402 234427
rect 311350 234363 311402 234369
rect 311254 233681 311306 233687
rect 311254 233623 311306 233629
rect 311158 233385 311210 233391
rect 311158 233327 311210 233333
rect 311062 228131 311114 228137
rect 311062 228073 311114 228079
rect 311266 227397 311294 233623
rect 311362 227545 311390 234363
rect 312226 231541 312254 239672
rect 312214 231535 312266 231541
rect 312214 231477 312266 231483
rect 311638 230499 311690 230505
rect 311638 230441 311690 230447
rect 311350 227539 311402 227545
rect 311350 227481 311402 227487
rect 311254 227391 311306 227397
rect 311254 227333 311306 227339
rect 311650 221482 311678 230441
rect 312310 225097 312362 225103
rect 312310 225039 312362 225045
rect 312322 221792 312350 225039
rect 312610 222735 312638 239672
rect 312706 234279 312734 239686
rect 313104 239672 313406 239700
rect 312694 234273 312746 234279
rect 312694 234215 312746 234221
rect 313078 230055 313130 230061
rect 313078 229997 313130 230003
rect 312598 222729 312650 222735
rect 312598 222671 312650 222677
rect 312322 221764 312398 221792
rect 312370 221482 312398 221764
rect 313090 221482 313118 229997
rect 313378 222957 313406 239672
rect 313474 228475 313502 239686
rect 313858 235907 313886 239686
rect 314208 239672 314462 239700
rect 314592 239672 314846 239700
rect 313942 235975 313994 235981
rect 313942 235917 313994 235923
rect 313846 235901 313898 235907
rect 313846 235843 313898 235849
rect 313846 233607 313898 233613
rect 313846 233549 313898 233555
rect 313460 228466 313516 228475
rect 313460 228401 313516 228410
rect 313858 228304 313886 233549
rect 313954 230875 313982 235917
rect 314434 234427 314462 239672
rect 314818 237313 314846 239672
rect 314806 237307 314858 237313
rect 314806 237249 314858 237255
rect 314422 234421 314474 234427
rect 314422 234363 314474 234369
rect 314518 231091 314570 231097
rect 314518 231033 314570 231039
rect 313942 230869 313994 230875
rect 313942 230811 313994 230817
rect 313858 228276 314078 228304
rect 313846 228205 313898 228211
rect 313846 228147 313898 228153
rect 313366 222951 313418 222957
rect 313366 222893 313418 222899
rect 313858 221482 313886 228147
rect 314050 228137 314078 228276
rect 314038 228131 314090 228137
rect 314038 228073 314090 228079
rect 314530 221792 314558 231033
rect 314914 228877 314942 239686
rect 315298 234797 315326 239686
rect 315286 234791 315338 234797
rect 315286 234733 315338 234739
rect 314902 228871 314954 228877
rect 314902 228813 314954 228819
rect 315382 227465 315434 227471
rect 315382 227407 315434 227413
rect 314530 221764 314606 221792
rect 314578 221482 314606 221764
rect 315394 221482 315422 227407
rect 315778 225621 315806 239686
rect 316176 239672 316382 239700
rect 316512 239672 316766 239700
rect 316896 239672 317150 239700
rect 316150 229907 316202 229913
rect 316150 229849 316202 229855
rect 315766 225615 315818 225621
rect 315766 225557 315818 225563
rect 316162 221482 316190 229849
rect 316354 223105 316382 239672
rect 316738 231435 316766 239672
rect 317122 237387 317150 239672
rect 317110 237381 317162 237387
rect 317110 237323 317162 237329
rect 317218 233465 317246 239686
rect 317602 237461 317630 239686
rect 317590 237455 317642 237461
rect 317590 237397 317642 237403
rect 317206 233459 317258 233465
rect 317206 233401 317258 233407
rect 316724 231426 316780 231435
rect 316724 231361 316780 231370
rect 317590 230573 317642 230579
rect 317590 230515 317642 230521
rect 316822 229759 316874 229765
rect 316822 229701 316874 229707
rect 316342 223099 316394 223105
rect 316342 223041 316394 223047
rect 316834 221792 316862 229701
rect 316834 221764 316910 221792
rect 316882 221482 316910 221764
rect 317602 221482 317630 230515
rect 317986 228951 318014 239686
rect 318384 239672 318590 239700
rect 318720 239672 318974 239700
rect 319200 239672 319454 239700
rect 318262 236049 318314 236055
rect 318262 235991 318314 235997
rect 317974 228945 318026 228951
rect 317974 228887 318026 228893
rect 318274 227471 318302 235991
rect 318358 235827 318410 235833
rect 318358 235769 318410 235775
rect 318370 230505 318398 235769
rect 318358 230499 318410 230505
rect 318358 230441 318410 230447
rect 318262 227465 318314 227471
rect 318262 227407 318314 227413
rect 318358 225245 318410 225251
rect 318358 225187 318410 225193
rect 318370 221482 318398 225187
rect 318562 223031 318590 239672
rect 318946 225515 318974 239672
rect 319126 229685 319178 229691
rect 319126 229627 319178 229633
rect 318932 225506 318988 225515
rect 318932 225441 318988 225450
rect 318550 223025 318602 223031
rect 318550 222967 318602 222973
rect 319138 221792 319166 229627
rect 319426 224585 319454 239672
rect 319522 231583 319550 239686
rect 319906 235981 319934 239686
rect 319894 235975 319946 235981
rect 319894 235917 319946 235923
rect 319606 233533 319658 233539
rect 319606 233475 319658 233481
rect 319508 231574 319564 231583
rect 319508 231509 319564 231518
rect 319618 227693 319646 233475
rect 320290 233317 320318 239686
rect 320640 239672 320894 239700
rect 321024 239672 321278 239700
rect 321408 239672 321662 239700
rect 320866 237535 320894 239672
rect 320854 237529 320906 237535
rect 320854 237471 320906 237477
rect 321046 234643 321098 234649
rect 321046 234585 321098 234591
rect 320758 234199 320810 234205
rect 320758 234141 320810 234147
rect 320278 233311 320330 233317
rect 320278 233253 320330 233259
rect 320662 231609 320714 231615
rect 320662 231551 320714 231557
rect 319606 227687 319658 227693
rect 319606 227629 319658 227635
rect 319894 227613 319946 227619
rect 319894 227555 319946 227561
rect 319414 224579 319466 224585
rect 319414 224521 319466 224527
rect 319138 221764 319214 221792
rect 319186 221482 319214 221764
rect 319906 221482 319934 227555
rect 320674 221482 320702 231551
rect 320770 230727 320798 234141
rect 320758 230721 320810 230727
rect 320758 230663 320810 230669
rect 321058 230579 321086 234585
rect 321046 230573 321098 230579
rect 321046 230515 321098 230521
rect 321250 230431 321278 239672
rect 321634 234871 321662 239672
rect 321622 234865 321674 234871
rect 321622 234807 321674 234813
rect 321238 230425 321290 230431
rect 321238 230367 321290 230373
rect 321334 225985 321386 225991
rect 321334 225927 321386 225933
rect 321346 221792 321374 225927
rect 321730 225663 321758 239686
rect 322128 239672 322334 239700
rect 322102 231165 322154 231171
rect 322102 231107 322154 231113
rect 321716 225654 321772 225663
rect 321716 225589 321772 225598
rect 321346 221764 321422 221792
rect 321394 221482 321422 221764
rect 322114 221482 322142 231107
rect 322306 224511 322334 239672
rect 322498 231731 322526 239686
rect 322944 239672 323198 239700
rect 323328 239672 323582 239700
rect 323712 239672 323966 239700
rect 322484 231722 322540 231731
rect 322484 231657 322540 231666
rect 322966 230351 323018 230357
rect 322966 230293 323018 230299
rect 322294 224505 322346 224511
rect 322294 224447 322346 224453
rect 322978 221496 323006 230293
rect 323170 224659 323198 239672
rect 323350 235679 323402 235685
rect 323350 235621 323402 235627
rect 323254 235013 323306 235019
rect 323254 234955 323306 234961
rect 323266 230653 323294 234955
rect 323362 230801 323390 235621
rect 323554 234649 323582 239672
rect 323938 238941 323966 239672
rect 323926 238935 323978 238941
rect 323926 238877 323978 238883
rect 323542 234643 323594 234649
rect 323542 234585 323594 234591
rect 323638 231017 323690 231023
rect 323638 230959 323690 230965
rect 323350 230795 323402 230801
rect 323350 230737 323402 230743
rect 323254 230647 323306 230653
rect 323254 230589 323306 230595
rect 323158 224653 323210 224659
rect 323158 224595 323210 224601
rect 322944 221468 323006 221496
rect 323650 221496 323678 230959
rect 324034 230209 324062 239686
rect 324418 239015 324446 239686
rect 324406 239009 324458 239015
rect 324406 238951 324458 238957
rect 324502 235161 324554 235167
rect 324502 235103 324554 235109
rect 324022 230203 324074 230209
rect 324022 230145 324074 230151
rect 324514 226065 324542 235103
rect 324802 233687 324830 239686
rect 325138 239404 325166 239686
rect 325536 239672 325790 239700
rect 325920 239672 326174 239700
rect 325090 239376 325166 239404
rect 324790 233681 324842 233687
rect 324790 233623 324842 233629
rect 324502 226059 324554 226065
rect 324502 226001 324554 226007
rect 324406 225689 324458 225695
rect 324406 225631 324458 225637
rect 323650 221468 323712 221496
rect 324418 221482 324446 225631
rect 325090 224437 325118 239376
rect 325174 231239 325226 231245
rect 325174 231181 325226 231187
rect 325078 224431 325130 224437
rect 325078 224373 325130 224379
rect 325186 221496 325214 231181
rect 325762 230357 325790 239672
rect 326146 235833 326174 239672
rect 326134 235827 326186 235833
rect 326134 235769 326186 235775
rect 326242 235685 326270 239686
rect 326722 238867 326750 239686
rect 326710 238861 326762 238867
rect 326710 238803 326762 238809
rect 326230 235679 326282 235685
rect 326230 235621 326282 235627
rect 326806 235605 326858 235611
rect 326806 235547 326858 235553
rect 326710 231683 326762 231689
rect 326710 231625 326762 231631
rect 325750 230351 325802 230357
rect 325750 230293 325802 230299
rect 325846 227983 325898 227989
rect 325846 227925 325898 227931
rect 325152 221468 325214 221496
rect 325858 221496 325886 227925
rect 325858 221468 325920 221496
rect 326722 221482 326750 231625
rect 326818 230949 326846 235547
rect 327106 231615 327134 239686
rect 327456 239672 327710 239700
rect 327840 239672 328094 239700
rect 327682 235167 327710 239672
rect 327670 235161 327722 235167
rect 327670 235103 327722 235109
rect 327094 231609 327146 231615
rect 327094 231551 327146 231557
rect 326806 230943 326858 230949
rect 326806 230885 326858 230891
rect 326806 230277 326858 230283
rect 326806 230219 326858 230225
rect 326818 227693 326846 230219
rect 326806 227687 326858 227693
rect 326806 227629 326858 227635
rect 327382 225837 327434 225843
rect 328066 225811 328094 239672
rect 328162 236174 328190 239686
rect 328162 236146 328286 236174
rect 328150 231757 328202 231763
rect 328150 231699 328202 231705
rect 327382 225779 327434 225785
rect 328052 225802 328108 225811
rect 327394 221792 327422 225779
rect 328052 225737 328108 225746
rect 327394 221764 327470 221792
rect 327442 221482 327470 221764
rect 328162 221482 328190 231699
rect 328258 224363 328286 236146
rect 328342 233829 328394 233835
rect 328342 233771 328394 233777
rect 328354 231097 328382 233771
rect 328342 231091 328394 231097
rect 328342 231033 328394 231039
rect 328546 230209 328574 239686
rect 328930 238793 328958 239686
rect 328918 238787 328970 238793
rect 328918 238729 328970 238735
rect 329314 233613 329342 239686
rect 329664 239672 329918 239700
rect 330048 239672 330302 239700
rect 329890 238719 329918 239672
rect 329878 238713 329930 238719
rect 329878 238655 329930 238661
rect 329302 233607 329354 233613
rect 329302 233549 329354 233555
rect 330274 233211 330302 239672
rect 330466 234205 330494 239686
rect 330454 234199 330506 234205
rect 330454 234141 330506 234147
rect 330260 233202 330316 233211
rect 330260 233137 330316 233146
rect 329590 230647 329642 230653
rect 329590 230589 329642 230595
rect 328534 230203 328586 230209
rect 328534 230145 328586 230151
rect 328918 228279 328970 228285
rect 328918 228221 328970 228227
rect 328246 224357 328298 224363
rect 328246 224299 328298 224305
rect 328930 221482 328958 228221
rect 329602 221792 329630 230589
rect 330850 227439 330878 239686
rect 331248 239672 331550 239700
rect 331414 235087 331466 235093
rect 331414 235029 331466 235035
rect 331222 233903 331274 233909
rect 331222 233845 331274 233851
rect 331234 231171 331262 233845
rect 331318 233163 331370 233169
rect 331318 233105 331370 233111
rect 331222 231165 331274 231171
rect 331222 231107 331274 231113
rect 330836 227430 330892 227439
rect 330836 227365 330892 227374
rect 331330 226972 331358 233105
rect 331234 226944 331358 226972
rect 330454 225911 330506 225917
rect 330454 225853 330506 225859
rect 329602 221764 329678 221792
rect 329650 221482 329678 221764
rect 330466 221482 330494 225853
rect 331234 221482 331262 226944
rect 331426 225917 331454 235029
rect 331414 225911 331466 225917
rect 331414 225853 331466 225859
rect 331522 224289 331550 239672
rect 331618 230135 331646 239686
rect 331968 239672 332222 239700
rect 332352 239672 332606 239700
rect 332194 233835 332222 239672
rect 332578 235611 332606 239672
rect 332674 238645 332702 239686
rect 332662 238639 332714 238645
rect 332662 238581 332714 238587
rect 332566 235605 332618 235611
rect 332566 235547 332618 235553
rect 332182 233829 332234 233835
rect 332182 233771 332234 233777
rect 331606 230129 331658 230135
rect 331606 230071 331658 230077
rect 331894 229981 331946 229987
rect 331894 229923 331946 229929
rect 331510 224283 331562 224289
rect 331510 224225 331562 224231
rect 331906 221792 331934 229923
rect 333058 228623 333086 239686
rect 333442 235019 333470 239686
rect 333430 235013 333482 235019
rect 333430 234955 333482 234961
rect 333044 228614 333100 228623
rect 333044 228549 333100 228558
rect 333826 227291 333854 239686
rect 334272 239672 334526 239700
rect 334656 239672 334910 239700
rect 334294 235531 334346 235537
rect 334294 235473 334346 235479
rect 334102 233755 334154 233761
rect 334102 233697 334154 233703
rect 334114 231245 334142 233697
rect 334198 233237 334250 233243
rect 334198 233179 334250 233185
rect 334102 231239 334154 231245
rect 334102 231181 334154 231187
rect 333812 227282 333868 227291
rect 333812 227217 333868 227226
rect 333526 225171 333578 225177
rect 333526 225113 333578 225119
rect 332662 223765 332714 223771
rect 332662 223707 332714 223713
rect 331906 221764 331982 221792
rect 331954 221482 331982 221764
rect 332674 221482 332702 223707
rect 333538 221482 333566 225113
rect 334210 221792 334238 233179
rect 334306 225991 334334 235473
rect 334294 225985 334346 225991
rect 334294 225927 334346 225933
rect 334498 224141 334526 239672
rect 334882 233063 334910 239672
rect 334978 235093 335006 239686
rect 334966 235087 335018 235093
rect 334966 235029 335018 235035
rect 335362 233539 335390 239686
rect 335746 238571 335774 239686
rect 336096 239672 336350 239700
rect 336480 239672 336734 239700
rect 335734 238565 335786 238571
rect 335734 238507 335786 238513
rect 335350 233533 335402 233539
rect 335350 233475 335402 233481
rect 334868 233054 334924 233063
rect 334868 232989 334924 232998
rect 336322 230061 336350 239672
rect 336706 238497 336734 239672
rect 336850 239404 336878 239686
rect 336850 239376 336926 239404
rect 336694 238491 336746 238497
rect 336694 238433 336746 238439
rect 336310 230055 336362 230061
rect 336310 229997 336362 230003
rect 334966 229463 335018 229469
rect 334966 229405 335018 229411
rect 334486 224135 334538 224141
rect 334486 224077 334538 224083
rect 334210 221764 334286 221792
rect 334258 221482 334286 221764
rect 334978 221482 335006 229405
rect 336898 227143 336926 239376
rect 336884 227134 336940 227143
rect 336884 227069 336940 227078
rect 336406 226725 336458 226731
rect 336406 226667 336458 226673
rect 335734 223839 335786 223845
rect 335734 223781 335786 223787
rect 335746 221482 335774 223781
rect 336418 221792 336446 226667
rect 337186 224067 337214 239686
rect 337270 232941 337322 232947
rect 337270 232883 337322 232889
rect 337174 224061 337226 224067
rect 337174 224003 337226 224009
rect 336418 221764 336494 221792
rect 336466 221482 336494 221764
rect 337282 221482 337310 232883
rect 337570 231689 337598 239686
rect 338050 236174 338078 239686
rect 338400 239672 338654 239700
rect 338784 239672 339038 239700
rect 339168 239672 339422 239700
rect 338050 236146 338174 236174
rect 338038 233089 338090 233095
rect 338038 233031 338090 233037
rect 337558 231683 337610 231689
rect 337558 231625 337610 231631
rect 338050 221482 338078 233031
rect 338146 224215 338174 236146
rect 338626 233761 338654 239672
rect 339010 238423 339038 239672
rect 338998 238417 339050 238423
rect 338998 238359 339050 238365
rect 339094 234125 339146 234131
rect 339094 234067 339146 234073
rect 338614 233755 338666 233761
rect 338614 233697 338666 233703
rect 339106 225695 339134 234067
rect 339394 228771 339422 239672
rect 339490 235389 339518 239686
rect 339478 235383 339530 235389
rect 339478 235325 339530 235331
rect 339766 233977 339818 233983
rect 339766 233919 339818 233925
rect 339380 228762 339436 228771
rect 339380 228697 339436 228706
rect 339478 226059 339530 226065
rect 339478 226001 339530 226007
rect 339094 225689 339146 225695
rect 339094 225631 339146 225637
rect 338134 224209 338186 224215
rect 338134 224151 338186 224157
rect 338710 223543 338762 223549
rect 338710 223485 338762 223491
rect 338722 221792 338750 223485
rect 338722 221764 338798 221792
rect 338770 221482 338798 221764
rect 339490 221482 339518 226001
rect 339778 225251 339806 233919
rect 339874 233909 339902 239686
rect 340272 239672 340478 239700
rect 340608 239672 340862 239700
rect 340992 239672 341246 239700
rect 341376 239672 341630 239700
rect 339862 233903 339914 233909
rect 339862 233845 339914 233851
rect 340246 232793 340298 232799
rect 340246 232735 340298 232741
rect 339766 225245 339818 225251
rect 339766 225187 339818 225193
rect 340258 221482 340286 232735
rect 340450 223993 340478 239672
rect 340834 233243 340862 239672
rect 341218 233983 341246 239672
rect 341398 234569 341450 234575
rect 341602 234543 341630 239672
rect 341794 238349 341822 239686
rect 341782 238343 341834 238349
rect 341782 238285 341834 238291
rect 341398 234511 341450 234517
rect 341588 234534 341644 234543
rect 341206 233977 341258 233983
rect 341206 233919 341258 233925
rect 340822 233237 340874 233243
rect 340822 233179 340874 233185
rect 341014 228057 341066 228063
rect 341014 227999 341066 228005
rect 340438 223987 340490 223993
rect 340438 223929 340490 223935
rect 341026 221792 341054 227999
rect 341410 227989 341438 234511
rect 341588 234469 341644 234478
rect 342178 230399 342206 239686
rect 342562 236023 342590 239686
rect 342912 239672 343070 239700
rect 343296 239672 343550 239700
rect 342548 236014 342604 236023
rect 342548 235949 342604 235958
rect 342646 233681 342698 233687
rect 342646 233623 342698 233629
rect 342164 230390 342220 230399
rect 342164 230325 342220 230334
rect 341398 227983 341450 227989
rect 341398 227925 341450 227931
rect 342550 225763 342602 225769
rect 342550 225705 342602 225711
rect 341782 223691 341834 223697
rect 341782 223633 341834 223639
rect 341026 221764 341102 221792
rect 341074 221482 341102 221764
rect 341794 221482 341822 223633
rect 342562 221482 342590 225705
rect 342658 225367 342686 233623
rect 343042 226995 343070 239672
rect 343522 233687 343550 239672
rect 343510 233681 343562 233687
rect 343510 233623 343562 233629
rect 343222 232719 343274 232725
rect 343222 232661 343274 232667
rect 343028 226986 343084 226995
rect 343028 226921 343084 226930
rect 342644 225358 342700 225367
rect 342644 225293 342700 225302
rect 343234 221792 343262 232661
rect 343618 223919 343646 239686
rect 343894 232571 343946 232577
rect 343894 232513 343946 232519
rect 343906 232355 343934 232513
rect 344002 232355 344030 239686
rect 344386 235135 344414 239686
rect 344180 235126 344236 235135
rect 344180 235061 344236 235070
rect 344372 235126 344428 235135
rect 344372 235061 344428 235070
rect 343894 232349 343946 232355
rect 343894 232291 343946 232297
rect 343990 232349 344042 232355
rect 343990 232291 344042 232297
rect 344194 228063 344222 235061
rect 344662 234051 344714 234057
rect 344662 233993 344714 233999
rect 344674 231023 344702 233993
rect 344662 231017 344714 231023
rect 344662 230959 344714 230965
rect 344182 228057 344234 228063
rect 344182 227999 344234 228005
rect 343990 227835 344042 227841
rect 343990 227777 344042 227783
rect 343606 223913 343658 223919
rect 343606 223855 343658 223861
rect 343234 221764 343310 221792
rect 343282 221482 343310 221764
rect 344002 221482 344030 227777
rect 344770 226847 344798 239686
rect 345120 239672 345374 239700
rect 345346 238275 345374 239672
rect 345538 239672 345600 239700
rect 345334 238269 345386 238275
rect 345334 238211 345386 238217
rect 345538 230251 345566 239672
rect 345718 235309 345770 235315
rect 345718 235251 345770 235257
rect 345524 230242 345580 230251
rect 345524 230177 345580 230186
rect 344756 226838 344812 226847
rect 344756 226773 344812 226782
rect 345730 225991 345758 235251
rect 345922 234575 345950 239686
rect 346320 239672 346622 239700
rect 345910 234569 345962 234575
rect 345910 234511 345962 234517
rect 346294 232793 346346 232799
rect 346294 232735 346346 232741
rect 345718 225985 345770 225991
rect 345718 225927 345770 225933
rect 345526 225911 345578 225917
rect 345526 225853 345578 225859
rect 344854 223617 344906 223623
rect 344854 223559 344906 223565
rect 344866 221482 344894 223559
rect 345538 221792 345566 225853
rect 345538 221764 345614 221792
rect 345586 221482 345614 221764
rect 346306 221482 346334 232735
rect 346594 223845 346622 239672
rect 346690 238201 346718 239686
rect 346678 238195 346730 238201
rect 346678 238137 346730 238143
rect 347074 233169 347102 239686
rect 347424 239672 347678 239700
rect 347808 239672 348062 239700
rect 347650 233803 347678 239672
rect 347636 233794 347692 233803
rect 347636 233729 347692 233738
rect 347062 233163 347114 233169
rect 347062 233105 347114 233111
rect 346966 232719 347018 232725
rect 346966 232661 347018 232667
rect 346978 232133 347006 232661
rect 346966 232127 347018 232133
rect 346966 232069 347018 232075
rect 346966 231757 347018 231763
rect 346966 231699 347018 231705
rect 346978 230875 347006 231699
rect 346966 230869 347018 230875
rect 346966 230811 347018 230817
rect 347062 229389 347114 229395
rect 347062 229331 347114 229337
rect 346582 223839 346634 223845
rect 346582 223781 346634 223787
rect 347074 221482 347102 229331
rect 348034 223771 348062 239672
rect 348022 223765 348074 223771
rect 348022 223707 348074 223713
rect 348130 223549 348158 239686
rect 348514 229987 348542 239686
rect 348898 235537 348926 239686
rect 349344 239672 349598 239700
rect 349728 239672 349982 239700
rect 350112 239672 350366 239700
rect 348886 235531 348938 235537
rect 348886 235473 348938 235479
rect 348694 235457 348746 235463
rect 348694 235399 348746 235405
rect 348502 229981 348554 229987
rect 348502 229923 348554 229929
rect 348598 227317 348650 227323
rect 348598 227259 348650 227265
rect 348118 223543 348170 223549
rect 348118 223485 348170 223491
rect 347734 223469 347786 223475
rect 347734 223411 347786 223417
rect 347746 221792 347774 223411
rect 347746 221764 347822 221792
rect 347794 221482 347822 221764
rect 348610 221482 348638 227259
rect 348706 224955 348734 235399
rect 349366 232497 349418 232503
rect 349366 232439 349418 232445
rect 348694 224949 348746 224955
rect 348694 224891 348746 224897
rect 349378 221482 349406 232439
rect 349570 223697 349598 239672
rect 349954 238127 349982 239672
rect 349942 238121 349994 238127
rect 349942 238063 349994 238069
rect 349748 234978 349804 234987
rect 349748 234913 349804 234922
rect 349762 225177 349790 234913
rect 350338 233095 350366 239672
rect 350326 233089 350378 233095
rect 350326 233031 350378 233037
rect 350518 232349 350570 232355
rect 350518 232291 350570 232297
rect 350530 232133 350558 232291
rect 350518 232127 350570 232133
rect 350518 232069 350570 232075
rect 350038 227761 350090 227767
rect 350038 227703 350090 227709
rect 349750 225171 349802 225177
rect 349750 225113 349802 225119
rect 349558 223691 349610 223697
rect 349558 223633 349610 223639
rect 350050 221792 350078 227703
rect 350818 223623 350846 239686
rect 350806 223617 350858 223623
rect 350806 223559 350858 223565
rect 351202 223475 351230 239686
rect 351552 239672 351806 239700
rect 351936 239672 352190 239700
rect 352320 239672 352574 239700
rect 351382 233903 351434 233909
rect 351382 233845 351434 233851
rect 351394 225959 351422 233845
rect 351778 229913 351806 239672
rect 352162 236129 352190 239672
rect 352150 236123 352202 236129
rect 352150 236065 352202 236071
rect 352342 232423 352394 232429
rect 352342 232365 352394 232371
rect 351766 229907 351818 229913
rect 351766 229849 351818 229855
rect 351574 227243 351626 227249
rect 351574 227185 351626 227191
rect 351380 225950 351436 225959
rect 351380 225885 351436 225894
rect 351190 223469 351242 223475
rect 351190 223411 351242 223417
rect 350806 223395 350858 223401
rect 350806 223337 350858 223343
rect 350050 221764 350126 221792
rect 350098 221482 350126 221764
rect 350818 221482 350846 223337
rect 351586 221482 351614 227185
rect 352354 221496 352382 232365
rect 352546 223401 352574 239672
rect 352738 237979 352766 239686
rect 352726 237973 352778 237979
rect 352726 237915 352778 237921
rect 353122 232947 353150 239686
rect 353506 238053 353534 239686
rect 353856 239672 354110 239700
rect 353494 238047 353546 238053
rect 353494 237989 353546 237995
rect 353110 232941 353162 232947
rect 353110 232883 353162 232889
rect 353110 227687 353162 227693
rect 353110 227629 353162 227635
rect 352534 223395 352586 223401
rect 352534 223337 352586 223343
rect 352354 221468 352416 221496
rect 353122 221482 353150 227629
rect 354082 223327 354110 239672
rect 354226 239404 354254 239686
rect 354624 239672 354878 239700
rect 354178 239376 354254 239404
rect 354178 224627 354206 239376
rect 354356 234830 354412 234839
rect 354356 234765 354412 234774
rect 354260 234682 354316 234691
rect 354260 234617 354316 234626
rect 354274 230653 354302 234617
rect 354262 230647 354314 230653
rect 354262 230589 354314 230595
rect 354370 225029 354398 234765
rect 354850 229765 354878 239672
rect 354946 235727 354974 239686
rect 355344 239672 355646 239700
rect 354932 235718 354988 235727
rect 354932 235653 354988 235662
rect 355318 232571 355370 232577
rect 355318 232513 355370 232519
rect 354838 229759 354890 229765
rect 354838 229701 354890 229707
rect 354550 226947 354602 226953
rect 354550 226889 354602 226895
rect 354358 225023 354410 225029
rect 354358 224965 354410 224971
rect 354164 224618 354220 224627
rect 354164 224553 354220 224562
rect 354070 223321 354122 223327
rect 354070 223263 354122 223269
rect 353878 223247 353930 223253
rect 353878 223189 353930 223195
rect 353890 221496 353918 223189
rect 353856 221468 353918 221496
rect 354562 221496 354590 226889
rect 354562 221468 354624 221496
rect 355330 221482 355358 232513
rect 355618 223253 355646 239672
rect 355714 237905 355742 239686
rect 356064 239672 356318 239700
rect 356544 239672 356798 239700
rect 355702 237899 355754 237905
rect 355702 237841 355754 237847
rect 356290 232799 356318 239672
rect 356770 234839 356798 239672
rect 356756 234830 356812 234839
rect 356756 234765 356812 234774
rect 356866 234691 356894 239686
rect 357264 239672 357566 239700
rect 356852 234682 356908 234691
rect 356852 234617 356908 234626
rect 356278 232793 356330 232799
rect 356278 232735 356330 232741
rect 356086 232645 356138 232651
rect 356086 232587 356138 232593
rect 355606 223247 355658 223253
rect 355606 223189 355658 223195
rect 356098 221792 356126 232587
rect 357538 224479 357566 239672
rect 357634 229395 357662 239686
rect 357718 237677 357770 237683
rect 357718 237619 357770 237625
rect 357622 229389 357674 229395
rect 357622 229331 357674 229337
rect 357730 228285 357758 237619
rect 358018 234131 358046 239686
rect 358368 239672 358622 239700
rect 358752 239672 359006 239700
rect 360022 239691 360074 239697
rect 358594 237831 358622 239672
rect 358582 237825 358634 237831
rect 358582 237767 358634 237773
rect 358390 234495 358442 234501
rect 358390 234437 358442 234443
rect 358006 234125 358058 234131
rect 358006 234067 358058 234073
rect 358294 232275 358346 232281
rect 358294 232217 358346 232223
rect 357718 228279 357770 228285
rect 357718 228221 357770 228227
rect 357622 227095 357674 227101
rect 357622 227037 357674 227043
rect 357524 224470 357580 224479
rect 357524 224405 357580 224414
rect 356854 222285 356906 222291
rect 356854 222227 356906 222233
rect 356098 221764 356174 221792
rect 356146 221482 356174 221764
rect 356866 221482 356894 222227
rect 357634 221482 357662 227037
rect 358306 221755 358334 232217
rect 358402 230875 358430 234437
rect 358390 230869 358442 230875
rect 358390 230811 358442 230817
rect 358978 229955 359006 239672
rect 359074 232915 359102 239686
rect 359060 232906 359116 232915
rect 359060 232841 359116 232850
rect 358964 229946 359020 229955
rect 358964 229881 359020 229890
rect 359158 227909 359210 227915
rect 359158 227851 359210 227857
rect 358306 221727 358382 221755
rect 358354 221482 358382 221727
rect 359170 221482 359198 227851
rect 359458 222999 359486 239686
rect 359842 236174 359870 239686
rect 359746 236146 359870 236174
rect 359746 224331 359774 236146
rect 360034 235907 360062 239691
rect 360022 235901 360074 235907
rect 360022 235843 360074 235849
rect 359828 228910 359884 228919
rect 359828 228845 359884 228854
rect 359842 226953 359870 228845
rect 359926 228279 359978 228285
rect 359926 228221 359978 228227
rect 359830 226947 359882 226953
rect 359830 226889 359882 226895
rect 359732 224322 359788 224331
rect 359732 224257 359788 224266
rect 359444 222990 359500 222999
rect 359444 222925 359500 222934
rect 359938 221482 359966 228221
rect 360322 224035 360350 239686
rect 360672 239672 360926 239700
rect 361056 239672 361310 239700
rect 360898 229691 360926 239672
rect 361282 233909 361310 239672
rect 361378 236174 361406 239686
rect 361762 237683 361790 239686
rect 361750 237677 361802 237683
rect 361750 237619 361802 237625
rect 361378 236146 361502 236174
rect 361270 233903 361322 233909
rect 361270 233845 361322 233851
rect 361366 232719 361418 232725
rect 361366 232661 361418 232667
rect 360886 229685 360938 229691
rect 360886 229627 360938 229633
rect 360598 227021 360650 227027
rect 360598 226963 360650 226969
rect 360308 224026 360364 224035
rect 360308 223961 360364 223970
rect 360610 221792 360638 226963
rect 360610 221764 360686 221792
rect 360658 221482 360686 221764
rect 361378 221482 361406 232661
rect 361474 224183 361502 236146
rect 361942 234939 361994 234945
rect 361942 234881 361994 234887
rect 361954 224807 361982 234881
rect 362146 232725 362174 239686
rect 362530 236055 362558 239686
rect 362880 239672 363134 239700
rect 363264 239672 363518 239700
rect 363106 237757 363134 239672
rect 363094 237751 363146 237757
rect 363094 237693 363146 237699
rect 362518 236049 362570 236055
rect 362518 235991 362570 235997
rect 362134 232719 362186 232725
rect 362134 232661 362186 232667
rect 362134 231757 362186 231763
rect 362134 231699 362186 231705
rect 361942 224801 361994 224807
rect 361942 224743 361994 224749
rect 361460 224174 361516 224183
rect 361460 224109 361516 224118
rect 362146 221482 362174 231699
rect 362806 229611 362858 229617
rect 362806 229553 362858 229559
rect 362818 224881 362846 229553
rect 362806 224875 362858 224881
rect 362806 224817 362858 224823
rect 363490 223887 363518 239672
rect 363586 230103 363614 239686
rect 363670 237603 363722 237609
rect 363670 237545 363722 237551
rect 363572 230094 363628 230103
rect 363572 230029 363628 230038
rect 363476 223878 363532 223887
rect 363476 223813 363532 223822
rect 363682 222273 363710 237545
rect 364066 235759 364094 239686
rect 364450 237609 364478 239686
rect 364800 239672 365054 239700
rect 365184 239672 365438 239700
rect 365568 239672 365726 239700
rect 364438 237603 364490 237609
rect 364438 237545 364490 237551
rect 364054 235753 364106 235759
rect 364054 235695 364106 235701
rect 365026 232577 365054 239672
rect 365410 232651 365438 239672
rect 365698 236174 365726 239672
rect 365698 236146 365822 236174
rect 365686 235235 365738 235241
rect 365686 235177 365738 235183
rect 365398 232645 365450 232651
rect 365398 232587 365450 232593
rect 365014 232571 365066 232577
rect 365014 232513 365066 232519
rect 364438 232201 364490 232207
rect 364438 232143 364490 232149
rect 364246 231313 364298 231319
rect 364246 231255 364298 231261
rect 364258 226879 364286 231255
rect 363766 226873 363818 226879
rect 363766 226815 363818 226821
rect 364246 226873 364298 226879
rect 364246 226815 364298 226821
rect 363010 222245 363710 222273
rect 363010 221792 363038 222245
rect 362962 221764 363038 221792
rect 362962 221482 362990 221764
rect 363778 221755 363806 226815
rect 363682 221727 363806 221755
rect 363682 221482 363710 221727
rect 364450 221482 364478 232143
rect 365110 230499 365162 230505
rect 365110 230441 365162 230447
rect 365122 221792 365150 230441
rect 365698 225917 365726 235177
rect 365794 229807 365822 236146
rect 365890 234057 365918 239686
rect 365878 234051 365930 234057
rect 365878 233993 365930 233999
rect 366274 232429 366302 239686
rect 366550 239675 366602 239681
rect 366550 239617 366602 239623
rect 366562 235981 366590 239617
rect 366550 235975 366602 235981
rect 366550 235917 366602 235923
rect 366262 232423 366314 232429
rect 366262 232365 366314 232371
rect 365780 229798 365836 229807
rect 365780 229733 365836 229742
rect 366658 229469 366686 239686
rect 367008 239672 367262 239700
rect 367392 239672 367646 239700
rect 367872 239672 368126 239700
rect 366742 236789 366794 236795
rect 366742 236731 366794 236737
rect 366646 229463 366698 229469
rect 366646 229405 366698 229411
rect 366754 228489 366782 236731
rect 367234 234247 367262 239672
rect 367220 234238 367276 234247
rect 367220 234173 367276 234182
rect 367126 232127 367178 232133
rect 367126 232069 367178 232075
rect 367138 231763 367166 232069
rect 367414 231979 367466 231985
rect 367414 231921 367466 231927
rect 367126 231757 367178 231763
rect 367126 231699 367178 231705
rect 365890 228461 366782 228489
rect 365686 225911 365738 225917
rect 365686 225853 365738 225859
rect 365122 221764 365198 221792
rect 365170 221482 365198 221764
rect 365890 221482 365918 228461
rect 366742 226799 366794 226805
rect 366742 226741 366794 226747
rect 366754 221482 366782 226741
rect 367426 221792 367454 231921
rect 367510 229315 367562 229321
rect 367510 229257 367562 229263
rect 367522 225103 367550 229257
rect 367510 225097 367562 225103
rect 367510 225039 367562 225045
rect 367618 223739 367646 239672
rect 368098 232207 368126 239672
rect 368194 232503 368222 239686
rect 368854 236863 368906 236869
rect 368854 236805 368906 236811
rect 368182 232497 368234 232503
rect 368182 232439 368234 232445
rect 368086 232201 368138 232207
rect 368086 232143 368138 232149
rect 368758 231091 368810 231097
rect 368758 231033 368810 231039
rect 368770 230727 368798 231033
rect 368566 230721 368618 230727
rect 368566 230663 368618 230669
rect 368758 230721 368810 230727
rect 368758 230663 368810 230669
rect 368182 230573 368234 230579
rect 368182 230515 368234 230521
rect 367604 223730 367660 223739
rect 367604 223665 367660 223674
rect 367426 221764 367502 221792
rect 367474 221482 367502 221764
rect 368194 221482 368222 230515
rect 368578 225843 368606 230663
rect 368866 227534 368894 236805
rect 368962 236319 368990 239686
rect 369312 239672 369566 239700
rect 369696 239672 369950 239700
rect 370080 239672 370334 239700
rect 368948 236310 369004 236319
rect 368948 236245 369004 236254
rect 369538 232133 369566 239672
rect 369526 232127 369578 232133
rect 369526 232069 369578 232075
rect 369922 229691 369950 239672
rect 370306 234099 370334 239672
rect 370402 236763 370430 239686
rect 370388 236754 370444 236763
rect 370388 236689 370444 236698
rect 370292 234090 370348 234099
rect 370292 234025 370348 234034
rect 370786 232767 370814 239686
rect 370772 232758 370828 232767
rect 370772 232693 370828 232702
rect 371170 232355 371198 239686
rect 371616 239672 371870 239700
rect 372000 239672 372254 239700
rect 371638 239453 371690 239459
rect 371638 239395 371690 239401
rect 371650 235907 371678 239395
rect 371842 235907 371870 239672
rect 372226 237059 372254 239672
rect 372212 237050 372268 237059
rect 372212 236985 372268 236994
rect 371638 235901 371690 235907
rect 371638 235843 371690 235849
rect 371830 235901 371882 235907
rect 371830 235843 371882 235849
rect 371158 232349 371210 232355
rect 371158 232291 371210 232297
rect 370390 232053 370442 232059
rect 370390 231995 370442 232001
rect 369910 229685 369962 229691
rect 369910 229627 369962 229633
rect 370402 227534 370430 231995
rect 372322 231985 372350 239686
rect 372706 232281 372734 239686
rect 372694 232275 372746 232281
rect 372694 232217 372746 232223
rect 372310 231979 372362 231985
rect 372310 231921 372362 231927
rect 371638 231387 371690 231393
rect 371638 231329 371690 231335
rect 371254 229241 371306 229247
rect 371254 229183 371306 229189
rect 368866 227506 368990 227534
rect 370402 227506 370526 227534
rect 368566 225837 368618 225843
rect 368566 225779 368618 225785
rect 368962 221482 368990 227506
rect 369622 227169 369674 227175
rect 369622 227111 369674 227117
rect 369634 221792 369662 227111
rect 369634 221764 369710 221792
rect 369682 221482 369710 221764
rect 370498 221482 370526 227506
rect 371266 221482 371294 229183
rect 371542 229167 371594 229173
rect 371542 229109 371594 229115
rect 371350 225763 371402 225769
rect 371350 225705 371402 225711
rect 371362 225103 371390 225705
rect 371350 225097 371402 225103
rect 371350 225039 371402 225045
rect 371446 225097 371498 225103
rect 371446 225039 371498 225045
rect 371458 224733 371486 225039
rect 371554 224733 371582 229109
rect 371650 226731 371678 231329
rect 373090 229659 373118 239686
rect 373474 236911 373502 239686
rect 373824 239672 374078 239700
rect 373460 236902 373516 236911
rect 373460 236837 373516 236846
rect 374050 231911 374078 239672
rect 374146 239672 374208 239700
rect 373462 231905 373514 231911
rect 373462 231847 373514 231853
rect 374038 231905 374090 231911
rect 374038 231847 374090 231853
rect 373076 229650 373132 229659
rect 373076 229585 373132 229594
rect 371638 226725 371690 226731
rect 371638 226667 371690 226673
rect 372694 225097 372746 225103
rect 372694 225039 372746 225045
rect 371446 224727 371498 224733
rect 371446 224669 371498 224675
rect 371542 224727 371594 224733
rect 371542 224669 371594 224675
rect 371926 222359 371978 222365
rect 371926 222301 371978 222307
rect 371938 221792 371966 222301
rect 371938 221764 372014 221792
rect 371986 221482 372014 221764
rect 372706 221482 372734 225039
rect 373474 221482 373502 231847
rect 374146 229321 374174 239672
rect 374530 235241 374558 239686
rect 374914 236615 374942 239686
rect 374900 236606 374956 236615
rect 374900 236541 374956 236550
rect 374518 235235 374570 235241
rect 374518 235177 374570 235183
rect 374710 234199 374762 234205
rect 374710 234141 374762 234147
rect 374614 233015 374666 233021
rect 374614 232957 374666 232963
rect 374134 229315 374186 229321
rect 374134 229257 374186 229263
rect 374518 229093 374570 229099
rect 374518 229035 374570 229041
rect 374422 229019 374474 229025
rect 374422 228961 374474 228967
rect 374434 225843 374462 228961
rect 374230 225837 374282 225843
rect 374230 225779 374282 225785
rect 374422 225837 374474 225843
rect 374422 225779 374474 225785
rect 374242 221774 374270 225779
rect 374530 225103 374558 229035
rect 374626 226805 374654 232957
rect 374614 226799 374666 226805
rect 374614 226741 374666 226747
rect 374518 225097 374570 225103
rect 374518 225039 374570 225045
rect 374722 222365 374750 234141
rect 375394 232619 375422 239686
rect 375380 232610 375436 232619
rect 375380 232545 375436 232554
rect 375778 232059 375806 239686
rect 376128 239672 376382 239700
rect 376512 239672 376766 239700
rect 376354 233951 376382 239672
rect 376738 236467 376766 239672
rect 376724 236458 376780 236467
rect 376724 236393 376780 236402
rect 376340 233942 376396 233951
rect 376340 233877 376396 233886
rect 375766 232053 375818 232059
rect 375766 231995 375818 232001
rect 376834 229173 376862 239686
rect 377110 230795 377162 230801
rect 377110 230737 377162 230743
rect 376822 229167 376874 229173
rect 376822 229109 376874 229115
rect 375766 227539 375818 227545
rect 377122 227534 377150 230737
rect 377218 229247 377246 239686
rect 377206 229241 377258 229247
rect 377206 229183 377258 229189
rect 377122 227506 377246 227534
rect 375766 227481 375818 227487
rect 374998 222433 375050 222439
rect 374998 222375 375050 222381
rect 374710 222359 374762 222365
rect 374710 222301 374762 222307
rect 374242 221746 374318 221774
rect 374290 221482 374318 221746
rect 375010 221482 375038 222375
rect 375778 221482 375806 227481
rect 376438 225763 376490 225769
rect 376438 225705 376490 225711
rect 376450 221792 376478 225705
rect 376450 221764 376526 221792
rect 376498 221482 376526 221764
rect 377218 221482 377246 227506
rect 377602 223591 377630 239686
rect 377782 236715 377834 236721
rect 377782 236657 377834 236663
rect 377794 236319 377822 236657
rect 377986 236319 378014 239686
rect 378336 239672 378590 239700
rect 378720 239672 378974 239700
rect 378454 239305 378506 239311
rect 378454 239247 378506 239253
rect 377780 236310 377836 236319
rect 377780 236245 377836 236254
rect 377972 236310 378028 236319
rect 377972 236245 378028 236254
rect 378466 233983 378494 239247
rect 378562 235852 378590 239672
rect 378562 235824 378878 235852
rect 378850 235759 378878 235824
rect 378838 235753 378890 235759
rect 378838 235695 378890 235701
rect 378550 234865 378602 234871
rect 378550 234807 378602 234813
rect 378562 234205 378590 234807
rect 378550 234199 378602 234205
rect 378550 234141 378602 234147
rect 378454 233977 378506 233983
rect 378454 233919 378506 233925
rect 378946 232471 378974 239672
rect 379138 234395 379166 239686
rect 379536 239672 379838 239700
rect 379124 234386 379180 234395
rect 379124 234321 379180 234330
rect 378932 232462 378988 232471
rect 378932 232397 378988 232406
rect 378562 229756 378782 229784
rect 378562 229691 378590 229756
rect 378550 229685 378602 229691
rect 378550 229627 378602 229633
rect 378646 229685 378698 229691
rect 378646 229627 378698 229633
rect 378658 229395 378686 229627
rect 378754 229395 378782 229756
rect 378646 229389 378698 229395
rect 378646 229331 378698 229337
rect 378742 229389 378794 229395
rect 378742 229331 378794 229337
rect 378742 226651 378794 226657
rect 378742 226593 378794 226599
rect 378070 226429 378122 226435
rect 378070 226371 378122 226377
rect 377588 223582 377644 223591
rect 377588 223517 377644 223526
rect 378082 221482 378110 226371
rect 378754 221792 378782 226593
rect 379510 224727 379562 224733
rect 379510 224669 379562 224675
rect 378754 221764 378830 221792
rect 378802 221482 378830 221764
rect 379522 221482 379550 224669
rect 379810 223295 379838 239672
rect 379906 229025 379934 239686
rect 380256 239672 380510 239700
rect 380640 239672 380894 239700
rect 381024 239672 381278 239700
rect 379990 231461 380042 231467
rect 379990 231403 380042 231409
rect 379894 229019 379946 229025
rect 379894 228961 379946 228967
rect 380002 226435 380030 231403
rect 380278 230943 380330 230949
rect 380278 230885 380330 230891
rect 380086 228501 380138 228507
rect 380086 228443 380138 228449
rect 379990 226429 380042 226435
rect 379990 226371 380042 226377
rect 380098 225769 380126 228443
rect 380086 225763 380138 225769
rect 380086 225705 380138 225711
rect 379796 223286 379852 223295
rect 379796 223221 379852 223230
rect 380290 221482 380318 230885
rect 380482 229099 380510 239672
rect 380866 239089 380894 239672
rect 380854 239083 380906 239089
rect 380854 239025 380906 239031
rect 380470 229093 380522 229099
rect 380470 229035 380522 229041
rect 381250 223443 381278 239672
rect 381346 229363 381374 239686
rect 381622 235235 381674 235241
rect 381622 235177 381674 235183
rect 381634 234945 381662 235177
rect 381622 234939 381674 234945
rect 381622 234881 381674 234887
rect 381730 232323 381758 239686
rect 382114 233983 382142 239686
rect 382560 239672 382814 239700
rect 382582 236863 382634 236869
rect 382582 236805 382634 236811
rect 382594 236763 382622 236805
rect 382786 236763 382814 239672
rect 382930 239404 382958 239686
rect 383328 239672 383582 239700
rect 383062 239527 383114 239533
rect 383062 239469 383114 239475
rect 382930 239376 383006 239404
rect 382580 236754 382636 236763
rect 382580 236689 382636 236698
rect 382772 236754 382828 236763
rect 382772 236689 382828 236698
rect 382774 234051 382826 234057
rect 382774 233993 382826 233999
rect 382102 233977 382154 233983
rect 382102 233919 382154 233925
rect 381716 232314 381772 232323
rect 381716 232249 381772 232258
rect 381332 229354 381388 229363
rect 381332 229289 381388 229298
rect 381718 228353 381770 228359
rect 381718 228295 381770 228301
rect 381730 226657 381758 228295
rect 381814 227465 381866 227471
rect 381814 227407 381866 227413
rect 381718 226651 381770 226657
rect 381718 226593 381770 226599
rect 381236 223434 381292 223443
rect 381236 223369 381292 223378
rect 381046 223173 381098 223179
rect 381046 223115 381098 223121
rect 381058 221496 381086 223115
rect 381058 221468 381120 221496
rect 381826 221482 381854 227407
rect 382678 225911 382730 225917
rect 382678 225853 382730 225859
rect 382690 225103 382718 225853
rect 382582 225097 382634 225103
rect 382582 225039 382634 225045
rect 382678 225097 382730 225103
rect 382678 225039 382730 225045
rect 382594 221496 382622 225039
rect 382786 222851 382814 233993
rect 382870 232867 382922 232873
rect 382870 232809 382922 232815
rect 382882 224733 382910 232809
rect 382978 231879 383006 239376
rect 383074 233835 383102 239469
rect 383062 233829 383114 233835
rect 383062 233771 383114 233777
rect 382964 231870 383020 231879
rect 382964 231805 383020 231814
rect 382966 229833 383018 229839
rect 382966 229775 383018 229781
rect 382978 225917 383006 229775
rect 383554 229511 383582 239672
rect 383650 234501 383678 239686
rect 384048 239672 384350 239700
rect 383638 234495 383690 234501
rect 383638 234437 383690 234443
rect 383540 229502 383596 229511
rect 383540 229437 383596 229446
rect 383254 228131 383306 228137
rect 383254 228073 383306 228079
rect 382966 225911 383018 225917
rect 382966 225853 383018 225859
rect 382870 224727 382922 224733
rect 382870 224669 382922 224675
rect 382772 222842 382828 222851
rect 382772 222777 382828 222786
rect 382560 221468 382622 221496
rect 383266 221496 383294 228073
rect 384022 227391 384074 227397
rect 384022 227333 384074 227339
rect 383266 221468 383328 221496
rect 384034 221482 384062 227333
rect 384322 223147 384350 239672
rect 384418 229215 384446 239686
rect 384768 239672 385022 239700
rect 385152 239672 385406 239700
rect 385536 239672 385790 239700
rect 384994 232175 385022 239672
rect 384980 232166 385036 232175
rect 384980 232101 385036 232110
rect 385378 232027 385406 239672
rect 385364 232018 385420 232027
rect 385364 231953 385420 231962
rect 384404 229206 384460 229215
rect 384404 229141 384460 229150
rect 385762 226509 385790 239672
rect 385858 235579 385886 239686
rect 386352 239672 386654 239700
rect 385942 236345 385994 236351
rect 385942 236287 385994 236293
rect 385954 236023 385982 236287
rect 385940 236014 385996 236023
rect 385940 235949 385996 235958
rect 385844 235570 385900 235579
rect 385844 235505 385900 235514
rect 385942 234199 385994 234205
rect 385942 234141 385994 234147
rect 385954 230949 385982 234141
rect 385942 230943 385994 230949
rect 385942 230885 385994 230891
rect 384790 226503 384842 226509
rect 384790 226445 384842 226451
rect 385750 226503 385802 226509
rect 385750 226445 385802 226451
rect 384308 223138 384364 223147
rect 384308 223073 384364 223082
rect 384802 221792 384830 226445
rect 386626 225843 386654 239672
rect 386722 235833 386750 239686
rect 387072 239672 387326 239700
rect 387456 239672 387710 239700
rect 387792 239672 388094 239700
rect 386710 235827 386762 235833
rect 386710 235769 386762 235775
rect 387298 226065 387326 239672
rect 387682 235283 387710 239672
rect 387956 236902 388012 236911
rect 387956 236837 388012 236846
rect 387970 236573 387998 236837
rect 387958 236567 388010 236573
rect 387958 236509 388010 236515
rect 387668 235274 387724 235283
rect 387668 235209 387724 235218
rect 387286 226059 387338 226065
rect 387286 226001 387338 226007
rect 388066 225991 388094 239672
rect 388162 227175 388190 239686
rect 388258 239672 388560 239700
rect 388944 239672 389150 239700
rect 389280 239672 389534 239700
rect 389664 239672 389918 239700
rect 388258 227397 388286 239672
rect 388724 237050 388780 237059
rect 388642 237008 388724 237036
rect 388342 236789 388394 236795
rect 388340 236754 388342 236763
rect 388394 236754 388396 236763
rect 388642 236721 388670 237008
rect 388724 236985 388780 236994
rect 388724 236902 388780 236911
rect 388724 236837 388726 236846
rect 388778 236837 388780 236846
rect 388726 236805 388778 236811
rect 389014 236789 389066 236795
rect 389014 236731 389066 236737
rect 388340 236689 388396 236698
rect 388630 236715 388682 236721
rect 388630 236657 388682 236663
rect 388630 236567 388682 236573
rect 388630 236509 388682 236515
rect 388642 236467 388670 236509
rect 388628 236458 388684 236467
rect 388628 236393 388684 236402
rect 389026 236319 389054 236731
rect 388820 236310 388876 236319
rect 388820 236245 388876 236254
rect 389012 236310 389068 236319
rect 389012 236245 389068 236254
rect 388834 236148 388862 236245
rect 389012 236162 389068 236171
rect 388834 236120 389012 236148
rect 389012 236097 389068 236106
rect 389122 229839 389150 239672
rect 389398 236789 389450 236795
rect 389398 236731 389450 236737
rect 389410 236023 389438 236731
rect 389396 236014 389452 236023
rect 389396 235949 389452 235958
rect 389110 229833 389162 229839
rect 389110 229775 389162 229781
rect 388246 227391 388298 227397
rect 388246 227333 388298 227339
rect 388150 227169 388202 227175
rect 388150 227111 388202 227117
rect 386998 225985 387050 225991
rect 386998 225927 387050 225933
rect 387766 225985 387818 225991
rect 387766 225927 387818 225933
rect 388054 225985 388106 225991
rect 388054 225927 388106 225933
rect 385558 225837 385610 225843
rect 385558 225779 385610 225785
rect 386614 225837 386666 225843
rect 386614 225779 386666 225785
rect 384802 221764 384878 221792
rect 384850 221482 384878 221764
rect 385570 221482 385598 225779
rect 386326 224727 386378 224733
rect 386326 224669 386378 224675
rect 386338 221482 386366 224669
rect 387010 221792 387038 225927
rect 387010 221764 387086 221792
rect 387058 221482 387086 221764
rect 387778 221482 387806 225927
rect 389506 225917 389534 239672
rect 389890 235019 389918 239672
rect 389878 235013 389930 235019
rect 389878 234955 389930 234961
rect 390082 227545 390110 239686
rect 390358 235161 390410 235167
rect 390358 235103 390410 235109
rect 390370 228137 390398 235103
rect 390358 228131 390410 228137
rect 390358 228073 390410 228079
rect 390070 227539 390122 227545
rect 390070 227481 390122 227487
rect 390070 226577 390122 226583
rect 390070 226519 390122 226525
rect 388726 225911 388778 225917
rect 388726 225853 388778 225859
rect 389494 225911 389546 225917
rect 389494 225853 389546 225859
rect 388738 225769 388766 225853
rect 388630 225763 388682 225769
rect 388630 225705 388682 225711
rect 388726 225763 388778 225769
rect 388726 225705 388778 225711
rect 389302 225763 389354 225769
rect 389302 225705 389354 225711
rect 388642 221482 388670 225705
rect 389314 221792 389342 225705
rect 389314 221764 389390 221792
rect 389362 221482 389390 221764
rect 390082 221482 390110 226519
rect 390466 224733 390494 239686
rect 390850 227471 390878 239686
rect 390838 227465 390890 227471
rect 390838 227407 390890 227413
rect 391234 227027 391262 239686
rect 391584 239672 391646 239700
rect 391968 239672 392222 239700
rect 391222 227021 391274 227027
rect 391222 226963 391274 226969
rect 391510 226799 391562 226805
rect 391510 226741 391562 226747
rect 390838 226355 390890 226361
rect 390838 226297 390890 226303
rect 390454 224727 390506 224733
rect 390454 224669 390506 224675
rect 390850 221482 390878 226297
rect 391522 221792 391550 226741
rect 391618 226699 391646 239672
rect 392194 235167 392222 239672
rect 392182 235161 392234 235167
rect 391796 235126 391852 235135
rect 392182 235103 392234 235109
rect 391796 235061 391852 235070
rect 391604 226690 391660 226699
rect 391604 226625 391660 226634
rect 391810 222439 391838 235061
rect 392290 227323 392318 239686
rect 392566 235901 392618 235907
rect 392564 235866 392566 235875
rect 392618 235866 392620 235875
rect 392564 235801 392620 235810
rect 392564 234386 392620 234395
rect 392564 234321 392620 234330
rect 392578 233655 392606 234321
rect 392564 233646 392620 233655
rect 392564 233581 392620 233590
rect 392374 228205 392426 228211
rect 392374 228147 392426 228153
rect 392278 227317 392330 227323
rect 392278 227259 392330 227265
rect 392086 226503 392138 226509
rect 392086 226445 392138 226451
rect 392098 225843 392126 226445
rect 392086 225837 392138 225843
rect 392086 225779 392138 225785
rect 391798 222433 391850 222439
rect 391798 222375 391850 222381
rect 391522 221764 391598 221792
rect 391570 221482 391598 221764
rect 392386 221482 392414 228147
rect 392674 227101 392702 239686
rect 392758 236049 392810 236055
rect 392758 235991 392810 235997
rect 392770 235852 392798 235991
rect 392770 235824 392990 235852
rect 392962 235759 392990 235824
rect 392854 235753 392906 235759
rect 392854 235695 392906 235701
rect 392950 235753 393002 235759
rect 392950 235695 393002 235701
rect 392866 235463 392894 235695
rect 392854 235457 392906 235463
rect 392854 235399 392906 235405
rect 393058 234691 393086 239686
rect 393140 235866 393196 235875
rect 393140 235801 393142 235810
rect 393194 235801 393196 235810
rect 393142 235769 393194 235775
rect 393442 234987 393470 239686
rect 393888 239672 394142 239700
rect 394272 239672 394526 239700
rect 393526 235087 393578 235093
rect 393526 235029 393578 235035
rect 393428 234978 393484 234987
rect 393428 234913 393484 234922
rect 392852 234682 392908 234691
rect 392852 234617 392908 234626
rect 393044 234682 393100 234691
rect 393044 234617 393100 234626
rect 392866 234395 392894 234617
rect 392852 234386 392908 234395
rect 392852 234321 392908 234330
rect 393538 228359 393566 235029
rect 393526 228353 393578 228359
rect 393526 228295 393578 228301
rect 392662 227095 392714 227101
rect 392662 227037 392714 227043
rect 393142 226947 393194 226953
rect 393142 226889 393194 226895
rect 393154 221482 393182 226889
rect 393814 226725 393866 226731
rect 393814 226667 393866 226673
rect 393826 221792 393854 226667
rect 394114 226403 394142 239672
rect 394498 226551 394526 239672
rect 394594 235093 394622 239686
rect 394978 235241 395006 239686
rect 395376 239672 395582 239700
rect 395712 239672 395870 239700
rect 396096 239672 396350 239700
rect 396480 239672 396638 239700
rect 395254 235383 395306 235389
rect 395254 235325 395306 235331
rect 394966 235235 395018 235241
rect 394966 235177 395018 235183
rect 394582 235087 394634 235093
rect 394582 235029 394634 235035
rect 394870 234125 394922 234131
rect 394870 234067 394922 234073
rect 394484 226542 394540 226551
rect 394484 226477 394540 226486
rect 394582 226429 394634 226435
rect 394100 226394 394156 226403
rect 394582 226371 394634 226377
rect 394100 226329 394156 226338
rect 393826 221764 393902 221792
rect 393874 221482 393902 221764
rect 394594 221482 394622 226371
rect 394882 223179 394910 234067
rect 395266 231319 395294 235325
rect 395254 231313 395306 231319
rect 395254 231255 395306 231261
rect 395350 231165 395402 231171
rect 395350 231107 395402 231113
rect 394870 223173 394922 223179
rect 394870 223115 394922 223121
rect 395362 221482 395390 231107
rect 395554 226953 395582 239672
rect 395734 234865 395786 234871
rect 395734 234807 395786 234813
rect 395746 231171 395774 234807
rect 395842 234205 395870 239672
rect 396322 235315 396350 239672
rect 396310 235309 396362 235315
rect 396310 235251 396362 235257
rect 396406 234791 396458 234797
rect 396406 234733 396458 234739
rect 396502 234791 396554 234797
rect 396502 234733 396554 234739
rect 395830 234199 395882 234205
rect 395830 234141 395882 234147
rect 395734 231165 395786 231171
rect 395734 231107 395786 231113
rect 396418 228211 396446 234733
rect 396514 234501 396542 234733
rect 396610 234501 396638 239672
rect 396694 239601 396746 239607
rect 396694 239543 396746 239549
rect 396706 235463 396734 239543
rect 396802 235463 396830 239686
rect 396694 235457 396746 235463
rect 396694 235399 396746 235405
rect 396790 235457 396842 235463
rect 396790 235399 396842 235405
rect 396502 234495 396554 234501
rect 396502 234437 396554 234443
rect 396598 234495 396650 234501
rect 396598 234437 396650 234443
rect 396982 229833 397034 229839
rect 396982 229775 397034 229781
rect 396406 228205 396458 228211
rect 396406 228147 396458 228153
rect 395542 226947 395594 226953
rect 395542 226889 395594 226895
rect 396118 226873 396170 226879
rect 396118 226815 396170 226821
rect 396130 221792 396158 226815
rect 396994 225695 397022 229775
rect 397186 226805 397214 239686
rect 397366 236271 397418 236277
rect 397366 236213 397418 236219
rect 397378 235537 397406 236213
rect 397366 235531 397418 235537
rect 397366 235473 397418 235479
rect 397666 226953 397694 239686
rect 398016 239672 398270 239700
rect 398400 239672 398558 239700
rect 398242 234871 398270 239672
rect 398422 239231 398474 239237
rect 398422 239173 398474 239179
rect 398434 235759 398462 239173
rect 398422 235753 398474 235759
rect 398422 235695 398474 235701
rect 398530 235389 398558 239672
rect 398626 239672 398784 239700
rect 398626 235759 398654 239672
rect 398996 237050 399052 237059
rect 398996 236985 399052 236994
rect 398708 236902 398764 236911
rect 399010 236888 399038 236985
rect 398764 236860 399038 236888
rect 398708 236837 398764 236846
rect 398614 235753 398666 235759
rect 398614 235695 398666 235701
rect 398518 235383 398570 235389
rect 398518 235325 398570 235331
rect 398806 234939 398858 234945
rect 398806 234881 398858 234887
rect 398230 234865 398282 234871
rect 398230 234807 398282 234813
rect 398818 233021 398846 234881
rect 398902 234717 398954 234723
rect 398902 234659 398954 234665
rect 398806 233015 398858 233021
rect 398806 232957 398858 232963
rect 398914 230505 398942 234659
rect 399106 234057 399134 239686
rect 399094 234051 399146 234057
rect 399094 233993 399146 233999
rect 398902 230499 398954 230505
rect 398902 230441 398954 230447
rect 399490 228919 399518 239686
rect 399874 235135 399902 239686
rect 400224 239672 400286 239700
rect 400608 239672 400862 239700
rect 400992 239672 401246 239700
rect 399860 235126 399916 235135
rect 399860 235061 399916 235070
rect 400258 234057 400286 239672
rect 400436 234830 400492 234839
rect 400436 234765 400492 234774
rect 400342 234569 400394 234575
rect 400342 234511 400394 234517
rect 400150 234051 400202 234057
rect 400150 233993 400202 233999
rect 400246 234051 400298 234057
rect 400246 233993 400298 233999
rect 399476 228910 399532 228919
rect 399476 228845 399532 228854
rect 398326 227983 398378 227989
rect 398326 227925 398378 227931
rect 397654 226947 397706 226953
rect 397654 226889 397706 226895
rect 397174 226799 397226 226805
rect 397174 226741 397226 226747
rect 397654 226651 397706 226657
rect 397654 226593 397706 226599
rect 396886 225689 396938 225695
rect 396886 225631 396938 225637
rect 396982 225689 397034 225695
rect 396982 225631 397034 225637
rect 396130 221764 396206 221792
rect 396178 221482 396206 221764
rect 396898 221482 396926 225631
rect 397666 221482 397694 226593
rect 398338 221792 398366 227925
rect 400162 225251 400190 233993
rect 400246 231831 400298 231837
rect 400246 231773 400298 231779
rect 399958 225245 400010 225251
rect 399958 225187 400010 225193
rect 400150 225245 400202 225251
rect 400150 225187 400202 225193
rect 399094 224949 399146 224955
rect 399094 224891 399146 224897
rect 398338 221764 398414 221792
rect 398386 221482 398414 221764
rect 399106 221482 399134 224891
rect 399970 221482 399998 225187
rect 400258 224752 400286 231773
rect 400354 231393 400382 234511
rect 400450 231467 400478 234765
rect 400726 233977 400778 233983
rect 400726 233919 400778 233925
rect 400738 233835 400766 233919
rect 400726 233829 400778 233835
rect 400726 233771 400778 233777
rect 400438 231461 400490 231467
rect 400438 231403 400490 231409
rect 400342 231387 400394 231393
rect 400342 231329 400394 231335
rect 400834 226731 400862 239672
rect 401218 235907 401246 239672
rect 401206 235901 401258 235907
rect 401410 235875 401438 239686
rect 401206 235843 401258 235849
rect 401396 235866 401452 235875
rect 401396 235801 401452 235810
rect 401794 234131 401822 239686
rect 401782 234125 401834 234131
rect 401782 234067 401834 234073
rect 401398 230721 401450 230727
rect 401398 230663 401450 230669
rect 400822 226725 400874 226731
rect 400822 226667 400874 226673
rect 400258 224724 400670 224752
rect 400642 221792 400670 224724
rect 400642 221764 400718 221792
rect 400690 221482 400718 221764
rect 401410 221482 401438 230663
rect 402178 226583 402206 239686
rect 402528 239672 402686 239700
rect 402912 239672 403166 239700
rect 402166 226577 402218 226583
rect 402166 226519 402218 226525
rect 402658 226435 402686 239672
rect 403138 236023 403166 239672
rect 403124 236014 403180 236023
rect 403124 235949 403180 235958
rect 403030 235457 403082 235463
rect 403030 235399 403082 235405
rect 403042 235241 403070 235399
rect 403030 235235 403082 235241
rect 403030 235177 403082 235183
rect 403126 235235 403178 235241
rect 403126 235177 403178 235183
rect 403138 235019 403166 235177
rect 403126 235013 403178 235019
rect 403126 234955 403178 234961
rect 403234 234205 403262 239686
rect 403316 235718 403372 235727
rect 403316 235653 403372 235662
rect 403126 234199 403178 234205
rect 403126 234141 403178 234147
rect 403222 234199 403274 234205
rect 403222 234141 403274 234147
rect 403138 229067 403166 234141
rect 403124 229058 403180 229067
rect 403124 228993 403180 229002
rect 403330 228507 403358 235653
rect 403618 235019 403646 239686
rect 404002 235431 404030 239686
rect 403988 235422 404044 235431
rect 403988 235357 404044 235366
rect 403606 235013 403658 235019
rect 403606 234955 403658 234961
rect 403318 228501 403370 228507
rect 403318 228443 403370 228449
rect 403702 227613 403754 227619
rect 403702 227555 403754 227561
rect 402646 226429 402698 226435
rect 402646 226371 402698 226377
rect 402838 226281 402890 226287
rect 402838 226223 402890 226229
rect 402166 224801 402218 224807
rect 402166 224743 402218 224749
rect 402178 221482 402206 224743
rect 402850 221792 402878 226223
rect 402850 221764 402926 221792
rect 402898 221482 402926 221764
rect 403714 221482 403742 227555
rect 404386 226509 404414 239686
rect 404736 239672 404990 239700
rect 405216 239672 405470 239700
rect 404470 230647 404522 230653
rect 404470 230589 404522 230595
rect 404374 226503 404426 226509
rect 404374 226445 404426 226451
rect 404482 221482 404510 230589
rect 404962 226361 404990 239672
rect 405046 234865 405098 234871
rect 405442 234839 405470 239672
rect 405538 235727 405566 239686
rect 405826 239672 405936 239700
rect 405524 235718 405580 235727
rect 405524 235653 405580 235662
rect 405046 234807 405098 234813
rect 405428 234830 405484 234839
rect 405058 231837 405086 234807
rect 405428 234765 405484 234774
rect 405716 234386 405772 234395
rect 405716 234321 405772 234330
rect 405046 231831 405098 231837
rect 405046 231773 405098 231779
rect 404950 226355 405002 226361
rect 404950 226297 405002 226303
rect 405142 224875 405194 224881
rect 405142 224817 405194 224823
rect 405154 221792 405182 224817
rect 405730 222703 405758 234321
rect 405826 226255 405854 239672
rect 406102 239379 406154 239385
rect 406102 239321 406154 239327
rect 406006 236863 406058 236869
rect 406006 236805 406058 236811
rect 405910 236567 405962 236573
rect 405910 236509 405962 236515
rect 405922 234247 405950 236509
rect 406018 236055 406046 236805
rect 406006 236049 406058 236055
rect 406006 235991 406058 235997
rect 406114 235833 406142 239321
rect 406306 236055 406334 239686
rect 406294 236049 406346 236055
rect 406294 235991 406346 235997
rect 406102 235827 406154 235833
rect 406102 235769 406154 235775
rect 406690 234945 406718 239686
rect 407040 239672 407294 239700
rect 407424 239672 407678 239700
rect 407158 236937 407210 236943
rect 407158 236879 407210 236885
rect 406678 234939 406730 234945
rect 406678 234881 406730 234887
rect 406870 234791 406922 234797
rect 406870 234733 406922 234739
rect 405908 234238 405964 234247
rect 405908 234173 405964 234182
rect 406882 229543 406910 234733
rect 406964 233646 407020 233655
rect 406964 233581 407020 233590
rect 406978 229839 407006 233581
rect 406966 229833 407018 229839
rect 406966 229775 407018 229781
rect 406774 229537 406826 229543
rect 406774 229479 406826 229485
rect 406870 229537 406922 229543
rect 406870 229479 406922 229485
rect 405812 226246 405868 226255
rect 405812 226181 405868 226190
rect 405910 225171 405962 225177
rect 405910 225113 405962 225119
rect 405716 222694 405772 222703
rect 405716 222629 405772 222638
rect 405154 221764 405230 221792
rect 405202 221482 405230 221764
rect 405922 221482 405950 225113
rect 406786 221482 406814 229479
rect 407170 221792 407198 236879
rect 407266 234247 407294 239672
rect 407252 234238 407308 234247
rect 407252 234173 407308 234182
rect 407650 226107 407678 239672
rect 407746 226287 407774 239686
rect 407926 234865 407978 234871
rect 407926 234807 407978 234813
rect 407938 234691 407966 234807
rect 408130 234691 408158 239686
rect 407924 234682 407980 234691
rect 407924 234617 407980 234626
rect 408116 234682 408172 234691
rect 408116 234617 408172 234626
rect 408022 234495 408074 234501
rect 408022 234437 408074 234443
rect 408034 234057 408062 234437
rect 408514 234395 408542 239686
rect 408960 239672 409214 239700
rect 409728 239672 409982 239700
rect 408692 237050 408748 237059
rect 408692 236985 408748 236994
rect 408884 237050 408940 237059
rect 409186 237036 409214 239672
rect 409186 237008 409310 237036
rect 408884 236985 408940 236994
rect 408706 236721 408734 236985
rect 408788 236754 408844 236763
rect 408694 236715 408746 236721
rect 408788 236689 408844 236698
rect 408694 236657 408746 236663
rect 408802 236647 408830 236689
rect 408790 236641 408842 236647
rect 408790 236583 408842 236589
rect 408898 236444 408926 236985
rect 408982 236937 409034 236943
rect 408980 236902 408982 236911
rect 409034 236902 409036 236911
rect 408980 236837 409036 236846
rect 409174 236863 409226 236869
rect 409174 236805 409226 236811
rect 408706 236416 408926 236444
rect 408706 236319 408734 236416
rect 409186 236319 409214 236805
rect 408692 236310 408748 236319
rect 408692 236245 408748 236254
rect 409172 236310 409228 236319
rect 409172 236245 409228 236254
rect 408788 236162 408844 236171
rect 408788 236097 408844 236106
rect 408802 235875 408830 236097
rect 408788 235866 408844 235875
rect 408788 235801 408844 235810
rect 408788 234978 408844 234987
rect 408788 234913 408844 234922
rect 408802 234871 408830 234913
rect 408790 234865 408842 234871
rect 408790 234807 408842 234813
rect 409282 234501 409310 237008
rect 409364 236902 409420 236911
rect 409364 236837 409420 236846
rect 409378 236795 409406 236837
rect 409366 236789 409418 236795
rect 409366 236731 409418 236737
rect 409954 234871 409982 239672
rect 410050 236129 410078 239686
rect 410038 236123 410090 236129
rect 410038 236065 410090 236071
rect 409942 234865 409994 234871
rect 409942 234807 409994 234813
rect 409270 234495 409322 234501
rect 409270 234437 409322 234443
rect 408500 234386 408556 234395
rect 408500 234321 408556 234330
rect 408022 234051 408074 234057
rect 408022 233993 408074 233999
rect 409654 231017 409706 231023
rect 409654 230959 409706 230965
rect 407734 226281 407786 226287
rect 407734 226223 407786 226229
rect 408982 226207 409034 226213
rect 408982 226149 409034 226155
rect 407636 226098 407692 226107
rect 407636 226033 407692 226042
rect 408214 225023 408266 225029
rect 408214 224965 408266 224971
rect 407170 221764 407534 221792
rect 407506 221482 407534 221764
rect 408226 221482 408254 224965
rect 408994 221482 409022 226149
rect 409666 221792 409694 230959
rect 410434 225177 410462 239686
rect 410818 234575 410846 239686
rect 411168 239672 411326 239700
rect 411190 237085 411242 237091
rect 411190 237027 411242 237033
rect 411202 236795 411230 237027
rect 411190 236789 411242 236795
rect 411190 236731 411242 236737
rect 410902 235827 410954 235833
rect 410902 235769 410954 235775
rect 410806 234569 410858 234575
rect 410806 234511 410858 234517
rect 410914 233465 410942 235769
rect 411298 234723 411326 239672
rect 411394 239672 411552 239700
rect 411936 239672 412190 239700
rect 411286 234717 411338 234723
rect 411286 234659 411338 234665
rect 410902 233459 410954 233465
rect 410902 233401 410954 233407
rect 410518 230499 410570 230505
rect 410518 230441 410570 230447
rect 410422 225171 410474 225177
rect 410422 225113 410474 225119
rect 409666 221764 409742 221792
rect 409714 221482 409742 221764
rect 410530 221482 410558 230441
rect 411394 226139 411422 239672
rect 411766 239157 411818 239163
rect 411766 239099 411818 239105
rect 411478 237159 411530 237165
rect 411478 237101 411530 237107
rect 411670 237159 411722 237165
rect 411670 237101 411722 237107
rect 411490 236869 411518 237101
rect 411574 237085 411626 237091
rect 411574 237027 411626 237033
rect 411478 236863 411530 236869
rect 411478 236805 411530 236811
rect 411478 236493 411530 236499
rect 411478 236435 411530 236441
rect 411490 233687 411518 236435
rect 411586 233803 411614 237027
rect 411682 235981 411710 237101
rect 411670 235975 411722 235981
rect 411670 235917 411722 235923
rect 411778 235907 411806 239099
rect 411766 235901 411818 235907
rect 411766 235843 411818 235849
rect 412162 234797 412190 239672
rect 412258 239607 412286 240685
rect 412340 240010 412396 240019
rect 412340 239945 412396 239954
rect 412246 239601 412298 239607
rect 412246 239543 412298 239549
rect 412354 239385 412382 239945
rect 412342 239379 412394 239385
rect 412342 239321 412394 239327
rect 412450 239089 412478 241425
rect 420308 241194 420364 241203
rect 420308 241129 420364 241138
rect 412724 240898 412780 240907
rect 412724 240833 412780 240842
rect 412628 240602 412684 240611
rect 412628 240537 412684 240546
rect 412532 240158 412588 240167
rect 412532 240093 412588 240102
rect 412438 239083 412490 239089
rect 412438 239025 412490 239031
rect 412546 236573 412574 240093
rect 412642 239163 412670 240537
rect 412630 239157 412682 239163
rect 412630 239099 412682 239105
rect 412738 237165 412766 240833
rect 413014 239971 413066 239977
rect 413014 239913 413066 239919
rect 412918 239601 412970 239607
rect 412918 239543 412970 239549
rect 412822 239379 412874 239385
rect 412822 239321 412874 239327
rect 412726 237159 412778 237165
rect 412726 237101 412778 237107
rect 412834 237091 412862 239321
rect 412822 237085 412874 237091
rect 412822 237027 412874 237033
rect 412534 236567 412586 236573
rect 412534 236509 412586 236515
rect 412930 236499 412958 239543
rect 412918 236493 412970 236499
rect 412918 236435 412970 236441
rect 413026 235833 413054 239913
rect 420322 239163 420350 241129
rect 566708 240750 566764 240759
rect 566708 240685 566764 240694
rect 544820 240306 544876 240315
rect 544820 240241 544876 240250
rect 541460 240158 541516 240167
rect 541460 240093 541516 240102
rect 442198 239971 442250 239977
rect 442198 239913 442250 239919
rect 434614 239749 434666 239755
rect 434614 239691 434666 239697
rect 420310 239157 420362 239163
rect 420310 239099 420362 239105
rect 413396 238974 413452 238983
rect 413396 238909 413452 238918
rect 413410 236647 413438 238909
rect 413684 238678 413740 238687
rect 413684 238613 413740 238622
rect 413698 236721 413726 238613
rect 413972 238382 414028 238391
rect 413972 238317 414028 238326
rect 413986 236943 414014 238317
rect 414260 238234 414316 238243
rect 414260 238169 414316 238178
rect 413974 236937 414026 236943
rect 413974 236879 414026 236885
rect 413686 236715 413738 236721
rect 413686 236657 413738 236663
rect 413398 236641 413450 236647
rect 413398 236583 413450 236589
rect 413014 235827 413066 235833
rect 413014 235769 413066 235775
rect 412150 234791 412202 234797
rect 412150 234733 412202 234739
rect 414274 233951 414302 238169
rect 414452 238086 414508 238095
rect 414452 238021 414508 238030
rect 414466 236319 414494 238021
rect 432406 237233 432458 237239
rect 432406 237175 432458 237181
rect 420310 237011 420362 237017
rect 420310 236953 420362 236959
rect 414550 236419 414602 236425
rect 414550 236361 414602 236367
rect 414452 236310 414508 236319
rect 414452 236245 414508 236254
rect 414260 233942 414316 233951
rect 414260 233877 414316 233886
rect 411766 233829 411818 233835
rect 411572 233794 411628 233803
rect 411766 233771 411818 233777
rect 411572 233729 411628 233738
rect 411478 233681 411530 233687
rect 411478 233623 411530 233629
rect 411778 232873 411806 233771
rect 414562 233391 414590 236361
rect 414644 236310 414700 236319
rect 414644 236245 414700 236254
rect 414658 236055 414686 236245
rect 414646 236049 414698 236055
rect 414646 235991 414698 235997
rect 416374 234347 416426 234353
rect 416374 234289 416426 234295
rect 414550 233385 414602 233391
rect 414550 233327 414602 233333
rect 411766 232867 411818 232873
rect 411766 232809 411818 232815
rect 415700 231130 415756 231139
rect 415700 231065 415756 231074
rect 413494 228427 413546 228433
rect 413494 228369 413546 228375
rect 412726 228057 412778 228063
rect 412726 227999 412778 228005
rect 411286 226133 411338 226139
rect 411286 226075 411338 226081
rect 411382 226133 411434 226139
rect 411382 226075 411434 226081
rect 411298 221496 411326 226075
rect 411958 225319 412010 225325
rect 411958 225261 412010 225267
rect 411264 221468 411326 221496
rect 411970 221496 411998 225261
rect 411970 221468 412032 221496
rect 412738 221482 412766 227999
rect 413506 221496 413534 228369
rect 415030 225393 415082 225399
rect 415030 225335 415082 225341
rect 414262 222507 414314 222513
rect 414262 222449 414314 222455
rect 413472 221468 413534 221496
rect 414274 221482 414302 222449
rect 415042 221482 415070 225335
rect 415714 221792 415742 231065
rect 416386 231023 416414 234289
rect 418294 234273 418346 234279
rect 418294 234215 418346 234221
rect 416470 231239 416522 231245
rect 416470 231181 416522 231187
rect 416374 231017 416426 231023
rect 416374 230959 416426 230965
rect 415714 221764 415790 221792
rect 415762 221482 415790 221764
rect 416482 221482 416510 231181
rect 418306 227619 418334 234215
rect 419542 230869 419594 230875
rect 419542 230811 419594 230817
rect 418774 228575 418826 228581
rect 418774 228517 418826 228523
rect 418294 227613 418346 227619
rect 418294 227555 418346 227561
rect 418006 225097 418058 225103
rect 418006 225039 418058 225045
rect 417238 222581 417290 222587
rect 417238 222523 417290 222529
rect 417250 221482 417278 222523
rect 418018 221792 418046 225039
rect 418018 221764 418094 221792
rect 418066 221482 418094 221764
rect 418786 221482 418814 228517
rect 419554 221482 419582 230811
rect 420322 221792 420350 236953
rect 426358 236863 426410 236869
rect 426358 236805 426410 236811
rect 423382 234421 423434 234427
rect 423382 234363 423434 234369
rect 423394 230505 423422 234363
rect 424724 231278 424780 231287
rect 424724 231213 424780 231222
rect 424054 231017 424106 231023
rect 424054 230959 424106 230965
rect 423382 230499 423434 230505
rect 423382 230441 423434 230447
rect 421846 228649 421898 228655
rect 421846 228591 421898 228597
rect 420982 225467 421034 225473
rect 420982 225409 421034 225415
rect 420274 221764 420350 221792
rect 420274 221482 420302 221764
rect 420994 221482 421022 225409
rect 421858 221482 421886 228591
rect 422518 222803 422570 222809
rect 422518 222745 422570 222751
rect 422530 221792 422558 222745
rect 423286 222655 423338 222661
rect 423286 222597 423338 222603
rect 422530 221764 422606 221792
rect 422578 221482 422606 221764
rect 423298 221482 423326 222597
rect 424066 221482 424094 230959
rect 424738 221792 424766 231213
rect 425590 228723 425642 228729
rect 425590 228665 425642 228671
rect 424738 221764 424814 221792
rect 424786 221482 424814 221764
rect 425602 221482 425630 228665
rect 426370 221482 426398 236805
rect 428662 236789 428714 236795
rect 428662 236731 428714 236737
rect 428276 234090 428332 234099
rect 428276 234025 428332 234034
rect 428290 228803 428318 234025
rect 427798 228797 427850 228803
rect 427798 228739 427850 228745
rect 428278 228797 428330 228803
rect 428278 228739 428330 228745
rect 427030 225541 427082 225547
rect 427030 225483 427082 225489
rect 427042 221792 427070 225483
rect 427042 221764 427118 221792
rect 427090 221482 427118 221764
rect 427810 221482 427838 228739
rect 428674 221482 428702 236731
rect 430102 236419 430154 236425
rect 430102 236361 430154 236367
rect 429334 222877 429386 222883
rect 429334 222819 429386 222825
rect 429346 221792 429374 222819
rect 429346 221764 429422 221792
rect 429394 221482 429422 221764
rect 430114 221482 430142 236361
rect 432022 233903 432074 233909
rect 432022 233845 432074 233851
rect 432034 228729 432062 233845
rect 432022 228723 432074 228729
rect 432022 228665 432074 228671
rect 430868 228318 430924 228327
rect 430868 228253 430924 228262
rect 430882 221482 430910 228253
rect 431542 222729 431594 222735
rect 431542 222671 431594 222677
rect 431554 221792 431582 222671
rect 431554 221764 431630 221792
rect 431602 221482 431630 221764
rect 432418 221482 432446 237175
rect 433846 231535 433898 231541
rect 433846 231477 433898 231483
rect 433174 227613 433226 227619
rect 433174 227555 433226 227561
rect 433186 221482 433214 227555
rect 433858 221792 433886 231477
rect 433858 221764 433934 221792
rect 433906 221482 433934 221764
rect 434626 221482 434654 239691
rect 441430 237381 441482 237387
rect 441430 237323 441482 237329
rect 438358 237307 438410 237313
rect 438358 237249 438410 237255
rect 434902 234643 434954 234649
rect 434902 234585 434954 234591
rect 434914 228655 434942 234585
rect 436150 230499 436202 230505
rect 436150 230441 436202 230447
rect 434902 228649 434954 228655
rect 434902 228591 434954 228597
rect 435382 222951 435434 222957
rect 435382 222893 435434 222899
rect 435394 221482 435422 222893
rect 436162 221792 436190 230441
rect 436916 228466 436972 228475
rect 436916 228401 436972 228410
rect 436162 221764 436238 221792
rect 436210 221482 436238 221764
rect 436930 221482 436958 228401
rect 437686 228205 437738 228211
rect 437686 228147 437738 228153
rect 437698 221482 437726 228147
rect 438370 221792 438398 237249
rect 441442 236174 441470 237323
rect 440770 236146 441470 236174
rect 439990 228871 440042 228877
rect 439990 228813 440042 228819
rect 439126 225615 439178 225621
rect 439126 225557 439178 225563
rect 438370 221764 438446 221792
rect 438418 221482 438446 221764
rect 439138 221482 439166 225557
rect 440002 221496 440030 228813
rect 440770 221792 440798 236146
rect 441430 223099 441482 223105
rect 441430 223041 441482 223047
rect 439968 221468 440030 221496
rect 440722 221764 440798 221792
rect 440722 221482 440750 221764
rect 441442 221482 441470 223041
rect 442210 221496 442238 239913
rect 508630 239823 508682 239829
rect 508630 239765 508682 239771
rect 446710 239675 446762 239681
rect 446710 239617 446762 239623
rect 444502 237455 444554 237461
rect 444502 237397 444554 237403
rect 442868 231426 442924 231435
rect 442868 231361 442924 231370
rect 442176 221468 442238 221496
rect 442882 221496 442910 231361
rect 443734 223025 443786 223031
rect 443734 222967 443786 222973
rect 442882 221468 442944 221496
rect 443746 221482 443774 222967
rect 444514 221792 444542 237397
rect 445942 228945 445994 228951
rect 445942 228887 445994 228893
rect 445172 225506 445228 225515
rect 445172 225441 445228 225450
rect 444466 221764 444542 221792
rect 444466 221482 444494 221764
rect 445186 221482 445214 225441
rect 445954 221482 445982 228887
rect 446722 221792 446750 239617
rect 495766 239601 495818 239607
rect 495766 239543 495818 239549
rect 470902 239527 470954 239533
rect 470902 239469 470954 239475
rect 458806 239453 458858 239459
rect 458806 239395 458858 239401
rect 455158 239009 455210 239015
rect 455158 238951 455210 238957
rect 455062 238935 455114 238941
rect 455062 238877 455114 238883
rect 449302 237529 449354 237535
rect 449302 237471 449354 237477
rect 449314 236174 449342 237471
rect 449314 236146 450494 236174
rect 449302 233607 449354 233613
rect 449302 233549 449354 233555
rect 448246 233311 448298 233317
rect 448246 233253 448298 233259
rect 447478 224579 447530 224585
rect 447478 224521 447530 224527
rect 446674 221764 446750 221792
rect 446674 221482 446702 221764
rect 447490 221482 447518 224521
rect 448258 221482 448286 233253
rect 448916 231574 448972 231583
rect 448916 231509 448972 231518
rect 448930 221792 448958 231509
rect 449314 228951 449342 233549
rect 449686 230943 449738 230949
rect 449686 230885 449738 230891
rect 449302 228945 449354 228951
rect 449302 228887 449354 228893
rect 448930 221764 449006 221792
rect 448978 221482 449006 221764
rect 449698 221482 449726 230885
rect 450466 221482 450494 236146
rect 451990 230425 452042 230431
rect 451990 230367 452042 230373
rect 451220 225654 451276 225663
rect 451220 225589 451276 225598
rect 451234 221792 451262 225589
rect 451234 221764 451310 221792
rect 451282 221482 451310 221764
rect 452002 221482 452030 230367
rect 454294 228649 454346 228655
rect 454294 228591 454346 228597
rect 452758 224653 452810 224659
rect 452758 224595 452810 224601
rect 452770 221482 452798 224595
rect 453430 224505 453482 224511
rect 453430 224447 453482 224453
rect 453442 221792 453470 224447
rect 453442 221764 453518 221792
rect 453490 221482 453518 221764
rect 454306 221482 454334 228591
rect 455074 228581 455102 238877
rect 455170 236174 455198 238951
rect 455170 236146 455774 236174
rect 455156 231722 455212 231731
rect 455156 231657 455212 231666
rect 455062 228575 455114 228581
rect 455062 228517 455114 228523
rect 455170 226232 455198 231657
rect 455074 226204 455198 226232
rect 455074 221482 455102 226204
rect 455746 221792 455774 236146
rect 458038 230277 458090 230283
rect 458038 230219 458090 230225
rect 456502 228575 456554 228581
rect 456502 228517 456554 228523
rect 455746 221764 455822 221792
rect 455794 221482 455822 221764
rect 456514 221482 456542 228517
rect 457268 225358 457324 225367
rect 457268 225293 457324 225302
rect 457282 221482 457310 225293
rect 458050 221792 458078 230219
rect 458050 221764 458126 221792
rect 458098 221482 458126 221764
rect 458818 221482 458846 239395
rect 462550 238861 462602 238867
rect 462550 238803 462602 238809
rect 460246 235679 460298 235685
rect 460246 235621 460298 235627
rect 459574 224431 459626 224437
rect 459574 224373 459626 224379
rect 459586 221482 459614 224373
rect 460258 221792 460286 235621
rect 461014 230351 461066 230357
rect 461014 230293 461066 230299
rect 460258 221764 460334 221792
rect 460306 221482 460334 221764
rect 461026 221482 461054 230293
rect 461878 228131 461930 228137
rect 461878 228073 461930 228079
rect 461890 221482 461918 228073
rect 462562 221792 462590 238803
rect 464758 238787 464810 238793
rect 464758 238729 464810 238735
rect 464566 233755 464618 233761
rect 464566 233697 464618 233703
rect 463606 233533 463658 233539
rect 463606 233475 463658 233481
rect 463618 230357 463646 233475
rect 464086 231609 464138 231615
rect 464086 231551 464138 231557
rect 463606 230351 463658 230357
rect 463606 230293 463658 230299
rect 463316 225802 463372 225811
rect 463316 225737 463372 225746
rect 462562 221764 462638 221792
rect 462610 221482 462638 221764
rect 463330 221482 463358 225737
rect 464098 221482 464126 231551
rect 464578 230283 464606 233697
rect 464566 230277 464618 230283
rect 464566 230219 464618 230225
rect 464770 221792 464798 238729
rect 468598 238713 468650 238719
rect 468598 238655 468650 238661
rect 467062 230203 467114 230209
rect 467062 230145 467114 230151
rect 466390 228945 466442 228951
rect 466390 228887 466442 228893
rect 465622 224357 465674 224363
rect 465622 224299 465674 224305
rect 464770 221764 464846 221792
rect 464818 221482 464846 221764
rect 465634 221482 465662 224299
rect 466402 221482 466430 228887
rect 467074 221792 467102 230145
rect 467830 222359 467882 222365
rect 467830 222301 467882 222307
rect 467074 221764 467150 221792
rect 467122 221482 467150 221764
rect 467842 221482 467870 222301
rect 468610 221482 468638 238655
rect 470132 233202 470188 233211
rect 470132 233137 470188 233146
rect 469364 227430 469420 227439
rect 469364 227365 469420 227374
rect 469378 221496 469406 227365
rect 469378 221468 469440 221496
rect 470146 221482 470174 233137
rect 470914 221496 470942 239469
rect 488278 239305 488330 239311
rect 488278 239247 488330 239253
rect 474646 238639 474698 238645
rect 474646 238581 474698 238587
rect 472342 235605 472394 235611
rect 472342 235547 472394 235553
rect 471574 224283 471626 224289
rect 471574 224225 471626 224231
rect 470880 221468 470942 221496
rect 471586 221496 471614 224225
rect 471586 221468 471648 221496
rect 472354 221482 472382 235547
rect 473878 231165 473930 231171
rect 473878 231107 473930 231113
rect 473110 230129 473162 230135
rect 473110 230071 473162 230077
rect 473122 221792 473150 230071
rect 473122 221764 473198 221792
rect 473170 221482 473198 221764
rect 473890 221482 473918 231107
rect 474658 221482 474686 238581
rect 480694 238565 480746 238571
rect 480694 238507 480746 238513
rect 479158 238491 479210 238497
rect 479158 238433 479210 238439
rect 479170 236174 479198 238433
rect 479170 236146 479966 236174
rect 475222 234051 475274 234057
rect 475222 233993 475274 233999
rect 475234 230209 475262 233993
rect 479254 233977 479306 233983
rect 479254 233919 479306 233925
rect 479156 233054 479212 233063
rect 479156 232989 479212 232998
rect 478390 230351 478442 230357
rect 478390 230293 478442 230299
rect 475222 230203 475274 230209
rect 475222 230145 475274 230151
rect 476180 228614 476236 228623
rect 476180 228549 476236 228558
rect 475316 227282 475372 227291
rect 475316 227217 475372 227226
rect 475330 221792 475358 227217
rect 475330 221764 475406 221792
rect 475378 221482 475406 221764
rect 476194 221482 476222 228549
rect 476950 228353 477002 228359
rect 476950 228295 477002 228301
rect 476962 221482 476990 228295
rect 477622 224135 477674 224141
rect 477622 224077 477674 224083
rect 477634 221792 477662 224077
rect 477634 221764 477710 221792
rect 477682 221482 477710 221764
rect 478402 221482 478430 230293
rect 479170 221482 479198 232989
rect 479266 230135 479294 233919
rect 479254 230129 479306 230135
rect 479254 230071 479306 230077
rect 479938 221792 479966 236146
rect 479938 221764 480014 221792
rect 479986 221482 480014 221764
rect 480706 221482 480734 238507
rect 486742 238417 486794 238423
rect 486742 238359 486794 238365
rect 486646 234125 486698 234131
rect 486646 234067 486698 234073
rect 485206 231683 485258 231689
rect 485206 231625 485258 231631
rect 484438 230277 484490 230283
rect 484438 230219 484490 230225
rect 482134 230055 482186 230061
rect 482134 229997 482186 230003
rect 481460 227134 481516 227143
rect 481460 227069 481516 227078
rect 481474 221482 481502 227069
rect 482146 221792 482174 229997
rect 482902 224209 482954 224215
rect 482902 224151 482954 224157
rect 482146 221764 482222 221792
rect 482194 221482 482222 221764
rect 482914 221482 482942 224151
rect 483766 224061 483818 224067
rect 483766 224003 483818 224009
rect 483778 221482 483806 224003
rect 484450 221792 484478 230219
rect 484450 221764 484526 221792
rect 484498 221482 484526 221764
rect 485218 221482 485246 231625
rect 485974 231313 486026 231319
rect 485974 231255 486026 231261
rect 485986 221482 486014 231255
rect 486658 230061 486686 234067
rect 486646 230055 486698 230061
rect 486646 229997 486698 230003
rect 486754 221792 486782 238359
rect 488290 236174 488318 239247
rect 492790 238343 492842 238349
rect 492790 238285 492842 238291
rect 492022 236345 492074 236351
rect 492022 236287 492074 236293
rect 488290 236146 488990 236174
rect 488276 228762 488332 228771
rect 488276 228697 488332 228706
rect 487508 225950 487564 225959
rect 487508 225885 487564 225894
rect 486706 221764 486782 221792
rect 486706 221482 486734 221764
rect 487522 221482 487550 225885
rect 488290 221482 488318 228697
rect 488962 221792 488990 236146
rect 490484 234534 490540 234543
rect 490484 234469 490540 234478
rect 489718 223987 489770 223993
rect 489718 223929 489770 223935
rect 488962 221764 489038 221792
rect 489010 221482 489038 221764
rect 489730 221482 489758 223929
rect 490498 221482 490526 234469
rect 491254 233237 491306 233243
rect 491254 233179 491306 233185
rect 491266 221792 491294 233179
rect 491266 221764 491342 221792
rect 491314 221482 491342 221764
rect 492034 221482 492062 236287
rect 492802 221482 492830 238285
rect 495380 234238 495436 234247
rect 495380 234173 495436 234182
rect 495394 233243 495422 234173
rect 495382 233237 495434 233243
rect 495382 233179 495434 233185
rect 495094 231757 495146 231763
rect 495094 231699 495146 231705
rect 494228 230390 494284 230399
rect 494228 230325 494284 230334
rect 493460 226986 493516 226995
rect 493460 226921 493516 226930
rect 493474 221792 493502 226921
rect 493474 221764 493550 221792
rect 493522 221482 493550 221764
rect 494242 221482 494270 230325
rect 495106 221482 495134 231699
rect 495778 221792 495806 239543
rect 502582 239379 502634 239385
rect 502582 239321 502634 239327
rect 500278 238269 500330 238275
rect 500278 238211 500330 238217
rect 498550 234199 498602 234205
rect 498550 234141 498602 234147
rect 498562 231763 498590 234141
rect 498550 231757 498602 231763
rect 498550 231699 498602 231705
rect 499606 231387 499658 231393
rect 499606 231329 499658 231335
rect 497972 230242 498028 230251
rect 497972 230177 498028 230186
rect 497302 223913 497354 223919
rect 497302 223855 497354 223861
rect 496534 222433 496586 222439
rect 496534 222375 496586 222381
rect 495778 221764 495854 221792
rect 495826 221482 495854 221764
rect 496546 221482 496574 222375
rect 497314 221482 497342 223855
rect 497986 221792 498014 230177
rect 498836 226838 498892 226847
rect 498836 226773 498892 226782
rect 497986 221764 498062 221792
rect 498034 221482 498062 221764
rect 498850 221482 498878 226773
rect 499618 221496 499646 231329
rect 499584 221468 499646 221496
rect 500290 221496 500318 238211
rect 501046 233163 501098 233169
rect 501046 233105 501098 233111
rect 500290 221468 500352 221496
rect 501058 221482 501086 233105
rect 501814 223839 501866 223845
rect 501814 223781 501866 223787
rect 501826 221792 501854 223781
rect 501826 221764 501902 221792
rect 501874 221482 501902 221764
rect 502594 221482 502622 239321
rect 503350 238195 503402 238201
rect 503350 238137 503402 238143
rect 503362 221482 503390 238137
rect 505654 236271 505706 236277
rect 505654 236213 505706 236219
rect 504022 229981 504074 229987
rect 504022 229923 504074 229929
rect 504034 221792 504062 229923
rect 504790 223765 504842 223771
rect 504790 223707 504842 223713
rect 504034 221764 504110 221792
rect 504082 221482 504110 221764
rect 504802 221482 504830 223707
rect 505666 221482 505694 236213
rect 507094 233089 507146 233095
rect 507094 233031 507146 233037
rect 506326 223543 506378 223549
rect 506326 223485 506378 223491
rect 506338 221792 506366 223485
rect 506338 221764 506414 221792
rect 506386 221482 506414 221764
rect 507106 221482 507134 233031
rect 507862 223691 507914 223697
rect 507862 223633 507914 223639
rect 507874 221482 507902 223633
rect 508642 221792 508670 239765
rect 532822 239231 532874 239237
rect 532822 239173 532874 239179
rect 509398 238121 509450 238127
rect 509398 238063 509450 238069
rect 508594 221764 508670 221792
rect 508594 221482 508622 221764
rect 509410 221482 509438 238063
rect 514678 238047 514730 238053
rect 514678 237989 514730 237995
rect 512758 237973 512810 237979
rect 512758 237915 512810 237921
rect 511606 236197 511658 236203
rect 511606 236139 511658 236145
rect 510166 229907 510218 229913
rect 510166 229849 510218 229855
rect 510178 221482 510206 229849
rect 510838 223617 510890 223623
rect 510838 223559 510890 223565
rect 510850 221792 510878 223559
rect 510850 221764 510926 221792
rect 510898 221482 510926 221764
rect 511618 221482 511646 236139
rect 512180 234386 512236 234395
rect 512180 234321 512236 234330
rect 512194 229913 512222 234321
rect 512182 229907 512234 229913
rect 512182 229849 512234 229855
rect 512374 223469 512426 223475
rect 512374 223411 512426 223417
rect 512386 221482 512414 223411
rect 512770 221773 512798 237915
rect 513058 233012 513278 233040
rect 513058 232799 513086 233012
rect 513250 232947 513278 233012
rect 513142 232941 513194 232947
rect 513142 232883 513194 232889
rect 513238 232941 513290 232947
rect 513238 232883 513290 232889
rect 513046 232793 513098 232799
rect 513046 232735 513098 232741
rect 513154 221792 513182 232883
rect 513910 223395 513962 223401
rect 513910 223337 513962 223343
rect 512758 221767 512810 221773
rect 513154 221764 513230 221792
rect 512758 221709 512810 221715
rect 513202 221482 513230 221764
rect 513922 221482 513950 223337
rect 514690 221482 514718 237989
rect 521494 237899 521546 237905
rect 521494 237841 521546 237847
rect 521206 234495 521258 234501
rect 521206 234437 521258 234443
rect 519190 232941 519242 232947
rect 519190 232883 519242 232889
rect 516118 229759 516170 229765
rect 516118 229701 516170 229707
rect 515398 221767 515450 221773
rect 515398 221709 515450 221715
rect 515410 221482 515438 221709
rect 516130 221482 516158 229701
rect 517654 228501 517706 228507
rect 517654 228443 517706 228449
rect 516982 223321 517034 223327
rect 516982 223263 517034 223269
rect 516994 221482 517022 223263
rect 517666 221792 517694 228443
rect 518420 224618 518476 224627
rect 518420 224553 518476 224562
rect 517666 221764 517742 221792
rect 517714 221482 517742 221764
rect 518434 221482 518462 224553
rect 519202 221482 519230 232883
rect 521218 232799 521246 234437
rect 521206 232793 521258 232799
rect 521206 232735 521258 232741
rect 520726 231461 520778 231467
rect 520726 231403 520778 231409
rect 519862 223247 519914 223253
rect 519862 223189 519914 223195
rect 519874 221792 519902 223189
rect 519874 221764 519950 221792
rect 519922 221482 519950 221764
rect 520738 221482 520766 231403
rect 521506 221482 521534 237841
rect 526006 237825 526058 237831
rect 526006 237767 526058 237773
rect 522646 234569 522698 234575
rect 522646 234511 522698 234517
rect 522658 229691 522686 234511
rect 525236 232906 525292 232915
rect 525236 232841 525292 232850
rect 522166 229685 522218 229691
rect 522166 229627 522218 229633
rect 522646 229685 522698 229691
rect 522646 229627 522698 229633
rect 522178 221792 522206 229627
rect 524468 224470 524524 224479
rect 524468 224405 524524 224414
rect 523798 223173 523850 223179
rect 523798 223115 523850 223121
rect 522932 222694 522988 222703
rect 522932 222629 522988 222638
rect 522178 221764 522254 221792
rect 522226 221482 522254 221764
rect 522946 221482 522974 222629
rect 523810 221482 523838 223115
rect 524482 221792 524510 224405
rect 524482 221764 524558 221792
rect 524530 221482 524558 221764
rect 525250 221482 525278 232841
rect 526018 221482 526046 237767
rect 528502 236123 528554 236129
rect 528502 236065 528554 236071
rect 528406 235753 528458 235759
rect 528406 235695 528458 235701
rect 527540 229946 527596 229955
rect 527540 229881 527596 229890
rect 526676 222990 526732 222999
rect 526676 222925 526732 222934
rect 526690 221792 526718 222925
rect 526690 221764 526766 221792
rect 526738 221482 526766 221764
rect 527554 221482 527582 229881
rect 528418 229765 528446 235695
rect 528406 229759 528458 229765
rect 528406 229701 528458 229707
rect 528514 229617 528542 236065
rect 531286 232719 531338 232725
rect 531286 232661 531338 232667
rect 528310 229611 528362 229617
rect 528310 229553 528362 229559
rect 528502 229611 528554 229617
rect 528502 229553 528554 229559
rect 528322 221496 528350 229553
rect 529750 228723 529802 228729
rect 529750 228665 529802 228671
rect 528980 224322 529036 224331
rect 528980 224257 529036 224266
rect 528288 221468 528350 221496
rect 528994 221496 529022 224257
rect 528994 221468 529056 221496
rect 529762 221482 529790 228665
rect 530516 224026 530572 224035
rect 530516 223961 530572 223970
rect 530530 221496 530558 223961
rect 530496 221468 530558 221496
rect 531298 221482 531326 232661
rect 532052 224174 532108 224183
rect 532052 224109 532108 224118
rect 532066 221482 532094 224109
rect 532834 221792 532862 239173
rect 538004 238086 538060 238095
rect 538004 238021 538060 238030
rect 535126 237751 535178 237757
rect 535126 237693 535178 237699
rect 533494 237677 533546 237683
rect 533494 237619 533546 237625
rect 532786 221764 532862 221792
rect 532786 221482 532814 221764
rect 533506 221482 533534 237619
rect 534260 230094 534316 230103
rect 534260 230029 534316 230038
rect 534274 221482 534302 230029
rect 535138 221792 535166 237693
rect 535798 237603 535850 237609
rect 535798 237545 535850 237551
rect 535810 228581 535838 237545
rect 538018 236174 538046 238021
rect 537922 236146 538046 236174
rect 541474 236174 541502 240093
rect 544340 238382 544396 238391
rect 544340 238317 544396 238326
rect 541474 236146 541790 236174
rect 537238 232645 537290 232651
rect 537238 232587 537290 232593
rect 535798 228575 535850 228581
rect 535798 228517 535850 228523
rect 535798 228427 535850 228433
rect 535798 228369 535850 228375
rect 535090 221764 535166 221792
rect 535090 221482 535118 221764
rect 535810 221482 535838 228369
rect 536564 223878 536620 223887
rect 536564 223813 536620 223822
rect 536578 221482 536606 223813
rect 537250 221792 537278 232587
rect 537922 228433 537950 236146
rect 539542 232571 539594 232577
rect 539542 232513 539594 232519
rect 538868 229798 538924 229807
rect 538868 229733 538924 229742
rect 538006 228575 538058 228581
rect 538006 228517 538058 228523
rect 537910 228427 537962 228433
rect 537910 228369 537962 228375
rect 537250 221764 537326 221792
rect 537298 221482 537326 221764
rect 538018 221482 538046 228517
rect 538882 221482 538910 229733
rect 539554 221792 539582 232513
rect 540310 229463 540362 229469
rect 540310 229405 540362 229411
rect 539554 221764 539630 221792
rect 539602 221482 539630 221764
rect 540322 221482 540350 229405
rect 541076 222842 541132 222851
rect 541076 222777 541132 222786
rect 541090 221482 541118 222777
rect 541762 221792 541790 236146
rect 543382 232497 543434 232503
rect 543382 232439 543434 232445
rect 542614 232423 542666 232429
rect 542614 232365 542666 232371
rect 541762 221764 541838 221792
rect 541810 221482 541838 221764
rect 542626 221482 542654 232365
rect 543394 221482 543422 232439
rect 544354 228581 544382 238317
rect 544342 228575 544394 228581
rect 544342 228517 544394 228523
rect 544052 223730 544108 223739
rect 544052 223665 544108 223674
rect 544066 221792 544094 223665
rect 544066 221764 544142 221792
rect 544114 221482 544142 221764
rect 544834 221482 544862 240241
rect 550868 240010 550924 240019
rect 550868 239945 550924 239954
rect 550196 238678 550252 238687
rect 550196 238613 550252 238622
rect 549430 232349 549482 232355
rect 549430 232291 549482 232297
rect 545590 232201 545642 232207
rect 545590 232143 545642 232149
rect 545602 221482 545630 232143
rect 548566 232127 548618 232133
rect 548566 232069 548618 232075
rect 546358 229389 546410 229395
rect 546358 229331 546410 229337
rect 546370 221792 546398 229331
rect 547894 228797 547946 228803
rect 547894 228739 547946 228745
rect 547126 228575 547178 228581
rect 547126 228517 547178 228523
rect 546370 221764 546446 221792
rect 546418 221482 546446 221764
rect 547138 221482 547166 228517
rect 547906 221482 547934 228739
rect 548578 221792 548606 232069
rect 548578 221764 548654 221792
rect 548626 221482 548654 221764
rect 549442 221482 549470 232291
rect 550210 221482 550238 238613
rect 550882 221792 550910 239945
rect 553940 238974 553996 238983
rect 553940 238909 553996 238918
rect 553954 236174 553982 238909
rect 559892 238234 559948 238243
rect 559892 238169 559948 238178
rect 559220 236606 559276 236615
rect 559220 236541 559276 236550
rect 557684 236458 557740 236467
rect 557684 236393 557740 236402
rect 553282 236146 553982 236174
rect 551636 232758 551692 232767
rect 551636 232693 551692 232702
rect 550882 221764 550958 221792
rect 550930 221482 550958 221764
rect 551650 221482 551678 232693
rect 552406 232275 552458 232281
rect 552406 232217 552458 232223
rect 552418 221482 552446 232217
rect 553282 221792 553310 236146
rect 557014 233015 557066 233021
rect 557014 232957 557066 232963
rect 554710 231979 554762 231985
rect 554710 231921 554762 231927
rect 553940 229650 553996 229659
rect 553940 229585 553996 229594
rect 553234 221764 553310 221792
rect 553234 221482 553262 221764
rect 553954 221482 553982 229585
rect 554722 221482 554750 231921
rect 555382 229315 555434 229321
rect 555382 229257 555434 229263
rect 555394 221792 555422 229257
rect 556150 228575 556202 228581
rect 556150 228517 556202 228523
rect 555394 221764 555470 221792
rect 555442 221482 555470 221764
rect 556162 221482 556190 228517
rect 557026 221496 557054 232957
rect 557590 231905 557642 231911
rect 557590 231847 557642 231853
rect 557602 221792 557630 231847
rect 557698 228581 557726 236393
rect 558454 232053 558506 232059
rect 558454 231995 558506 232001
rect 557686 228575 557738 228581
rect 557686 228517 557738 228523
rect 557602 221764 557726 221792
rect 556992 221468 557054 221496
rect 557698 221496 557726 221764
rect 557698 221468 557760 221496
rect 558466 221482 558494 231995
rect 559234 221496 559262 236541
rect 559200 221468 559262 221496
rect 559906 221496 559934 238169
rect 566036 236902 566092 236911
rect 566036 236837 566092 236846
rect 562196 236754 562252 236763
rect 562196 236689 562252 236698
rect 560756 232610 560812 232619
rect 560756 232545 560812 232554
rect 559906 221468 559968 221496
rect 560770 221482 560798 232545
rect 561430 229241 561482 229247
rect 561430 229183 561482 229189
rect 561442 221792 561470 229183
rect 561442 221764 561518 221792
rect 561490 221482 561518 221764
rect 562210 221482 562238 236689
rect 566050 236174 566078 236837
rect 565282 236146 566078 236174
rect 564500 232462 564556 232471
rect 564500 232397 564556 232406
rect 563638 229167 563690 229173
rect 563638 229109 563690 229115
rect 562964 223582 563020 223591
rect 562964 223517 563020 223526
rect 562978 221482 563006 223517
rect 563650 221792 563678 229109
rect 563650 221764 563726 221792
rect 563698 221482 563726 221764
rect 564514 221482 564542 232397
rect 565282 221482 565310 236146
rect 565942 229833 565994 229839
rect 565942 229775 565994 229781
rect 565954 221792 565982 229775
rect 565954 221764 566030 221792
rect 566002 221482 566030 221764
rect 566722 221482 566750 240685
rect 567394 228581 567422 241425
rect 581780 240898 581836 240907
rect 581780 240833 581836 240842
rect 573140 237050 573196 237059
rect 573140 236985 573196 236994
rect 573154 236174 573182 236985
rect 573154 236146 574334 236174
rect 572086 232867 572138 232873
rect 572086 232809 572138 232815
rect 570452 232314 570508 232323
rect 570452 232249 570508 232258
rect 567478 229093 567530 229099
rect 567478 229035 567530 229041
rect 567382 228575 567434 228581
rect 567382 228517 567434 228523
rect 567490 221482 567518 229035
rect 569782 229019 569834 229025
rect 569782 228961 569834 228967
rect 569014 228575 569066 228581
rect 569014 228517 569066 228523
rect 568244 223286 568300 223295
rect 568244 223221 568300 223230
rect 568258 221792 568286 223221
rect 568258 221764 568334 221792
rect 568306 221482 568334 221764
rect 569026 221482 569054 228517
rect 569794 221482 569822 228961
rect 570466 221792 570494 232249
rect 571316 223434 571372 223443
rect 571316 223369 571372 223378
rect 570466 221764 570542 221792
rect 570514 221482 570542 221764
rect 571330 221482 571358 223369
rect 572098 221482 572126 232809
rect 573524 229502 573580 229511
rect 573524 229437 573580 229446
rect 572756 229354 572812 229363
rect 572756 229289 572812 229298
rect 572770 221792 572798 229289
rect 572770 221764 572846 221792
rect 572818 221482 572846 221764
rect 573538 221482 573566 229437
rect 574306 221482 574334 236146
rect 580340 235570 580396 235579
rect 580340 235505 580396 235514
rect 576596 232166 576652 232175
rect 576596 232101 576652 232110
rect 575828 231870 575884 231879
rect 575828 231805 575884 231814
rect 575062 229537 575114 229543
rect 575062 229479 575114 229485
rect 575074 221792 575102 229479
rect 575074 221764 575150 221792
rect 575122 221482 575150 221764
rect 575842 221482 575870 231805
rect 576610 221482 576638 232101
rect 578036 232018 578092 232027
rect 578036 231953 578092 231962
rect 577268 223138 577324 223147
rect 577268 223073 577324 223082
rect 577282 221792 577310 223073
rect 577282 221764 577358 221792
rect 577330 221482 577358 221764
rect 578050 221482 578078 231953
rect 578900 229206 578956 229215
rect 578900 229141 578956 229150
rect 578914 221482 578942 229141
rect 579574 225837 579626 225843
rect 579574 225779 579626 225785
rect 579586 221792 579614 225779
rect 579586 221764 579662 221792
rect 579634 221482 579662 221764
rect 580354 221482 580382 235505
rect 581110 225763 581162 225769
rect 581110 225705 581162 225711
rect 581122 221482 581150 225705
rect 581794 221792 581822 240833
rect 599062 239157 599114 239163
rect 599062 239099 599114 239105
rect 593012 236162 593068 236171
rect 593012 236097 593068 236106
rect 591476 235866 591532 235875
rect 591476 235801 591532 235810
rect 588982 235531 589034 235537
rect 588982 235473 589034 235479
rect 588694 235457 588746 235463
rect 588694 235399 588746 235405
rect 583412 235274 583468 235283
rect 583412 235209 583468 235218
rect 587926 235235 587978 235241
rect 582646 226059 582698 226065
rect 582646 226001 582698 226007
rect 581794 221764 581870 221792
rect 581842 221482 581870 221764
rect 582658 221482 582686 226001
rect 583426 221482 583454 235209
rect 587926 235177 587978 235183
rect 585622 227391 585674 227397
rect 585622 227333 585674 227339
rect 584854 227169 584906 227175
rect 584854 227111 584906 227117
rect 584086 225985 584138 225991
rect 584086 225927 584138 225933
rect 584098 221792 584126 225927
rect 584098 221764 584174 221792
rect 584146 221482 584174 221764
rect 584866 221482 584894 227111
rect 585634 221482 585662 227333
rect 587158 225911 587210 225917
rect 587158 225853 587210 225859
rect 586390 225689 586442 225695
rect 586390 225631 586442 225637
rect 586402 221496 586430 225631
rect 586402 221468 586464 221496
rect 587170 221482 587198 225853
rect 587938 221496 587966 235177
rect 588598 227539 588650 227545
rect 588598 227481 588650 227487
rect 587904 221468 587966 221496
rect 588610 221496 588638 227481
rect 588706 225917 588734 235399
rect 588886 235309 588938 235315
rect 588886 235251 588938 235257
rect 588898 226657 588926 235251
rect 588886 226651 588938 226657
rect 588886 226593 588938 226599
rect 588694 225911 588746 225917
rect 588694 225853 588746 225859
rect 588994 225769 589022 235473
rect 590422 235383 590474 235389
rect 590422 235325 590474 235331
rect 590134 227465 590186 227471
rect 590134 227407 590186 227413
rect 588982 225763 589034 225769
rect 588982 225705 589034 225711
rect 589366 224727 589418 224733
rect 589366 224669 589418 224675
rect 588610 221468 588672 221496
rect 589378 221482 589406 224669
rect 590146 221792 590174 227407
rect 590434 225991 590462 235325
rect 590902 227021 590954 227027
rect 590902 226963 590954 226969
rect 590422 225985 590474 225991
rect 590422 225927 590474 225933
rect 590146 221764 590222 221792
rect 590194 221482 590222 221764
rect 590914 221482 590942 226963
rect 591490 226065 591518 235801
rect 592342 235161 592394 235167
rect 592342 235103 592394 235109
rect 591668 226690 591724 226699
rect 591668 226625 591724 226634
rect 591478 226059 591530 226065
rect 591478 226001 591530 226007
rect 591682 221482 591710 226625
rect 592354 221792 592382 235103
rect 593026 227471 593054 236097
rect 595892 236014 595948 236023
rect 595892 235949 595948 235958
rect 595412 235126 595468 235135
rect 595412 235061 595468 235070
rect 594644 234978 594700 234987
rect 594644 234913 594700 234922
rect 593014 227465 593066 227471
rect 593014 227407 593066 227413
rect 593110 227317 593162 227323
rect 593110 227259 593162 227265
rect 592354 221764 592430 221792
rect 592402 221482 592430 221764
rect 593122 221482 593150 227259
rect 593974 227095 594026 227101
rect 593974 227037 594026 227043
rect 593986 221482 594014 227037
rect 594658 221792 594686 234913
rect 594658 221764 594734 221792
rect 594706 221482 594734 221764
rect 595426 221482 595454 235061
rect 595906 227397 595934 235949
rect 597428 235718 597484 235727
rect 597428 235653 597484 235662
rect 596180 235422 596236 235431
rect 596180 235357 596236 235366
rect 596194 227545 596222 235357
rect 596182 227539 596234 227545
rect 596182 227481 596234 227487
rect 595894 227391 595946 227397
rect 595894 227333 595946 227339
rect 597442 227323 597470 235653
rect 597718 235087 597770 235093
rect 597718 235029 597770 235035
rect 597430 227317 597482 227323
rect 597430 227259 597482 227265
rect 596948 226542 597004 226551
rect 596948 226477 597004 226486
rect 596180 226394 596236 226403
rect 596180 226329 596236 226338
rect 596194 221482 596222 226329
rect 596962 221792 596990 226477
rect 596962 221764 597038 221792
rect 597010 221482 597038 221764
rect 597730 221482 597758 235029
rect 599074 227101 599102 239099
rect 599924 229058 599980 229067
rect 599924 228993 599980 229002
rect 599062 227095 599114 227101
rect 599062 227037 599114 227043
rect 599158 226873 599210 226879
rect 599158 226815 599210 226821
rect 598486 225911 598538 225917
rect 598486 225853 598538 225859
rect 598498 221482 598526 225853
rect 599170 221792 599198 226815
rect 599170 221764 599246 221792
rect 599218 221482 599246 221764
rect 599938 221482 599966 228993
rect 600418 226879 600446 241911
rect 601462 230203 601514 230209
rect 601462 230145 601514 230151
rect 600406 226873 600458 226879
rect 600406 226815 600458 226821
rect 600790 226651 600842 226657
rect 600790 226593 600842 226599
rect 600802 221482 600830 226593
rect 601474 221792 601502 230145
rect 603298 226805 603326 253455
rect 603382 250627 603434 250633
rect 603382 250569 603434 250575
rect 603394 226953 603422 250569
rect 603478 247815 603530 247821
rect 603478 247757 603530 247763
rect 603490 227249 603518 247757
rect 604534 231831 604586 231837
rect 604534 231773 604586 231779
rect 603478 227243 603530 227249
rect 603478 227185 603530 227191
rect 603670 227021 603722 227027
rect 603670 226963 603722 226969
rect 603382 226947 603434 226953
rect 603382 226889 603434 226895
rect 602998 226799 603050 226805
rect 602998 226741 603050 226747
rect 603286 226799 603338 226805
rect 603286 226741 603338 226747
rect 602230 225763 602282 225769
rect 602230 225705 602282 225711
rect 601474 221764 601550 221792
rect 601522 221482 601550 221764
rect 602242 221482 602270 225705
rect 603010 221482 603038 226741
rect 603682 221792 603710 226963
rect 603682 221764 603758 221792
rect 603730 221482 603758 221764
rect 604546 221482 604574 231773
rect 605974 229759 606026 229765
rect 605974 229701 606026 229707
rect 605302 225911 605354 225917
rect 605302 225853 605354 225859
rect 605314 221482 605342 225853
rect 605986 221792 606014 229701
rect 606178 226657 606206 262113
rect 606262 259285 606314 259291
rect 606262 259227 606314 259233
rect 606274 227027 606302 259227
rect 606358 256399 606410 256405
rect 606358 256341 606410 256347
rect 606370 227175 606398 256341
rect 629206 247741 629258 247747
rect 629206 247683 629258 247689
rect 610484 240602 610540 240611
rect 610484 240537 610540 240546
rect 609046 230129 609098 230135
rect 609046 230071 609098 230077
rect 607508 228910 607564 228919
rect 607508 228845 607564 228854
rect 606358 227169 606410 227175
rect 606358 227111 606410 227117
rect 606262 227021 606314 227027
rect 606262 226963 606314 226969
rect 606166 226651 606218 226657
rect 606166 226593 606218 226599
rect 606742 225245 606794 225251
rect 606742 225187 606794 225193
rect 605986 221764 606062 221792
rect 606034 221482 606062 221764
rect 606754 221482 606782 225187
rect 607522 221482 607550 228845
rect 608278 226059 608330 226065
rect 608278 226001 608330 226007
rect 608290 221792 608318 226001
rect 608290 221764 608366 221792
rect 608338 221482 608366 221764
rect 609058 221482 609086 230071
rect 609814 226725 609866 226731
rect 609814 226667 609866 226673
rect 609826 221482 609854 226667
rect 610498 221792 610526 240537
rect 627188 240454 627244 240463
rect 627188 240389 627244 240398
rect 621140 236310 621196 236319
rect 621140 236245 621196 236254
rect 615862 235013 615914 235019
rect 615862 234955 615914 234961
rect 614998 231757 615050 231763
rect 614998 231699 615050 231705
rect 612118 230055 612170 230061
rect 612118 229997 612170 230003
rect 611254 227465 611306 227471
rect 611254 227407 611306 227413
rect 610498 221764 610574 221792
rect 610546 221482 610574 221764
rect 611266 221482 611294 227407
rect 612130 221482 612158 229997
rect 614326 227391 614378 227397
rect 614326 227333 614378 227339
rect 612790 226577 612842 226583
rect 612790 226519 612842 226525
rect 612802 221792 612830 226519
rect 613558 226429 613610 226435
rect 613558 226371 613610 226377
rect 612802 221764 612878 221792
rect 612850 221482 612878 221764
rect 613570 221482 613598 226371
rect 614338 221482 614366 227333
rect 615010 221792 615038 231699
rect 615010 221764 615086 221792
rect 615058 221482 615086 221764
rect 615874 221482 615902 234955
rect 618836 234830 618892 234839
rect 618836 234765 618892 234774
rect 616630 227539 616682 227545
rect 616630 227481 616682 227487
rect 616642 221496 616670 227481
rect 617302 226503 617354 226509
rect 617302 226445 617354 226451
rect 616608 221468 616670 221496
rect 617314 221496 617342 226445
rect 618070 226355 618122 226361
rect 618070 226297 618122 226303
rect 617314 221468 617376 221496
rect 618082 221482 618110 226297
rect 618850 221792 618878 234765
rect 619606 227317 619658 227323
rect 619606 227259 619658 227265
rect 618850 221764 618926 221792
rect 618898 221482 618926 221764
rect 619618 221482 619646 227259
rect 620372 226246 620428 226255
rect 620372 226181 620428 226190
rect 620386 221482 620414 226181
rect 621154 221792 621182 236245
rect 621814 234939 621866 234945
rect 621814 234881 621866 234887
rect 621106 221764 621182 221792
rect 621106 221482 621134 221764
rect 621826 221482 621854 234881
rect 624884 234682 624940 234691
rect 624884 234617 624940 234626
rect 622678 233237 622730 233243
rect 622678 233179 622730 233185
rect 622690 221482 622718 233179
rect 624118 226281 624170 226287
rect 624118 226223 624170 226229
rect 623348 226098 623404 226107
rect 623348 226033 623404 226042
rect 623362 221792 623390 226033
rect 623362 221764 623438 221792
rect 623410 221482 623438 221764
rect 624130 221482 624158 226223
rect 624898 221482 624926 234617
rect 626422 232793 626474 232799
rect 626422 232735 626474 232741
rect 625558 229907 625610 229913
rect 625558 229849 625610 229855
rect 625570 221792 625598 229849
rect 625570 221764 625646 221792
rect 625618 221482 625646 221764
rect 626434 221482 626462 232735
rect 627202 221482 627230 240389
rect 627862 234865 627914 234871
rect 627862 234807 627914 234813
rect 627874 221792 627902 234807
rect 628630 229611 628682 229617
rect 628630 229553 628682 229559
rect 627874 221764 627950 221792
rect 627922 221482 627950 221764
rect 628642 221482 628670 229553
rect 629218 226435 629246 247683
rect 629302 244855 629354 244861
rect 629302 244797 629354 244803
rect 629314 227545 629342 244797
rect 632374 234791 632426 234797
rect 632374 234733 632426 234739
rect 630934 234717 630986 234723
rect 630934 234659 630986 234665
rect 630166 229685 630218 229691
rect 630166 229627 630218 229633
rect 629302 227539 629354 227545
rect 629302 227481 629354 227487
rect 629206 226429 629258 226435
rect 629206 226371 629258 226377
rect 629398 225171 629450 225177
rect 629398 225113 629450 225119
rect 629410 221482 629438 225113
rect 630178 221792 630206 229627
rect 630178 221764 630254 221792
rect 630226 221482 630254 221764
rect 630946 221482 630974 234659
rect 631702 226133 631754 226139
rect 631702 226075 631754 226081
rect 631714 221482 631742 226075
rect 632386 221792 632414 234733
rect 634006 227539 634058 227545
rect 634006 227481 634058 227487
rect 633142 227095 633194 227101
rect 633142 227037 633194 227043
rect 632386 221764 632462 221792
rect 632434 221482 632462 221764
rect 633154 221482 633182 227037
rect 634018 221482 634046 227481
rect 636214 227243 636266 227249
rect 636214 227185 636266 227191
rect 634678 226873 634730 226879
rect 634678 226815 634730 226821
rect 634690 221792 634718 226815
rect 635446 226429 635498 226435
rect 635446 226371 635498 226377
rect 634690 221764 634766 221792
rect 634738 221482 634766 221764
rect 635458 221482 635486 226371
rect 636226 221482 636254 227185
rect 638518 227169 638570 227175
rect 638518 227111 638570 227117
rect 636886 226947 636938 226953
rect 636886 226889 636938 226895
rect 636898 221792 636926 226889
rect 637750 226799 637802 226805
rect 637750 226741 637802 226747
rect 636898 221764 636974 221792
rect 636946 221482 636974 221764
rect 637762 221482 637790 226741
rect 638530 221482 638558 227111
rect 639190 227021 639242 227027
rect 639190 226963 639242 226969
rect 639202 221792 639230 226963
rect 639958 226651 640010 226657
rect 639958 226593 640010 226599
rect 639202 221764 639278 221792
rect 639250 221482 639278 221764
rect 639970 221482 639998 226593
rect 640148 212334 640204 212343
rect 640148 212269 640204 212278
rect 640162 211603 640190 212269
rect 640148 211594 640204 211603
rect 640148 211529 640204 211538
rect 190292 201382 190348 201391
rect 190292 201317 190348 201326
rect 190306 200577 190334 201317
rect 640148 200938 640204 200947
rect 640148 200873 640204 200882
rect 190292 200568 190348 200577
rect 190292 200503 190348 200512
rect 640162 200207 640190 200873
rect 640148 200198 640204 200207
rect 640148 200133 640204 200142
rect 187220 199162 187276 199171
rect 187220 199097 187276 199106
rect 185890 195826 186302 195854
rect 186070 185803 186122 185809
rect 186070 185745 186122 185751
rect 185974 182991 186026 182997
rect 185974 182933 186026 182939
rect 185780 182438 185836 182447
rect 185780 182373 185836 182382
rect 185602 175666 185726 175694
rect 185602 173271 185630 175666
rect 185588 173262 185644 173271
rect 185588 173197 185644 173206
rect 185986 136863 186014 182933
rect 186082 138343 186110 185745
rect 186166 182917 186218 182923
rect 186166 182859 186218 182865
rect 186068 138334 186124 138343
rect 186068 138269 186124 138278
rect 186178 137455 186206 182859
rect 186274 174751 186302 195826
rect 640244 185694 640300 185703
rect 640244 185629 640300 185638
rect 640258 184963 640286 185629
rect 640244 184954 640300 184963
rect 640244 184889 640300 184898
rect 645142 183139 645194 183145
rect 645142 183081 645194 183087
rect 645154 183039 645182 183081
rect 645140 183030 645196 183039
rect 645140 182965 645196 182974
rect 645142 179439 645194 179445
rect 645142 179381 645194 179387
rect 645154 179339 645182 179381
rect 645140 179330 645196 179339
rect 645140 179265 645196 179274
rect 186742 178403 186794 178409
rect 186742 178345 186794 178351
rect 186754 177711 186782 178345
rect 186740 177702 186796 177711
rect 186740 177637 186796 177646
rect 645142 174925 645194 174931
rect 645140 174890 645142 174899
rect 645194 174890 645196 174899
rect 645140 174825 645196 174834
rect 186260 174742 186316 174751
rect 186260 174677 186316 174686
rect 186262 174259 186314 174265
rect 186262 174201 186314 174207
rect 186164 137446 186220 137455
rect 186164 137381 186220 137390
rect 185972 136854 186028 136863
rect 185972 136789 186028 136798
rect 185492 135966 185548 135975
rect 185492 135901 185548 135910
rect 184534 135335 184586 135341
rect 184534 135277 184586 135283
rect 184438 135261 184490 135267
rect 184438 135203 184490 135209
rect 184342 135187 184394 135193
rect 184342 135129 184394 135135
rect 184354 134495 184382 135129
rect 184340 134486 184396 134495
rect 184340 134421 184396 134430
rect 184450 133755 184478 135203
rect 184436 133746 184492 133755
rect 184436 133681 184492 133690
rect 184546 133015 184574 135277
rect 186274 135235 186302 174201
rect 645142 171077 645194 171083
rect 645140 171042 645142 171051
rect 645194 171042 645196 171051
rect 645140 170977 645196 170986
rect 645142 168265 645194 168271
rect 645142 168207 645194 168213
rect 645154 167795 645182 168207
rect 645140 167786 645196 167795
rect 645140 167721 645196 167730
rect 645142 163381 645194 163387
rect 645140 163346 645142 163355
rect 645194 163346 645196 163355
rect 645140 163281 645196 163290
rect 645142 159755 645194 159761
rect 645142 159697 645194 159703
rect 645154 159507 645182 159697
rect 645140 159498 645196 159507
rect 645140 159433 645196 159442
rect 645142 156055 645194 156061
rect 645142 155997 645194 156003
rect 645154 155511 645182 155997
rect 645140 155502 645196 155511
rect 645140 155437 645196 155446
rect 645142 152577 645194 152583
rect 645140 152542 645142 152551
rect 645194 152542 645196 152551
rect 645140 152477 645196 152486
rect 645142 148211 645194 148217
rect 645142 148153 645194 148159
rect 645154 148111 645182 148153
rect 645140 148102 645196 148111
rect 645140 148037 645196 148046
rect 186742 146879 186794 146885
rect 186742 146821 186794 146827
rect 186754 145891 186782 146821
rect 186740 145882 186796 145891
rect 186740 145817 186796 145826
rect 186260 135226 186316 135235
rect 186260 135161 186316 135170
rect 185686 134003 185738 134009
rect 185686 133945 185738 133951
rect 185590 133929 185642 133935
rect 185590 133871 185642 133877
rect 184532 133006 184588 133015
rect 184532 132941 184588 132950
rect 183094 132449 183146 132455
rect 183094 132391 183146 132397
rect 184630 132449 184682 132455
rect 184630 132391 184682 132397
rect 184534 132375 184586 132381
rect 184534 132317 184586 132323
rect 184342 132301 184394 132307
rect 184342 132243 184394 132249
rect 184354 131535 184382 132243
rect 184438 132227 184490 132233
rect 184438 132169 184490 132175
rect 184340 131526 184396 131535
rect 184340 131461 184396 131470
rect 184450 129907 184478 132169
rect 184546 130647 184574 132317
rect 184642 132275 184670 132391
rect 184628 132266 184684 132275
rect 184628 132201 184684 132210
rect 184532 130638 184588 130647
rect 184532 130573 184588 130582
rect 184436 129898 184492 129907
rect 184436 129833 184492 129842
rect 184630 129563 184682 129569
rect 184630 129505 184682 129511
rect 184438 129489 184490 129495
rect 184438 129431 184490 129437
rect 184342 129341 184394 129347
rect 184342 129283 184394 129289
rect 184354 129167 184382 129283
rect 184340 129158 184396 129167
rect 184340 129093 184396 129102
rect 184450 128427 184478 129431
rect 184534 129415 184586 129421
rect 184534 129357 184586 129363
rect 184436 128418 184492 128427
rect 184436 128353 184492 128362
rect 184546 127687 184574 129357
rect 184532 127678 184588 127687
rect 184532 127613 184588 127622
rect 184642 126947 184670 129505
rect 184628 126938 184684 126947
rect 184628 126873 184684 126882
rect 184438 126677 184490 126683
rect 184438 126619 184490 126625
rect 184342 126529 184394 126535
rect 184342 126471 184394 126477
rect 184354 125467 184382 126471
rect 184450 126059 184478 126619
rect 184534 126603 184586 126609
rect 184534 126545 184586 126551
rect 184436 126050 184492 126059
rect 184436 125985 184492 125994
rect 184340 125458 184396 125467
rect 184340 125393 184396 125402
rect 184546 124579 184574 126545
rect 184532 124570 184588 124579
rect 184532 124505 184588 124514
rect 184342 123865 184394 123871
rect 184340 123830 184342 123839
rect 184394 123830 184396 123839
rect 184340 123765 184396 123774
rect 184438 123791 184490 123797
rect 184438 123733 184490 123739
rect 184342 123717 184394 123723
rect 184342 123659 184394 123665
rect 184354 122211 184382 123659
rect 184450 123099 184478 123733
rect 184534 123643 184586 123649
rect 184534 123585 184586 123591
rect 184436 123090 184492 123099
rect 184436 123025 184492 123034
rect 184340 122202 184396 122211
rect 184340 122137 184396 122146
rect 184546 121619 184574 123585
rect 184532 121610 184588 121619
rect 184532 121545 184588 121554
rect 184438 120979 184490 120985
rect 184438 120921 184490 120927
rect 184342 120757 184394 120763
rect 184450 120731 184478 120921
rect 184534 120905 184586 120911
rect 184534 120847 184586 120853
rect 184342 120699 184394 120705
rect 184436 120722 184492 120731
rect 184354 119251 184382 120699
rect 184436 120657 184492 120666
rect 184546 120139 184574 120847
rect 184630 120831 184682 120837
rect 184630 120773 184682 120779
rect 184532 120130 184588 120139
rect 184532 120065 184588 120074
rect 184340 119242 184396 119251
rect 184340 119177 184396 119186
rect 184642 118659 184670 120773
rect 184628 118650 184684 118659
rect 184628 118585 184684 118594
rect 182902 118167 182954 118173
rect 182902 118109 182954 118115
rect 182806 112321 182858 112327
rect 182806 112263 182858 112269
rect 180022 112247 180074 112253
rect 180022 112189 180074 112195
rect 180022 95079 180074 95085
rect 180022 95021 180074 95027
rect 179926 94635 179978 94641
rect 179926 94577 179978 94583
rect 168406 83461 168458 83467
rect 168406 83403 168458 83409
rect 162358 80501 162410 80507
rect 162358 80443 162410 80449
rect 180034 80433 180062 95021
rect 182914 94715 182942 118109
rect 184630 118093 184682 118099
rect 184630 118035 184682 118041
rect 184534 118019 184586 118025
rect 184534 117961 184586 117967
rect 184438 117945 184490 117951
rect 184438 117887 184490 117893
rect 184342 117871 184394 117877
rect 184342 117813 184394 117819
rect 184354 117771 184382 117813
rect 184340 117762 184396 117771
rect 184340 117697 184396 117706
rect 184450 117031 184478 117887
rect 184436 117022 184492 117031
rect 184436 116957 184492 116966
rect 184546 116291 184574 117961
rect 184532 116282 184588 116291
rect 184532 116217 184588 116226
rect 184642 115403 184670 118035
rect 184628 115394 184684 115403
rect 184628 115329 184684 115338
rect 184534 115207 184586 115213
rect 184534 115149 184586 115155
rect 184438 115133 184490 115139
rect 184438 115075 184490 115081
rect 184342 115059 184394 115065
rect 184342 115001 184394 115007
rect 184354 114811 184382 115001
rect 184340 114802 184396 114811
rect 184340 114737 184396 114746
rect 184450 113923 184478 115075
rect 184436 113914 184492 113923
rect 184436 113849 184492 113858
rect 184546 113183 184574 115149
rect 184532 113174 184588 113183
rect 184532 113109 184588 113118
rect 184342 112321 184394 112327
rect 184342 112263 184394 112269
rect 184354 111703 184382 112263
rect 184438 112247 184490 112253
rect 184438 112189 184490 112195
rect 184340 111694 184396 111703
rect 184340 111629 184396 111638
rect 184450 110963 184478 112189
rect 184534 112173 184586 112179
rect 184534 112115 184586 112121
rect 184436 110954 184492 110963
rect 184436 110889 184492 110898
rect 184546 110223 184574 112115
rect 184532 110214 184588 110223
rect 184532 110149 184588 110158
rect 184342 109435 184394 109441
rect 184342 109377 184394 109383
rect 184354 107115 184382 109377
rect 184438 109361 184490 109367
rect 184436 109326 184438 109335
rect 184490 109326 184492 109335
rect 184436 109261 184492 109270
rect 185602 108743 185630 133871
rect 185698 112443 185726 133945
rect 645718 129637 645770 129643
rect 645718 129579 645770 129585
rect 645730 129019 645758 129579
rect 645716 129010 645772 129019
rect 645716 128945 645772 128954
rect 646498 126905 646526 275317
rect 647362 269323 647390 278018
rect 648610 272135 648638 278018
rect 648596 272126 648652 272135
rect 648596 272061 648652 272070
rect 647348 269314 647404 269323
rect 647348 269249 647404 269258
rect 646580 267390 646636 267399
rect 646580 267325 646636 267334
rect 646486 126899 646538 126905
rect 646486 126841 646538 126847
rect 186166 123569 186218 123575
rect 186166 123511 186218 123517
rect 185684 112434 185740 112443
rect 185684 112369 185740 112378
rect 185588 108734 185644 108743
rect 185588 108669 185644 108678
rect 186178 107855 186206 123511
rect 646498 122063 646526 126841
rect 646594 126831 646622 267325
rect 646678 253513 646730 253519
rect 646678 253455 646730 253461
rect 646690 144263 646718 253455
rect 646774 207411 646826 207417
rect 646774 207353 646826 207359
rect 646676 144254 646732 144263
rect 646676 144189 646732 144198
rect 646786 141007 646814 207353
rect 649378 183145 649406 861106
rect 655222 792085 655274 792091
rect 655222 792027 655274 792033
rect 655030 783501 655082 783507
rect 655030 783443 655082 783449
rect 654358 780541 654410 780547
rect 654358 780483 654410 780489
rect 654370 773559 654398 780483
rect 655042 774743 655070 783443
rect 655124 777694 655180 777703
rect 655124 777629 655180 777638
rect 655028 774734 655084 774743
rect 655028 774669 655084 774678
rect 654356 773550 654412 773559
rect 654356 773485 654412 773494
rect 654070 737473 654122 737479
rect 654070 737415 654122 737421
rect 654082 728567 654110 737415
rect 654166 737399 654218 737405
rect 654166 737341 654218 737347
rect 654178 730195 654206 737341
rect 654164 730186 654220 730195
rect 654164 730121 654220 730130
rect 654068 728558 654124 728567
rect 654068 728493 654124 728502
rect 655138 714465 655166 777629
rect 655234 775779 655262 792027
rect 655412 778286 655468 778295
rect 655412 778221 655468 778230
rect 655220 775770 655276 775779
rect 655220 775705 655276 775714
rect 655316 734478 655372 734487
rect 655316 734413 655372 734422
rect 655220 731666 655276 731675
rect 655220 731601 655276 731610
rect 655126 714459 655178 714465
rect 655126 714401 655178 714407
rect 654358 702841 654410 702847
rect 654358 702783 654410 702789
rect 649462 702767 649514 702773
rect 649462 702709 649514 702715
rect 649366 183139 649418 183145
rect 649366 183081 649418 183087
rect 649474 179445 649502 702709
rect 654166 694331 654218 694337
rect 654166 694273 654218 694279
rect 654070 691371 654122 691377
rect 654070 691313 654122 691319
rect 654082 684611 654110 691313
rect 654178 685351 654206 694273
rect 654370 686979 654398 702783
rect 655124 689486 655180 689495
rect 655124 689421 655180 689430
rect 654356 686970 654412 686979
rect 654356 686905 654412 686914
rect 654164 685342 654220 685351
rect 654164 685277 654220 685286
rect 654068 684602 654124 684611
rect 654068 684537 654124 684546
rect 652246 666803 652298 666809
rect 652246 666745 652298 666751
rect 649750 666729 649802 666735
rect 649750 666671 649802 666677
rect 649558 654075 649610 654081
rect 649558 654017 649610 654023
rect 649462 179439 649514 179445
rect 649462 179381 649514 179387
rect 649570 174931 649598 654017
rect 649654 610711 649706 610717
rect 649654 610653 649706 610659
rect 649558 174925 649610 174931
rect 649558 174867 649610 174873
rect 649666 171083 649694 610653
rect 649762 263403 649790 666671
rect 649846 567421 649898 567427
rect 649846 567363 649898 567369
rect 649748 263394 649804 263403
rect 649748 263329 649804 263338
rect 649654 171077 649706 171083
rect 649654 171019 649706 171025
rect 649858 168271 649886 567363
rect 649942 521319 649994 521325
rect 649942 521261 649994 521267
rect 649846 168265 649898 168271
rect 649846 168207 649898 168213
rect 646870 164417 646922 164423
rect 646870 164359 646922 164365
rect 646772 140998 646828 141007
rect 646772 140933 646828 140942
rect 646582 126825 646634 126831
rect 646582 126767 646634 126773
rect 646594 123839 646622 126767
rect 646882 125763 646910 164359
rect 647062 164343 647114 164349
rect 647062 164285 647114 164291
rect 646966 164269 647018 164275
rect 646966 164211 647018 164217
rect 646978 127687 647006 164211
rect 647074 134791 647102 164285
rect 649954 163387 649982 521261
rect 650038 478177 650090 478183
rect 650038 478119 650090 478125
rect 649942 163381 649994 163387
rect 649942 163323 649994 163329
rect 650050 159761 650078 478119
rect 650134 388859 650186 388865
rect 650134 388801 650186 388807
rect 650038 159755 650090 159761
rect 650038 159697 650090 159703
rect 650146 156061 650174 388801
rect 650230 342757 650282 342763
rect 650230 342699 650282 342705
rect 650134 156055 650186 156061
rect 650134 155997 650186 156003
rect 650242 152583 650270 342699
rect 650326 299763 650378 299769
rect 650326 299705 650378 299711
rect 650230 152577 650282 152583
rect 650230 152519 650282 152525
rect 650338 148217 650366 299705
rect 652258 267251 652286 666745
rect 654166 656739 654218 656745
rect 654166 656681 654218 656687
rect 654178 640655 654206 656681
rect 654164 640646 654220 640655
rect 654164 640581 654220 640590
rect 655138 622261 655166 689421
rect 655234 665477 655262 731601
rect 655330 668215 655358 734413
rect 655426 714613 655454 778221
rect 655604 775918 655660 775927
rect 655604 775853 655660 775862
rect 655508 732702 655564 732711
rect 655508 732637 655564 732646
rect 655414 714607 655466 714613
rect 655414 714549 655466 714555
rect 655412 688450 655468 688459
rect 655412 688385 655468 688394
rect 655318 668209 655370 668215
rect 655318 668151 655370 668157
rect 655222 665471 655274 665477
rect 655222 665413 655274 665419
rect 655316 643014 655372 643023
rect 655316 642949 655372 642958
rect 655126 622255 655178 622261
rect 655126 622197 655178 622203
rect 655126 613523 655178 613529
rect 655126 613465 655178 613471
rect 653782 602053 653834 602059
rect 653782 601995 653834 602001
rect 653794 592999 653822 601995
rect 655138 595367 655166 613465
rect 655220 597874 655276 597883
rect 655220 597809 655276 597818
rect 655124 595358 655180 595367
rect 655124 595293 655180 595302
rect 653780 592990 653836 592999
rect 653780 592925 653836 592934
rect 654166 555877 654218 555883
rect 654166 555819 654218 555825
rect 654178 548599 654206 555819
rect 655124 553326 655180 553335
rect 655124 553261 655180 553270
rect 654164 548590 654220 548599
rect 654164 548525 654220 548534
rect 655138 489801 655166 553261
rect 655234 533017 655262 597809
rect 655330 579045 655358 642949
rect 655426 624999 655454 688385
rect 655522 668437 655550 732637
rect 655618 714761 655646 775853
rect 655702 748869 655754 748875
rect 655702 748811 655754 748817
rect 655714 731379 655742 748811
rect 670774 737547 670826 737553
rect 670774 737489 670826 737495
rect 655700 731370 655756 731379
rect 655700 731305 655756 731314
rect 655606 714755 655658 714761
rect 655606 714697 655658 714703
rect 669718 713127 669770 713133
rect 669718 713069 669770 713075
rect 669526 711943 669578 711949
rect 669526 711885 669578 711891
rect 655604 687118 655660 687127
rect 655604 687053 655660 687062
rect 655510 668431 655562 668437
rect 655510 668373 655562 668379
rect 655508 642422 655564 642431
rect 655508 642357 655564 642366
rect 655414 624993 655466 624999
rect 655414 624935 655466 624941
rect 655412 596690 655468 596699
rect 655412 596625 655468 596634
rect 655318 579039 655370 579045
rect 655318 578981 655370 578987
rect 655316 552142 655372 552151
rect 655316 552077 655372 552086
rect 655222 533011 655274 533017
rect 655222 532953 655274 532959
rect 655330 489949 655358 552077
rect 655426 533165 655454 596625
rect 655522 579193 655550 642357
rect 655618 622409 655646 687053
rect 668758 666803 668810 666809
rect 668758 666745 668810 666751
rect 668770 665551 668798 666745
rect 668758 665545 668810 665551
rect 668758 665487 668810 665493
rect 655798 648303 655850 648309
rect 655798 648245 655850 648251
rect 655700 640794 655756 640803
rect 655700 640729 655756 640738
rect 655606 622403 655658 622409
rect 655606 622345 655658 622351
rect 655604 595506 655660 595515
rect 655604 595441 655660 595450
rect 655510 579187 655562 579193
rect 655510 579129 655562 579135
rect 655508 551106 655564 551115
rect 655508 551041 655564 551050
rect 655414 533159 655466 533165
rect 655414 533101 655466 533107
rect 655522 490097 655550 551041
rect 655618 533313 655646 595441
rect 655714 579341 655742 640729
rect 655810 639175 655838 648245
rect 655990 645195 656042 645201
rect 655990 645137 656042 645143
rect 655796 639166 655852 639175
rect 655796 639101 655852 639110
rect 656002 638287 656030 645137
rect 655988 638278 656044 638287
rect 655988 638213 656044 638222
rect 655798 602127 655850 602133
rect 655798 602069 655850 602075
rect 655810 594183 655838 602069
rect 655796 594174 655852 594183
rect 655796 594109 655852 594118
rect 655702 579335 655754 579341
rect 655702 579277 655754 579283
rect 655702 567495 655754 567501
rect 655702 567437 655754 567443
rect 655714 550967 655742 567437
rect 656566 558837 656618 558843
rect 656566 558779 656618 558785
rect 655700 550958 655756 550967
rect 655700 550893 655756 550902
rect 656578 549783 656606 558779
rect 656564 549774 656620 549783
rect 656564 549709 656620 549718
rect 655606 533307 655658 533313
rect 655606 533249 655658 533255
rect 655510 490091 655562 490097
rect 655510 490033 655562 490039
rect 655318 489943 655370 489949
rect 655318 489885 655370 489891
rect 655126 489795 655178 489801
rect 655126 489737 655178 489743
rect 655126 400625 655178 400631
rect 655126 400567 655178 400573
rect 653782 381681 653834 381687
rect 653782 381623 653834 381629
rect 652342 381607 652394 381613
rect 652342 381549 652394 381555
rect 652354 270909 652382 381549
rect 653794 370999 653822 381623
rect 655138 373367 655166 400567
rect 655510 400551 655562 400557
rect 655510 400493 655562 400499
rect 655318 400477 655370 400483
rect 655318 400419 655370 400425
rect 655124 373358 655180 373367
rect 655124 373293 655180 373302
rect 655330 372183 655358 400419
rect 655522 374403 655550 400493
rect 655508 374394 655564 374403
rect 655508 374329 655564 374338
rect 655316 372174 655372 372183
rect 655316 372109 655372 372118
rect 653780 370990 653836 370999
rect 653780 370925 653836 370934
rect 655126 357187 655178 357193
rect 655126 357129 655178 357135
rect 654166 328327 654218 328333
rect 654166 328269 654218 328275
rect 654178 326303 654206 328269
rect 655138 328079 655166 357129
rect 655318 354375 655370 354381
rect 655318 354317 655370 354323
rect 655222 354301 655274 354307
rect 655222 354243 655274 354249
rect 655234 329855 655262 354243
rect 655220 329846 655276 329855
rect 655220 329781 655276 329790
rect 655124 328070 655180 328079
rect 655124 328005 655180 328014
rect 655330 327487 655358 354317
rect 666646 340685 666698 340691
rect 666646 340627 666698 340633
rect 666658 328333 666686 340627
rect 666646 328327 666698 328333
rect 666646 328269 666698 328275
rect 655316 327478 655372 327487
rect 655316 327413 655372 327422
rect 654164 326294 654220 326303
rect 654164 326229 654220 326238
rect 654262 311233 654314 311239
rect 654262 311175 654314 311181
rect 654166 311159 654218 311165
rect 654166 311101 654218 311107
rect 654070 311085 654122 311091
rect 654070 311027 654122 311033
rect 654082 302179 654110 311027
rect 654178 303363 654206 311101
rect 654164 303354 654220 303363
rect 654164 303289 654220 303298
rect 654068 302170 654124 302179
rect 654068 302105 654124 302114
rect 654274 300995 654302 311175
rect 654260 300986 654316 300995
rect 654260 300921 654316 300930
rect 654164 298766 654220 298775
rect 654164 298701 654220 298710
rect 654178 296703 654206 298701
rect 656468 297582 656524 297591
rect 656468 297517 656524 297526
rect 656084 296842 656140 296851
rect 656084 296777 656140 296786
rect 654164 296694 654220 296703
rect 654164 296629 654220 296638
rect 655892 294030 655948 294039
rect 655892 293965 655948 293974
rect 655796 290922 655852 290931
rect 655796 290857 655852 290866
rect 655604 289294 655660 289303
rect 655604 289229 655660 289238
rect 655412 288110 655468 288119
rect 655412 288045 655468 288054
rect 653780 284558 653836 284567
rect 653780 284493 653836 284502
rect 653794 284155 653822 284493
rect 653782 284149 653834 284155
rect 653782 284091 653834 284097
rect 655124 283374 655180 283383
rect 655124 283309 655180 283318
rect 654260 279822 654316 279831
rect 654260 279757 654316 279766
rect 654274 279493 654302 279757
rect 654262 279487 654314 279493
rect 654262 279429 654314 279435
rect 652342 270903 652394 270909
rect 652342 270845 652394 270851
rect 652244 267242 652300 267251
rect 652244 267177 652300 267186
rect 650326 148211 650378 148217
rect 650326 148153 650378 148159
rect 647060 134782 647116 134791
rect 647060 134717 647116 134726
rect 647828 130934 647884 130943
rect 647828 130869 647884 130878
rect 646964 127678 647020 127687
rect 646964 127613 647020 127622
rect 646868 125754 646924 125763
rect 646868 125689 646924 125698
rect 646580 123830 646636 123839
rect 646580 123765 646636 123774
rect 646484 122054 646540 122063
rect 646484 121989 646540 121998
rect 647842 118395 647870 130869
rect 655138 129865 655166 283309
rect 655316 282338 655372 282347
rect 655316 282273 655372 282282
rect 655220 281006 655276 281015
rect 655220 280941 655276 280950
rect 655234 130013 655262 280941
rect 655330 130161 655358 282273
rect 655426 175893 655454 288045
rect 655508 285742 655564 285751
rect 655508 285677 655564 285686
rect 655522 176041 655550 285677
rect 655618 201571 655646 289229
rect 655700 286926 655756 286935
rect 655700 286861 655756 286870
rect 655606 201565 655658 201571
rect 655606 201507 655658 201513
rect 655714 176189 655742 286861
rect 655810 219109 655838 290857
rect 655906 247673 655934 293965
rect 655988 292846 656044 292855
rect 655988 292781 656044 292790
rect 655894 247667 655946 247673
rect 655894 247609 655946 247615
rect 656002 221921 656030 292781
rect 656098 265137 656126 296777
rect 656180 291662 656236 291671
rect 656180 291597 656236 291606
rect 656086 265131 656138 265137
rect 656086 265073 656138 265079
rect 656194 222069 656222 291597
rect 656482 265285 656510 297517
rect 656564 295214 656620 295223
rect 656564 295149 656620 295158
rect 656578 265433 656606 295149
rect 658006 284149 658058 284155
rect 658006 284091 658058 284097
rect 656566 265427 656618 265433
rect 656566 265369 656618 265375
rect 656470 265279 656522 265285
rect 656470 265221 656522 265227
rect 656182 222063 656234 222069
rect 656182 222005 656234 222011
rect 655990 221915 656042 221921
rect 655990 221857 656042 221863
rect 655798 219103 655850 219109
rect 655798 219045 655850 219051
rect 655702 176183 655754 176189
rect 655702 176125 655754 176131
rect 655510 176035 655562 176041
rect 655510 175977 655562 175983
rect 655414 175887 655466 175893
rect 655414 175829 655466 175835
rect 658018 155543 658046 284091
rect 663766 279487 663818 279493
rect 663766 279429 663818 279435
rect 658006 155537 658058 155543
rect 658006 155479 658058 155485
rect 655318 130155 655370 130161
rect 655318 130097 655370 130103
rect 655222 130007 655274 130013
rect 655222 129949 655274 129955
rect 655126 129859 655178 129865
rect 655126 129801 655178 129807
rect 647924 119538 647980 119547
rect 647924 119473 647980 119482
rect 647830 118389 647882 118395
rect 647830 118331 647882 118337
rect 647938 118247 647966 119473
rect 647926 118241 647978 118247
rect 647926 118183 647978 118189
rect 645238 118167 645290 118173
rect 645238 118109 645290 118115
rect 645250 117623 645278 118109
rect 645236 117614 645292 117623
rect 645236 117549 645292 117558
rect 647924 115690 647980 115699
rect 647924 115625 647980 115634
rect 647938 115287 647966 115625
rect 647926 115281 647978 115287
rect 647926 115223 647978 115229
rect 663778 115213 663806 279429
rect 669538 275095 669566 711885
rect 669622 623217 669674 623223
rect 669622 623159 669674 623165
rect 669524 275086 669580 275095
rect 669524 275021 669580 275030
rect 669634 264915 669662 623159
rect 669730 275243 669758 713069
rect 670678 712683 670730 712689
rect 670678 712625 670730 712631
rect 670582 711573 670634 711579
rect 670582 711515 670634 711521
rect 670390 666063 670442 666069
rect 670390 666005 670442 666011
rect 670402 623223 670430 666005
rect 670594 665551 670622 711515
rect 670690 666735 670718 712625
rect 670678 666729 670730 666735
rect 670678 666671 670730 666677
rect 670582 665545 670634 665551
rect 670582 665487 670634 665493
rect 670678 665027 670730 665033
rect 670678 664969 670730 664975
rect 670582 644085 670634 644091
rect 670582 644027 670634 644033
rect 670486 642309 670538 642315
rect 670486 642251 670538 642257
rect 670390 623217 670442 623223
rect 670390 623159 670442 623165
rect 670198 622477 670250 622483
rect 670198 622419 670250 622425
rect 669814 619887 669866 619893
rect 669814 619829 669866 619835
rect 669716 275234 669772 275243
rect 669716 275169 669772 275178
rect 669826 264989 669854 619829
rect 670210 578894 670238 622419
rect 670294 621367 670346 621373
rect 670294 621309 670346 621315
rect 670114 578866 670238 578894
rect 670114 577491 670142 578866
rect 670102 577485 670154 577491
rect 670102 577427 670154 577433
rect 669910 576079 669962 576085
rect 669910 576021 669962 576027
rect 669922 277759 669950 576021
rect 670006 488167 670058 488173
rect 670006 488109 670058 488115
rect 669908 277750 669964 277759
rect 669908 277685 669964 277694
rect 670018 270655 670046 488109
rect 670114 277907 670142 577427
rect 670306 576603 670334 621309
rect 670294 576597 670346 576603
rect 670294 576539 670346 576545
rect 670306 576085 670334 576539
rect 670294 576079 670346 576085
rect 670294 576021 670346 576027
rect 670390 575931 670442 575937
rect 670390 575873 670442 575879
rect 670402 538574 670430 575873
rect 670498 571127 670526 642251
rect 670486 571121 670538 571127
rect 670486 571063 670538 571069
rect 670594 570609 670622 644027
rect 670690 621965 670718 664969
rect 670786 660519 670814 737489
rect 670882 711949 670910 890373
rect 670978 713133 671006 891409
rect 673270 782983 673322 782989
rect 673270 782925 673322 782931
rect 673174 778765 673226 778771
rect 673174 778707 673226 778713
rect 672598 734957 672650 734963
rect 672598 734899 672650 734905
rect 670966 713127 671018 713133
rect 670966 713069 671018 713075
rect 670870 711943 670922 711949
rect 670870 711885 670922 711891
rect 670966 693665 671018 693671
rect 670966 693607 671018 693613
rect 670774 660513 670826 660519
rect 670774 660455 670826 660461
rect 670870 648969 670922 648975
rect 670870 648911 670922 648917
rect 670774 648377 670826 648383
rect 670774 648319 670826 648325
rect 670678 621959 670730 621965
rect 670678 621901 670730 621907
rect 670690 619893 670718 621901
rect 670678 619887 670730 619893
rect 670678 619829 670730 619835
rect 670678 599315 670730 599321
rect 670678 599257 670730 599263
rect 670582 570603 670634 570609
rect 670582 570545 670634 570551
rect 670306 538546 670430 538574
rect 670306 531537 670334 538546
rect 670294 531531 670346 531537
rect 670294 531473 670346 531479
rect 670198 487131 670250 487137
rect 670198 487073 670250 487079
rect 670100 277898 670156 277907
rect 670100 277833 670156 277842
rect 670210 274355 670238 487073
rect 670306 278055 670334 531473
rect 670690 525987 670718 599257
rect 670786 571571 670814 648319
rect 670882 572311 670910 648911
rect 670978 617155 671006 693607
rect 672610 658669 672638 734899
rect 672982 734439 673034 734445
rect 672982 734381 673034 734387
rect 672886 732367 672938 732373
rect 672886 732309 672938 732315
rect 672790 713423 672842 713429
rect 672790 713365 672842 713371
rect 672694 687375 672746 687381
rect 672694 687317 672746 687323
rect 672598 658663 672650 658669
rect 672598 658605 672650 658611
rect 672598 623439 672650 623445
rect 672598 623381 672650 623387
rect 670966 617149 671018 617155
rect 670966 617091 671018 617097
rect 670966 603311 671018 603317
rect 670966 603253 671018 603259
rect 670870 572305 670922 572311
rect 670870 572247 670922 572253
rect 670774 571565 670826 571571
rect 670774 571507 670826 571513
rect 670870 551955 670922 551961
rect 670870 551897 670922 551903
rect 670678 525981 670730 525987
rect 670678 525923 670730 525929
rect 670882 481957 670910 551897
rect 670978 526727 671006 603253
rect 672610 578823 672638 623381
rect 672706 616563 672734 687317
rect 672802 667623 672830 713365
rect 672790 667617 672842 667623
rect 672790 667559 672842 667565
rect 672790 666803 672842 666809
rect 672790 666745 672842 666751
rect 672802 624037 672830 666745
rect 672898 660149 672926 732309
rect 672886 660143 672938 660149
rect 672886 660085 672938 660091
rect 672994 659779 673022 734381
rect 673078 734217 673130 734223
rect 673078 734159 673130 734165
rect 672982 659773 673034 659779
rect 672982 659715 673034 659721
rect 673090 658299 673118 734159
rect 673186 704919 673214 778707
rect 673282 705585 673310 782925
rect 673378 714243 673406 892371
rect 676052 891506 676108 891515
rect 676052 891441 676054 891450
rect 676106 891441 676108 891450
rect 676054 891409 676106 891415
rect 676052 890470 676108 890479
rect 676052 890405 676054 890414
rect 676106 890405 676108 890414
rect 676054 890373 676106 890379
rect 680276 890174 680332 890183
rect 680276 890109 680332 890118
rect 676244 889286 676300 889295
rect 676244 889221 676300 889230
rect 676052 887954 676108 887963
rect 676052 887889 676108 887898
rect 676066 887551 676094 887889
rect 674230 887545 674282 887551
rect 674230 887487 674282 887493
rect 676054 887545 676106 887551
rect 676054 887487 676106 887493
rect 674038 885103 674090 885109
rect 674038 885045 674090 885051
rect 674050 872751 674078 885045
rect 674134 881033 674186 881039
rect 674134 880975 674186 880981
rect 674038 872745 674090 872751
rect 674038 872687 674090 872693
rect 674146 868829 674174 880975
rect 674242 870605 674270 887487
rect 676052 887436 676108 887445
rect 676052 887371 676108 887380
rect 675094 887175 675146 887181
rect 675094 887117 675146 887123
rect 674902 884437 674954 884443
rect 674818 884385 674902 884388
rect 674818 884379 674954 884385
rect 674818 884360 674942 884379
rect 674614 883623 674666 883629
rect 674614 883565 674666 883571
rect 674422 881995 674474 882001
rect 674422 881937 674474 881943
rect 674326 881699 674378 881705
rect 674326 881641 674378 881647
rect 674338 876747 674366 881641
rect 674434 881039 674462 881937
rect 674422 881033 674474 881039
rect 674422 880975 674474 880981
rect 674422 880885 674474 880891
rect 674422 880827 674474 880833
rect 674326 876741 674378 876747
rect 674326 876683 674378 876689
rect 674230 870599 674282 870605
rect 674230 870541 674282 870547
rect 674134 868823 674186 868829
rect 674134 868765 674186 868771
rect 674434 865795 674462 880827
rect 674518 878665 674570 878671
rect 674518 878607 674570 878613
rect 674530 869791 674558 878607
rect 674626 870013 674654 883565
rect 674818 872844 674846 884360
rect 674902 884215 674954 884221
rect 674902 884157 674954 884163
rect 674914 872973 674942 884157
rect 675106 880891 675134 887117
rect 676066 887107 676094 887371
rect 676258 887181 676286 889221
rect 680084 888694 680140 888703
rect 680084 888629 680140 888638
rect 676246 887175 676298 887181
rect 676246 887117 676298 887123
rect 675190 887101 675242 887107
rect 675190 887043 675242 887049
rect 676054 887101 676106 887107
rect 676054 887043 676106 887049
rect 675094 880885 675146 880891
rect 675094 880827 675146 880833
rect 675094 880737 675146 880743
rect 675094 880679 675146 880685
rect 674998 879553 675050 879559
rect 674998 879495 675050 879501
rect 675010 873565 675038 879495
rect 675106 874971 675134 880679
rect 675202 878671 675230 887043
rect 679700 886770 679756 886779
rect 679700 886705 679756 886714
rect 676052 885512 676108 885521
rect 676052 885447 676108 885456
rect 676066 885109 676094 885447
rect 676054 885103 676106 885109
rect 676054 885045 676106 885051
rect 676052 884994 676108 885003
rect 676052 884929 676108 884938
rect 676066 884443 676094 884929
rect 676054 884437 676106 884443
rect 676054 884379 676106 884385
rect 676244 884254 676300 884263
rect 676244 884189 676246 884198
rect 676298 884189 676300 884198
rect 676246 884157 676298 884163
rect 676052 884032 676108 884041
rect 676052 883967 676108 883976
rect 676066 883629 676094 883967
rect 676054 883623 676106 883629
rect 676054 883565 676106 883571
rect 676052 883514 676108 883523
rect 676052 883449 676108 883458
rect 675286 882883 675338 882889
rect 675286 882825 675338 882831
rect 675190 878665 675242 878671
rect 675190 878607 675242 878613
rect 675190 878517 675242 878523
rect 675190 878459 675242 878465
rect 675094 874965 675146 874971
rect 675094 874907 675146 874913
rect 675202 874305 675230 878459
rect 675298 876840 675326 882825
rect 675766 882291 675818 882297
rect 675766 882233 675818 882239
rect 675478 881403 675530 881409
rect 675478 881345 675530 881351
rect 675490 878084 675518 881345
rect 675778 878375 675806 882233
rect 676066 882001 676094 883449
rect 679714 882889 679742 886705
rect 679892 886178 679948 886187
rect 679892 886113 679948 886122
rect 679702 882883 679754 882889
rect 679702 882825 679754 882831
rect 679796 882774 679852 882783
rect 679796 882709 679852 882718
rect 679810 882191 679838 882709
rect 679796 882182 679852 882191
rect 679796 882117 679852 882126
rect 676054 881995 676106 882001
rect 676054 881937 676106 881943
rect 679810 881483 679838 882117
rect 679798 881477 679850 881483
rect 679798 881419 679850 881425
rect 679906 878523 679934 886113
rect 679988 885734 680044 885743
rect 679988 885669 680044 885678
rect 680002 879559 680030 885669
rect 680098 882297 680126 888629
rect 680180 888250 680236 888259
rect 680180 888185 680236 888194
rect 680086 882291 680138 882297
rect 680086 882233 680138 882239
rect 680194 880743 680222 888185
rect 680290 881705 680318 890109
rect 685460 882182 685516 882191
rect 685460 882117 685516 882126
rect 685474 881747 685502 882117
rect 685460 881738 685516 881747
rect 680278 881699 680330 881705
rect 685460 881673 685516 881682
rect 680278 881641 680330 881647
rect 680182 880737 680234 880743
rect 680182 880679 680234 880685
rect 679990 879553 680042 879559
rect 679990 879495 680042 879501
rect 679894 878517 679946 878523
rect 679894 878459 679946 878465
rect 675766 878369 675818 878375
rect 675766 878311 675818 878317
rect 675766 877851 675818 877857
rect 675766 877793 675818 877799
rect 675778 877523 675806 877793
rect 675394 876840 675422 876900
rect 675298 876812 675422 876840
rect 675286 876741 675338 876747
rect 675286 876683 675338 876689
rect 675298 876248 675326 876683
rect 675298 876220 675408 876248
rect 675478 874965 675530 874971
rect 675478 874907 675530 874913
rect 675490 874384 675518 874907
rect 675190 874299 675242 874305
rect 675190 874241 675242 874247
rect 675478 874299 675530 874305
rect 675478 874241 675530 874247
rect 675490 873866 675518 874241
rect 674998 873559 675050 873565
rect 674998 873501 675050 873507
rect 675382 873559 675434 873565
rect 675382 873501 675434 873507
rect 675394 873200 675422 873501
rect 674902 872967 674954 872973
rect 674902 872909 674954 872915
rect 675382 872967 675434 872973
rect 675382 872909 675434 872915
rect 674818 872816 675230 872844
rect 674902 872745 674954 872751
rect 674902 872687 674954 872693
rect 674614 870007 674666 870013
rect 674614 869949 674666 869955
rect 674518 869785 674570 869791
rect 674518 869727 674570 869733
rect 674914 867423 674942 872687
rect 675094 872671 675146 872677
rect 675094 872613 675146 872619
rect 674998 869785 675050 869791
rect 674998 869727 675050 869733
rect 674902 867417 674954 867423
rect 674902 867359 674954 867365
rect 674422 865789 674474 865795
rect 674422 865731 674474 865737
rect 675010 863372 675038 869727
rect 675106 867693 675134 872613
rect 675202 868889 675230 872816
rect 675394 872534 675422 872909
rect 675478 870599 675530 870605
rect 675478 870541 675530 870547
rect 675490 870092 675518 870541
rect 675382 870007 675434 870013
rect 675382 869949 675434 869955
rect 675394 869500 675422 869949
rect 675202 868861 675408 868889
rect 675190 868823 675242 868829
rect 675190 868765 675242 868771
rect 675202 868256 675230 868765
rect 675202 868228 675408 868256
rect 675106 867665 675408 867693
rect 675478 867417 675530 867423
rect 675478 867359 675530 867365
rect 675490 867058 675518 867359
rect 675106 865825 675408 865853
rect 675106 864019 675134 865825
rect 675190 865789 675242 865795
rect 675190 865731 675242 865737
rect 675202 865222 675230 865731
rect 675202 865194 675408 865222
rect 675094 864013 675146 864019
rect 675094 863955 675146 863961
rect 675010 863344 675408 863372
rect 675382 792085 675434 792091
rect 675382 792027 675434 792033
rect 675394 788875 675422 792027
rect 675394 788063 675422 788322
rect 675380 788054 675436 788063
rect 675380 787989 675436 787998
rect 675682 787175 675710 787656
rect 675668 787166 675724 787175
rect 675668 787101 675724 787110
rect 675394 786731 675422 787035
rect 675380 786722 675436 786731
rect 675380 786657 675436 786666
rect 675394 784807 675422 785214
rect 675380 784798 675436 784807
rect 675380 784733 675436 784742
rect 675778 784215 675806 784622
rect 675764 784206 675820 784215
rect 675764 784141 675820 784150
rect 675298 783985 675408 784013
rect 674998 783501 675050 783507
rect 675298 783475 675326 783985
rect 674998 783443 675050 783449
rect 675284 783466 675340 783475
rect 675010 778919 675038 783443
rect 675284 783401 675340 783410
rect 675394 782989 675422 783364
rect 675382 782983 675434 782989
rect 675382 782925 675434 782931
rect 675490 780663 675518 780848
rect 675476 780654 675532 780663
rect 675476 780589 675532 780598
rect 675286 780541 675338 780547
rect 675286 780483 675338 780489
rect 674998 778913 675050 778919
rect 674998 778855 675050 778861
rect 675298 776644 675326 780483
rect 675778 779923 675806 780330
rect 675764 779914 675820 779923
rect 675764 779849 675820 779858
rect 675778 779183 675806 779664
rect 675764 779174 675820 779183
rect 675764 779109 675820 779118
rect 675382 778913 675434 778919
rect 675382 778855 675434 778861
rect 675394 778480 675422 778855
rect 675490 778771 675518 779031
rect 675478 778765 675530 778771
rect 675478 778707 675530 778713
rect 675778 777703 675806 777814
rect 675764 777694 675820 777703
rect 675764 777629 675820 777638
rect 675298 776616 675408 776644
rect 675778 775483 675806 775995
rect 675764 775474 675820 775483
rect 675764 775409 675820 775418
rect 675298 774141 675408 774169
rect 675298 773665 675326 774141
rect 674614 773659 674666 773665
rect 674614 773601 674666 773607
rect 675286 773659 675338 773665
rect 675286 773601 675338 773607
rect 674422 742801 674474 742807
rect 674422 742743 674474 742749
rect 674434 731948 674462 742743
rect 674518 737473 674570 737479
rect 674518 737415 674570 737421
rect 674530 732077 674558 737415
rect 674518 732071 674570 732077
rect 674518 732013 674570 732019
rect 674434 731920 674558 731948
rect 674422 730517 674474 730523
rect 674422 730459 674474 730465
rect 674134 728667 674186 728673
rect 674134 728609 674186 728615
rect 673366 714237 673418 714243
rect 673366 714179 673418 714185
rect 673270 705579 673322 705585
rect 673270 705521 673322 705527
rect 673174 704913 673226 704919
rect 673174 704855 673226 704861
rect 673174 689817 673226 689823
rect 673174 689759 673226 689765
rect 673078 658293 673130 658299
rect 673078 658235 673130 658241
rect 672982 644603 673034 644609
rect 672982 644545 673034 644551
rect 672886 643641 672938 643647
rect 672886 643583 672938 643589
rect 672790 624031 672842 624037
rect 672790 623973 672842 623979
rect 672694 616557 672746 616563
rect 672694 616499 672746 616505
rect 672790 598945 672842 598951
rect 672790 598887 672842 598893
rect 672694 597169 672746 597175
rect 672694 597111 672746 597117
rect 672598 578817 672650 578823
rect 672598 578759 672650 578765
rect 672502 577855 672554 577861
rect 672502 577797 672554 577803
rect 672514 533831 672542 577797
rect 672598 577115 672650 577121
rect 672598 577057 672650 577063
rect 672502 533825 672554 533831
rect 672502 533767 672554 533773
rect 672610 532721 672638 577057
rect 672406 532715 672458 532721
rect 672406 532657 672458 532663
rect 672598 532715 672650 532721
rect 672598 532657 672650 532663
rect 670966 526721 671018 526727
rect 670966 526663 671018 526669
rect 670870 481951 670922 481957
rect 670870 481893 670922 481899
rect 670484 308978 670540 308987
rect 670484 308913 670540 308922
rect 670498 278647 670526 308913
rect 670484 278638 670540 278647
rect 670484 278573 670540 278582
rect 670292 278046 670348 278055
rect 670292 277981 670348 277990
rect 672418 276279 672446 532657
rect 672706 526357 672734 597111
rect 672694 526351 672746 526357
rect 672694 526293 672746 526299
rect 672802 524507 672830 598887
rect 672898 569129 672926 643583
rect 672994 569647 673022 644545
rect 673186 615231 673214 689759
rect 673366 689373 673418 689379
rect 673366 689315 673418 689321
rect 673270 689151 673322 689157
rect 673270 689093 673322 689099
rect 673174 615225 673226 615231
rect 673174 615167 673226 615173
rect 673282 614491 673310 689093
rect 673378 615971 673406 689315
rect 674146 662369 674174 728609
rect 674326 685525 674378 685531
rect 674326 685467 674378 685473
rect 674230 683675 674282 683681
rect 674230 683617 674282 683623
rect 674134 662363 674186 662369
rect 674134 662305 674186 662311
rect 673846 648081 673898 648087
rect 673846 648023 673898 648029
rect 673366 615965 673418 615971
rect 673366 615907 673418 615913
rect 673270 614485 673322 614491
rect 673270 614427 673322 614433
rect 673270 606937 673322 606943
rect 673270 606879 673322 606885
rect 673078 601979 673130 601985
rect 673078 601921 673130 601927
rect 672982 569641 673034 569647
rect 672982 569583 673034 569589
rect 672886 569123 672938 569129
rect 672886 569065 672938 569071
rect 672886 553953 672938 553959
rect 672886 553895 672938 553901
rect 672790 524501 672842 524507
rect 672790 524443 672842 524449
rect 672898 481587 672926 553895
rect 673090 527467 673118 601921
rect 673174 599611 673226 599617
rect 673174 599553 673226 599559
rect 673078 527461 673130 527467
rect 673078 527403 673130 527409
rect 673186 524877 673214 599553
rect 673282 528059 673310 606879
rect 673366 603089 673418 603095
rect 673366 603031 673418 603037
rect 673270 528053 673322 528059
rect 673270 527995 673322 528001
rect 673378 525247 673406 603031
rect 673858 570239 673886 648023
rect 674242 618857 674270 683617
rect 674338 622039 674366 685467
rect 674434 665255 674462 730459
rect 674530 728567 674558 731920
rect 674516 728558 674572 728567
rect 674516 728493 674572 728502
rect 674626 711357 674654 773601
rect 674996 771922 675052 771931
rect 674996 771857 675052 771866
rect 674902 741469 674954 741475
rect 674902 741411 674954 741417
rect 674914 731675 674942 741411
rect 674900 731666 674956 731675
rect 674900 731601 674956 731610
rect 674614 711351 674666 711357
rect 674614 711293 674666 711299
rect 675010 708471 675038 771857
rect 675382 748869 675434 748875
rect 675382 748811 675434 748817
rect 675394 743848 675422 748811
rect 675202 743316 675408 743344
rect 675202 742807 675230 743316
rect 675190 742801 675242 742807
rect 675190 742743 675242 742749
rect 675298 742724 675422 742752
rect 675298 742678 675326 742724
rect 675202 742650 675326 742678
rect 675394 742664 675422 742724
rect 675202 741475 675230 742650
rect 675298 742021 675408 742049
rect 675190 741469 675242 741475
rect 675190 741411 675242 741417
rect 675298 741147 675326 742021
rect 675284 741138 675340 741147
rect 675284 741073 675340 741082
rect 675476 740398 675532 740407
rect 675476 740333 675532 740342
rect 675490 740222 675518 740333
rect 675284 739658 675340 739667
rect 675340 739616 675408 739644
rect 675284 739593 675340 739602
rect 675298 738985 675408 739013
rect 675298 737553 675326 738985
rect 675778 738039 675806 738372
rect 675764 738030 675820 738039
rect 675764 737965 675820 737974
rect 675286 737547 675338 737553
rect 675286 737489 675338 737495
rect 675286 737399 675338 737405
rect 675286 737341 675338 737347
rect 675298 736832 675326 737341
rect 675202 736804 675326 736832
rect 675202 733927 675230 736804
rect 675682 735523 675710 735856
rect 675668 735514 675724 735523
rect 675668 735449 675724 735458
rect 675394 734963 675422 735338
rect 675382 734957 675434 734963
rect 675382 734899 675434 734905
rect 675394 734445 675422 734672
rect 675382 734439 675434 734445
rect 675382 734381 675434 734387
rect 675382 734217 675434 734223
rect 675382 734159 675434 734165
rect 675394 734006 675422 734159
rect 675190 733921 675242 733927
rect 675190 733863 675242 733869
rect 675478 733921 675530 733927
rect 675478 733863 675530 733869
rect 675490 733488 675518 733863
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 679796 728114 679852 728123
rect 679796 728049 679852 728058
rect 676340 715534 676396 715543
rect 676340 715469 676396 715478
rect 676148 714942 676204 714951
rect 676148 714877 676204 714886
rect 676162 714613 676190 714877
rect 676244 714794 676300 714803
rect 676244 714729 676246 714738
rect 676298 714729 676300 714738
rect 676246 714697 676298 714703
rect 676150 714607 676202 714613
rect 676150 714549 676202 714555
rect 676354 714465 676382 715469
rect 676342 714459 676394 714465
rect 676342 714401 676394 714407
rect 676054 714237 676106 714243
rect 676052 714202 676054 714211
rect 676106 714202 676108 714211
rect 676052 714137 676108 714146
rect 676244 713462 676300 713471
rect 676244 713397 676246 713406
rect 676298 713397 676300 713406
rect 676246 713365 676298 713371
rect 676052 713166 676108 713175
rect 676052 713101 676054 713110
rect 676106 713101 676108 713110
rect 676054 713069 676106 713075
rect 676052 712722 676108 712731
rect 676052 712657 676054 712666
rect 676106 712657 676108 712666
rect 676054 712625 676106 712631
rect 676244 711982 676300 711991
rect 676244 711917 676246 711926
rect 676298 711917 676300 711926
rect 676246 711885 676298 711891
rect 676052 711612 676108 711621
rect 676052 711547 676054 711556
rect 676106 711547 676108 711556
rect 676054 711515 676106 711521
rect 676054 711351 676106 711357
rect 676054 711293 676106 711299
rect 676066 708587 676094 711293
rect 676052 708578 676108 708587
rect 676052 708513 676108 708522
rect 674998 708465 675050 708471
rect 674998 708407 675050 708413
rect 676054 708465 676106 708471
rect 676054 708407 676106 708413
rect 676066 708217 676094 708407
rect 676052 708208 676108 708217
rect 676052 708143 676108 708152
rect 679810 706959 679838 728049
rect 679796 706950 679852 706959
rect 679796 706885 679852 706894
rect 676052 705618 676108 705627
rect 676052 705553 676054 705562
rect 676106 705553 676108 705562
rect 676054 705521 676106 705527
rect 676246 704913 676298 704919
rect 676244 704878 676246 704887
rect 676298 704878 676300 704887
rect 676244 704813 676300 704822
rect 679988 704434 680044 704443
rect 679988 704369 680044 704378
rect 680002 703407 680030 704369
rect 679796 703398 679852 703407
rect 679796 703333 679852 703342
rect 679988 703398 680044 703407
rect 679988 703333 680044 703342
rect 679810 702963 679838 703333
rect 679796 702954 679852 702963
rect 679796 702889 679852 702898
rect 675382 702841 675434 702847
rect 675382 702783 675434 702789
rect 675394 698856 675422 702783
rect 680002 702773 680030 703333
rect 679990 702767 680042 702773
rect 679990 702709 680042 702715
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675778 697191 675806 697672
rect 675764 697182 675820 697191
rect 675764 697117 675820 697126
rect 675202 697043 675408 697049
rect 675188 697034 675408 697043
rect 675244 697021 675408 697034
rect 675188 696969 675244 696978
rect 675586 694823 675614 695195
rect 675572 694814 675628 694823
rect 675572 694749 675628 694758
rect 674998 694331 675050 694337
rect 674998 694273 675050 694279
rect 674902 692925 674954 692931
rect 674902 692867 674954 692873
rect 674614 690483 674666 690489
rect 674614 690425 674666 690431
rect 674422 665249 674474 665255
rect 674422 665191 674474 665197
rect 674326 622033 674378 622039
rect 674326 621975 674378 621981
rect 674626 619079 674654 690425
rect 674914 686535 674942 692867
rect 675010 688935 675038 694273
rect 675778 694231 675806 694638
rect 675764 694222 675820 694231
rect 675764 694157 675820 694166
rect 675490 693671 675518 693972
rect 675478 693665 675530 693671
rect 675478 693607 675530 693613
rect 675394 692931 675422 693380
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675190 691371 675242 691377
rect 675190 691313 675242 691319
rect 674998 688929 675050 688935
rect 674998 688871 675050 688877
rect 675202 687085 675230 691313
rect 675490 690489 675518 690864
rect 675478 690483 675530 690489
rect 675478 690425 675530 690431
rect 675394 689823 675422 690346
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675394 689379 675422 689680
rect 675382 689373 675434 689379
rect 675382 689315 675434 689321
rect 675382 689151 675434 689157
rect 675382 689093 675434 689099
rect 675394 689014 675422 689093
rect 675478 688929 675530 688935
rect 675478 688871 675530 688877
rect 675490 688496 675518 688871
rect 675490 687381 675518 687830
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 675190 687079 675242 687085
rect 675190 687021 675242 687027
rect 675478 687079 675530 687085
rect 675478 687021 675530 687027
rect 675490 686646 675518 687021
rect 674900 686526 674956 686535
rect 674900 686461 674956 686470
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 676244 668766 676300 668775
rect 676244 668701 676300 668710
rect 676258 668437 676286 668701
rect 676246 668431 676298 668437
rect 676246 668373 676298 668379
rect 676244 668322 676300 668331
rect 676244 668257 676300 668266
rect 676258 668215 676286 668257
rect 676246 668209 676298 668215
rect 676246 668151 676298 668157
rect 676052 668026 676108 668035
rect 676052 667961 676108 667970
rect 675958 667617 676010 667623
rect 675956 667582 675958 667591
rect 676010 667582 676012 667591
rect 675956 667517 676012 667526
rect 675956 666102 676012 666111
rect 675956 666037 675958 666046
rect 676010 666037 676012 666046
rect 675958 666005 676010 666011
rect 675958 665545 676010 665551
rect 675956 665510 675958 665519
rect 676010 665510 676012 665519
rect 676066 665477 676094 667961
rect 676244 666842 676300 666851
rect 676244 666777 676246 666786
rect 676298 666777 676300 666786
rect 676246 666745 676298 666751
rect 676150 666729 676202 666735
rect 676148 666694 676150 666703
rect 676202 666694 676204 666703
rect 676148 666629 676204 666638
rect 675956 665445 676012 665454
rect 676054 665471 676106 665477
rect 676054 665413 676106 665419
rect 676054 665249 676106 665255
rect 676054 665191 676106 665197
rect 675956 665066 676012 665075
rect 675956 665001 675958 665010
rect 676010 665001 676012 665010
rect 675958 664969 676010 664975
rect 676066 664039 676094 665191
rect 676052 664030 676108 664039
rect 676052 663965 676108 663974
rect 676054 662363 676106 662369
rect 676054 662305 676106 662311
rect 676066 662041 676094 662305
rect 676052 662032 676108 662041
rect 676052 661967 676108 661976
rect 676054 660513 676106 660519
rect 676052 660478 676054 660487
rect 676106 660478 676108 660487
rect 676052 660413 676108 660422
rect 676054 660143 676106 660149
rect 676052 660108 676054 660117
rect 676106 660108 676108 660117
rect 676052 660043 676108 660052
rect 676246 659773 676298 659779
rect 676244 659738 676246 659747
rect 676298 659738 676300 659747
rect 676244 659673 676300 659682
rect 676054 658663 676106 658669
rect 676052 658628 676054 658637
rect 676106 658628 676108 658637
rect 676052 658563 676108 658572
rect 676246 658293 676298 658299
rect 676244 658258 676246 658267
rect 676298 658258 676300 658267
rect 676244 658193 676300 658202
rect 679988 657370 680044 657379
rect 679988 657305 680044 657314
rect 680002 656787 680030 657305
rect 679796 656778 679852 656787
rect 675382 656739 675434 656745
rect 679796 656713 679852 656722
rect 679988 656778 680044 656787
rect 679988 656713 680044 656722
rect 675382 656681 675434 656687
rect 675394 653675 675422 656681
rect 679810 656343 679838 656713
rect 679796 656334 679852 656343
rect 679796 656269 679852 656278
rect 680002 654155 680030 656713
rect 679990 654149 680042 654155
rect 679990 654091 680042 654097
rect 675394 652643 675422 653124
rect 675380 652634 675436 652643
rect 675380 652569 675436 652578
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675394 651459 675422 651835
rect 675380 651450 675436 651459
rect 675380 651385 675436 651394
rect 675394 649683 675422 650016
rect 675380 649674 675436 649683
rect 675380 649609 675436 649618
rect 675298 649484 675422 649512
rect 675298 649438 675326 649484
rect 675202 649410 675326 649438
rect 675394 649424 675422 649484
rect 675202 648975 675230 649410
rect 675190 648969 675242 648975
rect 675190 648911 675242 648917
rect 675202 648785 675408 648813
rect 675202 648383 675230 648785
rect 675190 648377 675242 648383
rect 675190 648319 675242 648325
rect 674998 648303 675050 648309
rect 674998 648245 675050 648251
rect 675010 643721 675038 648245
rect 675202 648152 675408 648180
rect 675202 648087 675230 648152
rect 675190 648081 675242 648087
rect 675190 648023 675242 648029
rect 675682 645391 675710 645650
rect 675668 645382 675724 645391
rect 675668 645317 675724 645326
rect 675286 645195 675338 645201
rect 675286 645137 675338 645143
rect 674998 643715 675050 643721
rect 674998 643657 675050 643663
rect 675298 641446 675326 645137
rect 675394 644609 675422 645132
rect 675382 644603 675434 644609
rect 675382 644545 675434 644551
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675382 643715 675434 643721
rect 675382 643657 675434 643663
rect 675394 643282 675422 643657
rect 675490 643647 675518 643831
rect 675478 643641 675530 643647
rect 675478 643583 675530 643589
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675298 641418 675408 641446
rect 675298 640781 675408 640809
rect 675298 640063 675326 640781
rect 675284 640054 675340 640063
rect 675284 639989 675340 639998
rect 675778 638583 675806 638955
rect 675764 638574 675820 638583
rect 675764 638509 675820 638518
rect 678164 636650 678220 636659
rect 678164 636585 678220 636594
rect 676244 625106 676300 625115
rect 676244 625041 676300 625050
rect 676258 624999 676286 625041
rect 676246 624993 676298 624999
rect 676246 624935 676298 624941
rect 676148 624662 676204 624671
rect 676148 624597 676204 624606
rect 676054 624031 676106 624037
rect 676052 623996 676054 624005
rect 676106 623996 676108 624005
rect 676052 623931 676108 623940
rect 676052 623478 676108 623487
rect 676052 623413 676054 623422
rect 676106 623413 676108 623422
rect 676054 623381 676106 623387
rect 676052 622516 676108 622525
rect 676052 622451 676054 622460
rect 676106 622451 676108 622460
rect 676054 622419 676106 622425
rect 676162 622261 676190 624597
rect 676244 624218 676300 624227
rect 676244 624153 676300 624162
rect 676258 622409 676286 624153
rect 676342 623217 676394 623223
rect 676340 623182 676342 623191
rect 676394 623182 676396 623191
rect 676340 623117 676396 623126
rect 676246 622403 676298 622409
rect 676246 622345 676298 622351
rect 676150 622255 676202 622261
rect 676150 622197 676202 622203
rect 676246 622033 676298 622039
rect 676052 621998 676108 622007
rect 676246 621975 676298 621981
rect 676052 621933 676054 621942
rect 676106 621933 676108 621942
rect 676054 621901 676106 621907
rect 676052 621406 676108 621415
rect 676052 621341 676054 621350
rect 676106 621341 676108 621350
rect 676054 621309 676106 621315
rect 676258 620675 676286 621975
rect 676244 620666 676300 620675
rect 676244 620601 676300 620610
rect 674614 619073 674666 619079
rect 674614 619015 674666 619021
rect 676054 619073 676106 619079
rect 676054 619015 676106 619021
rect 676066 618973 676094 619015
rect 676052 618964 676108 618973
rect 676052 618899 676108 618908
rect 674230 618851 674282 618857
rect 674230 618793 674282 618799
rect 676246 618851 676298 618857
rect 676246 618793 676298 618799
rect 676258 618603 676286 618793
rect 676244 618594 676300 618603
rect 676244 618529 676300 618538
rect 678178 617715 678206 636585
rect 678164 617706 678220 617715
rect 678164 617641 678220 617650
rect 676246 617149 676298 617155
rect 676244 617114 676246 617123
rect 676298 617114 676300 617123
rect 676244 617049 676300 617058
rect 676054 616557 676106 616563
rect 676052 616522 676054 616531
rect 676106 616522 676108 616531
rect 676052 616457 676108 616466
rect 676054 615965 676106 615971
rect 676052 615930 676054 615939
rect 676106 615930 676108 615939
rect 676052 615865 676108 615874
rect 676246 615225 676298 615231
rect 676244 615190 676246 615199
rect 676298 615190 676300 615199
rect 676244 615125 676300 615134
rect 676054 614485 676106 614491
rect 676052 614450 676054 614459
rect 676106 614450 676108 614459
rect 676052 614385 676108 614394
rect 679988 613710 680044 613719
rect 679988 613645 680044 613654
rect 675382 613523 675434 613529
rect 675382 613465 675434 613471
rect 675394 608650 675422 613465
rect 680002 613275 680030 613645
rect 679796 613266 679852 613275
rect 679796 613201 679852 613210
rect 679988 613266 680044 613275
rect 679988 613201 680044 613210
rect 679810 612831 679838 613201
rect 679796 612822 679852 612831
rect 679796 612757 679852 612766
rect 680002 610717 680030 613201
rect 679990 610711 680042 610717
rect 679990 610653 680042 610659
rect 675202 608118 675408 608146
rect 675202 607799 675230 608118
rect 675188 607790 675244 607799
rect 675188 607725 675244 607734
rect 675202 607452 675408 607480
rect 675202 606943 675230 607452
rect 675190 606937 675242 606943
rect 675190 606879 675242 606885
rect 675202 606821 675408 606849
rect 675202 606023 675230 606821
rect 675188 606014 675244 606023
rect 675188 605949 675244 605958
rect 675298 604981 675408 605009
rect 675298 604839 675326 604981
rect 675284 604830 675340 604839
rect 675284 604765 675340 604774
rect 675298 604418 675408 604446
rect 674998 602127 675050 602133
rect 674998 602069 675050 602075
rect 674902 602053 674954 602059
rect 674902 601995 674954 602001
rect 674914 596879 674942 601995
rect 675010 598729 675038 602069
rect 675298 601985 675326 604418
rect 675394 603317 675422 603799
rect 675382 603311 675434 603317
rect 675382 603253 675434 603259
rect 675394 603095 675422 603174
rect 675382 603089 675434 603095
rect 675382 603031 675434 603037
rect 675286 601979 675338 601985
rect 675286 601921 675338 601927
rect 675490 600251 675518 600658
rect 675476 600242 675532 600251
rect 675476 600177 675532 600186
rect 675394 599617 675422 600140
rect 675382 599611 675434 599617
rect 675382 599553 675434 599559
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675382 598945 675434 598951
rect 675382 598887 675434 598893
rect 675394 598808 675422 598887
rect 674998 598723 675050 598729
rect 674998 598665 675050 598671
rect 675478 598723 675530 598729
rect 675478 598665 675530 598671
rect 675490 598290 675518 598665
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 674902 596873 674954 596879
rect 674902 596815 674954 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675778 593443 675806 593955
rect 675764 593434 675820 593443
rect 675764 593369 675820 593378
rect 676340 579818 676396 579827
rect 676340 579753 676396 579762
rect 676148 579374 676204 579383
rect 676148 579309 676204 579318
rect 676246 579335 676298 579341
rect 676162 579045 676190 579309
rect 676246 579277 676298 579283
rect 676258 579235 676286 579277
rect 676244 579226 676300 579235
rect 676354 579193 676382 579753
rect 676244 579161 676300 579170
rect 676342 579187 676394 579193
rect 676342 579129 676394 579135
rect 676150 579039 676202 579045
rect 676150 578981 676202 578987
rect 676246 578817 676298 578823
rect 676244 578782 676246 578791
rect 676298 578782 676300 578791
rect 676244 578717 676300 578726
rect 676244 577894 676300 577903
rect 676244 577829 676246 577838
rect 676298 577829 676300 577838
rect 676246 577797 676298 577803
rect 676052 577524 676108 577533
rect 676052 577459 676054 577468
rect 676106 577459 676108 577468
rect 676054 577427 676106 577433
rect 676052 577154 676108 577163
rect 676052 577089 676054 577098
rect 676106 577089 676108 577098
rect 676054 577057 676106 577063
rect 676054 576597 676106 576603
rect 676052 576562 676054 576571
rect 676106 576562 676108 576571
rect 676052 576497 676108 576506
rect 676052 575970 676108 575979
rect 676052 575905 676054 575914
rect 676106 575905 676108 575914
rect 676054 575873 676106 575879
rect 676246 572305 676298 572311
rect 676244 572270 676246 572279
rect 676298 572270 676300 572279
rect 676244 572205 676300 572214
rect 676054 571565 676106 571571
rect 676052 571530 676054 571539
rect 676106 571530 676108 571539
rect 676052 571465 676108 571474
rect 676054 571121 676106 571127
rect 676052 571086 676054 571095
rect 676106 571086 676108 571095
rect 676052 571021 676108 571030
rect 676054 570603 676106 570609
rect 676052 570568 676054 570577
rect 676106 570568 676108 570577
rect 676052 570503 676108 570512
rect 673846 570233 673898 570239
rect 676246 570233 676298 570239
rect 673846 570175 673898 570181
rect 676244 570198 676246 570207
rect 676298 570198 676300 570207
rect 676244 570133 676300 570142
rect 676054 569641 676106 569647
rect 676052 569606 676054 569615
rect 676106 569606 676108 569615
rect 676052 569541 676108 569550
rect 676054 569123 676106 569129
rect 676052 569088 676054 569097
rect 676106 569088 676108 569097
rect 676052 569023 676108 569032
rect 679988 568718 680044 568727
rect 679988 568653 680044 568662
rect 680002 567839 680030 568653
rect 679796 567830 679852 567839
rect 679796 567765 679852 567774
rect 679988 567830 680044 567839
rect 679988 567765 680044 567774
rect 675382 567495 675434 567501
rect 675382 567437 675434 567443
rect 675394 563475 675422 567437
rect 679810 567395 679838 567765
rect 680002 567427 680030 567765
rect 679990 567421 680042 567427
rect 679796 567386 679852 567395
rect 679990 567363 680042 567369
rect 679796 567321 679852 567330
rect 675188 562946 675244 562955
rect 675244 562904 675408 562932
rect 675188 562881 675244 562890
rect 675490 561771 675518 562252
rect 675476 561762 675532 561771
rect 675476 561697 675532 561706
rect 675394 561475 675422 561660
rect 675380 561466 675436 561475
rect 675380 561401 675436 561410
rect 675394 559583 675422 559810
rect 674422 559577 674474 559583
rect 674422 559519 674474 559525
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 673846 556025 673898 556031
rect 673846 555967 673898 555973
rect 673750 554397 673802 554403
rect 673750 554339 673802 554345
rect 673654 553361 673706 553367
rect 673654 553303 673706 553309
rect 673366 525241 673418 525247
rect 673366 525183 673418 525189
rect 673174 524871 673226 524877
rect 673174 524813 673226 524819
rect 672886 481581 672938 481587
rect 672886 481523 672938 481529
rect 673666 480107 673694 553303
rect 673762 480477 673790 554339
rect 673858 480847 673886 555967
rect 674326 548921 674378 548927
rect 674326 548863 674378 548869
rect 674230 548255 674282 548261
rect 674230 548197 674282 548203
rect 674242 483733 674270 548197
rect 674338 486619 674366 548863
rect 674326 486613 674378 486619
rect 674326 486555 674378 486561
rect 674434 486545 674462 559519
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 674998 558837 675050 558843
rect 674998 558779 675050 558785
rect 674614 558097 674666 558103
rect 674614 558039 674666 558045
rect 674422 486539 674474 486545
rect 674422 486481 674474 486487
rect 674626 483807 674654 558039
rect 674902 555063 674954 555069
rect 674902 555005 674954 555011
rect 674914 538574 674942 555005
rect 675010 553515 675038 558779
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675298 557946 675408 557974
rect 675298 556031 675326 557946
rect 675286 556025 675338 556031
rect 675286 555967 675338 555973
rect 675286 555877 675338 555883
rect 675286 555819 675338 555825
rect 674998 553509 675050 553515
rect 674998 553451 675050 553457
rect 675298 551240 675326 555819
rect 675490 555069 675518 555444
rect 675478 555063 675530 555069
rect 675478 555005 675530 555011
rect 675394 554403 675422 554926
rect 675382 554397 675434 554403
rect 675382 554339 675434 554345
rect 675490 553959 675518 554260
rect 675478 553953 675530 553959
rect 675478 553895 675530 553901
rect 675382 553509 675434 553515
rect 675382 553451 675434 553457
rect 675394 553076 675422 553451
rect 675490 553367 675518 553631
rect 675478 553361 675530 553367
rect 675478 553303 675530 553309
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675298 551212 675408 551240
rect 675298 550581 675408 550609
rect 675298 548927 675326 550581
rect 675286 548921 675338 548927
rect 675286 548863 675338 548869
rect 675298 548741 675408 548769
rect 675298 548261 675326 548741
rect 675286 548255 675338 548261
rect 675286 548197 675338 548203
rect 674818 538546 674942 538574
rect 674818 518414 674846 538546
rect 676148 534974 676204 534983
rect 676148 534909 676204 534918
rect 676052 534234 676108 534243
rect 676052 534169 676108 534178
rect 675958 533825 676010 533831
rect 675956 533790 675958 533799
rect 676010 533790 676012 533799
rect 675956 533725 676012 533734
rect 676066 533313 676094 534169
rect 676054 533307 676106 533313
rect 676054 533249 676106 533255
rect 676162 533165 676190 534909
rect 676244 534382 676300 534391
rect 676244 534317 676300 534326
rect 676150 533159 676202 533165
rect 676150 533101 676202 533107
rect 676258 533017 676286 534317
rect 676724 533050 676780 533059
rect 676246 533011 676298 533017
rect 676724 532985 676780 532994
rect 676246 532953 676298 532959
rect 676052 532754 676108 532763
rect 676052 532689 676054 532698
rect 676106 532689 676108 532698
rect 676054 532657 676106 532663
rect 676628 532014 676684 532023
rect 676628 531949 676684 531958
rect 676244 531570 676300 531579
rect 676244 531505 676246 531514
rect 676298 531505 676300 531514
rect 676246 531473 676298 531479
rect 676532 530978 676588 530987
rect 676532 530913 676588 530922
rect 676246 528053 676298 528059
rect 676244 528018 676246 528027
rect 676298 528018 676300 528027
rect 676244 527953 676300 527962
rect 676246 527461 676298 527467
rect 676244 527426 676246 527435
rect 676298 527426 676300 527435
rect 676244 527361 676300 527370
rect 676054 526721 676106 526727
rect 676052 526686 676054 526695
rect 676106 526686 676108 526695
rect 676052 526621 676108 526630
rect 676054 526351 676106 526357
rect 676052 526316 676054 526325
rect 676106 526316 676108 526325
rect 676052 526251 676108 526260
rect 676246 525981 676298 525987
rect 676244 525946 676246 525955
rect 676298 525946 676300 525955
rect 676244 525881 676300 525890
rect 676054 525241 676106 525247
rect 676052 525206 676054 525215
rect 676106 525206 676108 525215
rect 676052 525141 676108 525150
rect 676054 524871 676106 524877
rect 676052 524836 676054 524845
rect 676106 524836 676108 524845
rect 676052 524771 676108 524780
rect 676246 524501 676298 524507
rect 676244 524466 676246 524475
rect 676298 524466 676300 524475
rect 676244 524401 676300 524410
rect 674818 518386 674942 518414
rect 674914 486693 674942 518386
rect 676148 490574 676204 490583
rect 676148 490509 676204 490518
rect 676162 489949 676190 490509
rect 676340 490130 676396 490139
rect 676246 490091 676298 490097
rect 676340 490065 676396 490074
rect 676246 490033 676298 490039
rect 676258 489991 676286 490033
rect 676244 489982 676300 489991
rect 676150 489943 676202 489949
rect 676244 489917 676300 489926
rect 676150 489885 676202 489891
rect 676354 489801 676382 490065
rect 676342 489795 676394 489801
rect 676342 489737 676394 489743
rect 676052 488354 676108 488363
rect 676052 488289 676108 488298
rect 676066 488173 676094 488289
rect 676054 488167 676106 488173
rect 676054 488109 676106 488115
rect 675284 487910 675340 487919
rect 675284 487845 675340 487854
rect 674902 486687 674954 486693
rect 674902 486629 674954 486635
rect 674614 483801 674666 483807
rect 674614 483743 674666 483749
rect 674230 483727 674282 483733
rect 674230 483669 674282 483675
rect 673846 480841 673898 480847
rect 673846 480783 673898 480789
rect 673750 480471 673802 480477
rect 673750 480413 673802 480419
rect 673654 480101 673706 480107
rect 673654 480043 673706 480049
rect 675298 429195 675326 487845
rect 676244 487170 676300 487179
rect 676546 487137 676574 530913
rect 676642 488173 676670 531949
rect 676738 489251 676766 532985
rect 679796 523578 679852 523587
rect 679796 523513 679852 523522
rect 679810 522995 679838 523513
rect 679796 522986 679852 522995
rect 679796 522921 679852 522930
rect 685460 522986 685516 522995
rect 685460 522921 685516 522930
rect 679810 521325 679838 522921
rect 685474 522551 685502 522921
rect 685460 522542 685516 522551
rect 685460 522477 685516 522486
rect 679798 521319 679850 521325
rect 679798 521261 679850 521267
rect 676724 489242 676780 489251
rect 676724 489177 676780 489186
rect 676724 488650 676780 488659
rect 676724 488585 676780 488594
rect 676630 488167 676682 488173
rect 676630 488109 676682 488115
rect 676244 487105 676246 487114
rect 676298 487105 676300 487114
rect 676534 487131 676586 487137
rect 676246 487073 676298 487079
rect 676534 487073 676586 487079
rect 676054 486687 676106 486693
rect 676054 486629 676106 486635
rect 675958 486613 676010 486619
rect 675958 486555 676010 486561
rect 675970 485847 675998 486555
rect 675956 485838 676012 485847
rect 675956 485773 676012 485782
rect 676066 484367 676094 486629
rect 676246 486539 676298 486545
rect 676246 486481 676298 486487
rect 676258 485107 676286 486481
rect 676244 485098 676300 485107
rect 676244 485033 676300 485042
rect 676052 484358 676108 484367
rect 676052 484293 676108 484302
rect 676054 483801 676106 483807
rect 675956 483766 676012 483775
rect 676054 483743 676106 483749
rect 675956 483701 675958 483710
rect 676010 483701 676012 483710
rect 675958 483669 676010 483675
rect 676066 482295 676094 483743
rect 676052 482286 676108 482295
rect 676052 482221 676108 482230
rect 676054 481951 676106 481957
rect 676052 481916 676054 481925
rect 676106 481916 676108 481925
rect 676052 481851 676108 481860
rect 676246 481581 676298 481587
rect 676244 481546 676246 481555
rect 676298 481546 676300 481555
rect 676244 481481 676300 481490
rect 676054 480841 676106 480847
rect 676052 480806 676054 480815
rect 676106 480806 676108 480815
rect 676052 480741 676108 480750
rect 676054 480471 676106 480477
rect 676052 480436 676054 480445
rect 676106 480436 676108 480445
rect 676052 480371 676108 480380
rect 676246 480101 676298 480107
rect 676244 480066 676246 480075
rect 676298 480066 676300 480075
rect 676244 480001 676300 480010
rect 676630 479287 676682 479293
rect 676630 479229 676682 479235
rect 673846 429189 673898 429195
rect 673846 429131 673898 429137
rect 675286 429189 675338 429195
rect 675286 429131 675338 429137
rect 673366 400403 673418 400409
rect 673366 400345 673418 400351
rect 672502 400181 672554 400187
rect 672502 400123 672554 400129
rect 672514 277939 672542 400123
rect 673078 398035 673130 398041
rect 673078 397977 673130 397983
rect 673090 357134 673118 397977
rect 673174 395593 673226 395599
rect 673174 395535 673226 395541
rect 673186 372141 673214 395535
rect 673270 385899 673322 385905
rect 673270 385841 673322 385847
rect 673174 372135 673226 372141
rect 673174 372077 673226 372083
rect 672802 357106 673118 357134
rect 672598 354449 672650 354455
rect 672598 354391 672650 354397
rect 672502 277933 672554 277939
rect 672502 277875 672554 277881
rect 672404 276270 672460 276279
rect 672404 276205 672460 276214
rect 670196 274346 670252 274355
rect 670196 274281 670252 274290
rect 672610 273467 672638 354391
rect 672802 353937 672830 357106
rect 673282 354825 673310 385841
rect 673378 356231 673406 400345
rect 673858 400187 673886 429131
rect 676148 402366 676204 402375
rect 676148 402301 676204 402310
rect 676052 401626 676108 401635
rect 676052 401561 676108 401570
rect 676066 400483 676094 401561
rect 676162 400631 676190 402301
rect 676244 401774 676300 401783
rect 676244 401709 676300 401718
rect 676150 400625 676202 400631
rect 676150 400567 676202 400573
rect 676258 400557 676286 401709
rect 676246 400551 676298 400557
rect 676246 400493 676298 400499
rect 676054 400477 676106 400483
rect 676054 400419 676106 400425
rect 676244 400442 676300 400451
rect 676244 400377 676246 400386
rect 676298 400377 676300 400386
rect 676246 400345 676298 400351
rect 673846 400181 673898 400187
rect 676054 400181 676106 400187
rect 673846 400123 673898 400129
rect 676052 400146 676054 400155
rect 676106 400146 676108 400155
rect 676052 400081 676108 400090
rect 676052 399702 676108 399711
rect 676052 399637 676108 399646
rect 675956 398666 676012 398675
rect 675956 398601 676012 398610
rect 675970 398041 675998 398601
rect 675958 398035 676010 398041
rect 675958 397977 676010 397983
rect 675190 397961 675242 397967
rect 675190 397903 675242 397909
rect 674518 397739 674570 397745
rect 674518 397681 674570 397687
rect 674530 385905 674558 397681
rect 675202 397454 675230 397903
rect 676066 397745 676094 399637
rect 676642 399415 676670 479229
rect 676738 401043 676766 488585
rect 679700 486578 679756 486587
rect 679700 486513 679756 486522
rect 679714 479293 679742 486513
rect 679702 479287 679754 479293
rect 679702 479229 679754 479235
rect 679892 479178 679948 479187
rect 679892 479113 679948 479122
rect 679906 478595 679934 479113
rect 679700 478586 679756 478595
rect 679700 478521 679756 478530
rect 679892 478586 679948 478595
rect 679892 478521 679948 478530
rect 679714 478151 679742 478521
rect 679906 478183 679934 478521
rect 679894 478177 679946 478183
rect 679700 478142 679756 478151
rect 679894 478119 679946 478125
rect 679700 478077 679756 478086
rect 676724 401034 676780 401043
rect 676724 400969 676780 400978
rect 676628 399406 676684 399415
rect 676628 399341 676684 399350
rect 676642 397967 676670 399341
rect 676630 397961 676682 397967
rect 676630 397903 676682 397909
rect 676054 397739 676106 397745
rect 676054 397681 676106 397687
rect 675010 397426 675230 397454
rect 674518 385899 674570 385905
rect 674518 385841 674570 385847
rect 675010 381613 675038 397426
rect 676052 395632 676108 395641
rect 676052 395567 676054 395576
rect 676106 395567 676108 395576
rect 676054 395535 676106 395541
rect 679796 390970 679852 390979
rect 679796 390905 679852 390914
rect 679810 390387 679838 390905
rect 679796 390378 679852 390387
rect 679796 390313 679852 390322
rect 685460 390378 685516 390387
rect 685460 390313 685516 390322
rect 679810 388865 679838 390313
rect 685474 389943 685502 390313
rect 685460 389934 685516 389943
rect 685460 389869 685516 389878
rect 679798 388859 679850 388865
rect 679798 388801 679850 388807
rect 675106 386266 675408 386294
rect 675106 381687 675134 386266
rect 675188 385938 675244 385947
rect 675188 385873 675244 385882
rect 675202 385737 675230 385873
rect 675202 385709 675408 385737
rect 675764 385642 675820 385651
rect 675764 385577 675820 385586
rect 675778 385096 675806 385577
rect 675764 384902 675820 384911
rect 675764 384837 675820 384846
rect 675778 384430 675806 384837
rect 675764 382978 675820 382987
rect 675764 382913 675820 382922
rect 675778 382580 675806 382913
rect 675476 382386 675532 382395
rect 675476 382321 675532 382330
rect 675490 382062 675518 382321
rect 675764 381794 675820 381803
rect 675764 381729 675820 381738
rect 675094 381681 675146 381687
rect 675094 381623 675146 381629
rect 674998 381607 675050 381613
rect 674998 381549 675050 381555
rect 675778 381396 675806 381729
rect 675572 381202 675628 381211
rect 675572 381137 675628 381146
rect 675586 380730 675614 381137
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675764 378094 675820 378103
rect 675764 378029 675820 378038
rect 675778 377696 675806 378029
rect 675380 377206 675436 377215
rect 675380 377141 675436 377150
rect 675394 377075 675422 377141
rect 675476 376762 675532 376771
rect 675476 376697 675532 376706
rect 675490 376438 675518 376697
rect 675764 375726 675820 375735
rect 675764 375661 675820 375670
rect 675778 375254 675806 375661
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675382 372135 675434 372141
rect 675382 372077 675434 372083
rect 675394 371554 675422 372077
rect 676244 357226 676300 357235
rect 676244 357161 676246 357170
rect 676298 357161 676300 357170
rect 676246 357129 676298 357135
rect 676148 356782 676204 356791
rect 676148 356717 676204 356726
rect 676052 356412 676108 356421
rect 676052 356347 676108 356356
rect 673366 356225 673418 356231
rect 673366 356167 673418 356173
rect 675956 354858 676012 354867
rect 673270 354819 673322 354825
rect 675956 354793 675958 354802
rect 673270 354761 673322 354767
rect 676010 354793 676012 354802
rect 675958 354761 676010 354767
rect 673282 354455 673310 354761
rect 673270 354449 673322 354455
rect 673270 354391 673322 354397
rect 676066 354381 676094 356347
rect 676054 354375 676106 354381
rect 676054 354317 676106 354323
rect 676162 354307 676190 356717
rect 676246 356225 676298 356231
rect 676244 356190 676246 356199
rect 676298 356190 676300 356199
rect 676244 356125 676300 356134
rect 676150 354301 676202 354307
rect 676150 354243 676202 354249
rect 676052 353970 676108 353979
rect 672790 353931 672842 353937
rect 676052 353905 676054 353914
rect 672790 353873 672842 353879
rect 676106 353905 676108 353914
rect 676054 353873 676106 353879
rect 672802 273615 672830 353873
rect 676916 352194 676972 352203
rect 676916 352129 676972 352138
rect 675572 351898 675628 351907
rect 675572 351833 675628 351842
rect 674422 348677 674474 348683
rect 674422 348619 674474 348625
rect 674434 336621 674462 348619
rect 675286 348603 675338 348609
rect 675286 348545 675338 348551
rect 675190 348529 675242 348535
rect 675190 348471 675242 348477
rect 674806 347567 674858 347573
rect 674806 347509 674858 347515
rect 674422 336615 674474 336621
rect 674422 336557 674474 336563
rect 674818 332255 674846 347509
rect 674902 345791 674954 345797
rect 674902 345733 674954 345739
rect 674806 332249 674858 332255
rect 674806 332191 674858 332197
rect 674914 331811 674942 345733
rect 674998 345717 675050 345723
rect 674998 345659 675050 345665
rect 675010 332773 675038 345659
rect 675094 345643 675146 345649
rect 675094 345585 675146 345591
rect 675106 336103 675134 345585
rect 675202 337287 675230 348471
rect 675298 339896 675326 348545
rect 675586 348494 675614 351833
rect 676820 350270 676876 350279
rect 676820 350205 676876 350214
rect 676244 349826 676300 349835
rect 676244 349761 676300 349770
rect 676052 349530 676108 349539
rect 676052 349465 676108 349474
rect 675956 348938 676012 348947
rect 675956 348873 676012 348882
rect 675970 348683 675998 348873
rect 675958 348677 676010 348683
rect 675958 348619 676010 348625
rect 676066 348535 676094 349465
rect 676258 348609 676286 349761
rect 676246 348603 676298 348609
rect 676246 348545 676298 348551
rect 676054 348529 676106 348535
rect 675586 348466 675806 348494
rect 676054 348471 676106 348477
rect 675778 341431 675806 348466
rect 676052 347976 676108 347985
rect 676052 347911 676108 347920
rect 676066 347573 676094 347911
rect 676054 347567 676106 347573
rect 676054 347509 676106 347515
rect 676052 347458 676108 347467
rect 676052 347393 676108 347402
rect 676066 345649 676094 347393
rect 676244 346866 676300 346875
rect 676244 346801 676300 346810
rect 676148 346274 676204 346283
rect 676148 346209 676204 346218
rect 676162 345797 676190 346209
rect 676150 345791 676202 345797
rect 676150 345733 676202 345739
rect 676258 345723 676286 346801
rect 676246 345717 676298 345723
rect 676246 345659 676298 345665
rect 676054 345643 676106 345649
rect 676054 345585 676106 345591
rect 676834 343027 676862 350205
rect 676820 343018 676876 343027
rect 676820 342953 676876 342962
rect 676930 342879 676958 352129
rect 679700 345682 679756 345691
rect 679700 345617 679756 345626
rect 679714 345247 679742 345617
rect 679700 345238 679756 345247
rect 679700 345173 679756 345182
rect 685460 345238 685516 345247
rect 685460 345173 685516 345182
rect 676916 342870 676972 342879
rect 676916 342805 676972 342814
rect 679714 342763 679742 345173
rect 685474 344803 685502 345173
rect 685460 344794 685516 344803
rect 685460 344729 685516 344738
rect 679702 342757 679754 342763
rect 679702 342699 679754 342705
rect 675766 341425 675818 341431
rect 675766 341367 675818 341373
rect 675490 340691 675518 341066
rect 675766 340759 675818 340765
rect 675766 340701 675818 340707
rect 675478 340685 675530 340691
rect 675478 340627 675530 340633
rect 675778 340548 675806 340701
rect 675298 339868 675408 339896
rect 675764 339614 675820 339623
rect 675764 339549 675820 339558
rect 675778 339216 675806 339549
rect 675764 337838 675820 337847
rect 675764 337773 675820 337782
rect 675778 337395 675806 337773
rect 675190 337281 675242 337287
rect 675190 337223 675242 337229
rect 675478 337281 675530 337287
rect 675478 337223 675530 337229
rect 675490 336848 675518 337223
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675394 336182 675422 336557
rect 675094 336097 675146 336103
rect 675094 336039 675146 336045
rect 675382 336097 675434 336103
rect 675382 336039 675434 336045
rect 675394 335555 675422 336039
rect 675380 333546 675436 333555
rect 675380 333481 675436 333490
rect 675394 333074 675422 333481
rect 674998 332767 675050 332773
rect 674998 332709 675050 332715
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675478 332249 675530 332255
rect 675478 332191 675530 332197
rect 675490 331890 675518 332191
rect 674902 331805 674954 331811
rect 674902 331747 674954 331753
rect 675382 331805 675434 331811
rect 675382 331747 675434 331753
rect 675394 331224 675422 331747
rect 675572 330586 675628 330595
rect 675572 330521 675628 330530
rect 675586 330040 675614 330521
rect 675778 328079 675806 328190
rect 675764 328070 675820 328079
rect 675764 328005 675820 328014
rect 675764 326886 675820 326895
rect 675764 326821 675820 326830
rect 675778 326340 675806 326821
rect 676340 312234 676396 312243
rect 676340 312169 676396 312178
rect 676148 311642 676204 311651
rect 676148 311577 676204 311586
rect 676162 311165 676190 311577
rect 676246 311233 676298 311239
rect 676244 311198 676246 311207
rect 676298 311198 676300 311207
rect 676150 311159 676202 311165
rect 676244 311133 676300 311142
rect 676150 311101 676202 311107
rect 676354 311091 676382 312169
rect 676342 311085 676394 311091
rect 676342 311027 676394 311033
rect 676052 308016 676108 308025
rect 676052 307951 676108 307960
rect 676066 305393 676094 307951
rect 676244 306758 676300 306767
rect 676244 306693 676300 306702
rect 674614 305387 674666 305393
rect 674614 305329 674666 305335
rect 676054 305387 676106 305393
rect 676054 305329 676106 305335
rect 674230 302649 674282 302655
rect 674230 302591 674282 302597
rect 674242 291629 674270 302591
rect 674422 302575 674474 302581
rect 674422 302517 674474 302523
rect 674326 299689 674378 299695
rect 674326 299631 674378 299637
rect 674230 291623 674282 291629
rect 674230 291565 674282 291571
rect 674338 287781 674366 299631
rect 674434 292295 674462 302517
rect 674626 294811 674654 305329
rect 676258 305319 676286 306693
rect 676916 305722 676972 305731
rect 676916 305657 676972 305666
rect 675094 305313 675146 305319
rect 675094 305255 675146 305261
rect 676246 305313 676298 305319
rect 676246 305255 676298 305261
rect 674710 302501 674762 302507
rect 674710 302443 674762 302449
rect 674722 295477 674750 302443
rect 674902 302427 674954 302433
rect 674902 302369 674954 302375
rect 674710 295471 674762 295477
rect 674710 295413 674762 295419
rect 674614 294805 674666 294811
rect 674614 294747 674666 294753
rect 674422 292289 674474 292295
rect 674422 292231 674474 292237
rect 674914 291111 674942 302369
rect 674998 299615 675050 299621
rect 674998 299557 675050 299563
rect 674902 291105 674954 291111
rect 674902 291047 674954 291053
rect 674326 287775 674378 287781
rect 674326 287717 674378 287723
rect 675010 286819 675038 299557
rect 675106 295537 675134 305255
rect 676244 304834 676300 304843
rect 676244 304769 676300 304778
rect 676052 304464 676108 304473
rect 676052 304399 676108 304408
rect 675956 303946 676012 303955
rect 675956 303881 676012 303890
rect 675970 302655 675998 303881
rect 675958 302649 676010 302655
rect 675958 302591 676010 302597
rect 676066 302581 676094 304399
rect 676054 302575 676106 302581
rect 676054 302517 676106 302523
rect 676258 302507 676286 304769
rect 676820 303354 676876 303363
rect 676820 303289 676876 303298
rect 676246 302501 676298 302507
rect 676052 302466 676108 302475
rect 676246 302443 676298 302449
rect 676052 302401 676054 302410
rect 676106 302401 676108 302410
rect 676054 302369 676106 302375
rect 676052 302022 676108 302031
rect 676052 301957 676108 301966
rect 676066 299695 676094 301957
rect 676244 301282 676300 301291
rect 676244 301217 676300 301226
rect 676054 299689 676106 299695
rect 676054 299631 676106 299637
rect 676258 299621 676286 301217
rect 676246 299615 676298 299621
rect 676246 299557 676298 299563
rect 676834 299219 676862 303289
rect 676820 299210 676876 299219
rect 676820 299145 676876 299154
rect 676930 298775 676958 305657
rect 679988 300690 680044 300699
rect 679988 300625 680044 300634
rect 680002 300255 680030 300625
rect 679796 300246 679852 300255
rect 679796 300181 679852 300190
rect 679988 300246 680044 300255
rect 679988 300181 680044 300190
rect 679810 299811 679838 300181
rect 679796 299802 679852 299811
rect 680002 299769 680030 300181
rect 679796 299737 679852 299746
rect 679990 299763 680042 299769
rect 679990 299705 680042 299711
rect 676916 298766 676972 298775
rect 676916 298701 676972 298710
rect 675380 296694 675436 296703
rect 675380 296629 675436 296638
rect 675394 296074 675422 296629
rect 675106 295509 675408 295537
rect 675094 295471 675146 295477
rect 675094 295413 675146 295419
rect 675106 294904 675134 295413
rect 675106 294876 675408 294904
rect 675094 294805 675146 294811
rect 675094 294747 675146 294753
rect 675106 294238 675134 294747
rect 675106 294210 675408 294238
rect 675380 292846 675436 292855
rect 675380 292781 675436 292790
rect 675394 292374 675422 292781
rect 675478 292289 675530 292295
rect 675478 292231 675530 292237
rect 675490 291856 675518 292231
rect 675382 291623 675434 291629
rect 675382 291565 675434 291571
rect 675394 291190 675422 291565
rect 675382 291105 675434 291111
rect 675382 291047 675434 291053
rect 675394 290555 675422 291047
rect 675476 288554 675532 288563
rect 675476 288489 675532 288498
rect 675490 288082 675518 288489
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675476 287370 675532 287379
rect 675476 287305 675532 287314
rect 675490 286898 675518 287305
rect 674998 286813 675050 286819
rect 674998 286755 675050 286761
rect 675382 286813 675434 286819
rect 675382 286755 675434 286761
rect 675394 286232 675422 286755
rect 675668 285298 675724 285307
rect 675668 285233 675724 285242
rect 675682 285048 675710 285233
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675764 281894 675820 281903
rect 675764 281829 675820 281838
rect 675778 281348 675806 281829
rect 675284 278490 675340 278499
rect 675284 278425 675340 278434
rect 675298 276533 675326 278425
rect 675764 278342 675820 278351
rect 675764 278277 675820 278286
rect 675778 276681 675806 278277
rect 675766 276675 675818 276681
rect 675766 276617 675818 276623
rect 679798 276675 679850 276681
rect 679798 276617 679850 276623
rect 675286 276527 675338 276533
rect 675286 276469 675338 276475
rect 679702 276527 679754 276533
rect 679702 276469 679754 276475
rect 672788 273606 672844 273615
rect 672788 273541 672844 273550
rect 672596 273458 672652 273467
rect 672596 273393 672652 273402
rect 670004 270646 670060 270655
rect 670004 270581 670060 270590
rect 676340 267242 676396 267251
rect 676340 267177 676396 267186
rect 672788 267094 672844 267103
rect 672788 267029 672844 267038
rect 672596 266946 672652 266955
rect 672596 266881 672652 266890
rect 672404 266798 672460 266807
rect 672404 266733 672460 266742
rect 671828 266502 671884 266511
rect 671828 266437 671884 266446
rect 671842 265063 671870 266437
rect 671830 265057 671882 265063
rect 671830 264999 671882 265005
rect 669814 264983 669866 264989
rect 669814 264925 669866 264931
rect 669622 264909 669674 264915
rect 669622 264851 669674 264857
rect 668180 263542 668236 263551
rect 668180 263477 668236 263486
rect 665302 115281 665354 115287
rect 665302 115223 665354 115229
rect 663766 115207 663818 115213
rect 663766 115149 663818 115155
rect 665206 115207 665258 115213
rect 665206 115149 665258 115155
rect 646580 113174 646636 113183
rect 646580 113109 646636 113118
rect 186164 107846 186220 107855
rect 186164 107781 186220 107790
rect 184340 107106 184396 107115
rect 184340 107041 184396 107050
rect 184534 106549 184586 106555
rect 184534 106491 184586 106497
rect 184342 106475 184394 106481
rect 184342 106417 184394 106423
rect 184354 106375 184382 106417
rect 184340 106366 184396 106375
rect 184340 106301 184396 106310
rect 184438 106327 184490 106333
rect 184438 106269 184490 106275
rect 184450 104895 184478 106269
rect 184546 105635 184574 106491
rect 184630 106401 184682 106407
rect 184630 106343 184682 106349
rect 184532 105626 184588 105635
rect 184532 105561 184588 105570
rect 184436 104886 184492 104895
rect 184436 104821 184492 104830
rect 184642 104007 184670 106343
rect 645716 106070 645772 106079
rect 645716 106005 645772 106014
rect 184726 105143 184778 105149
rect 184726 105085 184778 105091
rect 184628 103998 184684 104007
rect 184628 103933 184684 103942
rect 184438 103663 184490 103669
rect 184438 103605 184490 103611
rect 184342 103589 184394 103595
rect 184342 103531 184394 103537
rect 184354 103415 184382 103531
rect 184340 103406 184396 103415
rect 184340 103341 184396 103350
rect 184450 102527 184478 103605
rect 184534 103515 184586 103521
rect 184534 103457 184586 103463
rect 184436 102518 184492 102527
rect 184436 102453 184492 102462
rect 184546 101047 184574 103457
rect 184738 101935 184766 105085
rect 645730 103743 645758 106005
rect 645718 103737 645770 103743
rect 645718 103679 645770 103685
rect 645140 102222 645196 102231
rect 645140 102157 645196 102166
rect 645154 102115 645182 102157
rect 645142 102109 645194 102115
rect 645142 102051 645194 102057
rect 184724 101926 184780 101935
rect 184724 101861 184780 101870
rect 184532 101038 184588 101047
rect 184532 100973 184588 100982
rect 184534 100777 184586 100783
rect 184534 100719 184586 100725
rect 184342 100629 184394 100635
rect 184342 100571 184394 100577
rect 184354 100307 184382 100571
rect 184438 100555 184490 100561
rect 184438 100497 184490 100503
rect 184340 100298 184396 100307
rect 184340 100233 184396 100242
rect 184450 99567 184478 100497
rect 184436 99558 184492 99567
rect 184436 99493 184492 99502
rect 184546 98679 184574 100719
rect 184630 100703 184682 100709
rect 184630 100645 184682 100651
rect 184532 98670 184588 98679
rect 184532 98605 184588 98614
rect 184642 98087 184670 100645
rect 184628 98078 184684 98087
rect 184246 98039 184298 98045
rect 184628 98013 184684 98022
rect 184246 97981 184298 97987
rect 182902 94709 182954 94715
rect 182902 94651 182954 94657
rect 184258 81955 184286 97981
rect 186166 97965 186218 97971
rect 186166 97907 186218 97913
rect 184342 97891 184394 97897
rect 184342 97833 184394 97839
rect 184354 97199 184382 97833
rect 184438 97817 184490 97823
rect 184438 97759 184490 97765
rect 184340 97190 184396 97199
rect 184340 97125 184396 97134
rect 184450 96459 184478 97759
rect 184534 97743 184586 97749
rect 184534 97685 184586 97691
rect 184436 96450 184492 96459
rect 184436 96385 184492 96394
rect 184546 95719 184574 97685
rect 184532 95710 184588 95719
rect 184532 95645 184588 95654
rect 184340 94970 184396 94979
rect 184340 94905 184342 94914
rect 184394 94905 184396 94914
rect 184342 94873 184394 94879
rect 184342 94783 184394 94789
rect 184342 94725 184394 94731
rect 184354 93499 184382 94725
rect 184630 94635 184682 94641
rect 184630 94577 184682 94583
rect 184340 93490 184396 93499
rect 184340 93425 184396 93434
rect 184642 92759 184670 94577
rect 184628 92750 184684 92759
rect 184628 92685 184684 92694
rect 184630 92119 184682 92125
rect 184630 92061 184682 92067
rect 184534 92045 184586 92051
rect 184534 91987 184586 91993
rect 184438 91971 184490 91977
rect 184438 91913 184490 91919
rect 184342 91897 184394 91903
rect 184340 91862 184342 91871
rect 184394 91862 184396 91871
rect 184340 91797 184396 91806
rect 184450 91131 184478 91913
rect 184436 91122 184492 91131
rect 184436 91057 184492 91066
rect 184546 90391 184574 91987
rect 184532 90382 184588 90391
rect 184532 90317 184588 90326
rect 184642 89651 184670 92061
rect 184628 89642 184684 89651
rect 184628 89577 184684 89586
rect 184630 89233 184682 89239
rect 184630 89175 184682 89181
rect 184534 89159 184586 89165
rect 184534 89101 184586 89107
rect 184438 89085 184490 89091
rect 184438 89027 184490 89033
rect 184342 89011 184394 89017
rect 184342 88953 184394 88959
rect 184354 88911 184382 88953
rect 184340 88902 184396 88911
rect 184340 88837 184396 88846
rect 184450 88171 184478 89027
rect 184436 88162 184492 88171
rect 184436 88097 184492 88106
rect 184546 87283 184574 89101
rect 184532 87274 184588 87283
rect 184532 87209 184588 87218
rect 184642 86691 184670 89175
rect 184628 86682 184684 86691
rect 184628 86617 184684 86626
rect 184438 86421 184490 86427
rect 184438 86363 184490 86369
rect 184342 86273 184394 86279
rect 184342 86215 184394 86221
rect 184354 85211 184382 86215
rect 184450 85803 184478 86363
rect 184534 86347 184586 86353
rect 184534 86289 184586 86295
rect 184436 85794 184492 85803
rect 184436 85729 184492 85738
rect 184340 85202 184396 85211
rect 184340 85137 184396 85146
rect 184546 84323 184574 86289
rect 184532 84314 184588 84323
rect 184532 84249 184588 84258
rect 184438 83535 184490 83541
rect 184438 83477 184490 83483
rect 184342 83461 184394 83467
rect 184340 83426 184342 83435
rect 184394 83426 184396 83435
rect 184340 83361 184396 83370
rect 184244 81946 184300 81955
rect 184244 81881 184300 81890
rect 184450 81363 184478 83477
rect 186178 82843 186206 97907
rect 645428 96006 645484 96015
rect 645428 95941 645430 95950
rect 645482 95941 645484 95950
rect 645430 95909 645482 95915
rect 186262 94709 186314 94715
rect 186262 94651 186314 94657
rect 186274 94239 186302 94651
rect 186260 94230 186316 94239
rect 186260 94165 186316 94174
rect 645526 92415 645578 92421
rect 645526 92357 645578 92363
rect 186164 82834 186220 82843
rect 186164 82769 186220 82778
rect 184436 81354 184492 81363
rect 184436 81289 184492 81298
rect 184438 80649 184490 80655
rect 184438 80591 184490 80597
rect 184342 80501 184394 80507
rect 184342 80443 184394 80449
rect 180022 80427 180074 80433
rect 180022 80369 180074 80375
rect 184354 78995 184382 80443
rect 184450 79883 184478 80591
rect 184534 80575 184586 80581
rect 184534 80517 184586 80523
rect 184436 79874 184492 79883
rect 184436 79809 184492 79818
rect 184340 78986 184396 78995
rect 184340 78921 184396 78930
rect 184546 78255 184574 80517
rect 184628 80466 184684 80475
rect 184628 80401 184630 80410
rect 184682 80401 184684 80410
rect 184630 80369 184682 80375
rect 645538 79439 645566 92357
rect 646486 92341 646538 92347
rect 646486 92283 646538 92289
rect 645908 88902 645964 88911
rect 645908 88837 645964 88846
rect 645922 87537 645950 88837
rect 645910 87531 645962 87537
rect 645910 87473 645962 87479
rect 645908 84462 645964 84471
rect 645908 84397 645964 84406
rect 645922 84207 645950 84397
rect 645910 84201 645962 84207
rect 645910 84143 645962 84149
rect 645524 79430 645580 79439
rect 645524 79365 645580 79374
rect 184532 78246 184588 78255
rect 184532 78181 184588 78190
rect 184342 77763 184394 77769
rect 184342 77705 184394 77711
rect 156406 77541 156458 77547
rect 184354 77515 184382 77705
rect 184438 77689 184490 77695
rect 184438 77631 184490 77637
rect 156406 77483 156458 77489
rect 184340 77506 184396 77515
rect 184340 77441 184396 77450
rect 184450 76775 184478 77631
rect 184534 77615 184586 77621
rect 184534 77557 184586 77563
rect 184436 76766 184492 76775
rect 184436 76701 184492 76710
rect 184546 76035 184574 77557
rect 184630 77541 184682 77547
rect 184630 77483 184682 77489
rect 184532 76026 184588 76035
rect 184532 75961 184588 75970
rect 184642 75147 184670 77483
rect 646006 76135 646058 76141
rect 646006 76077 646058 76083
rect 646018 75591 646046 76077
rect 646004 75582 646060 75591
rect 646004 75517 646060 75526
rect 184628 75138 184684 75147
rect 184628 75073 184684 75082
rect 184534 74877 184586 74883
rect 184534 74819 184586 74825
rect 184438 74729 184490 74735
rect 184438 74671 184490 74677
rect 154102 74655 154154 74661
rect 154102 74597 154154 74603
rect 184342 74655 184394 74661
rect 184342 74597 184394 74603
rect 184354 74407 184382 74597
rect 184340 74398 184396 74407
rect 184340 74333 184396 74342
rect 184450 72927 184478 74671
rect 184546 73667 184574 74819
rect 184630 74803 184682 74809
rect 184630 74745 184682 74751
rect 184532 73658 184588 73667
rect 184532 73593 184588 73602
rect 184436 72918 184492 72927
rect 184436 72853 184492 72862
rect 184642 72187 184670 74745
rect 184628 72178 184684 72187
rect 184628 72113 184684 72122
rect 184438 71991 184490 71997
rect 184438 71933 184490 71939
rect 149686 71917 149738 71923
rect 149686 71859 149738 71865
rect 149590 71843 149642 71849
rect 149590 71785 149642 71791
rect 184342 71843 184394 71849
rect 184342 71785 184394 71791
rect 149506 70952 149630 70980
rect 149492 70846 149548 70855
rect 149492 70781 149548 70790
rect 149396 69514 149452 69523
rect 149396 69449 149452 69458
rect 149302 68883 149354 68889
rect 149302 68825 149354 68831
rect 149204 68330 149260 68339
rect 149204 68265 149260 68274
rect 149110 66219 149162 66225
rect 149110 66161 149162 66167
rect 149014 65997 149066 66003
rect 149014 65939 149066 65945
rect 149218 63191 149246 68265
rect 149410 66151 149438 69449
rect 149398 66145 149450 66151
rect 149398 66087 149450 66093
rect 149506 66077 149534 70781
rect 149602 68963 149630 70952
rect 184354 70559 184382 71785
rect 184450 71447 184478 71933
rect 184534 71917 184586 71923
rect 184534 71859 184586 71865
rect 184436 71438 184492 71447
rect 184436 71373 184492 71382
rect 184340 70550 184396 70559
rect 184340 70485 184396 70494
rect 184546 69967 184574 71859
rect 184532 69958 184588 69967
rect 184532 69893 184588 69902
rect 184342 69105 184394 69111
rect 184340 69070 184342 69079
rect 184394 69070 184396 69079
rect 184340 69005 184396 69014
rect 184438 69031 184490 69037
rect 184438 68973 184490 68979
rect 149590 68957 149642 68963
rect 149590 68899 149642 68905
rect 184342 68957 184394 68963
rect 184342 68899 184394 68905
rect 184354 67599 184382 68899
rect 184450 68487 184478 68973
rect 184534 68883 184586 68889
rect 184534 68825 184586 68831
rect 184436 68478 184492 68487
rect 184436 68413 184492 68422
rect 184340 67590 184396 67599
rect 184340 67525 184396 67534
rect 149588 67146 149644 67155
rect 149588 67081 149644 67090
rect 149494 66071 149546 66077
rect 149494 66013 149546 66019
rect 149300 65370 149356 65379
rect 149300 65305 149356 65314
rect 149206 63185 149258 63191
rect 149206 63127 149258 63133
rect 149314 63117 149342 65305
rect 149396 64630 149452 64639
rect 149396 64565 149452 64574
rect 149410 63339 149438 64565
rect 149492 63446 149548 63455
rect 149492 63381 149548 63390
rect 149398 63333 149450 63339
rect 149398 63275 149450 63281
rect 149302 63111 149354 63117
rect 149302 63053 149354 63059
rect 149396 62262 149452 62271
rect 149396 62197 149452 62206
rect 149300 60634 149356 60643
rect 149300 60569 149356 60578
rect 149314 60305 149342 60569
rect 149410 60453 149438 62197
rect 149398 60447 149450 60453
rect 149398 60389 149450 60395
rect 149506 60379 149534 63381
rect 149602 63265 149630 67081
rect 184546 66859 184574 68825
rect 184532 66850 184588 66859
rect 184532 66785 184588 66794
rect 646004 66258 646060 66267
rect 184534 66219 184586 66225
rect 646004 66193 646006 66202
rect 184534 66161 184586 66167
rect 646058 66193 646060 66202
rect 646006 66161 646058 66167
rect 184340 66110 184396 66119
rect 184340 66045 184396 66054
rect 184438 66071 184490 66077
rect 184354 66003 184382 66045
rect 184438 66013 184490 66019
rect 184342 65997 184394 66003
rect 184342 65939 184394 65945
rect 184450 64639 184478 66013
rect 184546 65231 184574 66161
rect 184630 66145 184682 66151
rect 184630 66087 184682 66093
rect 184532 65222 184588 65231
rect 184532 65157 184588 65166
rect 184436 64630 184492 64639
rect 184436 64565 184492 64574
rect 184642 63751 184670 66087
rect 184628 63742 184684 63751
rect 184628 63677 184684 63686
rect 184630 63333 184682 63339
rect 184630 63275 184682 63281
rect 149590 63259 149642 63265
rect 149590 63201 149642 63207
rect 184534 63259 184586 63265
rect 184534 63201 184586 63207
rect 184342 63185 184394 63191
rect 184340 63150 184342 63159
rect 184394 63150 184396 63159
rect 184340 63085 184396 63094
rect 184438 63111 184490 63117
rect 184438 63053 184490 63059
rect 184450 61531 184478 63053
rect 184546 62271 184574 63201
rect 184532 62262 184588 62271
rect 184532 62197 184588 62206
rect 184436 61522 184492 61531
rect 184436 61457 184492 61466
rect 184642 60791 184670 63275
rect 184628 60782 184684 60791
rect 184628 60717 184684 60726
rect 184438 60447 184490 60453
rect 184438 60389 184490 60395
rect 149494 60373 149546 60379
rect 149494 60315 149546 60321
rect 184342 60373 184394 60379
rect 184342 60315 184394 60321
rect 149302 60299 149354 60305
rect 149302 60241 149354 60247
rect 184354 60051 184382 60315
rect 184340 60042 184396 60051
rect 184340 59977 184396 59986
rect 149396 59746 149452 59755
rect 149396 59681 149452 59690
rect 149410 59047 149438 59681
rect 184450 59311 184478 60389
rect 184534 60299 184586 60305
rect 184534 60241 184586 60247
rect 184436 59302 184492 59311
rect 184436 59237 184492 59246
rect 149398 59041 149450 59047
rect 149398 58983 149450 58989
rect 184342 59041 184394 59047
rect 184342 58983 184394 58989
rect 149396 58562 149452 58571
rect 149396 58497 149452 58506
rect 149410 57567 149438 58497
rect 184354 57683 184382 58983
rect 184546 58423 184574 60241
rect 646006 59115 646058 59121
rect 646006 59057 646058 59063
rect 646018 59015 646046 59057
rect 646004 59006 646060 59015
rect 646004 58941 646060 58950
rect 184532 58414 184588 58423
rect 184532 58349 184588 58358
rect 184340 57674 184396 57683
rect 184340 57609 184396 57618
rect 149398 57561 149450 57567
rect 149398 57503 149450 57509
rect 184342 57561 184394 57567
rect 184342 57503 184394 57509
rect 149492 57378 149548 57387
rect 149492 57313 149548 57322
rect 149398 56229 149450 56235
rect 149396 56194 149398 56203
rect 149450 56194 149452 56203
rect 149506 56161 149534 57313
rect 184354 56943 184382 57503
rect 184340 56934 184396 56943
rect 184340 56869 184396 56878
rect 184438 56229 184490 56235
rect 184340 56194 184396 56203
rect 149396 56129 149452 56138
rect 149494 56155 149546 56161
rect 184438 56171 184490 56177
rect 184340 56129 184342 56138
rect 149494 56097 149546 56103
rect 184394 56129 184396 56138
rect 184342 56097 184394 56103
rect 184450 55463 184478 56171
rect 184436 55454 184492 55463
rect 184436 55389 184492 55398
rect 149684 54862 149740 54871
rect 149684 54797 149740 54806
rect 149698 54681 149726 54797
rect 646498 54723 646526 92283
rect 646594 77695 646622 113109
rect 665218 112327 665246 115149
rect 665206 112321 665258 112327
rect 665206 112263 665258 112269
rect 647060 111398 647116 111407
rect 647060 111333 647116 111342
rect 646676 109474 646732 109483
rect 646676 109409 646732 109418
rect 646582 77689 646634 77695
rect 646582 77631 646634 77637
rect 646690 77621 646718 109409
rect 646772 107994 646828 108003
rect 646772 107929 646828 107938
rect 646786 92717 646814 107929
rect 646964 98078 647020 98087
rect 646964 98013 647020 98022
rect 646774 92711 646826 92717
rect 646774 92653 646826 92659
rect 646870 92267 646922 92273
rect 646870 92209 646922 92215
rect 646774 83609 646826 83615
rect 646774 83551 646826 83557
rect 646678 77615 646730 77621
rect 646678 77557 646730 77563
rect 646786 57091 646814 83551
rect 646882 68635 646910 92209
rect 646978 77769 647006 98013
rect 647074 87093 647102 111333
rect 665314 104895 665342 115223
rect 668194 106375 668222 263477
rect 670390 250701 670442 250707
rect 670390 250643 670442 250649
rect 670402 247673 670430 250643
rect 670390 247667 670442 247673
rect 670390 247609 670442 247615
rect 672418 174455 672446 266733
rect 672404 174446 672460 174455
rect 672404 174381 672460 174390
rect 672610 173567 672638 266881
rect 672802 218263 672830 267029
rect 672980 266650 673036 266659
rect 672980 266585 673036 266594
rect 676148 266650 676204 266659
rect 676148 266585 676204 266594
rect 672994 219299 673022 266585
rect 673460 266354 673516 266363
rect 673460 266289 673516 266298
rect 673270 265057 673322 265063
rect 673270 264999 673322 265005
rect 673282 259587 673310 264999
rect 673474 263403 673502 266289
rect 676162 265285 676190 266585
rect 676244 266206 676300 266215
rect 676244 266141 676300 266150
rect 676258 265433 676286 266141
rect 676246 265427 676298 265433
rect 676246 265369 676298 265375
rect 676150 265279 676202 265285
rect 676150 265221 676202 265227
rect 676354 265137 676382 267177
rect 679714 265179 679742 276469
rect 679700 265170 679756 265179
rect 676342 265131 676394 265137
rect 679700 265105 679756 265114
rect 676342 265073 676394 265079
rect 676246 265057 676298 265063
rect 676246 264999 676298 265005
rect 676258 264735 676286 264999
rect 676244 264726 676300 264735
rect 676244 264661 676300 264670
rect 679810 264291 679838 276617
rect 679796 264282 679852 264291
rect 679796 264217 679852 264226
rect 673460 263394 673516 263403
rect 673378 263352 673460 263380
rect 673270 259581 673322 259587
rect 673270 259523 673322 259529
rect 672980 219290 673036 219299
rect 672980 219225 673036 219234
rect 673378 218813 673406 263352
rect 673460 263329 673516 263338
rect 676244 262802 676300 262811
rect 676244 262737 676300 262746
rect 676258 262177 676286 262737
rect 676916 262210 676972 262219
rect 675190 262171 675242 262177
rect 675190 262113 675242 262119
rect 676246 262171 676298 262177
rect 676916 262145 676972 262154
rect 676246 262113 676298 262119
rect 674806 259951 674858 259957
rect 674806 259893 674858 259899
rect 673462 259581 673514 259587
rect 673462 259523 673514 259529
rect 673474 219923 673502 259523
rect 674710 259359 674762 259365
rect 674710 259301 674762 259307
rect 674614 256473 674666 256479
rect 674614 256415 674666 256421
rect 674626 242789 674654 256415
rect 674722 247694 674750 259301
rect 674818 247969 674846 259893
rect 674902 256399 674954 256405
rect 674902 256341 674954 256347
rect 674806 247963 674858 247969
rect 674806 247905 674858 247911
rect 674722 247666 674846 247694
rect 674818 247081 674846 247666
rect 674806 247075 674858 247081
rect 674806 247017 674858 247023
rect 674914 245897 674942 256341
rect 675202 249246 675230 262113
rect 676244 261322 676300 261331
rect 676244 261257 676300 261266
rect 676258 259957 676286 261257
rect 676820 260582 676876 260591
rect 676820 260517 676876 260526
rect 676246 259951 676298 259957
rect 676246 259893 676298 259899
rect 676244 259842 676300 259851
rect 676244 259777 676300 259786
rect 676052 259472 676108 259481
rect 676052 259407 676108 259416
rect 676066 259365 676094 259407
rect 676054 259359 676106 259365
rect 676054 259301 676106 259307
rect 676258 259291 676286 259777
rect 675286 259285 675338 259291
rect 675286 259227 675338 259233
rect 676246 259285 676298 259291
rect 676246 259227 676298 259233
rect 675298 250356 675326 259227
rect 676052 257474 676108 257483
rect 676052 257409 676108 257418
rect 675956 257030 676012 257039
rect 675956 256965 676012 256974
rect 675970 256479 675998 256965
rect 675958 256473 676010 256479
rect 675958 256415 676010 256421
rect 676066 256405 676094 257409
rect 676054 256399 676106 256405
rect 676054 256341 676106 256347
rect 676834 253339 676862 260517
rect 676820 253330 676876 253339
rect 676820 253265 676876 253274
rect 676930 253191 676958 262145
rect 679796 255698 679852 255707
rect 679796 255633 679852 255642
rect 679810 255263 679838 255633
rect 679796 255254 679852 255263
rect 679796 255189 679852 255198
rect 685556 255254 685612 255263
rect 685556 255189 685612 255198
rect 679810 253519 679838 255189
rect 685570 254819 685598 255189
rect 685556 254810 685612 254819
rect 685556 254745 685612 254754
rect 679798 253513 679850 253519
rect 679798 253455 679850 253461
rect 676916 253182 676972 253191
rect 676916 253117 676972 253126
rect 675394 250707 675422 251082
rect 675764 250814 675820 250823
rect 675764 250749 675820 250758
rect 675382 250701 675434 250707
rect 675382 250643 675434 250649
rect 675778 250523 675806 250749
rect 675298 250328 675518 250356
rect 675490 249898 675518 250328
rect 675202 249218 675408 249246
rect 675382 247963 675434 247969
rect 675382 247905 675434 247911
rect 675394 247382 675422 247905
rect 675478 247075 675530 247081
rect 675478 247017 675530 247023
rect 675490 246864 675518 247017
rect 675572 246670 675628 246679
rect 675572 246605 675628 246614
rect 675586 246198 675614 246605
rect 674902 245891 674954 245897
rect 674902 245833 674954 245839
rect 675382 245891 675434 245897
rect 675382 245833 675434 245839
rect 675394 245532 675422 245833
rect 675668 243562 675724 243571
rect 675668 243497 675724 243506
rect 675682 243090 675710 243497
rect 674614 242783 674666 242789
rect 674614 242725 674666 242731
rect 675382 242783 675434 242789
rect 675382 242725 675434 242731
rect 675394 242498 675422 242725
rect 675380 242082 675436 242091
rect 675380 242017 675436 242026
rect 675394 241875 675422 242017
rect 675476 241786 675532 241795
rect 675476 241721 675532 241730
rect 675490 241240 675518 241721
rect 675476 240602 675532 240611
rect 675476 240537 675532 240546
rect 675490 240056 675518 240537
rect 675764 238678 675820 238687
rect 675764 238613 675820 238622
rect 675778 238206 675806 238613
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 676244 222102 676300 222111
rect 676244 222037 676246 222046
rect 676298 222037 676300 222046
rect 676246 222005 676298 222011
rect 676244 221954 676300 221963
rect 676244 221889 676246 221898
rect 676298 221889 676300 221898
rect 676246 221857 676298 221863
rect 676052 221214 676108 221223
rect 676052 221149 676108 221158
rect 673462 219917 673514 219923
rect 673462 219859 673514 219865
rect 676066 219109 676094 221149
rect 676246 219917 676298 219923
rect 676244 219882 676246 219891
rect 676298 219882 676300 219891
rect 676244 219817 676300 219826
rect 676054 219103 676106 219109
rect 676054 219045 676106 219051
rect 673366 218807 673418 218813
rect 676054 218807 676106 218813
rect 673366 218749 673418 218755
rect 676052 218772 676054 218781
rect 676106 218772 676108 218781
rect 676052 218707 676108 218716
rect 672788 218254 672844 218263
rect 672788 218189 672844 218198
rect 677012 217070 677068 217079
rect 677012 217005 677068 217014
rect 675764 216774 675820 216783
rect 675764 216709 675820 216718
rect 675284 214850 675340 214859
rect 675284 214785 675340 214794
rect 674806 213257 674858 213263
rect 674806 213199 674858 213205
rect 674614 211925 674666 211931
rect 674614 211867 674666 211873
rect 674626 197057 674654 211867
rect 674710 210445 674762 210451
rect 674710 210387 674762 210393
rect 674614 197051 674666 197057
rect 674614 196993 674666 196999
rect 674722 196613 674750 210387
rect 674818 201349 674846 213199
rect 675094 213183 675146 213189
rect 675094 213125 675146 213131
rect 674902 210371 674954 210377
rect 674902 210313 674954 210319
rect 674806 201343 674858 201349
rect 674806 201285 674858 201291
rect 674914 197797 674942 210313
rect 674998 210297 675050 210303
rect 674998 210239 675050 210245
rect 675010 200905 675038 210239
rect 675106 205808 675134 213125
rect 675106 205780 675230 205808
rect 675094 205709 675146 205715
rect 675094 205651 675146 205657
rect 675106 201571 675134 205651
rect 675202 201941 675230 205780
rect 675298 204698 675326 214785
rect 675778 206159 675806 216709
rect 676916 214998 676972 215007
rect 676916 214933 676972 214942
rect 676244 214110 676300 214119
rect 676244 214045 676300 214054
rect 676052 213740 676108 213749
rect 676052 213675 676108 213684
rect 676066 213263 676094 213675
rect 676054 213257 676106 213263
rect 676054 213199 676106 213205
rect 676258 213189 676286 214045
rect 676246 213183 676298 213189
rect 676246 213125 676298 213131
rect 676820 213074 676876 213083
rect 676820 213009 676876 213018
rect 676052 212778 676108 212787
rect 676052 212713 676108 212722
rect 676066 211931 676094 212713
rect 676244 212038 676300 212047
rect 676244 211973 676300 211982
rect 676054 211925 676106 211931
rect 676054 211867 676106 211873
rect 676052 211816 676108 211825
rect 676052 211751 676108 211760
rect 675956 211298 676012 211307
rect 675956 211233 676012 211242
rect 675970 210451 675998 211233
rect 675958 210445 676010 210451
rect 675958 210387 676010 210393
rect 676066 210377 676094 211751
rect 676054 210371 676106 210377
rect 676054 210313 676106 210319
rect 676258 210303 676286 211973
rect 676246 210297 676298 210303
rect 676246 210239 676298 210245
rect 676834 207459 676862 213009
rect 676930 207607 676958 214933
rect 677026 207755 677054 217005
rect 679988 210558 680044 210567
rect 679988 210493 680044 210502
rect 680002 209975 680030 210493
rect 679796 209966 679852 209975
rect 679796 209901 679852 209910
rect 679988 209966 680044 209975
rect 679988 209901 680044 209910
rect 679810 209531 679838 209901
rect 679796 209522 679852 209531
rect 679796 209457 679852 209466
rect 677012 207746 677068 207755
rect 677012 207681 677068 207690
rect 676916 207598 676972 207607
rect 676916 207533 676972 207542
rect 676820 207450 676876 207459
rect 680002 207417 680030 209901
rect 676820 207385 676876 207394
rect 679990 207411 680042 207417
rect 679990 207353 680042 207359
rect 675766 206153 675818 206159
rect 675766 206095 675818 206101
rect 675490 205715 675518 205868
rect 675478 205709 675530 205715
rect 675478 205651 675530 205657
rect 675766 205635 675818 205641
rect 675766 205577 675818 205583
rect 675778 205350 675806 205577
rect 675298 204670 675408 204698
rect 675764 204490 675820 204499
rect 675764 204425 675820 204434
rect 675778 204018 675806 204425
rect 675668 202714 675724 202723
rect 675668 202649 675724 202658
rect 675682 202168 675710 202649
rect 675190 201935 675242 201941
rect 675190 201877 675242 201883
rect 675478 201935 675530 201941
rect 675478 201877 675530 201883
rect 675490 201650 675518 201877
rect 675094 201565 675146 201571
rect 675094 201507 675146 201513
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 674998 200899 675050 200905
rect 674998 200841 675050 200847
rect 675382 200899 675434 200905
rect 675382 200841 675434 200847
rect 675394 200355 675422 200841
rect 675572 198422 675628 198431
rect 675572 198357 675628 198366
rect 675586 197876 675614 198357
rect 674902 197791 674954 197797
rect 674902 197733 674954 197739
rect 675382 197791 675434 197797
rect 675382 197733 675434 197739
rect 675394 197319 675422 197733
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 674710 196607 674762 196613
rect 674710 196549 674762 196555
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675764 195314 675820 195323
rect 675764 195249 675820 195258
rect 675778 194842 675806 195249
rect 675764 193538 675820 193547
rect 675764 193473 675820 193482
rect 675778 192992 675806 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 676148 177406 676204 177415
rect 676148 177341 676204 177350
rect 676162 176189 676190 177341
rect 676340 176814 676396 176823
rect 676340 176749 676396 176758
rect 676244 176370 676300 176379
rect 676244 176305 676300 176314
rect 676150 176183 676202 176189
rect 676150 176125 676202 176131
rect 676258 176041 676286 176305
rect 676246 176035 676298 176041
rect 676246 175977 676298 175983
rect 676354 175893 676382 176749
rect 676342 175887 676394 175893
rect 676342 175829 676394 175835
rect 672596 173558 672652 173567
rect 672596 173493 672652 173502
rect 676916 172374 676972 172383
rect 676916 172309 676972 172318
rect 675572 172078 675628 172087
rect 675572 172013 675628 172022
rect 674806 170337 674858 170343
rect 674806 170279 674858 170285
rect 674710 166267 674762 166273
rect 674710 166209 674762 166215
rect 670390 160495 670442 160501
rect 670390 160437 670442 160443
rect 670402 155543 670430 160437
rect 670390 155537 670442 155543
rect 670390 155479 670442 155485
rect 674722 151473 674750 166209
rect 674818 157763 674846 170279
rect 675286 169967 675338 169973
rect 675286 169909 675338 169915
rect 674902 167747 674954 167753
rect 674902 167689 674954 167695
rect 674806 157757 674858 157763
rect 674806 157699 674858 157705
rect 674914 157097 674942 167689
rect 675190 167155 675242 167161
rect 675190 167097 675242 167103
rect 674998 167081 675050 167087
rect 675202 167054 675230 167097
rect 674998 167023 675050 167029
rect 675106 167026 675230 167054
rect 674902 157091 674954 157097
rect 674902 157033 674954 157039
rect 675010 155913 675038 167023
rect 675106 161294 675134 167026
rect 675106 161266 675230 161294
rect 675202 156579 675230 161266
rect 675298 159706 675326 169909
rect 675586 167054 675614 172013
rect 676052 171708 676108 171717
rect 676052 171643 676108 171652
rect 676066 170343 676094 171643
rect 676820 170450 676876 170459
rect 676820 170385 676876 170394
rect 676054 170337 676106 170343
rect 676054 170279 676106 170285
rect 676052 170228 676108 170237
rect 676052 170163 676108 170172
rect 676066 169973 676094 170163
rect 676054 169967 676106 169973
rect 676054 169909 676106 169915
rect 676052 169710 676108 169719
rect 676052 169645 676108 169654
rect 676066 167753 676094 169645
rect 676244 168970 676300 168979
rect 676244 168905 676300 168914
rect 676054 167747 676106 167753
rect 676054 167689 676106 167695
rect 676052 167638 676108 167647
rect 676052 167573 676108 167582
rect 676066 167087 676094 167573
rect 676258 167161 676286 168905
rect 676246 167155 676298 167161
rect 676246 167097 676298 167103
rect 676054 167081 676106 167087
rect 675586 167026 675710 167054
rect 675682 161167 675710 167026
rect 676054 167023 676106 167029
rect 676052 166676 676108 166685
rect 676052 166611 676108 166620
rect 676066 166273 676094 166611
rect 676054 166267 676106 166273
rect 676054 166209 676106 166215
rect 676052 166158 676108 166167
rect 676052 166093 676108 166102
rect 676066 164423 676094 166093
rect 676148 165418 676204 165427
rect 676148 165353 676204 165362
rect 676054 164417 676106 164423
rect 676054 164359 676106 164365
rect 676162 164275 676190 165353
rect 676244 164826 676300 164835
rect 676244 164761 676300 164770
rect 676258 164349 676286 164761
rect 676246 164343 676298 164349
rect 676246 164285 676298 164291
rect 676150 164269 676202 164275
rect 676150 164211 676202 164217
rect 676834 161431 676862 170385
rect 676930 161579 676958 172309
rect 676916 161570 676972 161579
rect 676916 161505 676972 161514
rect 676820 161422 676876 161431
rect 676820 161357 676876 161366
rect 675670 161161 675722 161167
rect 675670 161103 675722 161109
rect 675394 160501 675422 160876
rect 675670 160643 675722 160649
rect 675670 160585 675722 160591
rect 675382 160495 675434 160501
rect 675382 160437 675434 160443
rect 675682 160323 675710 160585
rect 675298 159678 675408 159706
rect 675764 159350 675820 159359
rect 675764 159285 675820 159294
rect 675778 159026 675806 159285
rect 675382 157757 675434 157763
rect 675382 157699 675434 157705
rect 675394 157176 675422 157699
rect 675478 157091 675530 157097
rect 675478 157033 675530 157039
rect 675490 156658 675518 157033
rect 675190 156573 675242 156579
rect 675190 156515 675242 156521
rect 675382 156573 675434 156579
rect 675382 156515 675434 156521
rect 675394 155992 675422 156515
rect 674998 155907 675050 155913
rect 674998 155849 675050 155855
rect 675382 155907 675434 155913
rect 675382 155849 675434 155855
rect 675394 155355 675422 155849
rect 675476 153430 675532 153439
rect 675476 153365 675532 153374
rect 675490 152884 675518 153365
rect 675380 152542 675436 152551
rect 675380 152477 675436 152486
rect 675394 152292 675422 152477
rect 675476 152246 675532 152255
rect 675476 152181 675532 152190
rect 675490 151700 675518 152181
rect 674710 151467 674762 151473
rect 674710 151409 674762 151415
rect 675382 151467 675434 151473
rect 675382 151409 675434 151415
rect 675394 151034 675422 151409
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675764 148546 675820 148555
rect 675764 148481 675820 148490
rect 675778 148000 675806 148481
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 676148 131822 676204 131831
rect 676148 131757 676204 131766
rect 676162 130161 676190 131757
rect 676340 131230 676396 131239
rect 676340 131165 676396 131174
rect 676244 130786 676300 130795
rect 676244 130721 676300 130730
rect 676150 130155 676202 130161
rect 676150 130097 676202 130103
rect 676258 130013 676286 130721
rect 676246 130007 676298 130013
rect 676246 129949 676298 129955
rect 676354 129865 676382 131165
rect 676342 129859 676394 129865
rect 676342 129801 676394 129807
rect 676244 129750 676300 129759
rect 676244 129685 676300 129694
rect 676258 129643 676286 129685
rect 676246 129637 676298 129643
rect 676246 129579 676298 129585
rect 676148 128862 676204 128871
rect 676148 128797 676204 128806
rect 676052 127604 676108 127613
rect 676052 127539 676108 127548
rect 676066 126757 676094 127539
rect 676162 126831 676190 128797
rect 676244 127826 676300 127835
rect 676244 127761 676300 127770
rect 676258 126905 676286 127761
rect 676246 126899 676298 126905
rect 676246 126841 676298 126847
rect 676150 126825 676202 126831
rect 676150 126767 676202 126773
rect 676916 126790 676972 126799
rect 674134 126751 674186 126757
rect 674134 126693 674186 126699
rect 676054 126751 676106 126757
rect 676916 126725 676972 126734
rect 676054 126693 676106 126699
rect 674038 124087 674090 124093
rect 674038 124029 674090 124035
rect 674050 111735 674078 124029
rect 674146 114177 674174 126693
rect 676244 126346 676300 126355
rect 676244 126281 676300 126290
rect 676052 126124 676108 126133
rect 676052 126059 676108 126068
rect 676066 124685 676094 126059
rect 674230 124679 674282 124685
rect 674230 124621 674282 124627
rect 676054 124679 676106 124685
rect 676054 124621 676106 124627
rect 674134 114171 674186 114177
rect 674134 114113 674186 114119
rect 674242 112549 674270 124621
rect 676052 124570 676108 124579
rect 676052 124505 676108 124514
rect 675956 124126 676012 124135
rect 675956 124061 675958 124070
rect 676010 124061 676012 124070
rect 675958 124029 676010 124035
rect 676066 124019 676094 124505
rect 674614 124013 674666 124019
rect 674614 123955 674666 123961
rect 676054 124013 676106 124019
rect 676054 123955 676106 123961
rect 674422 122163 674474 122169
rect 674422 122105 674474 122111
rect 674326 121127 674378 121133
rect 674326 121069 674378 121075
rect 674230 112543 674282 112549
rect 674230 112485 674282 112491
rect 674038 111729 674090 111735
rect 674038 111671 674090 111677
rect 674338 107369 674366 121069
rect 674434 111365 674462 122105
rect 674626 114843 674654 123955
rect 676258 123945 676286 126281
rect 676820 124866 676876 124875
rect 676820 124801 676876 124810
rect 675190 123939 675242 123945
rect 675190 123881 675242 123887
rect 676246 123939 676298 123945
rect 676246 123881 676298 123887
rect 674710 121201 674762 121207
rect 674710 121143 674762 121149
rect 674614 114837 674666 114843
rect 674614 114779 674666 114785
rect 674422 111359 674474 111365
rect 674422 111301 674474 111307
rect 674722 110699 674750 121143
rect 674806 121053 674858 121059
rect 674806 120995 674858 121001
rect 674710 110693 674762 110699
rect 674710 110635 674762 110641
rect 674326 107363 674378 107369
rect 674326 107305 674378 107311
rect 674818 106407 674846 120995
rect 675094 115429 675146 115435
rect 675094 115371 675146 115377
rect 675106 112327 675134 115371
rect 675202 115158 675230 123881
rect 676052 123534 676108 123543
rect 676052 123469 676108 123478
rect 676066 122169 676094 123469
rect 676054 122163 676106 122169
rect 676054 122105 676106 122111
rect 676052 122054 676108 122063
rect 676052 121989 676108 121998
rect 676066 121207 676094 121989
rect 676244 121462 676300 121471
rect 676244 121397 676300 121406
rect 676054 121201 676106 121207
rect 676054 121143 676106 121149
rect 676258 121133 676286 121397
rect 676246 121127 676298 121133
rect 676052 121092 676108 121101
rect 676246 121069 676298 121075
rect 676052 121027 676054 121036
rect 676106 121027 676108 121036
rect 676054 120995 676106 121001
rect 676052 120574 676108 120583
rect 676052 120509 676108 120518
rect 676066 118173 676094 120509
rect 676148 119834 676204 119843
rect 676148 119769 676204 119778
rect 676162 118247 676190 119769
rect 676244 119242 676300 119251
rect 676244 119177 676300 119186
rect 676258 118395 676286 119177
rect 676246 118389 676298 118395
rect 676246 118331 676298 118337
rect 676150 118241 676202 118247
rect 676150 118183 676202 118189
rect 676054 118167 676106 118173
rect 676054 118109 676106 118115
rect 676834 118067 676862 124801
rect 676820 118058 676876 118067
rect 676820 117993 676876 118002
rect 676930 117919 676958 126725
rect 676916 117910 676972 117919
rect 676916 117845 676972 117854
rect 675298 115648 675408 115676
rect 675298 115435 675326 115648
rect 675286 115429 675338 115435
rect 675286 115371 675338 115377
rect 675202 115130 675326 115158
rect 675298 115084 675326 115130
rect 675394 115084 675422 115144
rect 675298 115056 675422 115084
rect 675190 114837 675242 114843
rect 675190 114779 675242 114785
rect 675202 114492 675230 114779
rect 675202 114464 675408 114492
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675382 112543 675434 112549
rect 675382 112485 675434 112491
rect 675094 112321 675146 112327
rect 675094 112263 675146 112269
rect 675394 111995 675422 112485
rect 675382 111729 675434 111735
rect 675382 111671 675434 111677
rect 675394 111444 675422 111671
rect 675382 111359 675434 111365
rect 675382 111301 675434 111307
rect 675394 110778 675422 111301
rect 675382 110693 675434 110699
rect 675382 110635 675434 110641
rect 675394 110155 675422 110635
rect 675380 108142 675436 108151
rect 675380 108077 675436 108086
rect 675394 107670 675422 108077
rect 675382 107363 675434 107369
rect 675382 107305 675434 107311
rect 675394 107119 675422 107305
rect 675476 106662 675532 106671
rect 675476 106597 675532 106606
rect 675490 106486 675518 106597
rect 674806 106401 674858 106407
rect 668180 106366 668236 106375
rect 674806 106343 674858 106349
rect 675382 106401 675434 106407
rect 675382 106343 675434 106349
rect 668180 106301 668236 106310
rect 675394 105820 675422 106343
rect 668372 105182 668428 105191
rect 668372 105117 668428 105126
rect 675380 105182 675436 105191
rect 675380 105117 675436 105126
rect 665300 104886 665356 104895
rect 665300 104821 665356 104830
rect 647924 104146 647980 104155
rect 647924 104081 647980 104090
rect 647938 103817 647966 104081
rect 647926 103811 647978 103817
rect 647926 103753 647978 103759
rect 661174 103811 661226 103817
rect 661174 103753 661226 103759
rect 657526 103737 657578 103743
rect 657526 103679 657578 103685
rect 652438 102109 652490 102115
rect 652438 102051 652490 102057
rect 647924 99706 647980 99715
rect 647924 99641 647980 99650
rect 647938 97971 647966 99641
rect 647926 97965 647978 97971
rect 647926 97907 647978 97913
rect 647732 94082 647788 94091
rect 647732 94017 647788 94026
rect 647158 92193 647210 92199
rect 647158 92135 647210 92141
rect 647062 87087 647114 87093
rect 647062 87029 647114 87035
rect 646966 77763 647018 77769
rect 646966 77705 647018 77711
rect 647062 74951 647114 74957
rect 647062 74893 647114 74899
rect 646868 68626 646924 68635
rect 646868 68561 646924 68570
rect 647074 60347 647102 74893
rect 647170 71891 647198 92135
rect 647746 81617 647774 94017
rect 647828 92750 647884 92759
rect 647828 92685 647884 92694
rect 647842 81839 647870 92685
rect 650902 87531 650954 87537
rect 650902 87473 650954 87479
rect 647926 87309 647978 87315
rect 647926 87251 647978 87257
rect 647938 87135 647966 87251
rect 647924 87126 647980 87135
rect 647924 87061 647980 87070
rect 650914 86247 650942 87473
rect 650900 86238 650956 86247
rect 650900 86173 650956 86182
rect 652340 85350 652396 85359
rect 652340 85285 652396 85294
rect 651764 84314 651820 84323
rect 651764 84249 651820 84258
rect 651778 83615 651806 84249
rect 651766 83609 651818 83615
rect 651766 83551 651818 83557
rect 652244 83426 652300 83435
rect 652244 83361 652300 83370
rect 647924 82686 647980 82695
rect 647924 82621 647980 82630
rect 647938 81913 647966 82621
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647830 81833 647882 81839
rect 647830 81775 647882 81781
rect 647734 81611 647786 81617
rect 647734 81553 647786 81559
rect 647924 81058 647980 81067
rect 647924 80993 647980 81002
rect 647938 80803 647966 80993
rect 647926 80797 647978 80803
rect 647926 80739 647978 80745
rect 647926 77541 647978 77547
rect 647924 77506 647926 77515
rect 647978 77506 647980 77515
rect 647924 77441 647980 77450
rect 647924 73658 647980 73667
rect 647924 73593 647980 73602
rect 647938 72145 647966 73593
rect 647926 72139 647978 72145
rect 647926 72081 647978 72087
rect 647156 71882 647212 71891
rect 647156 71817 647212 71826
rect 647924 69662 647980 69671
rect 647924 69597 647980 69606
rect 647938 69481 647966 69597
rect 647926 69475 647978 69481
rect 647926 69417 647978 69423
rect 647924 64186 647980 64195
rect 647924 64121 647980 64130
rect 647938 63635 647966 64121
rect 647926 63629 647978 63635
rect 647926 63571 647978 63577
rect 647924 62262 647980 62271
rect 647924 62197 647980 62206
rect 647938 61045 647966 62197
rect 647926 61039 647978 61045
rect 647926 60981 647978 60987
rect 647060 60338 647116 60347
rect 647060 60273 647116 60282
rect 652258 59121 652286 83361
rect 652354 66225 652382 85285
rect 652450 82695 652478 102051
rect 653686 95967 653738 95973
rect 653686 95909 653738 95915
rect 653698 86987 653726 95909
rect 657538 88000 657566 103679
rect 660694 92341 660746 92347
rect 660694 92283 660746 92289
rect 659830 92267 659882 92273
rect 659830 92209 659882 92215
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 657538 87972 657792 88000
rect 658882 87986 658910 92135
rect 659348 90826 659404 90835
rect 659348 90761 659404 90770
rect 659362 88000 659390 90761
rect 659842 88000 659870 92209
rect 659362 87972 659616 88000
rect 659842 87972 660144 88000
rect 660706 87986 660734 92283
rect 661186 88000 661214 103753
rect 662518 97965 662570 97971
rect 662518 97907 662570 97913
rect 661750 92415 661802 92421
rect 661750 92357 661802 92363
rect 661762 88000 661790 92357
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 97907
rect 663094 92711 663146 92717
rect 663094 92653 663146 92659
rect 663106 87986 663134 92653
rect 658006 87309 658058 87315
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 653684 86978 653740 86987
rect 653684 86913 653740 86922
rect 663298 86395 663326 87029
rect 663284 86386 663340 86395
rect 663284 86321 663340 86330
rect 663284 84758 663340 84767
rect 663202 84716 663284 84744
rect 657046 84201 657098 84207
rect 657046 84143 657098 84149
rect 652436 82686 652492 82695
rect 652436 82621 652492 82630
rect 657058 81691 657086 84143
rect 657046 81685 657098 81691
rect 657046 81627 657098 81633
rect 658582 81685 658634 81691
rect 662420 81650 662476 81659
rect 658634 81633 658896 81636
rect 658582 81627 658896 81633
rect 658594 81608 658896 81627
rect 662420 81585 662422 81594
rect 662474 81585 662476 81594
rect 662422 81553 662474 81559
rect 656962 81016 657216 81044
rect 657538 81016 657792 81044
rect 656962 77547 656990 81016
rect 656950 77541 657002 77547
rect 656950 77483 657002 77489
rect 657538 76141 657566 81016
rect 658306 77769 658334 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658294 77763 658346 77769
rect 658294 77705 658346 77711
rect 659458 77695 659486 80665
rect 659446 77689 659498 77695
rect 659446 77631 659498 77637
rect 657526 76135 657578 76141
rect 657526 76077 657578 76083
rect 660130 74957 660158 81030
rect 660118 74951 660170 74957
rect 660118 74893 660170 74899
rect 660706 72145 660734 81030
rect 660886 81019 660938 81025
rect 661440 81016 661502 81044
rect 660886 80961 660938 80967
rect 660694 72139 660746 72145
rect 660694 72081 660746 72087
rect 652342 66219 652394 66225
rect 652342 66161 652394 66167
rect 652246 59115 652298 59121
rect 652246 59057 652298 59063
rect 646772 57082 646828 57091
rect 646772 57017 646828 57026
rect 184340 54714 184396 54723
rect 149686 54675 149738 54681
rect 184340 54649 184342 54658
rect 149686 54617 149738 54623
rect 184394 54649 184396 54658
rect 646484 54714 646540 54723
rect 646484 54649 646540 54658
rect 184342 54617 184394 54623
rect 184340 53974 184396 53983
rect 184340 53909 184396 53918
rect 149396 53826 149452 53835
rect 149396 53761 149452 53770
rect 149410 53275 149438 53761
rect 184354 53275 184382 53909
rect 149398 53269 149450 53275
rect 149398 53211 149450 53217
rect 184342 53269 184394 53275
rect 184342 53211 184394 53217
rect 145104 49788 145406 49816
rect 145378 47133 145406 49788
rect 199138 47133 199166 53650
rect 145366 47127 145418 47133
rect 145366 47069 145418 47075
rect 199126 47127 199178 47133
rect 199126 47069 199178 47075
rect 142114 46680 142416 46708
rect 142114 40219 142142 46680
rect 216418 41995 216446 53650
rect 233698 47725 233726 53650
rect 233686 47719 233738 47725
rect 233686 47661 233738 47667
rect 250978 47577 251006 53650
rect 268320 53636 268574 53664
rect 285600 53636 285854 53664
rect 268546 47651 268574 53636
rect 268534 47645 268586 47651
rect 268534 47587 268586 47593
rect 250966 47571 251018 47577
rect 250966 47513 251018 47519
rect 224566 44685 224618 44691
rect 224566 44627 224618 44633
rect 187604 41986 187660 41995
rect 187344 41944 187604 41972
rect 187604 41921 187660 41930
rect 216404 41986 216460 41995
rect 216404 41921 216460 41930
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 194324 41773 194380 41782
rect 224578 40515 224606 44627
rect 285826 43285 285854 53636
rect 302914 47799 302942 53650
rect 311062 47941 311114 47947
rect 311062 47883 311114 47889
rect 302902 47793 302954 47799
rect 302902 47735 302954 47741
rect 285814 43279 285866 43285
rect 285814 43221 285866 43227
rect 311074 42268 311102 47883
rect 320194 47873 320222 53650
rect 320182 47867 320234 47873
rect 320182 47809 320234 47815
rect 337474 46319 337502 53650
rect 354850 46319 354878 53650
rect 371938 53636 372192 53664
rect 389218 53636 389472 53664
rect 371938 47947 371966 53636
rect 371926 47941 371978 47947
rect 371926 47883 371978 47889
rect 324310 46313 324362 46319
rect 324310 46255 324362 46261
rect 337462 46313 337514 46319
rect 337462 46255 337514 46261
rect 345622 46313 345674 46319
rect 345622 46255 345674 46261
rect 354838 46313 354890 46319
rect 354838 46255 354890 46261
rect 310498 42240 311102 42268
rect 310498 42120 310526 42240
rect 310128 42092 310526 42120
rect 307222 42021 307274 42027
rect 307008 41969 307222 41972
rect 307008 41963 307274 41969
rect 311062 42021 311114 42027
rect 311062 41963 311114 41969
rect 307008 41944 307262 41963
rect 302900 41838 302956 41847
rect 302688 41796 302900 41824
rect 302900 41773 302956 41782
rect 224564 40506 224620 40515
rect 224564 40441 224620 40450
rect 142100 40210 142156 40219
rect 142100 40145 142156 40154
rect 311074 37259 311102 41963
rect 324322 37259 324350 46255
rect 345634 40515 345662 46255
rect 365314 42240 365726 42268
rect 365314 42120 365342 42240
rect 364944 42092 365342 42120
rect 362038 42021 362090 42027
rect 361776 41969 362038 41972
rect 361776 41963 362090 41969
rect 361776 41944 362078 41963
rect 357716 41838 357772 41847
rect 357456 41796 357716 41824
rect 365698 41824 365726 42240
rect 365974 42021 366026 42027
rect 365974 41963 366026 41969
rect 365698 41796 365918 41824
rect 357716 41773 357772 41782
rect 345620 40506 345676 40515
rect 345620 40441 345676 40450
rect 365890 37439 365918 41796
rect 365878 37433 365930 37439
rect 365878 37375 365930 37381
rect 365986 37365 366014 41963
rect 389218 37365 389246 53636
rect 406786 48021 406814 53650
rect 424066 48021 424094 53650
rect 434902 48163 434954 48169
rect 434902 48105 434954 48111
rect 394582 48015 394634 48021
rect 394582 47957 394634 47963
rect 406774 48015 406826 48021
rect 406774 47957 406826 47963
rect 411862 48015 411914 48021
rect 411862 47957 411914 47963
rect 424054 48015 424106 48021
rect 424054 47957 424106 47963
rect 426166 48015 426218 48021
rect 426166 47957 426218 47963
rect 394594 41847 394622 47957
rect 405526 47941 405578 47947
rect 405526 47883 405578 47889
rect 399862 42391 399914 42397
rect 399862 42333 399914 42339
rect 394580 41838 394636 41847
rect 394580 41773 394636 41782
rect 399874 37439 399902 42333
rect 405538 42106 405566 47883
rect 411874 42397 411902 47957
rect 426178 44955 426206 47957
rect 426164 44946 426220 44955
rect 426164 44881 426220 44890
rect 411862 42391 411914 42397
rect 411862 42333 411914 42339
rect 434914 41995 434942 48105
rect 441346 47947 441374 53650
rect 441334 47941 441386 47947
rect 441334 47883 441386 47889
rect 415220 41986 415276 41995
rect 415220 41921 415276 41930
rect 434900 41986 434956 41995
rect 434900 41921 434956 41930
rect 415234 41810 415262 41921
rect 416852 41838 416908 41847
rect 416592 41796 416852 41824
rect 416852 41773 416908 41782
rect 458626 40515 458654 53650
rect 475714 53636 475968 53664
rect 492994 53636 493248 53664
rect 510370 53636 510624 53664
rect 475714 48169 475742 53636
rect 475702 48163 475754 48169
rect 475702 48105 475754 48111
rect 460342 48089 460394 48095
rect 460342 48031 460394 48037
rect 460354 42106 460382 48031
rect 492994 48021 493022 53636
rect 510370 48095 510398 53636
rect 510358 48089 510410 48095
rect 510358 48031 510410 48037
rect 492982 48015 493034 48021
rect 492982 47957 493034 47963
rect 472246 47941 472298 47947
rect 472246 47883 472298 47889
rect 472258 44955 472286 47883
rect 523894 47793 523946 47799
rect 523894 47735 523946 47741
rect 475510 47719 475562 47725
rect 475510 47661 475562 47667
rect 505366 47719 505418 47725
rect 505366 47661 505418 47667
rect 472244 44946 472300 44955
rect 472244 44881 472300 44890
rect 470324 41838 470380 41847
rect 470160 41796 470324 41824
rect 471668 41838 471724 41847
rect 471408 41796 471668 41824
rect 470324 41773 470380 41782
rect 471668 41773 471724 41782
rect 458612 40506 458668 40515
rect 458612 40441 458668 40450
rect 475522 37439 475550 47661
rect 505378 40663 505406 47661
rect 517366 47645 517418 47651
rect 517366 47587 517418 47593
rect 517378 42143 517406 47587
rect 521206 47571 521258 47577
rect 521206 47513 521258 47519
rect 518722 43285 518834 43304
rect 518710 43279 518834 43285
rect 518762 43276 518834 43279
rect 518710 43221 518762 43227
rect 521218 42268 521246 47513
rect 523906 44025 523934 47735
rect 527938 47725 527966 53650
rect 529270 47867 529322 47873
rect 529270 47809 529322 47815
rect 527926 47719 527978 47725
rect 527926 47661 527978 47667
rect 523894 44019 523946 44025
rect 523894 43961 523946 43967
rect 525910 44019 525962 44025
rect 525910 43961 525962 43967
rect 521218 42240 521534 42268
rect 517364 42134 517420 42143
rect 517364 42069 517420 42078
rect 520340 42134 520396 42143
rect 521506 42120 521534 42240
rect 525922 42120 525950 43961
rect 520396 42092 520656 42120
rect 521506 42092 521856 42120
rect 525922 42092 526176 42120
rect 529282 42106 529310 47809
rect 520340 42069 520396 42078
rect 514882 41805 515136 41824
rect 514006 41799 514058 41805
rect 514006 41741 514058 41747
rect 514870 41799 515136 41805
rect 514922 41796 515136 41799
rect 514870 41741 514922 41747
rect 505364 40654 505420 40663
rect 505364 40589 505420 40598
rect 514018 37439 514046 41741
rect 545218 40515 545246 53650
rect 562498 47947 562526 53650
rect 579796 53602 579852 54402
rect 597092 53602 597148 54402
rect 614388 53602 614444 54402
rect 631684 53602 631740 54402
rect 562486 47941 562538 47947
rect 562486 47883 562538 47889
rect 660898 44691 660926 80961
rect 661474 69481 661502 81016
rect 661762 81016 662016 81044
rect 661762 77621 661790 81016
rect 662530 80803 662558 81030
rect 662518 80797 662570 80803
rect 662518 80739 662570 80745
rect 661750 77615 661802 77621
rect 661750 77557 661802 77563
rect 661462 69475 661514 69481
rect 661462 69417 661514 69423
rect 663202 63635 663230 84716
rect 663284 84693 663340 84702
rect 663476 84018 663532 84027
rect 663476 83953 663532 83962
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663190 63629 663242 63635
rect 663190 63571 663242 63577
rect 663490 61045 663518 83953
rect 668386 81025 668414 105117
rect 675394 104636 675422 105117
rect 675764 103258 675820 103267
rect 675764 103193 675820 103202
rect 675778 102786 675806 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 668374 81019 668426 81025
rect 668374 80961 668426 80967
rect 663478 61039 663530 61045
rect 663478 60981 663530 60987
rect 660886 44685 660938 44691
rect 660886 44627 660938 44633
rect 545204 40506 545260 40515
rect 545204 40441 545260 40450
rect 399862 37433 399914 37439
rect 399862 37375 399914 37381
rect 475510 37433 475562 37439
rect 475510 37375 475562 37381
rect 514006 37433 514058 37439
rect 514006 37375 514058 37381
rect 365974 37359 366026 37365
rect 365974 37301 366026 37307
rect 389206 37359 389258 37365
rect 389206 37301 389258 37307
rect 311060 37250 311116 37259
rect 311060 37185 311116 37194
rect 324308 37250 324364 37259
rect 324308 37185 324364 37194
<< via2 >>
rect 82292 1002319 82348 1002358
rect 82292 1002302 82294 1002319
rect 82294 1002302 82346 1002319
rect 82346 1002302 82348 1002319
rect 483668 1002319 483724 1002358
rect 483668 1002302 483670 1002319
rect 483670 1002302 483722 1002319
rect 483722 1002302 483724 1002319
rect 132404 997714 132460 997770
rect 184244 997714 184300 997770
rect 241172 997122 241228 997178
rect 80564 982914 80620 982970
rect 132404 982914 132460 982970
rect 184244 982914 184300 982970
rect 233204 982914 233260 982970
rect 240884 982953 240886 982970
rect 240886 982953 240938 982970
rect 240938 982953 240940 982970
rect 240884 982914 240940 982953
rect 241172 982914 241228 982970
rect 293108 997122 293164 997178
rect 285044 982914 285100 982970
rect 389588 983210 389644 983266
rect 292532 982953 292534 982970
rect 292534 982953 292586 982970
rect 292586 982953 292588 982970
rect 292532 982914 292588 982953
rect 293108 982914 293164 982970
rect 400340 997122 400396 997178
rect 535700 997714 535756 997770
rect 639380 997714 639436 997770
rect 394580 982914 394636 982970
rect 400340 982914 400396 982970
rect 486740 982914 486796 982970
rect 538580 982914 538636 982970
rect 639380 982914 639436 982970
rect 40148 961915 40204 961954
rect 40148 961898 40150 961915
rect 40150 961898 40202 961915
rect 40202 961898 40204 961915
rect 60020 961750 60076 961806
rect 653780 960457 653782 960474
rect 653782 960457 653834 960474
rect 653834 960457 653836 960474
rect 653780 960418 653836 960457
rect 679700 958494 679756 958550
rect 676148 894114 676204 894170
rect 676052 893374 676108 893430
rect 655220 867622 655276 867678
rect 655124 866438 655180 866494
rect 676244 893522 676300 893578
rect 676052 892429 676108 892468
rect 676052 892412 676054 892429
rect 676054 892412 676106 892429
rect 676106 892412 676108 892429
rect 655412 868806 655468 868862
rect 655316 865254 655372 865310
rect 654164 863922 654220 863978
rect 653780 862886 653836 862942
rect 41780 816653 41836 816692
rect 41780 816636 41782 816653
rect 41782 816636 41834 816653
rect 41834 816636 41836 816653
rect 41780 816135 41836 816174
rect 41780 816118 41782 816135
rect 41782 816118 41834 816135
rect 41834 816118 41836 816135
rect 41588 815395 41644 815434
rect 41588 815378 41590 815395
rect 41590 815378 41642 815395
rect 41642 815378 41644 815395
rect 41780 814655 41836 814694
rect 41780 814638 41782 814655
rect 41782 814638 41834 814655
rect 41834 814638 41836 814655
rect 41588 813471 41644 813510
rect 41588 813454 41590 813471
rect 41590 813454 41642 813471
rect 41642 813454 41644 813471
rect 41780 812583 41836 812622
rect 41780 812566 41782 812583
rect 41782 812566 41834 812583
rect 41834 812566 41836 812583
rect 41396 811974 41452 812030
rect 40244 811234 40300 811290
rect 28820 804426 28876 804482
rect 28820 803834 28876 803890
rect 40244 801318 40300 801374
rect 41972 811604 42028 811660
rect 41588 810494 41644 810550
rect 41684 809902 41740 809958
rect 41588 808439 41644 808478
rect 41588 808422 41590 808439
rect 41590 808422 41642 808439
rect 41642 808422 41644 808439
rect 41588 806959 41644 806998
rect 41588 806942 41590 806959
rect 41590 806942 41642 806959
rect 41642 806942 41644 806959
rect 41588 805462 41644 805518
rect 41492 803834 41548 803890
rect 41876 809606 41932 809662
rect 41780 807682 41836 807738
rect 41780 806202 41836 806258
rect 41684 800430 41740 800486
rect 42164 808126 42220 808182
rect 42068 806572 42124 806628
rect 41972 800282 42028 800338
rect 42164 800282 42220 800338
rect 41972 798062 42028 798118
rect 42836 795398 42892 795454
rect 41780 792882 41836 792938
rect 42836 791846 42892 791902
rect 42932 791698 42988 791754
rect 41588 774530 41644 774586
rect 41492 773938 41548 773994
rect 41780 773511 41836 773550
rect 41780 773494 41782 773511
rect 41782 773494 41834 773511
rect 41834 773494 41836 773511
rect 41780 772919 41836 772958
rect 41780 772902 41782 772919
rect 41782 772902 41834 772919
rect 41834 772902 41836 772919
rect 41780 772327 41836 772366
rect 41780 772310 41782 772327
rect 41782 772310 41834 772327
rect 41834 772310 41836 772327
rect 41780 771979 41782 771996
rect 41782 771979 41834 771996
rect 41834 771979 41836 771996
rect 41780 771940 41836 771979
rect 41780 771439 41836 771478
rect 41780 771422 41782 771439
rect 41782 771422 41834 771439
rect 41834 771422 41836 771439
rect 41588 770682 41644 770738
rect 41492 769646 41548 769702
rect 41588 768758 41644 768814
rect 38804 768018 38860 768074
rect 34484 765798 34540 765854
rect 28820 761210 28876 761266
rect 28820 760766 28876 760822
rect 34484 758842 34540 758898
rect 41684 768166 41740 768222
rect 41588 767278 41644 767334
rect 40340 766538 40396 766594
rect 38804 757510 38860 757566
rect 41300 765058 41356 765114
rect 41588 761654 41644 761710
rect 41588 760783 41644 760822
rect 41588 760766 41590 760783
rect 41590 760766 41642 760783
rect 41642 760766 41644 760783
rect 41972 766908 42028 766964
rect 41780 765445 41836 765484
rect 41780 765428 41782 765445
rect 41782 765428 41834 765445
rect 41834 765428 41836 765445
rect 41876 764466 41932 764522
rect 41780 763447 41836 763486
rect 41780 763430 41782 763447
rect 41782 763430 41834 763447
rect 41834 763430 41836 763447
rect 41780 762394 41836 762450
rect 42068 763874 42124 763930
rect 42164 762986 42220 763042
rect 43028 757954 43084 758010
rect 41972 757066 42028 757122
rect 42740 754698 42796 754754
rect 43124 757214 43180 757270
rect 42836 750406 42892 750462
rect 42836 747150 42892 747206
rect 42740 746854 42796 746910
rect 43028 751590 43084 751646
rect 41588 731462 41644 731518
rect 41684 731314 41740 731370
rect 41780 730443 41836 730482
rect 41780 730426 41782 730443
rect 41782 730426 41834 730443
rect 41834 730426 41836 730443
rect 41780 729925 41836 729964
rect 41780 729908 41782 729925
rect 41782 729908 41834 729925
rect 41834 729908 41836 729925
rect 41780 729407 41836 729446
rect 41780 729390 41782 729407
rect 41782 729390 41834 729407
rect 41834 729390 41836 729407
rect 41780 728985 41782 729002
rect 41782 728985 41834 729002
rect 41834 728985 41836 729002
rect 41780 728946 41836 728985
rect 41588 727614 41644 727670
rect 41780 728371 41836 728410
rect 41780 728354 41782 728371
rect 41782 728354 41834 728371
rect 41834 728354 41836 728371
rect 41780 727927 41836 727966
rect 41780 727910 41782 727927
rect 41782 727910 41834 727927
rect 41834 727910 41836 727927
rect 41780 726891 41836 726930
rect 41780 726874 41782 726891
rect 41782 726874 41834 726891
rect 41834 726874 41836 726891
rect 41684 726726 41740 726782
rect 41780 726003 41836 726042
rect 41780 725986 41782 726003
rect 41782 725986 41834 726003
rect 41834 725986 41836 726003
rect 41876 725394 41932 725450
rect 39764 724654 39820 724710
rect 34484 722730 34540 722786
rect 28820 718142 28876 718198
rect 28820 717698 28876 717754
rect 34484 715626 34540 715682
rect 41684 724062 41740 724118
rect 41588 721250 41644 721306
rect 41588 720675 41644 720714
rect 41588 720658 41590 720675
rect 41590 720658 41642 720675
rect 41642 720658 41644 720675
rect 41588 719770 41644 719826
rect 41588 719178 41644 719234
rect 41492 717715 41548 717754
rect 41492 717698 41494 717715
rect 41494 717698 41546 717715
rect 41546 717698 41548 717715
rect 39764 714886 39820 714942
rect 41780 723322 41836 723378
rect 41972 724506 42028 724562
rect 42164 722434 42220 722490
rect 42068 720362 42124 720418
rect 41972 713998 42028 714054
rect 42260 721842 42316 721898
rect 42164 714146 42220 714202
rect 42068 713850 42124 713906
rect 42740 715774 42796 715830
rect 42836 714442 42892 714498
rect 42932 711038 42988 711094
rect 42836 710742 42892 710798
rect 42164 707930 42220 707986
rect 42740 705118 42796 705174
rect 43028 708226 43084 708282
rect 42932 704082 42988 704138
rect 43124 707190 43180 707246
rect 41780 686857 41836 686896
rect 41780 686840 41782 686857
rect 41782 686840 41834 686857
rect 41834 686840 41836 686857
rect 41780 686339 41836 686378
rect 41780 686322 41782 686339
rect 41782 686322 41834 686339
rect 41834 686322 41836 686339
rect 41588 685599 41644 685638
rect 41588 685582 41590 685599
rect 41590 685582 41642 685599
rect 41642 685582 41644 685599
rect 41780 685325 41782 685342
rect 41782 685325 41834 685342
rect 41834 685325 41836 685342
rect 41780 685286 41836 685325
rect 41780 684859 41836 684898
rect 41780 684842 41782 684859
rect 41782 684842 41834 684859
rect 41834 684842 41836 684859
rect 41780 683845 41782 683862
rect 41782 683845 41834 683862
rect 41834 683845 41836 683862
rect 41780 683806 41836 683845
rect 43796 702010 43852 702066
rect 41588 682957 41590 682974
rect 41590 682957 41642 682974
rect 41642 682957 41644 682974
rect 41588 682918 41644 682957
rect 39764 682178 39820 682234
rect 37364 680698 37420 680754
rect 34484 678626 34540 678682
rect 23060 674482 23116 674538
rect 23060 674038 23116 674094
rect 41780 681808 41836 681864
rect 39860 681438 39916 681494
rect 41972 680254 42028 680310
rect 41780 679810 41836 679866
rect 40244 679070 40300 679126
rect 41684 676554 41740 676610
rect 41588 676127 41644 676166
rect 41588 676110 41590 676127
rect 41590 676110 41642 676127
rect 41642 676110 41644 676127
rect 41588 675666 41644 675722
rect 41588 674055 41644 674094
rect 41588 674038 41590 674055
rect 41590 674038 41642 674055
rect 41642 674038 41644 674055
rect 40244 673594 40300 673650
rect 39860 671078 39916 671134
rect 41684 670930 41740 670986
rect 41876 677886 41932 677942
rect 42260 678330 42316 678386
rect 42068 677294 42124 677350
rect 41876 670782 41932 670838
rect 42068 670634 42124 670690
rect 41876 666638 41932 666694
rect 42164 664714 42220 664770
rect 41780 660866 41836 660922
rect 42932 660274 42988 660330
rect 42836 659682 42892 659738
rect 41492 645030 41548 645086
rect 41684 644882 41740 644938
rect 41780 643715 41836 643754
rect 41780 643698 41782 643715
rect 41782 643698 41834 643715
rect 41834 643698 41836 643715
rect 41780 643123 41836 643162
rect 41780 643106 41782 643123
rect 41782 643106 41834 643123
rect 41834 643106 41836 643123
rect 41588 642383 41644 642422
rect 41588 642366 41590 642383
rect 41590 642366 41642 642383
rect 41642 642366 41644 642383
rect 41492 640886 41548 640942
rect 41780 642183 41782 642200
rect 41782 642183 41834 642200
rect 41834 642183 41836 642200
rect 41780 642144 41836 642183
rect 41780 641643 41836 641682
rect 41780 641626 41782 641643
rect 41782 641626 41834 641643
rect 41834 641626 41836 641643
rect 41780 640163 41836 640202
rect 41780 640146 41782 640163
rect 41782 640146 41834 640163
rect 41834 640146 41836 640163
rect 41684 639850 41740 639906
rect 37364 638962 37420 639018
rect 34388 636002 34444 636058
rect 23060 631414 23116 631470
rect 23060 630970 23116 631026
rect 34484 635410 34540 635466
rect 34388 628010 34444 628066
rect 40244 638222 40300 638278
rect 40148 637482 40204 637538
rect 41492 636890 41548 636946
rect 40244 627862 40300 627918
rect 41780 636594 41836 636650
rect 41588 633947 41644 633986
rect 41588 633930 41590 633947
rect 41590 633930 41642 633947
rect 41642 633930 41644 633947
rect 41588 630839 41644 630878
rect 41588 630822 41590 630839
rect 41590 630822 41642 630839
rect 41642 630822 41644 630839
rect 42068 635114 42124 635170
rect 41876 633190 41932 633246
rect 42836 634670 42892 634726
rect 42164 633634 42220 633690
rect 42260 632598 42316 632654
rect 42068 627418 42124 627474
rect 42164 625198 42220 625254
rect 42740 624754 42796 624810
rect 42836 617650 42892 617706
rect 42740 617206 42796 617262
rect 40340 602110 40396 602166
rect 41780 600499 41836 600538
rect 41780 600482 41782 600499
rect 41782 600482 41834 600499
rect 41834 600482 41836 600499
rect 41588 599759 41644 599798
rect 41588 599742 41590 599759
rect 41590 599742 41642 599759
rect 41642 599742 41644 599759
rect 41780 599389 41836 599428
rect 41780 599372 41782 599389
rect 41782 599372 41834 599389
rect 41834 599372 41836 599389
rect 41780 599019 41836 599058
rect 41780 599002 41782 599019
rect 41782 599002 41834 599019
rect 41834 599002 41836 599019
rect 41588 598279 41644 598318
rect 41588 598262 41590 598279
rect 41590 598262 41642 598279
rect 41642 598262 41644 598279
rect 40340 597670 40396 597726
rect 41588 596207 41644 596246
rect 41588 596190 41590 596207
rect 41590 596190 41642 596207
rect 41642 596190 41644 596207
rect 41492 595746 41548 595802
rect 34388 594710 34444 594766
rect 23060 588198 23116 588254
rect 23060 587754 23116 587810
rect 34484 592786 34540 592842
rect 34388 584794 34444 584850
rect 34484 584646 34540 584702
rect 41780 595450 41836 595506
rect 41684 594266 41740 594322
rect 41588 591306 41644 591362
rect 41588 589826 41644 589882
rect 41588 589234 41644 589290
rect 41588 587754 41644 587810
rect 42164 593970 42220 594026
rect 41780 593378 41836 593434
rect 41492 584498 41548 584554
rect 41684 584498 41740 584554
rect 41972 592490 42028 592546
rect 41876 590953 41932 590992
rect 41876 590936 41878 590953
rect 41878 590936 41930 590953
rect 41930 590936 41932 590953
rect 42068 591898 42124 591954
rect 41972 584646 42028 584702
rect 42356 590418 42412 590474
rect 41876 584202 41932 584258
rect 42836 578578 42892 578634
rect 42068 578134 42124 578190
rect 41780 573398 41836 573454
rect 43028 576802 43084 576858
rect 42932 573990 42988 574046
rect 43124 574434 43180 574490
rect 43028 544390 43084 544446
rect 41588 543075 41644 543114
rect 41588 543058 41590 543075
rect 41590 543058 41642 543075
rect 41642 543058 41644 543075
rect 41780 542705 41836 542744
rect 41780 542688 41782 542705
rect 41782 542688 41834 542705
rect 41834 542688 41836 542705
rect 41780 542187 41836 542226
rect 41780 542170 41782 542187
rect 41782 542170 41834 542187
rect 41834 542170 41836 542187
rect 41780 541765 41782 541782
rect 41782 541765 41834 541782
rect 41834 541765 41836 541782
rect 41780 541726 41836 541765
rect 41780 538174 41836 538230
rect 42740 536694 42796 536750
rect 41780 536250 41836 536306
rect 41972 534918 42028 534974
rect 41780 534178 41836 534234
rect 41780 533882 41836 533938
rect 43508 541134 43564 541190
rect 43412 540690 43468 540746
rect 43028 539210 43084 539266
rect 43124 538766 43180 538822
rect 43028 537286 43084 537342
rect 42932 536546 42988 536602
rect 42836 534622 42892 534678
rect 42740 533142 42796 533198
rect 42932 532698 42988 532754
rect 42836 530626 42892 530682
rect 41780 529590 41836 529646
rect 41684 525002 41740 525058
rect 41588 429263 41644 429302
rect 41588 429246 41590 429263
rect 41590 429246 41642 429263
rect 41642 429246 41644 429263
rect 41780 428967 41836 429006
rect 41780 428950 41782 428967
rect 41782 428950 41834 428967
rect 41834 428950 41836 428967
rect 41780 428375 41836 428414
rect 41780 428358 41782 428375
rect 41782 428358 41834 428375
rect 41834 428358 41836 428375
rect 41780 427953 41782 427970
rect 41782 427953 41834 427970
rect 41834 427953 41836 427970
rect 41780 427914 41836 427953
rect 41780 427413 41836 427452
rect 41780 427396 41782 427413
rect 41782 427396 41834 427413
rect 41834 427396 41836 427413
rect 41780 426895 41836 426934
rect 41780 426878 41782 426895
rect 41782 426878 41834 426895
rect 41834 426878 41836 426895
rect 25844 425546 25900 425602
rect 41780 425398 41836 425454
rect 41684 422142 41740 422198
rect 41588 420218 41644 420274
rect 25844 418738 25900 418794
rect 28820 417110 28876 417166
rect 41780 419922 41836 419978
rect 41780 418960 41836 419016
rect 41780 418442 41836 418498
rect 41780 416979 41836 417018
rect 41780 416962 41782 416979
rect 41782 416962 41834 416979
rect 41834 416962 41836 416979
rect 28820 416666 28876 416722
rect 41876 411190 41932 411246
rect 41876 406010 41932 406066
rect 42068 403790 42124 403846
rect 41780 403050 41836 403106
rect 41780 402606 41836 402662
rect 41780 401866 41836 401922
rect 41780 400090 41836 400146
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 41780 386491 41836 386530
rect 41780 386474 41782 386491
rect 41782 386474 41834 386491
rect 41834 386474 41836 386491
rect 41588 385751 41644 385790
rect 41588 385734 41590 385751
rect 41590 385734 41642 385751
rect 41642 385734 41644 385751
rect 41780 385381 41836 385420
rect 41780 385364 41782 385381
rect 41782 385364 41834 385381
rect 41834 385364 41836 385381
rect 41588 385181 41590 385198
rect 41590 385181 41642 385198
rect 41642 385181 41644 385198
rect 41588 385142 41644 385181
rect 41780 384419 41836 384458
rect 41780 384402 41782 384419
rect 41782 384402 41834 384419
rect 41834 384402 41836 384419
rect 34484 383662 34540 383718
rect 28724 381590 28780 381646
rect 43508 426434 43564 426490
rect 41780 383479 41782 383496
rect 41782 383479 41834 383496
rect 41834 383479 41836 383496
rect 41780 383440 41836 383479
rect 40244 382626 40300 382682
rect 23060 374190 23116 374246
rect 23060 373746 23116 373802
rect 39380 380702 39436 380758
rect 39284 379666 39340 379722
rect 39860 379666 39916 379722
rect 39764 378778 39820 378834
rect 39476 378186 39532 378242
rect 39668 377150 39724 377206
rect 39764 374190 39820 374246
rect 41780 376945 41836 376984
rect 41780 376928 41782 376945
rect 41782 376928 41834 376945
rect 41834 376928 41836 376945
rect 41780 375966 41836 376022
rect 41588 375226 41644 375282
rect 39860 373746 39916 373802
rect 39476 373154 39532 373210
rect 39380 372710 39436 372766
rect 28724 372414 28780 372470
rect 41876 373911 41932 373950
rect 41876 373894 41878 373911
rect 41878 373894 41930 373911
rect 41930 373894 41932 373911
rect 41780 368122 41836 368178
rect 41780 362794 41836 362850
rect 41972 360574 42028 360630
rect 41780 359834 41836 359890
rect 42068 359242 42124 359298
rect 41780 358798 41836 358854
rect 41876 356874 41932 356930
rect 41780 356134 41836 356190
rect 42164 355690 42220 355746
rect 41588 343275 41644 343314
rect 41588 343258 41590 343275
rect 41590 343258 41642 343275
rect 41642 343258 41644 343275
rect 41780 342905 41836 342944
rect 41780 342888 41782 342905
rect 41782 342888 41834 342905
rect 41834 342888 41836 342905
rect 41780 342387 41836 342426
rect 41780 342370 41782 342387
rect 41782 342370 41834 342387
rect 41834 342370 41836 342387
rect 41780 341965 41782 341982
rect 41782 341965 41834 341982
rect 41834 341965 41836 341982
rect 41780 341926 41836 341965
rect 41780 341425 41836 341464
rect 41780 341408 41782 341425
rect 41782 341408 41834 341425
rect 41834 341408 41836 341425
rect 41780 340907 41836 340946
rect 41780 340890 41782 340907
rect 41782 340890 41834 340907
rect 41834 340890 41836 340907
rect 41780 340485 41782 340502
rect 41782 340485 41834 340502
rect 41834 340485 41836 340502
rect 41780 340446 41836 340485
rect 41780 339871 41836 339910
rect 41780 339854 41782 339871
rect 41782 339854 41834 339871
rect 41834 339854 41836 339871
rect 41588 339745 41590 339762
rect 41590 339745 41642 339762
rect 41642 339745 41644 339762
rect 41588 339706 41644 339745
rect 28724 338670 28780 338726
rect 23060 331122 23116 331178
rect 23060 330678 23116 330734
rect 39284 337634 39340 337690
rect 41684 336154 41740 336210
rect 41588 334082 41644 334138
rect 39284 331122 39340 331178
rect 28724 329198 28780 329254
rect 41780 333934 41836 333990
rect 41780 332454 41836 332510
rect 41876 330991 41932 331030
rect 41876 330974 41878 330991
rect 41878 330974 41930 330991
rect 41930 330974 41932 330991
rect 41780 324906 41836 324962
rect 42164 320466 42220 320522
rect 41780 319726 41836 319782
rect 42164 317358 42220 317414
rect 41876 316766 41932 316822
rect 41780 316026 41836 316082
rect 41780 315582 41836 315638
rect 42068 313658 42124 313714
rect 41780 313066 41836 313122
rect 41780 312326 41836 312382
rect 41588 299894 41644 299950
rect 41780 299763 41836 299802
rect 41780 299746 41782 299763
rect 41782 299746 41834 299763
rect 41834 299746 41836 299763
rect 39668 299450 39724 299506
rect 28724 295454 28780 295510
rect 23060 287906 23116 287962
rect 23060 287462 23116 287518
rect 41780 298749 41782 298766
rect 41782 298749 41834 298766
rect 41834 298749 41836 298766
rect 41780 298710 41836 298749
rect 41780 298209 41836 298248
rect 41780 298192 41782 298209
rect 41782 298192 41834 298209
rect 41834 298192 41836 298209
rect 41780 297691 41836 297730
rect 41780 297674 41782 297691
rect 41782 297674 41834 297691
rect 41834 297674 41836 297691
rect 41876 297230 41932 297286
rect 41780 296729 41836 296768
rect 41780 296712 41782 296729
rect 41782 296712 41834 296729
rect 41834 296712 41836 296729
rect 39860 296490 39916 296546
rect 41684 292938 41740 292994
rect 41588 291014 41644 291070
rect 42452 290718 42508 290774
rect 41780 289756 41836 289812
rect 41780 289238 41836 289294
rect 28724 285094 28780 285150
rect 41876 287775 41932 287814
rect 41876 287758 41878 287775
rect 41878 287758 41930 287775
rect 41930 287758 41932 287775
rect 41876 281690 41932 281746
rect 42452 281542 42508 281598
rect 41972 277990 42028 278046
rect 42164 276510 42220 276566
rect 41780 274142 41836 274198
rect 41780 273550 41836 273606
rect 41780 272810 41836 272866
rect 41780 272218 41836 272274
rect 41780 270590 41836 270646
rect 41780 269998 41836 270054
rect 42164 269258 42220 269314
rect 23348 254754 23404 254810
rect 43316 263338 43372 263394
rect 41588 256826 41644 256882
rect 41780 256530 41836 256586
rect 41780 255977 41782 255994
rect 41782 255977 41834 255994
rect 41834 255977 41836 255994
rect 41780 255938 41836 255977
rect 41780 255533 41782 255550
rect 41782 255533 41834 255550
rect 41834 255533 41836 255550
rect 41780 255494 41836 255533
rect 41780 255067 41836 255106
rect 41780 255050 41782 255067
rect 41782 255050 41834 255067
rect 41834 255050 41836 255067
rect 23156 253866 23212 253922
rect 23540 253866 23596 253922
rect 23060 253274 23116 253330
rect 41780 250018 41836 250074
rect 41492 247798 41548 247854
rect 41588 247354 41644 247410
rect 41684 245874 41740 245930
rect 41684 245282 41740 245338
rect 41588 244877 41590 244894
rect 41590 244877 41642 244894
rect 41642 244877 41644 244894
rect 41588 244838 41644 244877
rect 41588 244246 41644 244302
rect 41876 246614 41932 246670
rect 41780 237882 41836 237938
rect 41780 233294 41836 233350
rect 41780 231074 41836 231130
rect 41780 230334 41836 230390
rect 41780 229594 41836 229650
rect 41780 229002 41836 229058
rect 41780 227374 41836 227430
rect 41876 226782 41932 226838
rect 41780 225894 41836 225950
rect 41780 213649 41782 213666
rect 41782 213649 41834 213666
rect 41834 213649 41836 213666
rect 41780 213610 41836 213649
rect 41780 213131 41782 213148
rect 41782 213131 41834 213148
rect 41834 213131 41836 213148
rect 41780 213092 41836 213131
rect 41588 212761 41590 212778
rect 41590 212761 41642 212778
rect 41642 212761 41644 212778
rect 41588 212722 41644 212761
rect 41780 212169 41782 212186
rect 41782 212169 41834 212186
rect 41834 212169 41836 212186
rect 41780 212130 41836 212169
rect 41780 211651 41782 211668
rect 41782 211651 41834 211668
rect 41834 211651 41836 211668
rect 41780 211612 41836 211651
rect 41588 211281 41590 211298
rect 41590 211281 41642 211298
rect 41642 211281 41644 211298
rect 41588 211242 41644 211281
rect 43508 267186 43564 267242
rect 41780 210689 41782 210706
rect 41782 210689 41834 210706
rect 41834 210689 41836 210706
rect 41780 210650 41836 210689
rect 41780 210097 41782 210114
rect 41782 210097 41834 210114
rect 41834 210097 41836 210114
rect 41780 210058 41836 210097
rect 57716 790810 57772 790866
rect 57620 789626 57676 789682
rect 58196 788442 58252 788498
rect 58388 787258 58444 787314
rect 59636 785482 59692 785538
rect 59156 784890 59212 784946
rect 44756 275326 44812 275382
rect 44660 267334 44716 267390
rect 58676 747594 58732 747650
rect 54740 745983 54796 746022
rect 54740 745966 54742 745983
rect 54742 745966 54794 745983
rect 54794 745966 54796 745983
rect 54644 745818 54700 745874
rect 59636 745670 59692 745726
rect 57620 745226 57676 745282
rect 58484 744042 58540 744098
rect 59636 742858 59692 742914
rect 59732 741674 59788 741730
rect 45044 278582 45100 278638
rect 44948 266446 45004 266502
rect 45908 658794 45964 658850
rect 45908 615578 45964 615634
rect 46196 572362 46252 572418
rect 46676 529294 46732 529350
rect 45236 426434 45292 426490
rect 45236 273254 45292 273310
rect 45140 266298 45196 266354
rect 41588 209801 41590 209818
rect 41590 209801 41642 209818
rect 41642 209801 41644 209818
rect 41588 209762 41644 209801
rect 25652 208874 25708 208930
rect 25556 207838 25612 207894
rect 25844 208282 25900 208338
rect 25748 206802 25804 206858
rect 25652 200882 25708 200938
rect 25556 199994 25612 200050
rect 34292 207394 34348 207450
rect 41876 206580 41932 206636
rect 41588 204286 41644 204342
rect 34292 201474 34348 201530
rect 25844 200882 25900 200938
rect 25748 199698 25804 199754
rect 41780 204138 41836 204194
rect 41780 203176 41836 203232
rect 41780 202658 41836 202714
rect 41780 201217 41782 201234
rect 41782 201217 41834 201234
rect 41834 201217 41836 201234
rect 41780 201178 41836 201217
rect 41972 202105 41974 202122
rect 41974 202105 42026 202122
rect 42026 202105 42028 202122
rect 41972 202066 42028 202105
rect 41972 201661 41974 201678
rect 41974 201661 42026 201678
rect 42026 201661 42028 201678
rect 41972 201622 42028 201661
rect 41780 195258 41836 195314
rect 45428 270590 45484 270646
rect 45716 276214 45772 276270
rect 59636 704378 59692 704434
rect 58772 702641 58774 702658
rect 58774 702641 58826 702658
rect 58826 702641 58828 702658
rect 58772 702602 58828 702641
rect 58676 700826 58732 700882
rect 59252 699642 59308 699698
rect 58868 698458 58924 698514
rect 59636 661162 59692 661218
rect 58772 659403 58828 659442
rect 58772 659386 58774 659403
rect 58774 659386 58826 659403
rect 58826 659386 58828 659403
rect 59156 657610 59212 657666
rect 58196 656426 58252 656482
rect 58388 655242 58444 655298
rect 58964 617946 59020 618002
rect 59636 616209 59638 616226
rect 59638 616209 59690 616226
rect 59690 616209 59692 616226
rect 59636 616170 59692 616209
rect 58964 614394 59020 614450
rect 59636 613210 59692 613266
rect 59540 612026 59596 612082
rect 58964 574730 59020 574786
rect 59636 572993 59638 573010
rect 59638 572993 59690 573010
rect 59690 572993 59692 573010
rect 59636 572954 59692 572993
rect 58964 571178 59020 571234
rect 59348 569994 59404 570050
rect 59540 568810 59596 568866
rect 57716 531662 57772 531718
rect 57620 530478 57676 530534
rect 59636 527535 59692 527574
rect 59636 527518 59638 527535
rect 59638 527518 59690 527535
rect 59690 527518 59692 527535
rect 59348 525890 59404 525946
rect 59636 525019 59692 525058
rect 59636 525002 59638 525019
rect 59638 525002 59690 525019
rect 59690 525002 59692 525019
rect 47828 263486 47884 263542
rect 58484 404086 58540 404142
rect 59348 402310 59404 402366
rect 57716 400534 57772 400590
rect 59636 399942 59692 399998
rect 59732 399350 59788 399406
rect 59540 398166 59596 398222
rect 58484 360870 58540 360926
rect 59156 359686 59212 359742
rect 57716 357466 57772 357522
rect 58388 356134 58444 356190
rect 59636 356726 59692 356782
rect 58484 354950 58540 355006
rect 41780 190078 41836 190134
rect 41876 187858 41932 187914
rect 41780 187118 41836 187174
rect 41780 186674 41836 186730
rect 41780 185786 41836 185842
rect 42164 184158 42220 184214
rect 41876 183566 41932 183622
rect 42068 182826 42124 182882
rect 58484 317654 58540 317710
rect 59156 316470 59212 316526
rect 59060 314102 59116 314158
rect 59636 313510 59692 313566
rect 59732 312918 59788 312974
rect 59540 311734 59596 311790
rect 50612 275178 50668 275234
rect 50420 275030 50476 275086
rect 59252 295158 59308 295214
rect 59636 292790 59692 292846
rect 58196 292642 58252 292698
rect 60308 293974 60364 294030
rect 60212 291458 60268 291514
rect 57620 284502 57676 284558
rect 58580 283318 58636 283374
rect 59540 289238 59596 289294
rect 59156 288071 59212 288110
rect 59156 288054 59158 288071
rect 59158 288054 59210 288071
rect 59210 288054 59212 288071
rect 59252 286870 59308 286926
rect 58964 285686 59020 285742
rect 58388 280950 58444 281006
rect 58580 279766 58636 279822
rect 59636 282430 59692 282486
rect 61940 278434 61996 278490
rect 62132 278286 62188 278342
rect 62036 266890 62092 266946
rect 61844 266742 61900 266798
rect 62324 602110 62380 602166
rect 62324 278138 62380 278194
rect 62516 547202 62572 547258
rect 62708 544390 62764 544446
rect 62612 277990 62668 278046
rect 62900 277842 62956 277898
rect 62996 277694 63052 277750
rect 62708 273550 62764 273606
rect 62516 273402 62572 273458
rect 70580 272070 70636 272126
rect 69428 269554 69484 269610
rect 67028 269406 67084 269462
rect 72980 272218 73036 272274
rect 71732 269258 71788 269314
rect 78836 272366 78892 272422
rect 77588 269702 77644 269758
rect 62420 267038 62476 267094
rect 62228 266594 62284 266650
rect 88340 272514 88396 272570
rect 91892 272662 91948 272718
rect 139124 269850 139180 269906
rect 148340 244542 148396 244598
rect 148244 239658 148300 239714
rect 147668 232258 147724 232314
rect 146900 229890 146956 229946
rect 147668 218938 147724 218994
rect 147284 217771 147340 217810
rect 147284 217754 147286 217771
rect 147286 217754 147338 217771
rect 147338 217754 147340 217771
rect 147380 214794 147436 214850
rect 147572 214054 147628 214110
rect 146900 212887 146956 212926
rect 146900 212870 146902 212887
rect 146902 212870 146954 212887
rect 146954 212870 146956 212887
rect 147380 211686 147436 211742
rect 147380 210371 147436 210410
rect 147380 210354 147382 210371
rect 147382 210354 147434 210371
rect 147434 210354 147436 210371
rect 146900 209170 146956 209226
rect 146996 207986 147052 208042
rect 147092 206358 147148 206414
rect 147668 204434 147724 204490
rect 147476 199550 147532 199606
rect 147284 195850 147340 195906
rect 147284 190966 147340 191022
rect 147668 175130 147724 175186
rect 148532 243358 148588 243414
rect 148436 234774 148492 234830
rect 148724 242026 148780 242082
rect 148628 236698 148684 236754
rect 149012 240842 149068 240898
rect 148820 238474 148876 238530
rect 148724 170246 148780 170302
rect 148916 233590 148972 233646
rect 148916 173946 148972 174002
rect 148724 166250 148780 166306
rect 148532 165510 148588 165566
rect 148340 164326 148396 164382
rect 148244 161810 148300 161866
rect 146900 159442 146956 159498
rect 147092 139906 147148 139962
rect 147188 130303 147244 130342
rect 147188 130286 147190 130303
rect 147190 130286 147242 130303
rect 147242 130286 147244 130303
rect 148436 160626 148492 160682
rect 148148 125402 148204 125458
rect 147668 108399 147724 108438
rect 147668 108382 147670 108399
rect 147670 108382 147722 108399
rect 147722 108382 147724 108399
rect 146996 107198 147052 107254
rect 148628 163142 148684 163198
rect 148820 155742 148876 155798
rect 149108 235958 149164 236014
rect 149396 231091 149452 231130
rect 149396 231074 149398 231091
rect 149398 231074 149450 231091
rect 149450 231074 149452 231091
rect 149396 228114 149452 228170
rect 149300 227374 149356 227430
rect 149396 226338 149452 226394
rect 149492 225154 149548 225210
rect 149492 223822 149548 223878
rect 149396 222638 149452 222694
rect 149492 221454 149548 221510
rect 149396 219678 149452 219734
rect 149396 216570 149452 216626
rect 149396 205618 149452 205674
rect 149492 203250 149548 203306
rect 149396 201639 149452 201678
rect 149396 201622 149398 201639
rect 149398 201622 149450 201639
rect 149450 201622 149452 201639
rect 149396 200734 149452 200790
rect 149300 198366 149356 198422
rect 149396 197034 149452 197090
rect 149492 194666 149548 194722
rect 149396 193334 149452 193390
rect 149396 192150 149452 192206
rect 149396 189782 149452 189838
rect 149300 187414 149356 187470
rect 149204 186230 149260 186286
rect 149588 188006 149644 188062
rect 149396 184454 149452 184510
rect 149492 183714 149548 183770
rect 149396 182530 149452 182586
rect 149492 181346 149548 181402
rect 149300 179570 149356 179626
rect 149396 178830 149452 178886
rect 149492 177646 149548 177702
rect 149396 176462 149452 176518
rect 149204 170986 149260 171042
rect 149012 168026 149068 168082
rect 148532 129102 148588 129158
rect 149588 172762 149644 172818
rect 149492 169062 149548 169118
rect 148820 141255 148876 141294
rect 148820 141238 148822 141255
rect 148822 141238 148874 141255
rect 148874 141238 148876 141255
rect 149300 157666 149356 157722
rect 149204 153078 149260 153134
rect 149204 152042 149260 152098
rect 149204 149861 149206 149878
rect 149206 149861 149258 149878
rect 149258 149861 149260 149878
rect 149204 149822 149260 149861
rect 149204 147306 149260 147362
rect 149204 144494 149260 144550
rect 149204 142422 149260 142478
rect 149204 138722 149260 138778
rect 149204 135910 149260 135966
rect 148820 132654 148876 132710
rect 148532 115190 148588 115246
rect 148244 111934 148300 111990
rect 148436 110898 148492 110954
rect 148340 104682 148396 104738
rect 148532 106014 148588 106070
rect 148628 102314 148684 102370
rect 148916 130878 148972 130934
rect 149492 135022 149548 135078
rect 149396 133838 149452 133894
rect 149684 156926 149740 156982
rect 149684 154558 149740 154614
rect 149684 150858 149740 150914
rect 149684 148490 149740 148546
rect 149684 146122 149740 146178
rect 149684 143606 149740 143662
rect 149684 137538 149740 137594
rect 149108 127918 149164 127974
rect 149012 122442 149068 122498
rect 149588 126586 149644 126642
rect 149300 124218 149356 124274
rect 149204 121702 149260 121758
rect 149396 120518 149452 120574
rect 149492 119334 149548 119390
rect 149396 118167 149452 118206
rect 149396 118150 149398 118167
rect 149398 118150 149450 118167
rect 149450 118150 149452 118167
rect 149396 116818 149452 116874
rect 149492 115634 149548 115690
rect 149396 115190 149452 115246
rect 149492 114450 149548 114506
rect 149396 113118 149452 113174
rect 149396 109583 149452 109622
rect 149396 109566 149398 109583
rect 149398 109566 149450 109583
rect 149450 109566 149452 109583
rect 149588 103498 149644 103554
rect 149396 100851 149452 100890
rect 149396 100834 149398 100851
rect 149398 100834 149450 100851
rect 149450 100834 149452 100851
rect 149492 99798 149548 99854
rect 149396 98614 149452 98670
rect 149492 97430 149548 97486
rect 149396 95654 149452 95710
rect 149492 93730 149548 93786
rect 149396 92546 149452 92602
rect 149204 91362 149260 91418
rect 148724 86495 148780 86534
rect 148724 86478 148726 86495
rect 148726 86478 148778 86495
rect 148778 86478 148780 86495
rect 148436 85294 148492 85350
rect 147092 84110 147148 84166
rect 148244 81594 148300 81650
rect 149108 82334 149164 82390
rect 148820 77894 148876 77950
rect 149300 90178 149356 90234
rect 149396 88994 149452 89050
rect 149492 87366 149548 87422
rect 149684 94914 149740 94970
rect 149588 80410 149644 80466
rect 149204 76710 149260 76766
rect 149012 73010 149068 73066
rect 149108 71974 149164 72030
rect 149396 75526 149452 75582
rect 149300 73750 149356 73806
rect 149684 79226 149740 79282
rect 184340 219530 184396 219586
rect 184340 218829 184342 218846
rect 184342 218829 184394 218846
rect 184394 218829 184396 218846
rect 184340 218790 184396 218829
rect 184340 199698 184396 199754
rect 184244 197626 184300 197682
rect 192596 269406 192652 269462
rect 194420 272218 194476 272274
rect 196628 272366 196684 272422
rect 193748 272070 193804 272126
rect 193076 269554 193132 269610
rect 194228 269258 194284 269314
rect 196148 269702 196204 269758
rect 199220 272514 199276 272570
rect 200468 272662 200524 272718
rect 208148 268074 208204 268130
rect 213332 269850 213388 269906
rect 214292 268074 214348 268130
rect 341684 274438 341740 274494
rect 347636 274586 347692 274642
rect 350228 274734 350284 274790
rect 353396 274882 353452 274938
rect 370100 271626 370156 271682
rect 369620 271478 369676 271534
rect 367892 270442 367948 270498
rect 368372 269110 368428 269166
rect 374324 268814 374380 268870
rect 375572 271774 375628 271830
rect 377012 270294 377068 270350
rect 379028 276066 379084 276122
rect 378644 271922 378700 271978
rect 383444 275918 383500 275974
rect 382964 273106 383020 273162
rect 382388 270738 382444 270794
rect 385556 270146 385612 270202
rect 388724 270738 388780 270794
rect 388436 269998 388492 270054
rect 390356 275770 390412 275826
rect 390164 272958 390220 273014
rect 391508 269850 391564 269906
rect 392756 272810 392812 272866
rect 393908 276658 393964 276714
rect 396692 276510 396748 276566
rect 397076 268962 397132 269018
rect 398900 275622 398956 275678
rect 398708 272662 398764 272718
rect 402548 276806 402604 276862
rect 403028 269702 403084 269758
rect 404180 272514 404236 272570
rect 405620 269554 405676 269610
rect 407828 275474 407884 275530
rect 407252 272366 407308 272422
rect 408884 273254 408940 273310
rect 410900 272218 410956 272274
rect 410420 269406 410476 269462
rect 411764 272070 411820 272126
rect 411572 269258 411628 269314
rect 474836 274438 474892 274494
rect 489044 274586 489100 274642
rect 496052 274734 496108 274790
rect 503156 274882 503212 274938
rect 508244 268814 508300 268870
rect 526964 276806 527020 276862
rect 532820 268962 532876 269018
rect 539828 270442 539884 270498
rect 540980 269110 541036 269166
rect 544532 271626 544588 271682
rect 543380 271478 543436 271534
rect 558740 271774 558796 271830
rect 566996 276066 567052 276122
rect 565844 271922 565900 271978
rect 562292 270294 562348 270350
rect 577652 275918 577708 275974
rect 576500 273106 576556 273162
rect 583604 270146 583660 270202
rect 595412 275770 595468 275826
rect 594164 272958 594220 273014
rect 590612 269998 590668 270054
rect 597716 269850 597772 269906
rect 601268 272810 601324 272866
rect 603668 276658 603724 276714
rect 610772 276510 610828 276566
rect 616628 275622 616684 275678
rect 615476 272662 615532 272718
rect 626132 269702 626188 269758
rect 629684 272514 629740 272570
rect 633236 269554 633292 269610
rect 637940 275474 637996 275530
rect 636788 272366 636844 272422
rect 646484 275326 646540 275382
rect 646196 272218 646252 272274
rect 645044 269406 645100 269462
rect 420404 262171 420460 262210
rect 420404 262154 420406 262171
rect 420406 262154 420458 262171
rect 420458 262154 420460 262171
rect 420404 259786 420460 259842
rect 191540 259342 191596 259398
rect 185492 198218 185548 198274
rect 184436 196738 184492 196794
rect 184340 195998 184396 196054
rect 184340 195258 184396 195314
rect 184436 194370 184492 194426
rect 184532 193778 184588 193834
rect 184436 192890 184492 192946
rect 184340 192298 184396 192354
rect 184532 191410 184588 191466
rect 184628 190670 184684 190726
rect 184340 189969 184342 189986
rect 184342 189969 184394 189986
rect 184394 189969 184396 189986
rect 184340 189930 184396 189969
rect 184532 189190 184588 189246
rect 184436 188450 184492 188506
rect 184340 187562 184396 187618
rect 184340 186822 184396 186878
rect 184436 186082 184492 186138
rect 184628 185342 184684 185398
rect 184532 184602 184588 184658
rect 184340 183862 184396 183918
rect 184436 183122 184492 183178
rect 184532 181494 184588 181550
rect 184340 180754 184396 180810
rect 184436 180014 184492 180070
rect 184628 179274 184684 179330
rect 184532 178534 184588 178590
rect 184340 177054 184396 177110
rect 184436 176166 184492 176222
rect 184340 175591 184396 175630
rect 184340 175574 184342 175591
rect 184342 175574 184394 175591
rect 184394 175574 184396 175591
rect 184436 173946 184492 174002
rect 184340 172466 184396 172522
rect 184532 171726 184588 171782
rect 184628 170838 184684 170894
rect 184436 170246 184492 170302
rect 184340 169358 184396 169414
rect 184436 168618 184492 168674
rect 184628 167878 184684 167934
rect 184532 167138 184588 167194
rect 184340 166398 184396 166454
rect 184436 165658 184492 165714
rect 184532 164770 184588 164826
rect 184340 164047 184396 164086
rect 184340 164030 184342 164047
rect 184342 164030 184394 164047
rect 184394 164030 184396 164047
rect 184340 163290 184396 163346
rect 185300 162550 185356 162606
rect 184436 161810 184492 161866
rect 184340 160922 184396 160978
rect 184436 160330 184492 160386
rect 184532 159442 184588 159498
rect 184628 158850 184684 158906
rect 184340 156482 184396 156538
rect 184532 157962 184588 158018
rect 184628 157370 184684 157426
rect 184436 155594 184492 155650
rect 184340 155002 184396 155058
rect 184436 154114 184492 154170
rect 184532 153522 184588 153578
rect 184628 152634 184684 152690
rect 184340 151894 184396 151950
rect 184532 151154 184588 151210
rect 184436 150414 184492 150470
rect 184340 149713 184342 149730
rect 184342 149713 184394 149730
rect 184394 149713 184396 149730
rect 184340 149674 184396 149713
rect 184436 148934 184492 148990
rect 184340 148046 184396 148102
rect 184532 147306 184588 147362
rect 184340 145086 184396 145142
rect 185396 146566 185452 146622
rect 184436 144346 184492 144402
rect 184340 142718 184396 142774
rect 184436 142126 184492 142182
rect 184628 143606 184684 143662
rect 184532 141238 184588 141294
rect 184340 140498 184396 140554
rect 184436 139758 184492 139814
rect 184532 138870 184588 138926
rect 186068 213462 186124 213518
rect 186260 214942 186316 214998
rect 186452 210502 186508 210558
rect 186356 207246 186412 207302
rect 186836 221010 186892 221066
rect 187124 243358 187180 243414
rect 187028 220270 187084 220326
rect 186932 218050 186988 218106
rect 186740 216422 186796 216478
rect 187028 211982 187084 212038
rect 186644 209022 186700 209078
rect 186548 205174 186604 205230
rect 186164 204286 186220 204342
rect 185972 202806 186028 202862
rect 190196 251646 190252 251702
rect 420404 256974 420460 257030
rect 420404 255198 420460 255254
rect 420404 252830 420460 252886
rect 420308 250462 420364 250518
rect 420404 248094 420460 248150
rect 420404 245282 420460 245338
rect 420308 243506 420364 243562
rect 412436 241434 412492 241490
rect 567380 241434 567436 241490
rect 412244 240694 412300 240750
rect 412148 240398 412204 240454
rect 412052 240250 412108 240306
rect 292148 228854 292204 228910
rect 299348 234922 299404 234978
rect 299444 234774 299500 234830
rect 298964 234626 299020 234682
rect 301652 235070 301708 235126
rect 302900 231074 302956 231130
rect 307604 231222 307660 231278
rect 310676 228262 310732 228318
rect 313460 228410 313516 228466
rect 316724 231370 316780 231426
rect 318932 225450 318988 225506
rect 319508 231518 319564 231574
rect 321716 225598 321772 225654
rect 322484 231666 322540 231722
rect 328052 225746 328108 225802
rect 330260 233146 330316 233202
rect 330836 227374 330892 227430
rect 333044 228558 333100 228614
rect 333812 227226 333868 227282
rect 334868 232998 334924 233054
rect 336884 227078 336940 227134
rect 339380 228706 339436 228762
rect 341588 234478 341644 234534
rect 342548 235958 342604 236014
rect 342164 230334 342220 230390
rect 343028 226930 343084 226986
rect 342644 225302 342700 225358
rect 344180 235070 344236 235126
rect 344372 235070 344428 235126
rect 345524 230186 345580 230242
rect 344756 226782 344812 226838
rect 347636 233738 347692 233794
rect 349748 234922 349804 234978
rect 351380 225894 351436 225950
rect 354356 234774 354412 234830
rect 354260 234626 354316 234682
rect 354932 235662 354988 235718
rect 354164 224562 354220 224618
rect 356756 234774 356812 234830
rect 356852 234626 356908 234682
rect 357524 224414 357580 224470
rect 359060 232850 359116 232906
rect 358964 229890 359020 229946
rect 359828 228854 359884 228910
rect 359732 224266 359788 224322
rect 359444 222934 359500 222990
rect 360308 223970 360364 224026
rect 361460 224118 361516 224174
rect 363572 230038 363628 230094
rect 363476 223822 363532 223878
rect 365780 229742 365836 229798
rect 367220 234182 367276 234238
rect 367604 223674 367660 223730
rect 368948 236254 369004 236310
rect 370388 236698 370444 236754
rect 370292 234034 370348 234090
rect 370772 232702 370828 232758
rect 372212 236994 372268 237050
rect 373460 236846 373516 236902
rect 373076 229594 373132 229650
rect 374900 236550 374956 236606
rect 375380 232554 375436 232610
rect 376724 236402 376780 236458
rect 376340 233886 376396 233942
rect 377780 236254 377836 236310
rect 377972 236254 378028 236310
rect 379124 234330 379180 234386
rect 378932 232406 378988 232462
rect 377588 223526 377644 223582
rect 379796 223230 379852 223286
rect 382580 236698 382636 236754
rect 382772 236698 382828 236754
rect 381716 232258 381772 232314
rect 381332 229298 381388 229354
rect 381236 223378 381292 223434
rect 382964 231814 383020 231870
rect 383540 229446 383596 229502
rect 382772 222786 382828 222842
rect 384980 232110 385036 232166
rect 385364 231962 385420 232018
rect 384404 229150 384460 229206
rect 385940 235958 385996 236014
rect 385844 235514 385900 235570
rect 384308 223082 384364 223138
rect 387956 236846 388012 236902
rect 387668 235218 387724 235274
rect 388340 236737 388342 236754
rect 388342 236737 388394 236754
rect 388394 236737 388396 236754
rect 388340 236698 388396 236737
rect 388724 236994 388780 237050
rect 388724 236863 388780 236902
rect 388724 236846 388726 236863
rect 388726 236846 388778 236863
rect 388778 236846 388780 236863
rect 388628 236402 388684 236458
rect 388820 236254 388876 236310
rect 389012 236254 389068 236310
rect 389012 236106 389068 236162
rect 389396 235958 389452 236014
rect 391796 235070 391852 235126
rect 391604 226634 391660 226690
rect 392564 235849 392566 235866
rect 392566 235849 392618 235866
rect 392618 235849 392620 235866
rect 392564 235810 392620 235849
rect 392564 234330 392620 234386
rect 392564 233590 392620 233646
rect 393140 235827 393196 235866
rect 393140 235810 393142 235827
rect 393142 235810 393194 235827
rect 393194 235810 393196 235827
rect 393428 234922 393484 234978
rect 392852 234626 392908 234682
rect 393044 234626 393100 234682
rect 392852 234330 392908 234386
rect 394484 226486 394540 226542
rect 394100 226338 394156 226394
rect 398996 236994 399052 237050
rect 398708 236846 398764 236902
rect 399860 235070 399916 235126
rect 400436 234774 400492 234830
rect 399476 228854 399532 228910
rect 401396 235810 401452 235866
rect 403124 235958 403180 236014
rect 403316 235662 403372 235718
rect 403124 229002 403180 229058
rect 403988 235366 404044 235422
rect 405524 235662 405580 235718
rect 405428 234774 405484 234830
rect 405716 234330 405772 234386
rect 405908 234182 405964 234238
rect 406964 233590 407020 233646
rect 405812 226190 405868 226246
rect 405716 222638 405772 222694
rect 407252 234182 407308 234238
rect 407924 234626 407980 234682
rect 408116 234626 408172 234682
rect 408692 236994 408748 237050
rect 408884 236994 408940 237050
rect 408788 236698 408844 236754
rect 408980 236885 408982 236902
rect 408982 236885 409034 236902
rect 409034 236885 409036 236902
rect 408980 236846 409036 236885
rect 408692 236254 408748 236310
rect 409172 236254 409228 236310
rect 408788 236106 408844 236162
rect 408788 235810 408844 235866
rect 408788 234922 408844 234978
rect 409364 236846 409420 236902
rect 408500 234330 408556 234386
rect 407636 226042 407692 226098
rect 412340 239954 412396 240010
rect 420308 241138 420364 241194
rect 412724 240842 412780 240898
rect 412628 240546 412684 240602
rect 412532 240102 412588 240158
rect 566708 240694 566764 240750
rect 544820 240250 544876 240306
rect 541460 240102 541516 240158
rect 413396 238918 413452 238974
rect 413684 238622 413740 238678
rect 413972 238326 414028 238382
rect 414260 238178 414316 238234
rect 414452 238030 414508 238086
rect 414452 236254 414508 236310
rect 414260 233886 414316 233942
rect 411572 233738 411628 233794
rect 414644 236254 414700 236310
rect 415700 231074 415756 231130
rect 424724 231222 424780 231278
rect 428276 234034 428332 234090
rect 430868 228262 430924 228318
rect 436916 228410 436972 228466
rect 442868 231370 442924 231426
rect 445172 225450 445228 225506
rect 448916 231518 448972 231574
rect 451220 225598 451276 225654
rect 455156 231666 455212 231722
rect 457268 225302 457324 225358
rect 463316 225746 463372 225802
rect 470132 233146 470188 233202
rect 469364 227374 469420 227430
rect 479156 232998 479212 233054
rect 476180 228558 476236 228614
rect 475316 227226 475372 227282
rect 481460 227078 481516 227134
rect 488276 228706 488332 228762
rect 487508 225894 487564 225950
rect 490484 234478 490540 234534
rect 495380 234182 495436 234238
rect 494228 230334 494284 230390
rect 493460 226930 493516 226986
rect 497972 230186 498028 230242
rect 498836 226782 498892 226838
rect 512180 234330 512236 234386
rect 518420 224562 518476 224618
rect 525236 232850 525292 232906
rect 524468 224414 524524 224470
rect 522932 222638 522988 222694
rect 527540 229890 527596 229946
rect 526676 222934 526732 222990
rect 528980 224266 529036 224322
rect 530516 223970 530572 224026
rect 532052 224118 532108 224174
rect 538004 238030 538060 238086
rect 534260 230038 534316 230094
rect 544340 238326 544396 238382
rect 536564 223822 536620 223878
rect 538868 229742 538924 229798
rect 541076 222786 541132 222842
rect 544052 223674 544108 223730
rect 550868 239954 550924 240010
rect 550196 238622 550252 238678
rect 553940 238918 553996 238974
rect 559892 238178 559948 238234
rect 559220 236550 559276 236606
rect 557684 236402 557740 236458
rect 551636 232702 551692 232758
rect 553940 229594 553996 229650
rect 566036 236846 566092 236902
rect 562196 236698 562252 236754
rect 560756 232554 560812 232610
rect 564500 232406 564556 232462
rect 562964 223526 563020 223582
rect 581780 240842 581836 240898
rect 573140 236994 573196 237050
rect 570452 232258 570508 232314
rect 568244 223230 568300 223286
rect 571316 223378 571372 223434
rect 573524 229446 573580 229502
rect 572756 229298 572812 229354
rect 580340 235514 580396 235570
rect 576596 232110 576652 232166
rect 575828 231814 575884 231870
rect 578036 231962 578092 232018
rect 577268 223082 577324 223138
rect 578900 229150 578956 229206
rect 593012 236106 593068 236162
rect 591476 235810 591532 235866
rect 583412 235218 583468 235274
rect 591668 226634 591724 226690
rect 595892 235958 595948 236014
rect 595412 235070 595468 235126
rect 594644 234922 594700 234978
rect 597428 235662 597484 235718
rect 596180 235366 596236 235422
rect 596948 226486 597004 226542
rect 596180 226338 596236 226394
rect 599924 229002 599980 229058
rect 610484 240546 610540 240602
rect 607508 228854 607564 228910
rect 627188 240398 627244 240454
rect 621140 236254 621196 236310
rect 618836 234774 618892 234830
rect 620372 226190 620428 226246
rect 624884 234626 624940 234682
rect 623348 226042 623404 226098
rect 640148 212278 640204 212334
rect 640148 211538 640204 211594
rect 190292 201326 190348 201382
rect 640148 200882 640204 200938
rect 190292 200512 190348 200568
rect 640148 200142 640204 200198
rect 187220 199106 187276 199162
rect 185780 182382 185836 182438
rect 185588 173206 185644 173262
rect 186068 138278 186124 138334
rect 640244 185638 640300 185694
rect 640244 184898 640300 184954
rect 645140 182974 645196 183030
rect 645140 179274 645196 179330
rect 186740 177646 186796 177702
rect 645140 174873 645142 174890
rect 645142 174873 645194 174890
rect 645194 174873 645196 174890
rect 645140 174834 645196 174873
rect 186260 174686 186316 174742
rect 186164 137390 186220 137446
rect 185972 136798 186028 136854
rect 185492 135910 185548 135966
rect 184340 134430 184396 134486
rect 184436 133690 184492 133746
rect 645140 171025 645142 171042
rect 645142 171025 645194 171042
rect 645194 171025 645196 171042
rect 645140 170986 645196 171025
rect 645140 167730 645196 167786
rect 645140 163329 645142 163346
rect 645142 163329 645194 163346
rect 645194 163329 645196 163346
rect 645140 163290 645196 163329
rect 645140 159442 645196 159498
rect 645140 155446 645196 155502
rect 645140 152525 645142 152542
rect 645142 152525 645194 152542
rect 645194 152525 645196 152542
rect 645140 152486 645196 152525
rect 645140 148046 645196 148102
rect 186740 145826 186796 145882
rect 186260 135170 186316 135226
rect 184532 132950 184588 133006
rect 184340 131470 184396 131526
rect 184628 132210 184684 132266
rect 184532 130582 184588 130638
rect 184436 129842 184492 129898
rect 184340 129102 184396 129158
rect 184436 128362 184492 128418
rect 184532 127622 184588 127678
rect 184628 126882 184684 126938
rect 184436 125994 184492 126050
rect 184340 125402 184396 125458
rect 184532 124514 184588 124570
rect 184340 123813 184342 123830
rect 184342 123813 184394 123830
rect 184394 123813 184396 123830
rect 184340 123774 184396 123813
rect 184436 123034 184492 123090
rect 184340 122146 184396 122202
rect 184532 121554 184588 121610
rect 184436 120666 184492 120722
rect 184532 120074 184588 120130
rect 184340 119186 184396 119242
rect 184628 118594 184684 118650
rect 184340 117706 184396 117762
rect 184436 116966 184492 117022
rect 184532 116226 184588 116282
rect 184628 115338 184684 115394
rect 184340 114746 184396 114802
rect 184436 113858 184492 113914
rect 184532 113118 184588 113174
rect 184340 111638 184396 111694
rect 184436 110898 184492 110954
rect 184532 110158 184588 110214
rect 184436 109309 184438 109326
rect 184438 109309 184490 109326
rect 184490 109309 184492 109326
rect 184436 109270 184492 109309
rect 645716 128954 645772 129010
rect 648596 272070 648652 272126
rect 647348 269258 647404 269314
rect 646580 267334 646636 267390
rect 185684 112378 185740 112434
rect 185588 108678 185644 108734
rect 646676 144198 646732 144254
rect 655124 777638 655180 777694
rect 655028 774678 655084 774734
rect 654356 773494 654412 773550
rect 654164 730130 654220 730186
rect 654068 728502 654124 728558
rect 655412 778230 655468 778286
rect 655220 775714 655276 775770
rect 655316 734422 655372 734478
rect 655220 731610 655276 731666
rect 655124 689430 655180 689486
rect 654356 686914 654412 686970
rect 654164 685286 654220 685342
rect 654068 684546 654124 684602
rect 649748 263338 649804 263394
rect 646772 140942 646828 140998
rect 654164 640590 654220 640646
rect 655604 775862 655660 775918
rect 655508 732646 655564 732702
rect 655412 688394 655468 688450
rect 655316 642958 655372 643014
rect 655220 597818 655276 597874
rect 655124 595302 655180 595358
rect 653780 592934 653836 592990
rect 655124 553270 655180 553326
rect 654164 548534 654220 548590
rect 655700 731314 655756 731370
rect 655604 687062 655660 687118
rect 655508 642366 655564 642422
rect 655412 596634 655468 596690
rect 655316 552086 655372 552142
rect 655700 640738 655756 640794
rect 655604 595450 655660 595506
rect 655508 551050 655564 551106
rect 655796 639110 655852 639166
rect 655988 638222 656044 638278
rect 655796 594118 655852 594174
rect 655700 550902 655756 550958
rect 656564 549718 656620 549774
rect 655124 373302 655180 373358
rect 655508 374338 655564 374394
rect 655316 372118 655372 372174
rect 653780 370934 653836 370990
rect 655220 329790 655276 329846
rect 655124 328014 655180 328070
rect 655316 327422 655372 327478
rect 654164 326238 654220 326294
rect 654164 303298 654220 303354
rect 654068 302114 654124 302170
rect 654260 300930 654316 300986
rect 654164 298710 654220 298766
rect 656468 297526 656524 297582
rect 656084 296786 656140 296842
rect 654164 296638 654220 296694
rect 655892 293974 655948 294030
rect 655796 290866 655852 290922
rect 655604 289238 655660 289294
rect 655412 288054 655468 288110
rect 653780 284502 653836 284558
rect 655124 283318 655180 283374
rect 654260 279766 654316 279822
rect 652244 267186 652300 267242
rect 647060 134726 647116 134782
rect 647828 130878 647884 130934
rect 646964 127622 647020 127678
rect 646868 125698 646924 125754
rect 646580 123774 646636 123830
rect 646484 121998 646540 122054
rect 655316 282282 655372 282338
rect 655220 280950 655276 281006
rect 655508 285686 655564 285742
rect 655700 286870 655756 286926
rect 655988 292790 656044 292846
rect 656180 291606 656236 291662
rect 656564 295158 656620 295214
rect 647924 119482 647980 119538
rect 645236 117558 645292 117614
rect 647924 115634 647980 115690
rect 669524 275030 669580 275086
rect 669716 275178 669772 275234
rect 669908 277694 669964 277750
rect 670100 277842 670156 277898
rect 676052 891467 676108 891506
rect 676052 891450 676054 891467
rect 676054 891450 676106 891467
rect 676106 891450 676108 891467
rect 676052 890431 676108 890470
rect 676052 890414 676054 890431
rect 676054 890414 676106 890431
rect 676106 890414 676108 890431
rect 680276 890118 680332 890174
rect 676244 889230 676300 889286
rect 676052 887898 676108 887954
rect 676052 887380 676108 887436
rect 680084 888638 680140 888694
rect 679700 886714 679756 886770
rect 676052 885456 676108 885512
rect 676052 884938 676108 884994
rect 676244 884215 676300 884254
rect 676244 884198 676246 884215
rect 676246 884198 676298 884215
rect 676298 884198 676300 884215
rect 676052 883976 676108 884032
rect 676052 883458 676108 883514
rect 679892 886122 679948 886178
rect 679796 882718 679852 882774
rect 679796 882126 679852 882182
rect 679988 885678 680044 885734
rect 680180 888194 680236 888250
rect 685460 882126 685516 882182
rect 685460 881682 685516 881738
rect 675380 787998 675436 788054
rect 675668 787110 675724 787166
rect 675380 786666 675436 786722
rect 675380 784742 675436 784798
rect 675764 784150 675820 784206
rect 675284 783410 675340 783466
rect 675476 780598 675532 780654
rect 675764 779858 675820 779914
rect 675764 779118 675820 779174
rect 675764 777638 675820 777694
rect 675764 775418 675820 775474
rect 670484 308922 670540 308978
rect 670484 278582 670540 278638
rect 670292 277990 670348 278046
rect 674516 728502 674572 728558
rect 674996 771866 675052 771922
rect 674900 731610 674956 731666
rect 675284 741082 675340 741138
rect 675476 740342 675532 740398
rect 675284 739602 675340 739658
rect 675764 737974 675820 738030
rect 675668 735458 675724 735514
rect 679796 728058 679852 728114
rect 676340 715478 676396 715534
rect 676148 714886 676204 714942
rect 676244 714755 676300 714794
rect 676244 714738 676246 714755
rect 676246 714738 676298 714755
rect 676298 714738 676300 714755
rect 676052 714185 676054 714202
rect 676054 714185 676106 714202
rect 676106 714185 676108 714202
rect 676052 714146 676108 714185
rect 676244 713423 676300 713462
rect 676244 713406 676246 713423
rect 676246 713406 676298 713423
rect 676298 713406 676300 713423
rect 676052 713127 676108 713166
rect 676052 713110 676054 713127
rect 676054 713110 676106 713127
rect 676106 713110 676108 713127
rect 676052 712683 676108 712722
rect 676052 712666 676054 712683
rect 676054 712666 676106 712683
rect 676106 712666 676108 712683
rect 676244 711943 676300 711982
rect 676244 711926 676246 711943
rect 676246 711926 676298 711943
rect 676298 711926 676300 711943
rect 676052 711573 676108 711612
rect 676052 711556 676054 711573
rect 676054 711556 676106 711573
rect 676106 711556 676108 711573
rect 676052 708522 676108 708578
rect 676052 708152 676108 708208
rect 679796 706894 679852 706950
rect 676052 705579 676108 705618
rect 676052 705562 676054 705579
rect 676054 705562 676106 705579
rect 676106 705562 676108 705579
rect 676244 704861 676246 704878
rect 676246 704861 676298 704878
rect 676298 704861 676300 704878
rect 676244 704822 676300 704861
rect 679988 704378 680044 704434
rect 679796 703342 679852 703398
rect 679988 703342 680044 703398
rect 679796 702898 679852 702954
rect 675380 697866 675436 697922
rect 675764 697126 675820 697182
rect 675188 696978 675244 697034
rect 675572 694758 675628 694814
rect 675764 694166 675820 694222
rect 674900 686470 674956 686526
rect 676244 668710 676300 668766
rect 676244 668266 676300 668322
rect 676052 667970 676108 668026
rect 675956 667565 675958 667582
rect 675958 667565 676010 667582
rect 676010 667565 676012 667582
rect 675956 667526 676012 667565
rect 675956 666063 676012 666102
rect 675956 666046 675958 666063
rect 675958 666046 676010 666063
rect 676010 666046 676012 666063
rect 675956 665493 675958 665510
rect 675958 665493 676010 665510
rect 676010 665493 676012 665510
rect 675956 665454 676012 665493
rect 676244 666803 676300 666842
rect 676244 666786 676246 666803
rect 676246 666786 676298 666803
rect 676298 666786 676300 666803
rect 676148 666677 676150 666694
rect 676150 666677 676202 666694
rect 676202 666677 676204 666694
rect 676148 666638 676204 666677
rect 675956 665027 676012 665066
rect 675956 665010 675958 665027
rect 675958 665010 676010 665027
rect 676010 665010 676012 665027
rect 676052 663974 676108 664030
rect 676052 661976 676108 662032
rect 676052 660461 676054 660478
rect 676054 660461 676106 660478
rect 676106 660461 676108 660478
rect 676052 660422 676108 660461
rect 676052 660091 676054 660108
rect 676054 660091 676106 660108
rect 676106 660091 676108 660108
rect 676052 660052 676108 660091
rect 676244 659721 676246 659738
rect 676246 659721 676298 659738
rect 676298 659721 676300 659738
rect 676244 659682 676300 659721
rect 676052 658611 676054 658628
rect 676054 658611 676106 658628
rect 676106 658611 676108 658628
rect 676052 658572 676108 658611
rect 676244 658241 676246 658258
rect 676246 658241 676298 658258
rect 676298 658241 676300 658258
rect 676244 658202 676300 658241
rect 679988 657314 680044 657370
rect 679796 656722 679852 656778
rect 679988 656722 680044 656778
rect 679796 656278 679852 656334
rect 675380 652578 675436 652634
rect 675476 652134 675532 652190
rect 675380 651394 675436 651450
rect 675380 649618 675436 649674
rect 675668 645326 675724 645382
rect 675284 639998 675340 640054
rect 675764 638518 675820 638574
rect 678164 636594 678220 636650
rect 676244 625050 676300 625106
rect 676148 624606 676204 624662
rect 676052 623979 676054 623996
rect 676054 623979 676106 623996
rect 676106 623979 676108 623996
rect 676052 623940 676108 623979
rect 676052 623439 676108 623478
rect 676052 623422 676054 623439
rect 676054 623422 676106 623439
rect 676106 623422 676108 623439
rect 676052 622477 676108 622516
rect 676052 622460 676054 622477
rect 676054 622460 676106 622477
rect 676106 622460 676108 622477
rect 676244 624162 676300 624218
rect 676340 623165 676342 623182
rect 676342 623165 676394 623182
rect 676394 623165 676396 623182
rect 676340 623126 676396 623165
rect 676052 621959 676108 621998
rect 676052 621942 676054 621959
rect 676054 621942 676106 621959
rect 676106 621942 676108 621959
rect 676052 621367 676108 621406
rect 676052 621350 676054 621367
rect 676054 621350 676106 621367
rect 676106 621350 676108 621367
rect 676244 620610 676300 620666
rect 676052 618908 676108 618964
rect 676244 618538 676300 618594
rect 678164 617650 678220 617706
rect 676244 617097 676246 617114
rect 676246 617097 676298 617114
rect 676298 617097 676300 617114
rect 676244 617058 676300 617097
rect 676052 616505 676054 616522
rect 676054 616505 676106 616522
rect 676106 616505 676108 616522
rect 676052 616466 676108 616505
rect 676052 615913 676054 615930
rect 676054 615913 676106 615930
rect 676106 615913 676108 615930
rect 676052 615874 676108 615913
rect 676244 615173 676246 615190
rect 676246 615173 676298 615190
rect 676298 615173 676300 615190
rect 676244 615134 676300 615173
rect 676052 614433 676054 614450
rect 676054 614433 676106 614450
rect 676106 614433 676108 614450
rect 676052 614394 676108 614433
rect 679988 613654 680044 613710
rect 679796 613210 679852 613266
rect 679988 613210 680044 613266
rect 679796 612766 679852 612822
rect 675188 607734 675244 607790
rect 675188 605958 675244 606014
rect 675284 604774 675340 604830
rect 675476 600186 675532 600242
rect 675764 595302 675820 595358
rect 675764 593378 675820 593434
rect 676340 579762 676396 579818
rect 676148 579318 676204 579374
rect 676244 579170 676300 579226
rect 676244 578765 676246 578782
rect 676246 578765 676298 578782
rect 676298 578765 676300 578782
rect 676244 578726 676300 578765
rect 676244 577855 676300 577894
rect 676244 577838 676246 577855
rect 676246 577838 676298 577855
rect 676298 577838 676300 577855
rect 676052 577485 676108 577524
rect 676052 577468 676054 577485
rect 676054 577468 676106 577485
rect 676106 577468 676108 577485
rect 676052 577115 676108 577154
rect 676052 577098 676054 577115
rect 676054 577098 676106 577115
rect 676106 577098 676108 577115
rect 676052 576545 676054 576562
rect 676054 576545 676106 576562
rect 676106 576545 676108 576562
rect 676052 576506 676108 576545
rect 676052 575931 676108 575970
rect 676052 575914 676054 575931
rect 676054 575914 676106 575931
rect 676106 575914 676108 575931
rect 676244 572253 676246 572270
rect 676246 572253 676298 572270
rect 676298 572253 676300 572270
rect 676244 572214 676300 572253
rect 676052 571513 676054 571530
rect 676054 571513 676106 571530
rect 676106 571513 676108 571530
rect 676052 571474 676108 571513
rect 676052 571069 676054 571086
rect 676054 571069 676106 571086
rect 676106 571069 676108 571086
rect 676052 571030 676108 571069
rect 676052 570551 676054 570568
rect 676054 570551 676106 570568
rect 676106 570551 676108 570568
rect 676052 570512 676108 570551
rect 676244 570181 676246 570198
rect 676246 570181 676298 570198
rect 676298 570181 676300 570198
rect 676244 570142 676300 570181
rect 676052 569589 676054 569606
rect 676054 569589 676106 569606
rect 676106 569589 676108 569606
rect 676052 569550 676108 569589
rect 676052 569071 676054 569088
rect 676054 569071 676106 569088
rect 676106 569071 676108 569088
rect 676052 569032 676108 569071
rect 679988 568662 680044 568718
rect 679796 567774 679852 567830
rect 679988 567774 680044 567830
rect 679796 567330 679852 567386
rect 675188 562890 675244 562946
rect 675476 561706 675532 561762
rect 675380 561410 675436 561466
rect 675476 558894 675532 558950
rect 676148 534918 676204 534974
rect 676052 534178 676108 534234
rect 675956 533773 675958 533790
rect 675958 533773 676010 533790
rect 676010 533773 676012 533790
rect 675956 533734 676012 533773
rect 676244 534326 676300 534382
rect 676724 532994 676780 533050
rect 676052 532715 676108 532754
rect 676052 532698 676054 532715
rect 676054 532698 676106 532715
rect 676106 532698 676108 532715
rect 676628 531958 676684 532014
rect 676244 531531 676300 531570
rect 676244 531514 676246 531531
rect 676246 531514 676298 531531
rect 676298 531514 676300 531531
rect 676532 530922 676588 530978
rect 676244 528001 676246 528018
rect 676246 528001 676298 528018
rect 676298 528001 676300 528018
rect 676244 527962 676300 528001
rect 676244 527409 676246 527426
rect 676246 527409 676298 527426
rect 676298 527409 676300 527426
rect 676244 527370 676300 527409
rect 676052 526669 676054 526686
rect 676054 526669 676106 526686
rect 676106 526669 676108 526686
rect 676052 526630 676108 526669
rect 676052 526299 676054 526316
rect 676054 526299 676106 526316
rect 676106 526299 676108 526316
rect 676052 526260 676108 526299
rect 676244 525929 676246 525946
rect 676246 525929 676298 525946
rect 676298 525929 676300 525946
rect 676244 525890 676300 525929
rect 676052 525189 676054 525206
rect 676054 525189 676106 525206
rect 676106 525189 676108 525206
rect 676052 525150 676108 525189
rect 676052 524819 676054 524836
rect 676054 524819 676106 524836
rect 676106 524819 676108 524836
rect 676052 524780 676108 524819
rect 676244 524449 676246 524466
rect 676246 524449 676298 524466
rect 676298 524449 676300 524466
rect 676244 524410 676300 524449
rect 676148 490518 676204 490574
rect 676340 490074 676396 490130
rect 676244 489926 676300 489982
rect 676052 488298 676108 488354
rect 675284 487854 675340 487910
rect 676244 487131 676300 487170
rect 679796 523522 679852 523578
rect 679796 522930 679852 522986
rect 685460 522930 685516 522986
rect 685460 522486 685516 522542
rect 676724 489186 676780 489242
rect 676724 488594 676780 488650
rect 676244 487114 676246 487131
rect 676246 487114 676298 487131
rect 676298 487114 676300 487131
rect 675956 485782 676012 485838
rect 676244 485042 676300 485098
rect 676052 484302 676108 484358
rect 675956 483727 676012 483766
rect 675956 483710 675958 483727
rect 675958 483710 676010 483727
rect 676010 483710 676012 483727
rect 676052 482230 676108 482286
rect 676052 481899 676054 481916
rect 676054 481899 676106 481916
rect 676106 481899 676108 481916
rect 676052 481860 676108 481899
rect 676244 481529 676246 481546
rect 676246 481529 676298 481546
rect 676298 481529 676300 481546
rect 676244 481490 676300 481529
rect 676052 480789 676054 480806
rect 676054 480789 676106 480806
rect 676106 480789 676108 480806
rect 676052 480750 676108 480789
rect 676052 480419 676054 480436
rect 676054 480419 676106 480436
rect 676106 480419 676108 480436
rect 676052 480380 676108 480419
rect 676244 480049 676246 480066
rect 676246 480049 676298 480066
rect 676298 480049 676300 480066
rect 676244 480010 676300 480049
rect 672404 276214 672460 276270
rect 670196 274290 670252 274346
rect 676148 402310 676204 402366
rect 676052 401570 676108 401626
rect 676244 401718 676300 401774
rect 676244 400403 676300 400442
rect 676244 400386 676246 400403
rect 676246 400386 676298 400403
rect 676298 400386 676300 400403
rect 676052 400129 676054 400146
rect 676054 400129 676106 400146
rect 676106 400129 676108 400146
rect 676052 400090 676108 400129
rect 676052 399646 676108 399702
rect 675956 398610 676012 398666
rect 679700 486522 679756 486578
rect 679892 479122 679948 479178
rect 679700 478530 679756 478586
rect 679892 478530 679948 478586
rect 679700 478086 679756 478142
rect 676724 400978 676780 401034
rect 676628 399350 676684 399406
rect 676052 395593 676108 395632
rect 676052 395576 676054 395593
rect 676054 395576 676106 395593
rect 676106 395576 676108 395593
rect 679796 390914 679852 390970
rect 679796 390322 679852 390378
rect 685460 390322 685516 390378
rect 685460 389878 685516 389934
rect 675188 385882 675244 385938
rect 675764 385586 675820 385642
rect 675764 384846 675820 384902
rect 675764 382922 675820 382978
rect 675476 382330 675532 382386
rect 675764 381738 675820 381794
rect 675572 381146 675628 381202
rect 675476 378778 675532 378834
rect 675764 378038 675820 378094
rect 675380 377150 675436 377206
rect 675476 376706 675532 376762
rect 675764 375670 675820 375726
rect 675476 373894 675532 373950
rect 676244 357187 676300 357226
rect 676244 357170 676246 357187
rect 676246 357170 676298 357187
rect 676298 357170 676300 357187
rect 676148 356726 676204 356782
rect 676052 356356 676108 356412
rect 675956 354819 676012 354858
rect 675956 354802 675958 354819
rect 675958 354802 676010 354819
rect 676010 354802 676012 354819
rect 676244 356173 676246 356190
rect 676246 356173 676298 356190
rect 676298 356173 676300 356190
rect 676244 356134 676300 356173
rect 676052 353931 676108 353970
rect 676052 353914 676054 353931
rect 676054 353914 676106 353931
rect 676106 353914 676108 353931
rect 676916 352138 676972 352194
rect 675572 351842 675628 351898
rect 676820 350214 676876 350270
rect 676244 349770 676300 349826
rect 676052 349474 676108 349530
rect 675956 348882 676012 348938
rect 676052 347920 676108 347976
rect 676052 347402 676108 347458
rect 676244 346810 676300 346866
rect 676148 346218 676204 346274
rect 676820 342962 676876 343018
rect 679700 345626 679756 345682
rect 679700 345182 679756 345238
rect 685460 345182 685516 345238
rect 676916 342814 676972 342870
rect 685460 344738 685516 344794
rect 675764 339558 675820 339614
rect 675764 337782 675820 337838
rect 675380 333490 675436 333546
rect 675572 330530 675628 330586
rect 675764 328014 675820 328070
rect 675764 326830 675820 326886
rect 676340 312178 676396 312234
rect 676148 311586 676204 311642
rect 676244 311181 676246 311198
rect 676246 311181 676298 311198
rect 676298 311181 676300 311198
rect 676244 311142 676300 311181
rect 676052 307960 676108 308016
rect 676244 306702 676300 306758
rect 676916 305666 676972 305722
rect 676244 304778 676300 304834
rect 676052 304408 676108 304464
rect 675956 303890 676012 303946
rect 676820 303298 676876 303354
rect 676052 302427 676108 302466
rect 676052 302410 676054 302427
rect 676054 302410 676106 302427
rect 676106 302410 676108 302427
rect 676052 301966 676108 302022
rect 676244 301226 676300 301282
rect 676820 299154 676876 299210
rect 679988 300634 680044 300690
rect 679796 300190 679852 300246
rect 679988 300190 680044 300246
rect 679796 299746 679852 299802
rect 676916 298710 676972 298766
rect 675380 296638 675436 296694
rect 675380 292790 675436 292846
rect 675476 288498 675532 288554
rect 675476 287314 675532 287370
rect 675668 285242 675724 285298
rect 675380 283614 675436 283670
rect 675764 281838 675820 281894
rect 675284 278434 675340 278490
rect 675764 278286 675820 278342
rect 672788 273550 672844 273606
rect 672596 273402 672652 273458
rect 670004 270590 670060 270646
rect 676340 267186 676396 267242
rect 672788 267038 672844 267094
rect 672596 266890 672652 266946
rect 672404 266742 672460 266798
rect 671828 266446 671884 266502
rect 668180 263486 668236 263542
rect 646580 113118 646636 113174
rect 186164 107790 186220 107846
rect 184340 107050 184396 107106
rect 184340 106310 184396 106366
rect 184532 105570 184588 105626
rect 184436 104830 184492 104886
rect 645716 106014 645772 106070
rect 184628 103942 184684 103998
rect 184340 103350 184396 103406
rect 184436 102462 184492 102518
rect 645140 102166 645196 102222
rect 184724 101870 184780 101926
rect 184532 100982 184588 101038
rect 184340 100242 184396 100298
rect 184436 99502 184492 99558
rect 184532 98614 184588 98670
rect 184628 98022 184684 98078
rect 184340 97134 184396 97190
rect 184436 96394 184492 96450
rect 184532 95654 184588 95710
rect 184340 94931 184396 94970
rect 184340 94914 184342 94931
rect 184342 94914 184394 94931
rect 184394 94914 184396 94931
rect 184340 93434 184396 93490
rect 184628 92694 184684 92750
rect 184340 91845 184342 91862
rect 184342 91845 184394 91862
rect 184394 91845 184396 91862
rect 184340 91806 184396 91845
rect 184436 91066 184492 91122
rect 184532 90326 184588 90382
rect 184628 89586 184684 89642
rect 184340 88846 184396 88902
rect 184436 88106 184492 88162
rect 184532 87218 184588 87274
rect 184628 86626 184684 86682
rect 184436 85738 184492 85794
rect 184340 85146 184396 85202
rect 184532 84258 184588 84314
rect 184340 83409 184342 83426
rect 184342 83409 184394 83426
rect 184394 83409 184396 83426
rect 184340 83370 184396 83409
rect 184244 81890 184300 81946
rect 645428 95967 645484 96006
rect 645428 95950 645430 95967
rect 645430 95950 645482 95967
rect 645482 95950 645484 95967
rect 186260 94174 186316 94230
rect 186164 82778 186220 82834
rect 184436 81298 184492 81354
rect 184436 79818 184492 79874
rect 184340 78930 184396 78986
rect 184628 80427 184684 80466
rect 184628 80410 184630 80427
rect 184630 80410 184682 80427
rect 184682 80410 184684 80427
rect 645908 88846 645964 88902
rect 645908 84406 645964 84462
rect 645524 79374 645580 79430
rect 184532 78190 184588 78246
rect 184340 77450 184396 77506
rect 184436 76710 184492 76766
rect 184532 75970 184588 76026
rect 646004 75526 646060 75582
rect 184628 75082 184684 75138
rect 184340 74342 184396 74398
rect 184532 73602 184588 73658
rect 184436 72862 184492 72918
rect 184628 72122 184684 72178
rect 149492 70790 149548 70846
rect 149396 69458 149452 69514
rect 149204 68274 149260 68330
rect 184436 71382 184492 71438
rect 184340 70494 184396 70550
rect 184532 69902 184588 69958
rect 184340 69053 184342 69070
rect 184342 69053 184394 69070
rect 184394 69053 184396 69070
rect 184340 69014 184396 69053
rect 184436 68422 184492 68478
rect 184340 67534 184396 67590
rect 149588 67090 149644 67146
rect 149300 65314 149356 65370
rect 149396 64574 149452 64630
rect 149492 63390 149548 63446
rect 149396 62206 149452 62262
rect 149300 60578 149356 60634
rect 184532 66794 184588 66850
rect 646004 66219 646060 66258
rect 646004 66202 646006 66219
rect 646006 66202 646058 66219
rect 646058 66202 646060 66219
rect 184340 66054 184396 66110
rect 184532 65166 184588 65222
rect 184436 64574 184492 64630
rect 184628 63686 184684 63742
rect 184340 63133 184342 63150
rect 184342 63133 184394 63150
rect 184394 63133 184396 63150
rect 184340 63094 184396 63133
rect 184532 62206 184588 62262
rect 184436 61466 184492 61522
rect 184628 60726 184684 60782
rect 184340 59986 184396 60042
rect 149396 59690 149452 59746
rect 184436 59246 184492 59302
rect 149396 58506 149452 58562
rect 646004 58950 646060 59006
rect 184532 58358 184588 58414
rect 184340 57618 184396 57674
rect 149492 57322 149548 57378
rect 149396 56177 149398 56194
rect 149398 56177 149450 56194
rect 149450 56177 149452 56194
rect 149396 56138 149452 56177
rect 184340 56878 184396 56934
rect 184340 56155 184396 56194
rect 184340 56138 184342 56155
rect 184342 56138 184394 56155
rect 184394 56138 184396 56155
rect 184436 55398 184492 55454
rect 149684 54806 149740 54862
rect 647060 111342 647116 111398
rect 646676 109418 646732 109474
rect 646772 107938 646828 107994
rect 646964 98022 647020 98078
rect 672404 174390 672460 174446
rect 672980 266594 673036 266650
rect 676148 266594 676204 266650
rect 673460 266298 673516 266354
rect 676244 266150 676300 266206
rect 679700 265114 679756 265170
rect 676244 264670 676300 264726
rect 679796 264226 679852 264282
rect 672980 219234 673036 219290
rect 673460 263338 673516 263394
rect 676244 262746 676300 262802
rect 676916 262154 676972 262210
rect 676244 261266 676300 261322
rect 676820 260526 676876 260582
rect 676244 259786 676300 259842
rect 676052 259416 676108 259472
rect 676052 257418 676108 257474
rect 675956 256974 676012 257030
rect 676820 253274 676876 253330
rect 679796 255642 679852 255698
rect 679796 255198 679852 255254
rect 685556 255198 685612 255254
rect 685556 254754 685612 254810
rect 676916 253126 676972 253182
rect 675764 250758 675820 250814
rect 675572 246614 675628 246670
rect 675668 243506 675724 243562
rect 675380 242026 675436 242082
rect 675476 241730 675532 241786
rect 675476 240546 675532 240602
rect 675764 238622 675820 238678
rect 675764 236846 675820 236902
rect 676244 222063 676300 222102
rect 676244 222046 676246 222063
rect 676246 222046 676298 222063
rect 676298 222046 676300 222063
rect 676244 221915 676300 221954
rect 676244 221898 676246 221915
rect 676246 221898 676298 221915
rect 676298 221898 676300 221915
rect 676052 221158 676108 221214
rect 676244 219865 676246 219882
rect 676246 219865 676298 219882
rect 676298 219865 676300 219882
rect 676244 219826 676300 219865
rect 676052 218755 676054 218772
rect 676054 218755 676106 218772
rect 676106 218755 676108 218772
rect 676052 218716 676108 218755
rect 672788 218198 672844 218254
rect 677012 217014 677068 217070
rect 675764 216718 675820 216774
rect 675284 214794 675340 214850
rect 676916 214942 676972 214998
rect 676244 214054 676300 214110
rect 676052 213684 676108 213740
rect 676820 213018 676876 213074
rect 676052 212722 676108 212778
rect 676244 211982 676300 212038
rect 676052 211760 676108 211816
rect 675956 211242 676012 211298
rect 679988 210502 680044 210558
rect 679796 209910 679852 209966
rect 679988 209910 680044 209966
rect 679796 209466 679852 209522
rect 677012 207690 677068 207746
rect 676916 207542 676972 207598
rect 676820 207394 676876 207450
rect 675764 204434 675820 204490
rect 675668 202658 675724 202714
rect 675572 198366 675628 198422
rect 675764 195258 675820 195314
rect 675764 193482 675820 193538
rect 675764 191558 675820 191614
rect 676148 177350 676204 177406
rect 676340 176758 676396 176814
rect 676244 176314 676300 176370
rect 672596 173502 672652 173558
rect 676916 172318 676972 172374
rect 675572 172022 675628 172078
rect 676052 171652 676108 171708
rect 676820 170394 676876 170450
rect 676052 170172 676108 170228
rect 676052 169654 676108 169710
rect 676244 168914 676300 168970
rect 676052 167582 676108 167638
rect 676052 166620 676108 166676
rect 676052 166102 676108 166158
rect 676148 165362 676204 165418
rect 676244 164770 676300 164826
rect 676916 161514 676972 161570
rect 676820 161366 676876 161422
rect 675764 159294 675820 159350
rect 675476 153374 675532 153430
rect 675380 152486 675436 152542
rect 675476 152190 675532 152246
rect 675476 150266 675532 150322
rect 675764 148490 675820 148546
rect 675764 146566 675820 146622
rect 676148 131766 676204 131822
rect 676340 131174 676396 131230
rect 676244 130730 676300 130786
rect 676244 129694 676300 129750
rect 676148 128806 676204 128862
rect 676052 127548 676108 127604
rect 676244 127770 676300 127826
rect 676916 126734 676972 126790
rect 676244 126290 676300 126346
rect 676052 126068 676108 126124
rect 676052 124514 676108 124570
rect 675956 124087 676012 124126
rect 675956 124070 675958 124087
rect 675958 124070 676010 124087
rect 676010 124070 676012 124087
rect 676820 124810 676876 124866
rect 676052 123478 676108 123534
rect 676052 121998 676108 122054
rect 676244 121406 676300 121462
rect 676052 121053 676108 121092
rect 676052 121036 676054 121053
rect 676054 121036 676106 121053
rect 676106 121036 676108 121053
rect 676052 120518 676108 120574
rect 676148 119778 676204 119834
rect 676244 119186 676300 119242
rect 676820 118002 676876 118058
rect 676916 117854 676972 117910
rect 675380 108086 675436 108142
rect 675476 106606 675532 106662
rect 668180 106310 668236 106366
rect 668372 105126 668428 105182
rect 675380 105126 675436 105182
rect 665300 104830 665356 104886
rect 647924 104090 647980 104146
rect 647924 99650 647980 99706
rect 647732 94026 647788 94082
rect 646868 68570 646924 68626
rect 647828 92694 647884 92750
rect 647924 87070 647980 87126
rect 650900 86182 650956 86238
rect 652340 85294 652396 85350
rect 651764 84258 651820 84314
rect 652244 83370 652300 83426
rect 647924 82630 647980 82686
rect 647924 81002 647980 81058
rect 647924 77489 647926 77506
rect 647926 77489 647978 77506
rect 647978 77489 647980 77506
rect 647924 77450 647980 77489
rect 647924 73602 647980 73658
rect 647156 71826 647212 71882
rect 647924 69606 647980 69662
rect 647924 64130 647980 64186
rect 647924 62206 647980 62262
rect 647060 60282 647116 60338
rect 659348 90770 659404 90826
rect 653684 86922 653740 86978
rect 663284 86330 663340 86386
rect 652436 82630 652492 82686
rect 662420 81611 662476 81650
rect 662420 81594 662422 81611
rect 662422 81594 662474 81611
rect 662474 81594 662476 81611
rect 646772 57026 646828 57082
rect 184340 54675 184396 54714
rect 184340 54658 184342 54675
rect 184342 54658 184394 54675
rect 184394 54658 184396 54675
rect 646484 54658 646540 54714
rect 184340 53918 184396 53974
rect 149396 53770 149452 53826
rect 187604 41930 187660 41986
rect 216404 41930 216460 41986
rect 194324 41782 194380 41838
rect 302900 41782 302956 41838
rect 224564 40450 224620 40506
rect 142100 40154 142156 40210
rect 357716 41782 357772 41838
rect 345620 40450 345676 40506
rect 394580 41782 394636 41838
rect 426164 44890 426220 44946
rect 415220 41930 415276 41986
rect 434900 41930 434956 41986
rect 416852 41782 416908 41838
rect 472244 44890 472300 44946
rect 470324 41782 470380 41838
rect 471668 41782 471724 41838
rect 458612 40450 458668 40506
rect 517364 42078 517420 42134
rect 520340 42078 520396 42134
rect 505364 40598 505420 40654
rect 663284 84702 663340 84758
rect 663476 83962 663532 84018
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 675764 103202 675820 103258
rect 675764 101426 675820 101482
rect 545204 40450 545260 40506
rect 311060 37194 311116 37250
rect 324308 37194 324364 37250
<< metal3 >>
rect 82287 1002360 82353 1002363
rect 82272 1002358 82353 1002360
rect 82272 1002302 82292 1002358
rect 82348 1002302 82353 1002358
rect 82272 1002300 82353 1002302
rect 82287 1002297 82353 1002300
rect 483663 1002360 483729 1002363
rect 483663 1002358 483744 1002360
rect 483663 1002302 483668 1002358
rect 483724 1002302 483744 1002358
rect 483663 1002300 483744 1002302
rect 483663 1002297 483729 1002300
rect 132399 997772 132465 997775
rect 184239 997772 184305 997775
rect 535695 997772 535761 997775
rect 639375 997772 639441 997775
rect 132399 997770 133728 997772
rect 132399 997714 132404 997770
rect 132460 997714 133728 997770
rect 132399 997712 133728 997714
rect 184239 997770 184992 997772
rect 184239 997714 184244 997770
rect 184300 997714 184992 997770
rect 535008 997770 535761 997772
rect 184239 997712 184992 997714
rect 132399 997709 132465 997712
rect 184239 997709 184305 997712
rect 241218 997183 241278 997742
rect 241167 997178 241278 997183
rect 241167 997122 241172 997178
rect 241228 997122 241278 997178
rect 241167 997120 241278 997122
rect 293058 997183 293118 997742
rect 400386 997183 400446 997742
rect 535008 997714 535700 997770
rect 535756 997714 535761 997770
rect 535008 997712 535761 997714
rect 636768 997770 639441 997772
rect 636768 997714 639380 997770
rect 639436 997714 639441 997770
rect 636768 997712 639441 997714
rect 535695 997709 535761 997712
rect 639375 997709 639441 997712
rect 293058 997178 293169 997183
rect 293058 997122 293108 997178
rect 293164 997122 293169 997178
rect 293058 997120 293169 997122
rect 241167 997117 241233 997120
rect 293103 997117 293169 997120
rect 400335 997178 400446 997183
rect 400335 997122 400340 997178
rect 400396 997122 400446 997178
rect 400335 997120 400446 997122
rect 400335 997117 400401 997120
rect 389583 983268 389649 983271
rect 389583 983266 389694 983268
rect 389583 983210 389588 983266
rect 389644 983210 389694 983266
rect 389583 983205 389694 983210
rect 80559 982972 80625 982975
rect 132399 982972 132465 982975
rect 184239 982972 184305 982975
rect 233199 982972 233265 982975
rect 240879 982972 240945 982975
rect 80559 982970 81726 982972
rect 80559 982914 80564 982970
rect 80620 982914 81726 982970
rect 80559 982912 81726 982914
rect 80559 982909 80625 982912
rect 81666 982646 81726 982912
rect 132399 982970 133566 982972
rect 132399 982914 132404 982970
rect 132460 982914 133566 982970
rect 132399 982912 133566 982914
rect 132399 982909 132465 982912
rect 133506 982646 133566 982912
rect 184239 982970 185598 982972
rect 184239 982914 184244 982970
rect 184300 982914 185598 982970
rect 184239 982912 185598 982914
rect 184239 982909 184305 982912
rect 185538 982646 185598 982912
rect 233199 982970 236286 982972
rect 233199 982914 233204 982970
rect 233260 982914 236286 982970
rect 233199 982912 236286 982914
rect 233199 982909 233265 982912
rect 236226 982646 236286 982912
rect 240834 982970 240945 982972
rect 240834 982914 240884 982970
rect 240940 982914 240945 982970
rect 240834 982909 240945 982914
rect 241167 982972 241233 982975
rect 285039 982972 285105 982975
rect 292527 982972 292593 982975
rect 293103 982972 293169 982975
rect 241167 982970 241278 982972
rect 241167 982914 241172 982970
rect 241228 982914 241278 982970
rect 241167 982909 241278 982914
rect 285039 982970 288126 982972
rect 285039 982914 285044 982970
rect 285100 982914 288126 982970
rect 285039 982912 288126 982914
rect 285039 982909 285105 982912
rect 240834 982646 240894 982909
rect 241218 982646 241278 982909
rect 288066 982646 288126 982912
rect 292482 982970 292593 982972
rect 292482 982914 292532 982970
rect 292588 982914 292593 982970
rect 292482 982909 292593 982914
rect 293058 982970 293169 982972
rect 293058 982914 293108 982970
rect 293164 982914 293169 982970
rect 293058 982909 293169 982914
rect 292482 982646 292542 982909
rect 293058 982646 293118 982909
rect 389634 982646 389694 983205
rect 394575 982972 394641 982975
rect 400335 982972 400401 982975
rect 486735 982972 486801 982975
rect 538575 982972 538641 982975
rect 639375 982972 639441 982975
rect 394242 982970 394641 982972
rect 394242 982914 394580 982970
rect 394636 982914 394641 982970
rect 394242 982912 394641 982914
rect 394242 982646 394302 982912
rect 394575 982909 394641 982912
rect 399426 982970 400401 982972
rect 399426 982914 400340 982970
rect 400396 982914 400401 982970
rect 399426 982912 400401 982914
rect 399426 982646 399486 982912
rect 400335 982909 400401 982912
rect 483522 982970 486801 982972
rect 483522 982914 486740 982970
rect 486796 982914 486801 982970
rect 483522 982912 486801 982914
rect 483522 982646 483582 982912
rect 486735 982909 486801 982912
rect 535554 982970 538641 982972
rect 535554 982914 538580 982970
rect 538636 982914 538641 982970
rect 535554 982912 538641 982914
rect 535554 982646 535614 982912
rect 538575 982909 538641 982912
rect 636738 982970 639441 982972
rect 636738 982914 639380 982970
rect 639436 982914 639441 982970
rect 636738 982912 639441 982914
rect 636738 982646 636798 982912
rect 639375 982909 639441 982912
rect 40143 961956 40209 961959
rect 39840 961954 40209 961956
rect 39840 961898 40148 961954
rect 40204 961898 40209 961954
rect 39840 961896 40209 961898
rect 40143 961893 40209 961896
rect 60015 961808 60081 961811
rect 60015 961806 65376 961808
rect 60015 961750 60020 961806
rect 60076 961750 65376 961806
rect 60015 961748 65376 961750
rect 60015 961745 60081 961748
rect 653775 960476 653841 960479
rect 649248 960474 653841 960476
rect 649248 960418 653780 960474
rect 653836 960418 653841 960474
rect 649248 960416 653841 960418
rect 653775 960413 653841 960416
rect 679746 958555 679806 958670
rect 679695 958550 679806 958555
rect 679695 958494 679700 958550
rect 679756 958494 679806 958550
rect 679695 958492 679806 958494
rect 679695 958489 679761 958492
rect 676143 894172 676209 894175
rect 676290 894172 676350 894438
rect 676143 894170 676350 894172
rect 676143 894114 676148 894170
rect 676204 894114 676350 894170
rect 676143 894112 676350 894114
rect 676143 894109 676209 894112
rect 676290 893583 676350 893920
rect 676239 893578 676350 893583
rect 676239 893522 676244 893578
rect 676300 893522 676350 893578
rect 676239 893520 676350 893522
rect 676239 893517 676305 893520
rect 676047 893432 676113 893435
rect 676047 893430 676320 893432
rect 676047 893374 676052 893430
rect 676108 893374 676320 893430
rect 676047 893372 676320 893374
rect 676047 893369 676113 893372
rect 676047 892470 676113 892473
rect 676047 892468 676320 892470
rect 676047 892412 676052 892468
rect 676108 892412 676320 892468
rect 676047 892410 676320 892412
rect 676047 892407 676113 892410
rect 676047 891508 676113 891511
rect 676047 891506 676320 891508
rect 676047 891450 676052 891506
rect 676108 891450 676320 891506
rect 676047 891448 676320 891450
rect 676047 891445 676113 891448
rect 676047 890472 676113 890475
rect 676047 890470 676320 890472
rect 676047 890414 676052 890470
rect 676108 890414 676320 890470
rect 676047 890412 676320 890414
rect 676047 890409 676113 890412
rect 680271 890176 680337 890179
rect 680271 890174 680382 890176
rect 680271 890118 680276 890174
rect 680332 890118 680382 890174
rect 680271 890113 680382 890118
rect 680322 889998 680382 890113
rect 676290 889291 676350 889406
rect 676239 889286 676350 889291
rect 676239 889230 676244 889286
rect 676300 889230 676350 889286
rect 676239 889228 676350 889230
rect 676239 889225 676305 889228
rect 680130 888699 680190 888888
rect 680079 888694 680190 888699
rect 680079 888638 680084 888694
rect 680140 888638 680190 888694
rect 680079 888636 680190 888638
rect 680079 888633 680145 888636
rect 680130 888255 680190 888518
rect 680130 888250 680241 888255
rect 680130 888194 680180 888250
rect 680236 888194 680241 888250
rect 680130 888192 680241 888194
rect 680175 888189 680241 888192
rect 676047 887956 676113 887959
rect 676047 887954 676320 887956
rect 676047 887898 676052 887954
rect 676108 887898 676320 887954
rect 676047 887896 676320 887898
rect 676047 887893 676113 887896
rect 676047 887438 676113 887441
rect 676047 887436 676320 887438
rect 676047 887380 676052 887436
rect 676108 887380 676320 887436
rect 676047 887378 676320 887380
rect 676047 887375 676113 887378
rect 679746 886775 679806 887038
rect 679695 886770 679806 886775
rect 679695 886714 679700 886770
rect 679756 886714 679806 886770
rect 679695 886712 679806 886714
rect 679695 886709 679761 886712
rect 679938 886183 679998 886446
rect 679887 886178 679998 886183
rect 679887 886122 679892 886178
rect 679948 886122 679998 886178
rect 679887 886120 679998 886122
rect 679887 886117 679953 886120
rect 679938 885739 679998 885854
rect 679938 885734 680049 885739
rect 679938 885678 679988 885734
rect 680044 885678 680049 885734
rect 679938 885676 680049 885678
rect 679983 885673 680049 885676
rect 676047 885514 676113 885517
rect 676047 885512 676320 885514
rect 676047 885456 676052 885512
rect 676108 885456 676320 885512
rect 676047 885454 676320 885456
rect 676047 885451 676113 885454
rect 676047 884996 676113 884999
rect 676047 884994 676320 884996
rect 676047 884938 676052 884994
rect 676108 884938 676320 884994
rect 676047 884936 676320 884938
rect 676047 884933 676113 884936
rect 676290 884259 676350 884374
rect 676239 884254 676350 884259
rect 676239 884198 676244 884254
rect 676300 884198 676350 884254
rect 676239 884196 676350 884198
rect 676239 884193 676305 884196
rect 676047 884034 676113 884037
rect 676047 884032 676320 884034
rect 676047 883976 676052 884032
rect 676108 883976 676320 884032
rect 676047 883974 676320 883976
rect 676047 883971 676113 883974
rect 676047 883516 676113 883519
rect 676047 883514 676320 883516
rect 676047 883458 676052 883514
rect 676108 883458 676320 883514
rect 676047 883456 676320 883458
rect 676047 883453 676113 883456
rect 679746 882779 679806 882894
rect 679746 882774 679857 882779
rect 679746 882718 679796 882774
rect 679852 882718 679857 882774
rect 679746 882716 679857 882718
rect 679791 882713 679857 882716
rect 685506 882187 685566 882450
rect 679791 882184 679857 882187
rect 679746 882182 679857 882184
rect 679746 882126 679796 882182
rect 679852 882126 679857 882182
rect 679746 882121 679857 882126
rect 685455 882182 685566 882187
rect 685455 882126 685460 882182
rect 685516 882126 685566 882182
rect 685455 882124 685566 882126
rect 685455 882121 685521 882124
rect 679746 882006 679806 882121
rect 685455 881740 685521 881743
rect 685455 881738 685566 881740
rect 685455 881682 685460 881738
rect 685516 881682 685566 881738
rect 685455 881677 685566 881682
rect 685506 881414 685566 881677
rect 655407 868864 655473 868867
rect 649986 868862 655473 868864
rect 649986 868806 655412 868862
rect 655468 868806 655473 868862
rect 649986 868804 655473 868806
rect 649986 868246 650046 868804
rect 655407 868801 655473 868804
rect 655215 867680 655281 867683
rect 649986 867678 655281 867680
rect 649986 867622 655220 867678
rect 655276 867622 655281 867678
rect 649986 867620 655281 867622
rect 649986 867064 650046 867620
rect 655215 867617 655281 867620
rect 655119 866496 655185 866499
rect 649986 866494 655185 866496
rect 649986 866438 655124 866494
rect 655180 866438 655185 866494
rect 649986 866436 655185 866438
rect 649986 865882 650046 866436
rect 655119 866433 655185 866436
rect 655311 865312 655377 865315
rect 649986 865310 655377 865312
rect 649986 865254 655316 865310
rect 655372 865254 655377 865310
rect 649986 865252 655377 865254
rect 649986 864700 650046 865252
rect 655311 865249 655377 865252
rect 654159 863980 654225 863983
rect 649986 863978 654225 863980
rect 649986 863922 654164 863978
rect 654220 863922 654225 863978
rect 649986 863920 654225 863922
rect 649986 863518 650046 863920
rect 654159 863917 654225 863920
rect 653775 862944 653841 862947
rect 649986 862942 653841 862944
rect 649986 862886 653780 862942
rect 653836 862886 653841 862942
rect 649986 862884 653841 862886
rect 649986 862336 650046 862884
rect 653775 862881 653841 862884
rect 41775 816694 41841 816697
rect 41568 816692 41841 816694
rect 41568 816636 41780 816692
rect 41836 816636 41841 816692
rect 41568 816634 41841 816636
rect 41775 816631 41841 816634
rect 41775 816176 41841 816179
rect 41568 816174 41841 816176
rect 41568 816118 41780 816174
rect 41836 816118 41841 816174
rect 41568 816116 41841 816118
rect 41775 816113 41841 816116
rect 41538 815439 41598 815554
rect 41538 815434 41649 815439
rect 41538 815378 41588 815434
rect 41644 815378 41649 815434
rect 41538 815376 41649 815378
rect 41583 815373 41649 815376
rect 41775 814696 41841 814699
rect 41568 814694 41841 814696
rect 41568 814638 41780 814694
rect 41836 814638 41841 814694
rect 41568 814636 41841 814638
rect 41775 814633 41841 814636
rect 40386 813958 40446 814074
rect 40378 813894 40384 813958
rect 40448 813894 40454 813958
rect 41538 813515 41598 813630
rect 41538 813510 41649 813515
rect 41538 813454 41588 813510
rect 41644 813454 41649 813510
rect 41538 813452 41649 813454
rect 41583 813449 41649 813452
rect 40578 812774 40638 813186
rect 40570 812710 40576 812774
rect 40640 812710 40646 812774
rect 41775 812624 41841 812627
rect 41568 812622 41841 812624
rect 41568 812566 41780 812622
rect 41836 812566 41841 812622
rect 41568 812564 41841 812566
rect 41775 812561 41841 812564
rect 41346 812035 41406 812150
rect 41346 812030 41457 812035
rect 41346 811974 41396 812030
rect 41452 811974 41457 812030
rect 41346 811972 41457 811974
rect 41391 811969 41457 811972
rect 41967 811662 42033 811665
rect 41568 811660 42033 811662
rect 41568 811604 41972 811660
rect 42028 811604 42033 811660
rect 41568 811602 42033 811604
rect 41967 811599 42033 811602
rect 40239 811292 40305 811295
rect 40194 811290 40305 811292
rect 40194 811234 40244 811290
rect 40300 811234 40305 811290
rect 40194 811229 40305 811234
rect 40194 811114 40254 811229
rect 41538 810555 41598 810670
rect 41538 810550 41649 810555
rect 41538 810494 41588 810550
rect 41644 810494 41649 810550
rect 41538 810492 41649 810494
rect 41583 810489 41649 810492
rect 41538 809960 41598 810152
rect 41679 809960 41745 809963
rect 41538 809958 41745 809960
rect 41538 809902 41684 809958
rect 41740 809902 41745 809958
rect 41538 809900 41745 809902
rect 41679 809897 41745 809900
rect 41871 809664 41937 809667
rect 41568 809662 41937 809664
rect 41568 809606 41876 809662
rect 41932 809606 41937 809662
rect 41568 809604 41937 809606
rect 41871 809601 41937 809604
rect 41538 808926 41598 809190
rect 41530 808862 41536 808926
rect 41600 808862 41606 808926
rect 41538 808483 41598 808598
rect 41538 808478 41649 808483
rect 41538 808422 41588 808478
rect 41644 808422 41649 808478
rect 41538 808420 41649 808422
rect 41583 808417 41649 808420
rect 42159 808184 42225 808187
rect 41568 808182 42225 808184
rect 41568 808126 42164 808182
rect 42220 808126 42225 808182
rect 41568 808124 42225 808126
rect 42159 808121 42225 808124
rect 41775 807740 41841 807743
rect 41568 807738 41841 807740
rect 41568 807682 41780 807738
rect 41836 807682 41841 807738
rect 41568 807680 41841 807682
rect 41775 807677 41841 807680
rect 41538 807003 41598 807118
rect 41538 806998 41649 807003
rect 41538 806942 41588 806998
rect 41644 806942 41649 806998
rect 41538 806940 41649 806942
rect 41583 806937 41649 806940
rect 42063 806630 42129 806633
rect 41568 806628 42129 806630
rect 41568 806572 42068 806628
rect 42124 806572 42129 806628
rect 41568 806570 42129 806572
rect 42063 806567 42129 806570
rect 41775 806260 41841 806263
rect 41568 806258 41841 806260
rect 41568 806202 41780 806258
rect 41836 806202 41841 806258
rect 41568 806200 41841 806202
rect 41775 806197 41841 806200
rect 41538 805523 41598 805638
rect 41538 805518 41649 805523
rect 41538 805462 41588 805518
rect 41644 805462 41649 805518
rect 41538 805460 41649 805462
rect 41583 805457 41649 805460
rect 41538 804928 41598 805120
rect 41538 804868 41790 804928
rect 28866 804487 28926 804750
rect 28815 804482 28926 804487
rect 41730 804484 41790 804868
rect 28815 804426 28820 804482
rect 28876 804426 28926 804482
rect 28815 804424 28926 804426
rect 41538 804424 41790 804484
rect 28815 804421 28881 804424
rect 41538 803895 41598 804424
rect 28815 803892 28881 803895
rect 28815 803890 28926 803892
rect 28815 803834 28820 803890
rect 28876 803834 28926 803890
rect 28815 803829 28926 803834
rect 41487 803890 41598 803895
rect 41487 803834 41492 803890
rect 41548 803834 41598 803890
rect 41487 803832 41598 803834
rect 41487 803829 41553 803832
rect 28866 803566 28926 803829
rect 40239 801376 40305 801379
rect 41146 801376 41152 801378
rect 40239 801374 41152 801376
rect 40239 801318 40244 801374
rect 40300 801318 41152 801374
rect 40239 801316 41152 801318
rect 40239 801313 40305 801316
rect 41146 801314 41152 801316
rect 41216 801314 41222 801378
rect 41679 800490 41745 800491
rect 41679 800488 41728 800490
rect 41636 800486 41728 800488
rect 41636 800430 41684 800486
rect 41636 800428 41728 800430
rect 41679 800426 41728 800428
rect 41792 800426 41798 800490
rect 41679 800425 41745 800426
rect 41967 800342 42033 800343
rect 41914 800278 41920 800342
rect 41984 800340 42033 800342
rect 42159 800340 42225 800343
rect 42298 800340 42304 800342
rect 41984 800338 42076 800340
rect 42028 800282 42076 800338
rect 41984 800280 42076 800282
rect 42159 800338 42304 800340
rect 42159 800282 42164 800338
rect 42220 800282 42304 800338
rect 42159 800280 42304 800282
rect 41984 800278 42033 800280
rect 41967 800277 42033 800278
rect 42159 800277 42225 800280
rect 42298 800278 42304 800280
rect 42368 800278 42374 800342
rect 41967 798122 42033 798123
rect 41914 798120 41920 798122
rect 41876 798060 41920 798120
rect 41984 798118 42033 798122
rect 42028 798062 42033 798118
rect 41914 798058 41920 798060
rect 41984 798058 42033 798062
rect 41967 798057 42033 798058
rect 42298 795394 42304 795458
rect 42368 795456 42374 795458
rect 42831 795456 42897 795459
rect 42368 795454 42897 795456
rect 42368 795398 42836 795454
rect 42892 795398 42897 795454
rect 42368 795396 42897 795398
rect 42368 795394 42374 795396
rect 42831 795393 42897 795396
rect 41775 792942 41841 792943
rect 41722 792940 41728 792942
rect 41684 792880 41728 792940
rect 41792 792938 41841 792942
rect 41836 792882 41841 792938
rect 41722 792878 41728 792880
rect 41792 792878 41841 792882
rect 41775 792877 41841 792878
rect 41530 791842 41536 791906
rect 41600 791904 41606 791906
rect 42831 791904 42897 791907
rect 41600 791902 42897 791904
rect 41600 791846 42836 791902
rect 42892 791846 42897 791902
rect 41600 791844 42897 791846
rect 41600 791842 41606 791844
rect 42831 791841 42897 791844
rect 41146 791694 41152 791758
rect 41216 791756 41222 791758
rect 42927 791756 42993 791759
rect 41216 791754 42993 791756
rect 41216 791698 42932 791754
rect 42988 791698 42993 791754
rect 41216 791696 42993 791698
rect 41216 791694 41222 791696
rect 42927 791693 42993 791696
rect 57711 790868 57777 790871
rect 57711 790866 64638 790868
rect 57711 790810 57716 790866
rect 57772 790810 64638 790866
rect 57711 790808 64638 790810
rect 57711 790805 57777 790808
rect 64578 790304 64638 790808
rect 57615 789684 57681 789687
rect 57615 789682 64638 789684
rect 57615 789626 57620 789682
rect 57676 789626 64638 789682
rect 57615 789624 64638 789626
rect 57615 789621 57681 789624
rect 64578 789122 64638 789624
rect 58191 788500 58257 788503
rect 58191 788498 64638 788500
rect 58191 788442 58196 788498
rect 58252 788442 64638 788498
rect 58191 788440 64638 788442
rect 58191 788437 58257 788440
rect 64578 787940 64638 788440
rect 675130 787994 675136 788058
rect 675200 788056 675206 788058
rect 675375 788056 675441 788059
rect 675200 788054 675441 788056
rect 675200 787998 675380 788054
rect 675436 787998 675441 788054
rect 675200 787996 675441 787998
rect 675200 787994 675206 787996
rect 675375 787993 675441 787996
rect 58383 787316 58449 787319
rect 58383 787314 64638 787316
rect 58383 787258 58388 787314
rect 58444 787258 64638 787314
rect 58383 787256 64638 787258
rect 58383 787253 58449 787256
rect 64578 786758 64638 787256
rect 675663 787170 675729 787171
rect 675663 787166 675712 787170
rect 675776 787168 675782 787170
rect 675663 787110 675668 787166
rect 675663 787106 675712 787110
rect 675776 787108 675820 787168
rect 675776 787106 675782 787108
rect 675663 787105 675729 787106
rect 674170 786662 674176 786726
rect 674240 786724 674246 786726
rect 675375 786724 675441 786727
rect 674240 786722 675441 786724
rect 674240 786666 675380 786722
rect 675436 786666 675441 786722
rect 674240 786664 675441 786666
rect 674240 786662 674246 786664
rect 675375 786661 675441 786664
rect 59631 785540 59697 785543
rect 64578 785540 64638 785576
rect 59631 785538 64638 785540
rect 59631 785482 59636 785538
rect 59692 785482 64638 785538
rect 59631 785480 64638 785482
rect 59631 785477 59697 785480
rect 59151 784948 59217 784951
rect 59151 784946 64638 784948
rect 59151 784890 59156 784946
rect 59212 784890 64638 784946
rect 59151 784888 64638 784890
rect 59151 784885 59217 784888
rect 64578 784394 64638 784888
rect 675375 784802 675441 784803
rect 675322 784800 675328 784802
rect 675284 784740 675328 784800
rect 675392 784798 675441 784802
rect 675436 784742 675441 784798
rect 675322 784738 675328 784740
rect 675392 784738 675441 784742
rect 675375 784737 675441 784738
rect 675759 784208 675825 784211
rect 676090 784208 676096 784210
rect 675759 784206 676096 784208
rect 675759 784150 675764 784206
rect 675820 784150 676096 784206
rect 675759 784148 676096 784150
rect 675759 784145 675825 784148
rect 676090 784146 676096 784148
rect 676160 784146 676166 784210
rect 673978 783406 673984 783470
rect 674048 783468 674054 783470
rect 675279 783468 675345 783471
rect 674048 783466 675345 783468
rect 674048 783410 675284 783466
rect 675340 783410 675345 783466
rect 674048 783408 675345 783410
rect 674048 783406 674054 783408
rect 675279 783405 675345 783408
rect 675471 780658 675537 780659
rect 675471 780654 675520 780658
rect 675584 780656 675590 780658
rect 675471 780598 675476 780654
rect 675471 780594 675520 780598
rect 675584 780596 675628 780656
rect 675584 780594 675590 780596
rect 675471 780593 675537 780594
rect 675759 779916 675825 779919
rect 676282 779916 676288 779918
rect 675759 779914 676288 779916
rect 675759 779858 675764 779914
rect 675820 779858 676288 779914
rect 675759 779856 676288 779858
rect 675759 779853 675825 779856
rect 676282 779854 676288 779856
rect 676352 779854 676358 779918
rect 675759 779176 675825 779179
rect 676474 779176 676480 779178
rect 675759 779174 676480 779176
rect 675759 779118 675764 779174
rect 675820 779118 676480 779174
rect 675759 779116 676480 779118
rect 675759 779113 675825 779116
rect 676474 779114 676480 779116
rect 676544 779114 676550 779178
rect 649986 778288 650046 778824
rect 655407 778288 655473 778291
rect 649986 778286 655473 778288
rect 649986 778230 655412 778286
rect 655468 778230 655473 778286
rect 649986 778228 655473 778230
rect 655407 778225 655473 778228
rect 655119 777696 655185 777699
rect 649986 777694 655185 777696
rect 649986 777638 655124 777694
rect 655180 777638 655185 777694
rect 649986 777636 655185 777638
rect 655119 777633 655185 777636
rect 675759 777696 675825 777699
rect 676666 777696 676672 777698
rect 675759 777694 676672 777696
rect 675759 777638 675764 777694
rect 675820 777638 676672 777694
rect 675759 777636 676672 777638
rect 675759 777633 675825 777636
rect 676666 777634 676672 777636
rect 676736 777634 676742 777698
rect 649986 775920 650046 776460
rect 655599 775920 655665 775923
rect 649986 775918 655665 775920
rect 649986 775862 655604 775918
rect 655660 775862 655665 775918
rect 649986 775860 655665 775862
rect 655599 775857 655665 775860
rect 655215 775772 655281 775775
rect 649986 775770 655281 775772
rect 649986 775714 655220 775770
rect 655276 775714 655281 775770
rect 649986 775712 655281 775714
rect 649986 775278 650046 775712
rect 655215 775709 655281 775712
rect 675759 775476 675825 775479
rect 675898 775476 675904 775478
rect 675759 775474 675904 775476
rect 675759 775418 675764 775474
rect 675820 775418 675904 775474
rect 675759 775416 675904 775418
rect 675759 775413 675825 775416
rect 675898 775414 675904 775416
rect 675968 775414 675974 775478
rect 655023 774736 655089 774739
rect 649986 774734 655089 774736
rect 649986 774678 655028 774734
rect 655084 774678 655089 774734
rect 649986 774676 655089 774678
rect 40378 774526 40384 774590
rect 40448 774588 40454 774590
rect 41583 774588 41649 774591
rect 40448 774586 41649 774588
rect 40448 774530 41588 774586
rect 41644 774530 41649 774586
rect 40448 774528 41649 774530
rect 40448 774526 40454 774528
rect 41583 774525 41649 774528
rect 649986 774096 650046 774676
rect 655023 774673 655089 774676
rect 40570 773934 40576 773998
rect 40640 773996 40646 773998
rect 41487 773996 41553 773999
rect 40640 773994 41553 773996
rect 40640 773938 41492 773994
rect 41548 773938 41553 773994
rect 40640 773936 41553 773938
rect 40640 773934 40646 773936
rect 41487 773933 41553 773936
rect 41775 773552 41841 773555
rect 654351 773552 654417 773555
rect 41568 773550 41841 773552
rect 41568 773494 41780 773550
rect 41836 773494 41841 773550
rect 41568 773492 41841 773494
rect 41775 773489 41841 773492
rect 649986 773550 654417 773552
rect 649986 773494 654356 773550
rect 654412 773494 654417 773550
rect 649986 773492 654417 773494
rect 41775 772960 41841 772963
rect 41568 772958 41841 772960
rect 41568 772902 41780 772958
rect 41836 772902 41841 772958
rect 649986 772914 650046 773492
rect 654351 773489 654417 773492
rect 41568 772900 41841 772902
rect 41775 772897 41841 772900
rect 41775 772368 41841 772371
rect 41568 772366 41841 772368
rect 41568 772310 41780 772366
rect 41836 772310 41841 772366
rect 41568 772308 41841 772310
rect 41775 772305 41841 772308
rect 41775 771998 41841 772001
rect 41568 771996 41841 771998
rect 41568 771940 41780 771996
rect 41836 771940 41841 771996
rect 41568 771938 41841 771940
rect 41775 771935 41841 771938
rect 674991 771924 675057 771927
rect 675706 771924 675712 771926
rect 674991 771922 675712 771924
rect 674991 771866 674996 771922
rect 675052 771866 675712 771922
rect 674991 771864 675712 771866
rect 674991 771861 675057 771864
rect 675706 771862 675712 771864
rect 675776 771862 675782 771926
rect 41775 771480 41841 771483
rect 41568 771478 41841 771480
rect 41568 771422 41780 771478
rect 41836 771422 41841 771478
rect 41568 771420 41841 771422
rect 41775 771417 41841 771420
rect 40386 770742 40446 770858
rect 40378 770678 40384 770742
rect 40448 770678 40454 770742
rect 41583 770740 41649 770743
rect 41538 770738 41649 770740
rect 41538 770682 41588 770738
rect 41644 770682 41649 770738
rect 41538 770677 41649 770682
rect 41538 770488 41598 770677
rect 40578 769706 40638 769970
rect 40570 769642 40576 769706
rect 40640 769642 40646 769706
rect 41487 769704 41553 769707
rect 41487 769702 41598 769704
rect 41487 769646 41492 769702
rect 41548 769646 41598 769702
rect 41487 769641 41598 769646
rect 41538 769378 41598 769641
rect 41538 768819 41598 768934
rect 41538 768814 41649 768819
rect 41538 768758 41588 768814
rect 41644 768758 41649 768814
rect 41538 768756 41649 768758
rect 41583 768753 41649 768756
rect 41538 768224 41598 768490
rect 41679 768224 41745 768227
rect 41538 768222 41745 768224
rect 41538 768166 41684 768222
rect 41740 768166 41745 768222
rect 41538 768164 41745 768166
rect 41679 768161 41745 768164
rect 38799 768076 38865 768079
rect 38799 768074 38910 768076
rect 38799 768018 38804 768074
rect 38860 768018 38910 768074
rect 38799 768013 38910 768018
rect 38850 767898 38910 768013
rect 41538 767339 41598 767454
rect 41538 767334 41649 767339
rect 41538 767278 41588 767334
rect 41644 767278 41649 767334
rect 41538 767276 41649 767278
rect 41583 767273 41649 767276
rect 41967 766966 42033 766969
rect 41568 766964 42033 766966
rect 41568 766908 41972 766964
rect 42028 766908 42033 766964
rect 41568 766906 42033 766908
rect 41967 766903 42033 766906
rect 40335 766596 40401 766599
rect 40335 766594 40446 766596
rect 40335 766538 40340 766594
rect 40396 766538 40446 766594
rect 40335 766533 40446 766538
rect 40386 766418 40446 766533
rect 34434 765859 34494 765974
rect 34434 765854 34545 765859
rect 34434 765798 34484 765854
rect 34540 765798 34545 765854
rect 34434 765796 34545 765798
rect 34479 765793 34545 765796
rect 41775 765486 41841 765489
rect 41568 765484 41841 765486
rect 41568 765428 41780 765484
rect 41836 765428 41841 765484
rect 41568 765426 41841 765428
rect 41775 765423 41841 765426
rect 41295 765116 41361 765119
rect 41295 765114 41406 765116
rect 41295 765058 41300 765114
rect 41356 765058 41406 765114
rect 41295 765053 41406 765058
rect 41346 764938 41406 765053
rect 41871 764524 41937 764527
rect 41568 764522 41937 764524
rect 41568 764466 41876 764522
rect 41932 764466 41937 764522
rect 41568 764464 41937 764466
rect 41871 764461 41937 764464
rect 42063 763932 42129 763935
rect 41568 763930 42129 763932
rect 41568 763874 42068 763930
rect 42124 763874 42129 763930
rect 41568 763872 42129 763874
rect 42063 763869 42129 763872
rect 41775 763488 41841 763491
rect 41568 763486 41841 763488
rect 41568 763430 41780 763486
rect 41836 763430 41841 763486
rect 41568 763428 41841 763430
rect 41775 763425 41841 763428
rect 42159 763044 42225 763047
rect 41568 763042 42225 763044
rect 41568 762986 42164 763042
rect 42220 762986 42225 763042
rect 41568 762984 42225 762986
rect 42159 762981 42225 762984
rect 41775 762452 41841 762455
rect 41568 762450 41841 762452
rect 41568 762394 41780 762450
rect 41836 762394 41841 762450
rect 41568 762392 41841 762394
rect 41775 762389 41841 762392
rect 41538 761715 41598 761904
rect 41538 761710 41649 761715
rect 41538 761654 41588 761710
rect 41644 761654 41649 761710
rect 41538 761652 41649 761654
rect 41583 761649 41649 761652
rect 28866 761271 28926 761534
rect 28815 761266 28926 761271
rect 28815 761210 28820 761266
rect 28876 761210 28926 761266
rect 28815 761208 28926 761210
rect 28815 761205 28881 761208
rect 41538 760827 41598 760942
rect 28815 760824 28881 760827
rect 28815 760822 28926 760824
rect 28815 760766 28820 760822
rect 28876 760766 28926 760822
rect 28815 760761 28926 760766
rect 41538 760822 41649 760827
rect 41538 760766 41588 760822
rect 41644 760766 41649 760822
rect 41538 760764 41649 760766
rect 41583 760761 41649 760764
rect 28866 760424 28926 760761
rect 34479 758900 34545 758903
rect 40762 758900 40768 758902
rect 34479 758898 40768 758900
rect 34479 758842 34484 758898
rect 34540 758842 40768 758898
rect 34479 758840 40768 758842
rect 34479 758837 34545 758840
rect 40762 758838 40768 758840
rect 40832 758838 40838 758902
rect 43023 758014 43089 758015
rect 43023 758010 43072 758014
rect 43136 758012 43142 758014
rect 43023 757954 43028 758010
rect 43023 757950 43072 757954
rect 43136 757952 43180 758012
rect 43136 757950 43142 757952
rect 43023 757949 43089 757950
rect 38799 757568 38865 757571
rect 40954 757568 40960 757570
rect 38799 757566 40960 757568
rect 38799 757510 38804 757566
rect 38860 757510 40960 757566
rect 38799 757508 40960 757510
rect 38799 757505 38865 757508
rect 40954 757506 40960 757508
rect 41024 757506 41030 757570
rect 42874 757210 42880 757274
rect 42944 757272 42950 757274
rect 43119 757272 43185 757275
rect 42944 757270 43185 757272
rect 42944 757214 43124 757270
rect 43180 757214 43185 757270
rect 42944 757212 43185 757214
rect 42944 757210 42950 757212
rect 43119 757209 43185 757212
rect 41967 757124 42033 757127
rect 42106 757124 42112 757126
rect 41967 757122 42112 757124
rect 41967 757066 41972 757122
rect 42028 757066 42112 757122
rect 41967 757064 42112 757066
rect 41967 757061 42033 757064
rect 42106 757062 42112 757064
rect 42176 757062 42182 757126
rect 42106 754694 42112 754758
rect 42176 754756 42182 754758
rect 42735 754756 42801 754759
rect 42176 754754 42801 754756
rect 42176 754698 42740 754754
rect 42796 754698 42801 754754
rect 42176 754696 42801 754698
rect 42176 754694 42182 754696
rect 42735 754693 42801 754696
rect 42874 751586 42880 751650
rect 42944 751648 42950 751650
rect 43023 751648 43089 751651
rect 42944 751646 43089 751648
rect 42944 751590 43028 751646
rect 43084 751590 43089 751646
rect 42944 751588 43089 751590
rect 42944 751586 42950 751588
rect 43023 751585 43089 751588
rect 42831 750464 42897 750467
rect 43066 750464 43072 750466
rect 42831 750462 43072 750464
rect 42831 750406 42836 750462
rect 42892 750406 43072 750462
rect 42831 750404 43072 750406
rect 42831 750401 42897 750404
rect 43066 750402 43072 750404
rect 43136 750402 43142 750466
rect 58671 747652 58737 747655
rect 58671 747650 64638 747652
rect 58671 747594 58676 747650
rect 58732 747594 64638 747650
rect 58671 747592 64638 747594
rect 58671 747589 58737 747592
rect 40762 747146 40768 747210
rect 40832 747208 40838 747210
rect 42831 747208 42897 747211
rect 40832 747206 42897 747208
rect 40832 747150 42836 747206
rect 42892 747150 42897 747206
rect 40832 747148 42897 747150
rect 40832 747146 40838 747148
rect 42831 747145 42897 747148
rect 64578 747082 64638 747592
rect 40954 746850 40960 746914
rect 41024 746912 41030 746914
rect 42735 746912 42801 746915
rect 41024 746910 42801 746912
rect 41024 746854 42740 746910
rect 42796 746854 42801 746910
rect 41024 746852 42801 746854
rect 41024 746850 41030 746852
rect 42735 746849 42801 746852
rect 54735 746024 54801 746027
rect 54690 746022 54801 746024
rect 54690 745966 54740 746022
rect 54796 745966 54801 746022
rect 54690 745961 54801 745966
rect 54690 745879 54750 745961
rect 54639 745874 54750 745879
rect 54639 745818 54644 745874
rect 54700 745818 54750 745874
rect 54639 745816 54750 745818
rect 54639 745813 54705 745816
rect 59631 745728 59697 745731
rect 64578 745728 64638 745900
rect 676282 745814 676288 745878
rect 676352 745876 676358 745878
rect 677434 745876 677440 745878
rect 676352 745816 677440 745876
rect 676352 745814 676358 745816
rect 677434 745814 677440 745816
rect 677504 745814 677510 745878
rect 59631 745726 64638 745728
rect 59631 745670 59636 745726
rect 59692 745670 64638 745726
rect 59631 745668 64638 745670
rect 59631 745665 59697 745668
rect 57615 745284 57681 745287
rect 57615 745282 64638 745284
rect 57615 745226 57620 745282
rect 57676 745226 64638 745282
rect 57615 745224 64638 745226
rect 57615 745221 57681 745224
rect 64578 744718 64638 745224
rect 58479 744100 58545 744103
rect 58479 744098 64638 744100
rect 58479 744042 58484 744098
rect 58540 744042 64638 744098
rect 58479 744040 64638 744042
rect 58479 744037 58545 744040
rect 64578 743536 64638 744040
rect 59631 742916 59697 742919
rect 59631 742914 64638 742916
rect 59631 742858 59636 742914
rect 59692 742858 64638 742914
rect 59631 742856 64638 742858
rect 59631 742853 59697 742856
rect 64578 742354 64638 742856
rect 59727 741732 59793 741735
rect 59727 741730 64638 741732
rect 59727 741674 59732 741730
rect 59788 741674 64638 741730
rect 59727 741672 64638 741674
rect 59727 741669 59793 741672
rect 64578 741172 64638 741672
rect 674362 741078 674368 741142
rect 674432 741140 674438 741142
rect 675279 741140 675345 741143
rect 674432 741138 675345 741140
rect 674432 741082 675284 741138
rect 675340 741082 675345 741138
rect 674432 741080 675345 741082
rect 674432 741078 674438 741080
rect 675279 741077 675345 741080
rect 674938 740338 674944 740402
rect 675008 740400 675014 740402
rect 675471 740400 675537 740403
rect 675008 740398 675537 740400
rect 675008 740342 675476 740398
rect 675532 740342 675537 740398
rect 675008 740340 675537 740342
rect 675008 740338 675014 740340
rect 675471 740337 675537 740340
rect 674554 739598 674560 739662
rect 674624 739660 674630 739662
rect 675279 739660 675345 739663
rect 674624 739658 675345 739660
rect 674624 739602 675284 739658
rect 675340 739602 675345 739658
rect 674624 739600 675345 739602
rect 674624 739598 674630 739600
rect 675279 739597 675345 739600
rect 675759 738032 675825 738035
rect 676858 738032 676864 738034
rect 675759 738030 676864 738032
rect 675759 737974 675764 738030
rect 675820 737974 676864 738030
rect 675759 737972 676864 737974
rect 675759 737969 675825 737972
rect 676858 737970 676864 737972
rect 676928 737970 676934 738034
rect 675663 735518 675729 735519
rect 675663 735514 675712 735518
rect 675776 735516 675782 735518
rect 675663 735458 675668 735514
rect 675663 735454 675712 735458
rect 675776 735456 675820 735516
rect 675776 735454 675782 735456
rect 675663 735453 675729 735454
rect 655311 734480 655377 734483
rect 649986 734478 655377 734480
rect 649986 734422 655316 734478
rect 655372 734422 655377 734478
rect 649986 734420 655377 734422
rect 649986 734402 650046 734420
rect 655311 734417 655377 734420
rect 649986 732704 650046 733220
rect 676474 732938 676480 733002
rect 676544 733000 676550 733002
rect 677050 733000 677056 733002
rect 676544 732940 677056 733000
rect 676544 732938 676550 732940
rect 677050 732938 677056 732940
rect 677120 732938 677126 733002
rect 655503 732704 655569 732707
rect 649986 732702 655569 732704
rect 649986 732646 655508 732702
rect 655564 732646 655569 732702
rect 649986 732644 655569 732646
rect 655503 732641 655569 732644
rect 676858 732494 676864 732558
rect 676928 732494 676934 732558
rect 676866 732114 676926 732494
rect 676858 732050 676864 732114
rect 676928 732050 676934 732114
rect 649986 731668 650046 732038
rect 655215 731668 655281 731671
rect 649986 731666 655281 731668
rect 649986 731610 655220 731666
rect 655276 731610 655281 731666
rect 649986 731608 655281 731610
rect 655215 731605 655281 731608
rect 674746 731606 674752 731670
rect 674816 731668 674822 731670
rect 674895 731668 674961 731671
rect 674816 731666 674961 731668
rect 674816 731610 674900 731666
rect 674956 731610 674961 731666
rect 674816 731608 674961 731610
rect 674816 731606 674822 731608
rect 674895 731605 674961 731608
rect 40378 731458 40384 731522
rect 40448 731520 40454 731522
rect 41583 731520 41649 731523
rect 40448 731518 41649 731520
rect 40448 731462 41588 731518
rect 41644 731462 41649 731518
rect 40448 731460 41649 731462
rect 40448 731458 40454 731460
rect 41583 731457 41649 731460
rect 40570 731310 40576 731374
rect 40640 731372 40646 731374
rect 41679 731372 41745 731375
rect 655695 731372 655761 731375
rect 40640 731370 41745 731372
rect 40640 731314 41684 731370
rect 41740 731314 41745 731370
rect 40640 731312 41745 731314
rect 40640 731310 40646 731312
rect 41679 731309 41745 731312
rect 649986 731370 655761 731372
rect 649986 731314 655700 731370
rect 655756 731314 655761 731370
rect 649986 731312 655761 731314
rect 649986 730856 650046 731312
rect 655695 731309 655761 731312
rect 41775 730484 41841 730487
rect 41568 730482 41841 730484
rect 41568 730426 41780 730482
rect 41836 730426 41841 730482
rect 41568 730424 41841 730426
rect 41775 730421 41841 730424
rect 654159 730188 654225 730191
rect 649986 730186 654225 730188
rect 649986 730130 654164 730186
rect 654220 730130 654225 730186
rect 649986 730128 654225 730130
rect 41775 729966 41841 729969
rect 41568 729964 41841 729966
rect 41568 729908 41780 729964
rect 41836 729908 41841 729964
rect 41568 729906 41841 729908
rect 41775 729903 41841 729906
rect 649986 729674 650046 730128
rect 654159 730125 654225 730128
rect 41775 729448 41841 729451
rect 41568 729446 41841 729448
rect 41568 729390 41780 729446
rect 41836 729390 41841 729446
rect 41568 729388 41841 729390
rect 41775 729385 41841 729388
rect 41775 729004 41841 729007
rect 41568 729002 41841 729004
rect 41568 728946 41780 729002
rect 41836 728946 41841 729002
rect 41568 728944 41841 728946
rect 41775 728941 41841 728944
rect 654063 728560 654129 728563
rect 649986 728558 654129 728560
rect 649986 728502 654068 728558
rect 654124 728502 654129 728558
rect 649986 728500 654129 728502
rect 649986 728492 650046 728500
rect 654063 728497 654129 728500
rect 674511 728560 674577 728563
rect 676282 728560 676288 728562
rect 674511 728558 676288 728560
rect 674511 728502 674516 728558
rect 674572 728502 676288 728558
rect 674511 728500 676288 728502
rect 674511 728497 674577 728500
rect 676282 728498 676288 728500
rect 676352 728498 676358 728562
rect 41775 728412 41841 728415
rect 41568 728410 41841 728412
rect 41568 728354 41780 728410
rect 41836 728354 41841 728410
rect 41568 728352 41841 728354
rect 41775 728349 41841 728352
rect 676666 728054 676672 728118
rect 676736 728116 676742 728118
rect 679791 728116 679857 728119
rect 676736 728114 679857 728116
rect 676736 728058 679796 728114
rect 679852 728058 679857 728114
rect 676736 728056 679857 728058
rect 676736 728054 676742 728056
rect 679791 728053 679857 728056
rect 41775 727968 41841 727971
rect 41568 727966 41841 727968
rect 41568 727910 41780 727966
rect 41836 727910 41841 727966
rect 41568 727908 41841 727910
rect 41775 727905 41841 727908
rect 41583 727672 41649 727675
rect 41538 727670 41649 727672
rect 41538 727614 41588 727670
rect 41644 727614 41649 727670
rect 41538 727609 41649 727614
rect 41538 727494 41598 727609
rect 41775 726932 41841 726935
rect 41568 726930 41841 726932
rect 41568 726874 41780 726930
rect 41836 726874 41841 726930
rect 41568 726872 41841 726874
rect 41775 726869 41841 726872
rect 41679 726784 41745 726787
rect 41538 726782 41745 726784
rect 41538 726726 41684 726782
rect 41740 726726 41745 726782
rect 41538 726724 41745 726726
rect 41538 726384 41598 726724
rect 41679 726721 41745 726724
rect 41775 726044 41841 726047
rect 41568 726042 41841 726044
rect 41568 725986 41780 726042
rect 41836 725986 41841 726042
rect 41568 725984 41841 725986
rect 41775 725981 41841 725984
rect 41871 725452 41937 725455
rect 41568 725450 41937 725452
rect 41568 725394 41876 725450
rect 41932 725394 41937 725450
rect 41568 725392 41937 725394
rect 41871 725389 41937 725392
rect 39810 724715 39870 724904
rect 39759 724710 39870 724715
rect 39759 724654 39764 724710
rect 39820 724654 39870 724710
rect 39759 724652 39870 724654
rect 39759 724649 39825 724652
rect 41967 724564 42033 724567
rect 41568 724562 42033 724564
rect 41568 724506 41972 724562
rect 42028 724506 42033 724562
rect 41568 724504 42033 724506
rect 41967 724501 42033 724504
rect 41679 724120 41745 724123
rect 41538 724118 41745 724120
rect 41538 724062 41684 724118
rect 41740 724062 41745 724118
rect 41538 724060 41745 724062
rect 41538 723942 41598 724060
rect 41679 724057 41745 724060
rect 41775 723380 41841 723383
rect 41568 723378 41841 723380
rect 41568 723322 41780 723378
rect 41836 723322 41841 723378
rect 41568 723320 41841 723322
rect 41775 723317 41841 723320
rect 34434 722791 34494 722980
rect 34434 722786 34545 722791
rect 34434 722730 34484 722786
rect 34540 722730 34545 722786
rect 34434 722728 34545 722730
rect 34479 722725 34545 722728
rect 42159 722492 42225 722495
rect 41568 722490 42225 722492
rect 41568 722434 42164 722490
rect 42220 722434 42225 722490
rect 41568 722432 42225 722434
rect 42159 722429 42225 722432
rect 42255 721900 42321 721903
rect 41568 721898 42321 721900
rect 41568 721842 42260 721898
rect 42316 721842 42321 721898
rect 41568 721840 42321 721842
rect 42255 721837 42321 721840
rect 41538 721311 41598 721500
rect 41538 721306 41649 721311
rect 41538 721250 41588 721306
rect 41644 721250 41649 721306
rect 41538 721248 41649 721250
rect 41583 721245 41649 721248
rect 41538 720719 41598 720982
rect 41538 720714 41649 720719
rect 41538 720658 41588 720714
rect 41644 720658 41649 720714
rect 41538 720656 41649 720658
rect 41583 720653 41649 720656
rect 42063 720420 42129 720423
rect 41568 720418 42129 720420
rect 41568 720362 42068 720418
rect 42124 720362 42129 720418
rect 41568 720360 42129 720362
rect 42063 720357 42129 720360
rect 41538 719831 41598 719946
rect 41538 719826 41649 719831
rect 41538 719770 41588 719826
rect 41644 719770 41649 719826
rect 41538 719768 41649 719770
rect 41583 719765 41649 719768
rect 41538 719239 41598 719502
rect 41538 719234 41649 719239
rect 41538 719178 41588 719234
rect 41644 719178 41649 719234
rect 41538 719176 41649 719178
rect 41583 719173 41649 719176
rect 41568 718880 41790 718940
rect 28866 718203 28926 718466
rect 41730 718348 41790 718880
rect 28815 718198 28926 718203
rect 28815 718142 28820 718198
rect 28876 718142 28926 718198
rect 28815 718140 28926 718142
rect 41538 718288 41790 718348
rect 28815 718137 28881 718140
rect 41538 717759 41598 718288
rect 28815 717756 28881 717759
rect 28815 717754 28926 717756
rect 28815 717698 28820 717754
rect 28876 717698 28926 717754
rect 28815 717693 28926 717698
rect 41487 717754 41598 717759
rect 41487 717698 41492 717754
rect 41548 717698 41598 717754
rect 41487 717696 41598 717698
rect 41487 717693 41553 717696
rect 28866 717430 28926 717693
rect 42735 715834 42801 715835
rect 42682 715832 42688 715834
rect 42644 715772 42688 715832
rect 42752 715830 42801 715834
rect 42796 715774 42801 715830
rect 42682 715770 42688 715772
rect 42752 715770 42801 715774
rect 42735 715769 42801 715770
rect 34479 715684 34545 715687
rect 40378 715684 40384 715686
rect 34479 715682 40384 715684
rect 34479 715626 34484 715682
rect 34540 715626 40384 715682
rect 34479 715624 40384 715626
rect 34479 715621 34545 715624
rect 40378 715622 40384 715624
rect 40448 715622 40454 715686
rect 676290 715539 676350 715654
rect 676290 715534 676401 715539
rect 676290 715478 676340 715534
rect 676396 715478 676401 715534
rect 676290 715476 676401 715478
rect 676335 715473 676401 715476
rect 39759 714944 39825 714947
rect 41338 714944 41344 714946
rect 39759 714942 41344 714944
rect 39759 714886 39764 714942
rect 39820 714886 41344 714942
rect 39759 714884 41344 714886
rect 39759 714881 39825 714884
rect 41338 714882 41344 714884
rect 41408 714882 41414 714946
rect 676143 714944 676209 714947
rect 676290 714944 676350 715136
rect 676143 714942 676350 714944
rect 676143 714886 676148 714942
rect 676204 714886 676350 714942
rect 676143 714884 676350 714886
rect 676143 714881 676209 714884
rect 676239 714796 676305 714799
rect 676239 714794 676350 714796
rect 676239 714738 676244 714794
rect 676300 714738 676350 714794
rect 676239 714733 676350 714738
rect 676290 714618 676350 714733
rect 42831 714502 42897 714503
rect 42831 714498 42880 714502
rect 42944 714500 42950 714502
rect 42831 714442 42836 714498
rect 42831 714438 42880 714442
rect 42944 714440 42988 714500
rect 42944 714438 42950 714440
rect 42831 714437 42897 714438
rect 42159 714206 42225 714207
rect 42106 714204 42112 714206
rect 42068 714144 42112 714204
rect 42176 714202 42225 714206
rect 42220 714146 42225 714202
rect 42106 714142 42112 714144
rect 42176 714142 42225 714146
rect 42159 714141 42225 714142
rect 676047 714204 676113 714207
rect 676047 714202 676320 714204
rect 676047 714146 676052 714202
rect 676108 714146 676320 714202
rect 676047 714144 676320 714146
rect 676047 714141 676113 714144
rect 41967 714056 42033 714059
rect 42490 714056 42496 714058
rect 41967 714054 42496 714056
rect 41967 713998 41972 714054
rect 42028 713998 42496 714054
rect 41967 713996 42496 713998
rect 41967 713993 42033 713996
rect 42490 713994 42496 713996
rect 42560 713994 42566 714058
rect 42063 713908 42129 713911
rect 42298 713908 42304 713910
rect 42063 713906 42304 713908
rect 42063 713850 42068 713906
rect 42124 713850 42304 713906
rect 42063 713848 42304 713850
rect 42063 713845 42129 713848
rect 42298 713846 42304 713848
rect 42368 713846 42374 713910
rect 676290 713467 676350 713582
rect 676239 713462 676350 713467
rect 676239 713406 676244 713462
rect 676300 713406 676350 713462
rect 676239 713404 676350 713406
rect 676239 713401 676305 713404
rect 676047 713168 676113 713171
rect 676047 713166 676320 713168
rect 676047 713110 676052 713166
rect 676108 713110 676320 713166
rect 676047 713108 676320 713110
rect 676047 713105 676113 713108
rect 676047 712724 676113 712727
rect 676047 712722 676320 712724
rect 676047 712666 676052 712722
rect 676108 712666 676320 712722
rect 676047 712664 676320 712666
rect 676047 712661 676113 712664
rect 676290 711987 676350 712102
rect 676239 711982 676350 711987
rect 676239 711926 676244 711982
rect 676300 711926 676350 711982
rect 676239 711924 676350 711926
rect 676239 711921 676305 711924
rect 676047 711614 676113 711617
rect 676047 711612 676320 711614
rect 676047 711556 676052 711612
rect 676108 711556 676320 711612
rect 676047 711554 676320 711556
rect 676047 711551 676113 711554
rect 674170 711182 674176 711246
rect 674240 711244 674246 711246
rect 674240 711184 676320 711244
rect 674240 711182 674246 711184
rect 42298 711034 42304 711098
rect 42368 711096 42374 711098
rect 42927 711096 42993 711099
rect 42368 711094 42993 711096
rect 42368 711038 42932 711094
rect 42988 711038 42993 711094
rect 42368 711036 42993 711038
rect 42368 711034 42374 711036
rect 42927 711033 42993 711036
rect 42490 710738 42496 710802
rect 42560 710800 42566 710802
rect 42831 710800 42897 710803
rect 42560 710798 42897 710800
rect 42560 710742 42836 710798
rect 42892 710742 42897 710798
rect 42560 710740 42897 710742
rect 42560 710738 42566 710740
rect 42831 710737 42897 710740
rect 675898 710590 675904 710654
rect 675968 710652 675974 710654
rect 675968 710592 676320 710652
rect 675968 710590 675974 710592
rect 675130 710442 675136 710506
rect 675200 710504 675206 710506
rect 675200 710444 676350 710504
rect 675200 710442 675206 710444
rect 676290 710104 676350 710444
rect 675322 709702 675328 709766
rect 675392 709764 675398 709766
rect 675392 709704 676320 709764
rect 675392 709702 675398 709704
rect 675514 709110 675520 709174
rect 675584 709172 675590 709174
rect 675584 709112 676320 709172
rect 675584 709110 675590 709112
rect 676047 708580 676113 708583
rect 676047 708578 676320 708580
rect 676047 708522 676052 708578
rect 676108 708522 676320 708578
rect 676047 708520 676320 708522
rect 676047 708517 676113 708520
rect 42874 708222 42880 708286
rect 42944 708284 42950 708286
rect 43023 708284 43089 708287
rect 42944 708282 43089 708284
rect 42944 708226 43028 708282
rect 43084 708226 43089 708282
rect 42944 708224 43089 708226
rect 42944 708222 42950 708224
rect 43023 708221 43089 708224
rect 676047 708210 676113 708213
rect 676047 708208 676320 708210
rect 676047 708152 676052 708208
rect 676108 708152 676320 708208
rect 676047 708150 676320 708152
rect 676047 708147 676113 708150
rect 42159 707990 42225 707991
rect 42106 707988 42112 707990
rect 42068 707928 42112 707988
rect 42176 707986 42225 707990
rect 42220 707930 42225 707986
rect 42106 707926 42112 707928
rect 42176 707926 42225 707930
rect 676090 707926 676096 707990
rect 676160 707988 676166 707990
rect 676160 707928 676350 707988
rect 676160 707926 676166 707928
rect 42159 707925 42225 707926
rect 676290 707662 676350 707928
rect 42682 707186 42688 707250
rect 42752 707248 42758 707250
rect 43119 707248 43185 707251
rect 42752 707246 43185 707248
rect 42752 707190 43124 707246
rect 43180 707190 43185 707246
rect 42752 707188 43185 707190
rect 42752 707186 42758 707188
rect 43119 707185 43185 707188
rect 673978 707038 673984 707102
rect 674048 707100 674054 707102
rect 674048 707040 676320 707100
rect 674048 707038 674054 707040
rect 679791 706952 679857 706955
rect 679746 706950 679857 706952
rect 679746 706894 679796 706950
rect 679852 706894 679857 706950
rect 679746 706889 679857 706894
rect 679746 706700 679806 706889
rect 677242 706446 677248 706510
rect 677312 706446 677318 706510
rect 677250 706182 677310 706446
rect 676047 705620 676113 705623
rect 676047 705618 676320 705620
rect 676047 705562 676052 705618
rect 676108 705562 676320 705618
rect 676047 705560 676320 705562
rect 676047 705557 676113 705560
rect 677434 705410 677440 705474
rect 677504 705410 677510 705474
rect 41338 705114 41344 705178
rect 41408 705176 41414 705178
rect 42735 705176 42801 705179
rect 41408 705174 42801 705176
rect 41408 705118 42740 705174
rect 42796 705118 42801 705174
rect 677442 705146 677502 705410
rect 41408 705116 42801 705118
rect 41408 705114 41414 705116
rect 42735 705113 42801 705116
rect 676239 704880 676305 704883
rect 676239 704878 676350 704880
rect 676239 704822 676244 704878
rect 676300 704822 676350 704878
rect 676239 704817 676350 704822
rect 676290 704702 676350 704817
rect 59631 704436 59697 704439
rect 679983 704436 680049 704439
rect 59631 704434 64638 704436
rect 59631 704378 59636 704434
rect 59692 704378 64638 704434
rect 59631 704376 64638 704378
rect 59631 704373 59697 704376
rect 40378 704078 40384 704142
rect 40448 704140 40454 704142
rect 42927 704140 42993 704143
rect 40448 704138 42993 704140
rect 40448 704082 42932 704138
rect 42988 704082 42993 704138
rect 40448 704080 42993 704082
rect 40448 704078 40454 704080
rect 42927 704077 42993 704080
rect 64578 703860 64638 704376
rect 679938 704434 680049 704436
rect 679938 704378 679988 704434
rect 680044 704378 680049 704434
rect 679938 704373 680049 704378
rect 679938 704110 679998 704373
rect 679746 703403 679806 703666
rect 679746 703398 679857 703403
rect 679983 703400 680049 703403
rect 679746 703342 679796 703398
rect 679852 703342 679857 703398
rect 679746 703340 679857 703342
rect 679791 703337 679857 703340
rect 679938 703398 680049 703400
rect 679938 703342 679988 703398
rect 680044 703342 680049 703398
rect 679938 703337 680049 703342
rect 679938 703148 679998 703337
rect 679791 702956 679857 702959
rect 679746 702954 679857 702956
rect 679746 702898 679796 702954
rect 679852 702898 679857 702954
rect 679746 702893 679857 702898
rect 58767 702660 58833 702663
rect 64578 702660 64638 702678
rect 58767 702658 64638 702660
rect 58767 702602 58772 702658
rect 58828 702602 64638 702658
rect 679746 702630 679806 702893
rect 58767 702600 64638 702602
rect 58767 702597 58833 702600
rect 43791 702068 43857 702071
rect 43791 702066 64638 702068
rect 43791 702010 43796 702066
rect 43852 702010 64638 702066
rect 43791 702008 64638 702010
rect 43791 702005 43857 702008
rect 64578 701496 64638 702008
rect 58671 700884 58737 700887
rect 58671 700882 64638 700884
rect 58671 700826 58676 700882
rect 58732 700826 64638 700882
rect 58671 700824 64638 700826
rect 58671 700821 58737 700824
rect 64578 700314 64638 700824
rect 59247 699700 59313 699703
rect 59247 699698 64638 699700
rect 59247 699642 59252 699698
rect 59308 699642 64638 699698
rect 59247 699640 64638 699642
rect 59247 699637 59313 699640
rect 64578 699132 64638 699640
rect 58863 698516 58929 698519
rect 58863 698514 64638 698516
rect 58863 698458 58868 698514
rect 58924 698458 64638 698514
rect 58863 698456 64638 698458
rect 58863 698453 58929 698456
rect 64578 697950 64638 698456
rect 675130 697862 675136 697926
rect 675200 697924 675206 697926
rect 675375 697924 675441 697927
rect 675200 697922 675441 697924
rect 675200 697866 675380 697922
rect 675436 697866 675441 697922
rect 675200 697864 675441 697866
rect 675200 697862 675206 697864
rect 675375 697861 675441 697864
rect 675759 697184 675825 697187
rect 675898 697184 675904 697186
rect 675759 697182 675904 697184
rect 675759 697126 675764 697182
rect 675820 697126 675904 697182
rect 675759 697124 675904 697126
rect 675759 697121 675825 697124
rect 675898 697122 675904 697124
rect 675968 697122 675974 697186
rect 674170 696974 674176 697038
rect 674240 697036 674246 697038
rect 675183 697036 675249 697039
rect 674240 697034 675249 697036
rect 674240 696978 675188 697034
rect 675244 696978 675249 697034
rect 674240 696976 675249 696978
rect 674240 696974 674246 696976
rect 675183 696973 675249 696976
rect 675567 694818 675633 694819
rect 675514 694816 675520 694818
rect 675476 694756 675520 694816
rect 675584 694814 675633 694818
rect 675628 694758 675633 694814
rect 675514 694754 675520 694756
rect 675584 694754 675633 694758
rect 675567 694753 675633 694754
rect 675759 694224 675825 694227
rect 676666 694224 676672 694226
rect 675759 694222 676672 694224
rect 675759 694166 675764 694222
rect 675820 694166 676672 694222
rect 675759 694164 676672 694166
rect 675759 694161 675825 694164
rect 676666 694162 676672 694164
rect 676736 694162 676742 694226
rect 649986 689488 650046 689980
rect 655119 689488 655185 689491
rect 649986 689486 655185 689488
rect 649986 689430 655124 689486
rect 655180 689430 655185 689486
rect 649986 689428 655185 689430
rect 655119 689425 655185 689428
rect 649986 688452 650046 688798
rect 655407 688452 655473 688455
rect 649986 688450 655473 688452
rect 649986 688394 655412 688450
rect 655468 688394 655473 688450
rect 649986 688392 655473 688394
rect 655407 688389 655473 688392
rect 649986 687120 650046 687616
rect 655599 687120 655665 687123
rect 649986 687118 655665 687120
rect 649986 687062 655604 687118
rect 655660 687062 655665 687118
rect 649986 687060 655665 687062
rect 655599 687057 655665 687060
rect 654351 686972 654417 686975
rect 649986 686970 654417 686972
rect 649986 686914 654356 686970
rect 654412 686914 654417 686970
rect 649986 686912 654417 686914
rect 41775 686898 41841 686901
rect 41568 686896 41841 686898
rect 41568 686840 41780 686896
rect 41836 686840 41841 686896
rect 41568 686838 41841 686840
rect 41775 686835 41841 686838
rect 649986 686434 650046 686912
rect 654351 686909 654417 686912
rect 674895 686528 674961 686531
rect 677050 686528 677056 686530
rect 674895 686526 677056 686528
rect 674895 686470 674900 686526
rect 674956 686470 677056 686526
rect 674895 686468 677056 686470
rect 674895 686465 674961 686468
rect 677050 686466 677056 686468
rect 677120 686466 677126 686530
rect 41775 686380 41841 686383
rect 41568 686378 41841 686380
rect 41568 686322 41780 686378
rect 41836 686322 41841 686378
rect 41568 686320 41841 686322
rect 41775 686317 41841 686320
rect 41538 685643 41598 685758
rect 41538 685638 41649 685643
rect 41538 685582 41588 685638
rect 41644 685582 41649 685638
rect 41538 685580 41649 685582
rect 41583 685577 41649 685580
rect 41775 685344 41841 685347
rect 654159 685344 654225 685347
rect 41568 685342 41841 685344
rect 41568 685286 41780 685342
rect 41836 685286 41841 685342
rect 41568 685284 41841 685286
rect 41775 685281 41841 685284
rect 649986 685342 654225 685344
rect 649986 685286 654164 685342
rect 654220 685286 654225 685342
rect 649986 685284 654225 685286
rect 649986 685252 650046 685284
rect 654159 685281 654225 685284
rect 41775 684900 41841 684903
rect 41568 684898 41841 684900
rect 41568 684842 41780 684898
rect 41836 684842 41841 684898
rect 41568 684840 41841 684842
rect 41775 684837 41841 684840
rect 654063 684604 654129 684607
rect 649986 684602 654129 684604
rect 649986 684546 654068 684602
rect 654124 684546 654129 684602
rect 649986 684544 654129 684546
rect 40578 684162 40638 684278
rect 40570 684098 40576 684162
rect 40640 684098 40646 684162
rect 649986 684070 650046 684544
rect 654063 684541 654129 684544
rect 41775 683864 41841 683867
rect 41568 683862 41841 683864
rect 41568 683806 41780 683862
rect 41836 683806 41841 683862
rect 41568 683804 41841 683806
rect 41775 683801 41841 683804
rect 40386 682978 40446 683390
rect 40378 682914 40384 682978
rect 40448 682914 40454 682978
rect 41583 682976 41649 682979
rect 41538 682974 41649 682976
rect 41538 682918 41588 682974
rect 41644 682918 41649 682974
rect 41538 682913 41649 682918
rect 41538 682798 41598 682913
rect 39810 682239 39870 682354
rect 39759 682234 39870 682239
rect 39759 682178 39764 682234
rect 39820 682178 39870 682234
rect 39759 682176 39870 682178
rect 39759 682173 39825 682176
rect 41775 681866 41841 681869
rect 41568 681864 41841 681866
rect 41568 681808 41780 681864
rect 41836 681808 41841 681864
rect 41568 681806 41841 681808
rect 41775 681803 41841 681806
rect 39855 681496 39921 681499
rect 39810 681494 39921 681496
rect 39810 681438 39860 681494
rect 39916 681438 39921 681494
rect 39810 681433 39921 681438
rect 39810 681318 39870 681433
rect 37314 680759 37374 680874
rect 37314 680754 37425 680759
rect 37314 680698 37364 680754
rect 37420 680698 37425 680754
rect 37314 680696 37425 680698
rect 37359 680693 37425 680696
rect 41967 680312 42033 680315
rect 41568 680310 42033 680312
rect 41568 680254 41972 680310
rect 42028 680254 42033 680310
rect 41568 680252 42033 680254
rect 41967 680249 42033 680252
rect 41775 679868 41841 679871
rect 41568 679866 41841 679868
rect 41568 679810 41780 679866
rect 41836 679810 41841 679866
rect 41568 679808 41841 679810
rect 41775 679805 41841 679808
rect 40194 679131 40254 679394
rect 40194 679126 40305 679131
rect 40194 679070 40244 679126
rect 40300 679070 40305 679126
rect 40194 679068 40305 679070
rect 40239 679065 40305 679068
rect 34434 678687 34494 678802
rect 34434 678682 34545 678687
rect 34434 678626 34484 678682
rect 34540 678626 34545 678682
rect 34434 678624 34545 678626
rect 34479 678621 34545 678624
rect 42255 678388 42321 678391
rect 41568 678386 42321 678388
rect 41568 678330 42260 678386
rect 42316 678330 42321 678386
rect 41568 678328 42321 678330
rect 42255 678325 42321 678328
rect 41871 677944 41937 677947
rect 41568 677942 41937 677944
rect 41568 677886 41876 677942
rect 41932 677886 41937 677942
rect 41568 677884 41937 677886
rect 41871 677881 41937 677884
rect 42063 677352 42129 677355
rect 41568 677350 42129 677352
rect 41568 677294 42068 677350
rect 42124 677294 42129 677350
rect 41568 677292 42129 677294
rect 42063 677289 42129 677292
rect 41538 676612 41598 676804
rect 41679 676612 41745 676615
rect 41538 676610 41745 676612
rect 41538 676554 41684 676610
rect 41740 676554 41745 676610
rect 41538 676552 41745 676554
rect 41679 676549 41745 676552
rect 41538 676171 41598 676434
rect 41538 676166 41649 676171
rect 41538 676110 41588 676166
rect 41644 676110 41649 676166
rect 41538 676108 41649 676110
rect 41583 676105 41649 676108
rect 41538 675727 41598 675842
rect 41538 675722 41649 675727
rect 41538 675666 41588 675722
rect 41644 675666 41649 675722
rect 41538 675664 41649 675666
rect 41583 675661 41649 675664
rect 41538 675132 41598 675250
rect 41538 675072 41790 675132
rect 23106 674543 23166 674954
rect 41730 674688 41790 675072
rect 23055 674538 23166 674543
rect 23055 674482 23060 674538
rect 23116 674482 23166 674538
rect 23055 674480 23166 674482
rect 41538 674628 41790 674688
rect 23055 674477 23121 674480
rect 41538 674099 41598 674628
rect 23055 674096 23121 674099
rect 23055 674094 23166 674096
rect 23055 674038 23060 674094
rect 23116 674038 23166 674094
rect 23055 674033 23166 674038
rect 41538 674094 41649 674099
rect 41538 674038 41588 674094
rect 41644 674038 41649 674094
rect 41538 674036 41649 674038
rect 41583 674033 41649 674036
rect 23106 673770 23166 674033
rect 40239 673652 40305 673655
rect 41530 673652 41536 673654
rect 40239 673650 41536 673652
rect 40239 673594 40244 673650
rect 40300 673594 41536 673650
rect 40239 673592 41536 673594
rect 40239 673589 40305 673592
rect 41530 673590 41536 673592
rect 41600 673590 41606 673654
rect 39855 671136 39921 671139
rect 41338 671136 41344 671138
rect 39855 671134 41344 671136
rect 39855 671078 39860 671134
rect 39916 671078 41344 671134
rect 39855 671076 41344 671078
rect 39855 671073 39921 671076
rect 41338 671074 41344 671076
rect 41408 671074 41414 671138
rect 41679 670990 41745 670991
rect 41679 670988 41728 670990
rect 41636 670986 41728 670988
rect 41636 670930 41684 670986
rect 41636 670928 41728 670930
rect 41679 670926 41728 670928
rect 41792 670926 41798 670990
rect 41679 670925 41745 670926
rect 41871 670842 41937 670843
rect 41871 670840 41920 670842
rect 41828 670838 41920 670840
rect 41828 670782 41876 670838
rect 41828 670780 41920 670782
rect 41871 670778 41920 670780
rect 41984 670778 41990 670842
rect 41871 670777 41937 670778
rect 42063 670694 42129 670695
rect 42063 670692 42112 670694
rect 42020 670690 42112 670692
rect 42020 670634 42068 670690
rect 42020 670632 42112 670634
rect 42063 670630 42112 670632
rect 42176 670630 42182 670694
rect 42063 670629 42129 670630
rect 676290 668771 676350 669034
rect 676239 668766 676350 668771
rect 676239 668710 676244 668766
rect 676300 668710 676350 668766
rect 676239 668708 676350 668710
rect 676239 668705 676305 668708
rect 676290 668327 676350 668516
rect 676239 668322 676350 668327
rect 676239 668266 676244 668322
rect 676300 668266 676350 668322
rect 676239 668264 676350 668266
rect 676239 668261 676305 668264
rect 676047 668028 676113 668031
rect 676047 668026 676320 668028
rect 676047 667970 676052 668026
rect 676108 667970 676320 668026
rect 676047 667968 676320 667970
rect 676047 667965 676113 667968
rect 675951 667584 676017 667587
rect 675951 667582 676320 667584
rect 675951 667526 675956 667582
rect 676012 667526 676320 667582
rect 675951 667524 676320 667526
rect 675951 667521 676017 667524
rect 676290 666847 676350 667036
rect 676239 666842 676350 666847
rect 676239 666786 676244 666842
rect 676300 666786 676350 666842
rect 676239 666784 676350 666786
rect 676239 666781 676305 666784
rect 41871 666698 41937 666699
rect 41871 666694 41920 666698
rect 41984 666696 41990 666698
rect 676143 666696 676209 666699
rect 41871 666638 41876 666694
rect 41871 666634 41920 666638
rect 41984 666636 42028 666696
rect 676143 666694 676350 666696
rect 676143 666638 676148 666694
rect 676204 666638 676350 666694
rect 676143 666636 676350 666638
rect 41984 666634 41990 666636
rect 41871 666633 41937 666634
rect 676143 666633 676209 666636
rect 676290 666518 676350 666636
rect 675951 666104 676017 666107
rect 675951 666102 676320 666104
rect 675951 666046 675956 666102
rect 676012 666046 676320 666102
rect 675951 666044 676320 666046
rect 675951 666041 676017 666044
rect 675951 665512 676017 665515
rect 675951 665510 676320 665512
rect 675951 665454 675956 665510
rect 676012 665454 676320 665510
rect 675951 665452 676320 665454
rect 675951 665449 676017 665452
rect 675951 665068 676017 665071
rect 675951 665066 676320 665068
rect 675951 665010 675956 665066
rect 676012 665010 676320 665066
rect 675951 665008 676320 665010
rect 675951 665005 676017 665008
rect 42159 664774 42225 664775
rect 42106 664772 42112 664774
rect 42068 664712 42112 664772
rect 42176 664770 42225 664774
rect 42220 664714 42225 664770
rect 42106 664710 42112 664712
rect 42176 664710 42225 664714
rect 42159 664709 42225 664710
rect 674362 664562 674368 664626
rect 674432 664624 674438 664626
rect 674432 664564 676320 664624
rect 674432 664562 674438 664564
rect 676047 664032 676113 664035
rect 676047 664030 676320 664032
rect 676047 663974 676052 664030
rect 676108 663974 676320 664030
rect 676047 663972 676320 663974
rect 676047 663969 676113 663972
rect 676282 663822 676288 663886
rect 676352 663822 676358 663886
rect 676290 663484 676350 663822
rect 674938 663082 674944 663146
rect 675008 663144 675014 663146
rect 675008 663084 676320 663144
rect 675008 663082 675014 663084
rect 675706 662490 675712 662554
rect 675776 662552 675782 662554
rect 675776 662492 676320 662552
rect 675776 662490 675782 662492
rect 676047 662034 676113 662037
rect 676047 662032 676320 662034
rect 676047 661976 676052 662032
rect 676108 661976 676320 662032
rect 676047 661974 676320 661976
rect 676047 661971 676113 661974
rect 674746 661602 674752 661666
rect 674816 661664 674822 661666
rect 674816 661604 676320 661664
rect 674816 661602 674822 661604
rect 59631 661220 59697 661223
rect 59631 661218 64638 661220
rect 59631 661162 59636 661218
rect 59692 661162 64638 661218
rect 59631 661160 64638 661162
rect 59631 661157 59697 661160
rect 41775 660926 41841 660927
rect 41722 660924 41728 660926
rect 41684 660864 41728 660924
rect 41792 660922 41841 660926
rect 41836 660866 41841 660922
rect 41722 660862 41728 660864
rect 41792 660862 41841 660866
rect 41775 660861 41841 660862
rect 64578 660638 64638 661160
rect 674554 661010 674560 661074
rect 674624 661072 674630 661074
rect 674624 661012 676320 661072
rect 674624 661010 674630 661012
rect 676047 660480 676113 660483
rect 676047 660478 676320 660480
rect 676047 660422 676052 660478
rect 676108 660422 676320 660478
rect 676047 660420 676320 660422
rect 676047 660417 676113 660420
rect 41338 660270 41344 660334
rect 41408 660332 41414 660334
rect 42927 660332 42993 660335
rect 41408 660330 42993 660332
rect 41408 660274 42932 660330
rect 42988 660274 42993 660330
rect 41408 660272 42993 660274
rect 41408 660270 41414 660272
rect 42927 660269 42993 660272
rect 676047 660110 676113 660113
rect 676047 660108 676320 660110
rect 676047 660052 676052 660108
rect 676108 660052 676320 660108
rect 676047 660050 676320 660052
rect 676047 660047 676113 660050
rect 41530 659678 41536 659742
rect 41600 659740 41606 659742
rect 42831 659740 42897 659743
rect 41600 659738 42897 659740
rect 41600 659682 42836 659738
rect 42892 659682 42897 659738
rect 41600 659680 42897 659682
rect 41600 659678 41606 659680
rect 42831 659677 42897 659680
rect 676239 659740 676305 659743
rect 676239 659738 676350 659740
rect 676239 659682 676244 659738
rect 676300 659682 676350 659738
rect 676239 659677 676350 659682
rect 676290 659562 676350 659677
rect 58767 659444 58833 659447
rect 64578 659444 64638 659456
rect 58767 659442 64638 659444
rect 58767 659386 58772 659442
rect 58828 659386 64638 659442
rect 58767 659384 64638 659386
rect 58767 659381 58833 659384
rect 676858 659234 676864 659298
rect 676928 659234 676934 659298
rect 676866 658970 676926 659234
rect 45903 658852 45969 658855
rect 45903 658850 64638 658852
rect 45903 658794 45908 658850
rect 45964 658794 64638 658850
rect 45903 658792 64638 658794
rect 45903 658789 45969 658792
rect 64578 658274 64638 658792
rect 676047 658630 676113 658633
rect 676047 658628 676320 658630
rect 676047 658572 676052 658628
rect 676108 658572 676320 658628
rect 676047 658570 676320 658572
rect 676047 658567 676113 658570
rect 676239 658260 676305 658263
rect 676239 658258 676350 658260
rect 676239 658202 676244 658258
rect 676300 658202 676350 658258
rect 676239 658197 676350 658202
rect 676290 658082 676350 658197
rect 59151 657668 59217 657671
rect 59151 657666 64638 657668
rect 59151 657610 59156 657666
rect 59212 657610 64638 657666
rect 59151 657608 64638 657610
rect 59151 657605 59217 657608
rect 64578 657092 64638 657608
rect 679938 657375 679998 657490
rect 679938 657370 680049 657375
rect 679938 657314 679988 657370
rect 680044 657314 680049 657370
rect 679938 657312 680049 657314
rect 679983 657309 680049 657312
rect 679746 656783 679806 657046
rect 679746 656778 679857 656783
rect 679983 656780 680049 656783
rect 679746 656722 679796 656778
rect 679852 656722 679857 656778
rect 679746 656720 679857 656722
rect 679791 656717 679857 656720
rect 679938 656778 680049 656780
rect 679938 656722 679988 656778
rect 680044 656722 680049 656778
rect 679938 656717 680049 656722
rect 679938 656602 679998 656717
rect 58191 656484 58257 656487
rect 58191 656482 64638 656484
rect 58191 656426 58196 656482
rect 58252 656426 64638 656482
rect 58191 656424 64638 656426
rect 58191 656421 58257 656424
rect 64578 655910 64638 656424
rect 679791 656336 679857 656339
rect 679746 656334 679857 656336
rect 679746 656278 679796 656334
rect 679852 656278 679857 656334
rect 679746 656273 679857 656278
rect 679746 656010 679806 656273
rect 58383 655300 58449 655303
rect 58383 655298 64638 655300
rect 58383 655242 58388 655298
rect 58444 655242 64638 655298
rect 58383 655240 64638 655242
rect 58383 655237 58449 655240
rect 64578 654728 64638 655240
rect 674938 652574 674944 652638
rect 675008 652636 675014 652638
rect 675375 652636 675441 652639
rect 675008 652634 675441 652636
rect 675008 652578 675380 652634
rect 675436 652578 675441 652634
rect 675008 652576 675441 652578
rect 675008 652574 675014 652576
rect 675375 652573 675441 652576
rect 674362 652130 674368 652194
rect 674432 652192 674438 652194
rect 675471 652192 675537 652195
rect 674432 652190 675537 652192
rect 674432 652134 675476 652190
rect 675532 652134 675537 652190
rect 674432 652132 675537 652134
rect 674432 652130 674438 652132
rect 675471 652129 675537 652132
rect 674746 651390 674752 651454
rect 674816 651452 674822 651454
rect 675375 651452 675441 651455
rect 674816 651450 675441 651452
rect 674816 651394 675380 651450
rect 675436 651394 675441 651450
rect 674816 651392 675441 651394
rect 674816 651390 674822 651392
rect 675375 651389 675441 651392
rect 675375 649678 675441 649679
rect 675322 649676 675328 649678
rect 675284 649616 675328 649676
rect 675392 649674 675441 649678
rect 675436 649618 675441 649674
rect 675322 649614 675328 649616
rect 675392 649614 675441 649618
rect 675375 649613 675441 649614
rect 675663 645386 675729 645387
rect 675663 645382 675712 645386
rect 675776 645384 675782 645386
rect 675663 645326 675668 645382
rect 675663 645322 675712 645326
rect 675776 645324 675820 645384
rect 675776 645322 675782 645324
rect 675663 645321 675729 645322
rect 40570 645026 40576 645090
rect 40640 645088 40646 645090
rect 41487 645088 41553 645091
rect 40640 645086 41553 645088
rect 40640 645030 41492 645086
rect 41548 645030 41553 645086
rect 40640 645028 41553 645030
rect 40640 645026 40646 645028
rect 41487 645025 41553 645028
rect 40378 644878 40384 644942
rect 40448 644940 40454 644942
rect 41679 644940 41745 644943
rect 40448 644938 41745 644940
rect 40448 644882 41684 644938
rect 41740 644882 41745 644938
rect 40448 644880 41745 644882
rect 40448 644878 40454 644880
rect 41679 644877 41745 644880
rect 41775 643756 41841 643759
rect 41568 643754 41841 643756
rect 41568 643698 41780 643754
rect 41836 643698 41841 643754
rect 41568 643696 41841 643698
rect 41775 643693 41841 643696
rect 41775 643164 41841 643167
rect 41568 643162 41841 643164
rect 41568 643106 41780 643162
rect 41836 643106 41841 643162
rect 41568 643104 41841 643106
rect 41775 643101 41841 643104
rect 649986 643016 650046 643558
rect 655311 643016 655377 643019
rect 649986 643014 655377 643016
rect 649986 642958 655316 643014
rect 655372 642958 655377 643014
rect 649986 642956 655377 642958
rect 655311 642953 655377 642956
rect 41538 642427 41598 642542
rect 41538 642422 41649 642427
rect 655503 642424 655569 642427
rect 41538 642366 41588 642422
rect 41644 642366 41649 642422
rect 41538 642364 41649 642366
rect 649986 642422 655569 642424
rect 649986 642366 655508 642422
rect 655564 642366 655569 642422
rect 649986 642364 655569 642366
rect 41583 642361 41649 642364
rect 655503 642361 655569 642364
rect 41775 642202 41841 642205
rect 41568 642200 41841 642202
rect 41568 642144 41780 642200
rect 41836 642144 41841 642200
rect 41568 642142 41841 642144
rect 41775 642139 41841 642142
rect 41775 641684 41841 641687
rect 41568 641682 41841 641684
rect 41568 641626 41780 641682
rect 41836 641626 41841 641682
rect 41568 641624 41841 641626
rect 41775 641621 41841 641624
rect 41722 641092 41728 641094
rect 41568 641032 41728 641092
rect 41722 641030 41728 641032
rect 41792 641030 41798 641094
rect 41487 640944 41553 640947
rect 41487 640942 41598 640944
rect 41487 640886 41492 640942
rect 41548 640886 41598 640942
rect 41487 640881 41598 640886
rect 41538 640618 41598 640881
rect 649986 640796 650046 641194
rect 655695 640796 655761 640799
rect 649986 640794 655761 640796
rect 649986 640738 655700 640794
rect 655756 640738 655761 640794
rect 649986 640736 655761 640738
rect 655695 640733 655761 640736
rect 654159 640648 654225 640651
rect 649986 640646 654225 640648
rect 649986 640590 654164 640646
rect 654220 640590 654225 640646
rect 649986 640588 654225 640590
rect 41775 640204 41841 640207
rect 41568 640202 41841 640204
rect 41568 640146 41780 640202
rect 41836 640146 41841 640202
rect 41568 640144 41841 640146
rect 41775 640141 41841 640144
rect 649986 640012 650046 640588
rect 654159 640585 654225 640588
rect 673978 639994 673984 640058
rect 674048 640056 674054 640058
rect 675279 640056 675345 640059
rect 674048 640054 675345 640056
rect 674048 639998 675284 640054
rect 675340 639998 675345 640054
rect 674048 639996 675345 639998
rect 674048 639994 674054 639996
rect 675279 639993 675345 639996
rect 41679 639908 41745 639911
rect 41538 639906 41745 639908
rect 41538 639850 41684 639906
rect 41740 639850 41745 639906
rect 41538 639848 41745 639850
rect 41538 639582 41598 639848
rect 41679 639845 41745 639848
rect 655791 639168 655857 639171
rect 649986 639166 655857 639168
rect 37314 639023 37374 639138
rect 649986 639110 655796 639166
rect 655852 639110 655857 639166
rect 649986 639108 655857 639110
rect 37314 639018 37425 639023
rect 37314 638962 37364 639018
rect 37420 638962 37425 639018
rect 37314 638960 37425 638962
rect 37359 638957 37425 638960
rect 649986 638830 650046 639108
rect 655791 639105 655857 639108
rect 40239 638280 40305 638283
rect 41538 638282 41598 638694
rect 675759 638576 675825 638579
rect 676090 638576 676096 638578
rect 675759 638574 676096 638576
rect 675759 638518 675764 638574
rect 675820 638518 676096 638574
rect 675759 638516 676096 638518
rect 675759 638513 675825 638516
rect 676090 638514 676096 638516
rect 676160 638514 676166 638578
rect 40194 638278 40305 638280
rect 40194 638222 40244 638278
rect 40300 638222 40305 638278
rect 40194 638217 40305 638222
rect 41530 638218 41536 638282
rect 41600 638218 41606 638282
rect 655983 638280 656049 638283
rect 649986 638278 656049 638280
rect 649986 638222 655988 638278
rect 656044 638222 656049 638278
rect 649986 638220 656049 638222
rect 40194 638102 40254 638217
rect 40194 637543 40254 637658
rect 649986 637648 650046 638220
rect 655983 638217 656049 638220
rect 40143 637538 40254 637543
rect 40143 637482 40148 637538
rect 40204 637482 40254 637538
rect 40143 637480 40254 637482
rect 40143 637477 40209 637480
rect 41538 636951 41598 637140
rect 41487 636946 41598 636951
rect 41487 636890 41492 636946
rect 41548 636890 41598 636946
rect 41487 636888 41598 636890
rect 41487 636885 41553 636888
rect 41775 636652 41841 636655
rect 41568 636650 41841 636652
rect 41568 636594 41780 636650
rect 41836 636594 41841 636650
rect 41568 636592 41841 636594
rect 41775 636589 41841 636592
rect 676666 636590 676672 636654
rect 676736 636652 676742 636654
rect 678159 636652 678225 636655
rect 676736 636650 678225 636652
rect 676736 636594 678164 636650
rect 678220 636594 678225 636650
rect 676736 636592 678225 636594
rect 676736 636590 676742 636592
rect 678159 636589 678225 636592
rect 34434 636063 34494 636178
rect 34383 636058 34494 636063
rect 34383 636002 34388 636058
rect 34444 636002 34494 636058
rect 34383 636000 34494 636002
rect 34383 635997 34449 636000
rect 34434 635471 34494 635586
rect 34434 635466 34545 635471
rect 34434 635410 34484 635466
rect 34540 635410 34545 635466
rect 34434 635408 34545 635410
rect 34479 635405 34545 635408
rect 42063 635172 42129 635175
rect 41568 635170 42129 635172
rect 41568 635114 42068 635170
rect 42124 635114 42129 635170
rect 41568 635112 42129 635114
rect 42063 635109 42129 635112
rect 42831 634728 42897 634731
rect 41568 634726 42897 634728
rect 41568 634670 42836 634726
rect 42892 634670 42897 634726
rect 41568 634668 42897 634670
rect 42831 634665 42897 634668
rect 41538 633991 41598 634106
rect 41538 633986 41649 633991
rect 41538 633930 41588 633986
rect 41644 633930 41649 633986
rect 41538 633928 41649 633930
rect 41583 633925 41649 633928
rect 42159 633692 42225 633695
rect 41568 633690 42225 633692
rect 41568 633634 42164 633690
rect 42220 633634 42225 633690
rect 41568 633632 42225 633634
rect 42159 633629 42225 633632
rect 41871 633248 41937 633251
rect 41568 633246 41937 633248
rect 41568 633190 41876 633246
rect 41932 633190 41937 633246
rect 41568 633188 41937 633190
rect 41871 633185 41937 633188
rect 42255 632656 42321 632659
rect 41568 632654 42321 632656
rect 41568 632598 42260 632654
rect 42316 632598 42321 632654
rect 41568 632596 42321 632598
rect 42255 632593 42321 632596
rect 41538 631916 41598 632108
rect 41538 631856 41790 631916
rect 23106 631475 23166 631738
rect 23055 631470 23166 631475
rect 41730 631472 41790 631856
rect 23055 631414 23060 631470
rect 23116 631414 23166 631470
rect 23055 631412 23166 631414
rect 41538 631412 41790 631472
rect 23055 631409 23121 631412
rect 23055 631028 23121 631031
rect 23055 631026 23166 631028
rect 23055 630970 23060 631026
rect 23116 630970 23166 631026
rect 23055 630965 23166 630970
rect 23106 630554 23166 630965
rect 41538 630883 41598 631412
rect 41538 630878 41649 630883
rect 41538 630822 41588 630878
rect 41644 630822 41649 630878
rect 41538 630820 41649 630822
rect 41583 630817 41649 630820
rect 34383 628068 34449 628071
rect 40378 628068 40384 628070
rect 34383 628066 40384 628068
rect 34383 628010 34388 628066
rect 34444 628010 40384 628066
rect 34383 628008 40384 628010
rect 34383 628005 34449 628008
rect 40378 628006 40384 628008
rect 40448 628006 40454 628070
rect 40239 627920 40305 627923
rect 40762 627920 40768 627922
rect 40239 627918 40768 627920
rect 40239 627862 40244 627918
rect 40300 627862 40768 627918
rect 40239 627860 40768 627862
rect 40239 627857 40305 627860
rect 40762 627858 40768 627860
rect 40832 627858 40838 627922
rect 42063 627476 42129 627479
rect 42298 627476 42304 627478
rect 42063 627474 42304 627476
rect 42063 627418 42068 627474
rect 42124 627418 42304 627474
rect 42063 627416 42304 627418
rect 42063 627413 42129 627416
rect 42298 627414 42304 627416
rect 42368 627414 42374 627478
rect 41530 625194 41536 625258
rect 41600 625256 41606 625258
rect 42159 625256 42225 625259
rect 41600 625254 42225 625256
rect 41600 625198 42164 625254
rect 42220 625198 42225 625254
rect 41600 625196 42225 625198
rect 41600 625194 41606 625196
rect 42159 625193 42225 625196
rect 676290 625111 676350 625522
rect 676239 625106 676350 625111
rect 676239 625050 676244 625106
rect 676300 625050 676350 625106
rect 676239 625048 676350 625050
rect 676239 625045 676305 625048
rect 42298 624750 42304 624814
rect 42368 624812 42374 624814
rect 42735 624812 42801 624815
rect 42368 624810 42801 624812
rect 42368 624754 42740 624810
rect 42796 624754 42801 624810
rect 42368 624752 42801 624754
rect 42368 624750 42374 624752
rect 42735 624749 42801 624752
rect 676143 624664 676209 624667
rect 676290 624664 676350 624930
rect 676143 624662 676350 624664
rect 676143 624606 676148 624662
rect 676204 624606 676350 624662
rect 676143 624604 676350 624606
rect 676143 624601 676209 624604
rect 676290 624223 676350 624338
rect 676239 624218 676350 624223
rect 676239 624162 676244 624218
rect 676300 624162 676350 624218
rect 676239 624160 676350 624162
rect 676239 624157 676305 624160
rect 676047 623998 676113 624001
rect 676047 623996 676320 623998
rect 676047 623940 676052 623996
rect 676108 623940 676320 623996
rect 676047 623938 676320 623940
rect 676047 623935 676113 623938
rect 676047 623480 676113 623483
rect 676047 623478 676320 623480
rect 676047 623422 676052 623478
rect 676108 623422 676320 623478
rect 676047 623420 676320 623422
rect 676047 623417 676113 623420
rect 676335 623184 676401 623187
rect 676290 623182 676401 623184
rect 676290 623126 676340 623182
rect 676396 623126 676401 623182
rect 676290 623121 676401 623126
rect 676290 622858 676350 623121
rect 676047 622518 676113 622521
rect 676047 622516 676320 622518
rect 676047 622460 676052 622516
rect 676108 622460 676320 622516
rect 676047 622458 676320 622460
rect 676047 622455 676113 622458
rect 676047 622000 676113 622003
rect 676047 621998 676320 622000
rect 676047 621942 676052 621998
rect 676108 621942 676320 621998
rect 676047 621940 676320 621942
rect 676047 621937 676113 621940
rect 676047 621408 676113 621411
rect 676047 621406 676320 621408
rect 676047 621350 676052 621406
rect 676108 621350 676320 621406
rect 676047 621348 676320 621350
rect 676047 621345 676113 621348
rect 674170 620902 674176 620966
rect 674240 620964 674246 620966
rect 674240 620904 676320 620964
rect 674240 620902 674246 620904
rect 676239 620668 676305 620671
rect 676239 620666 676350 620668
rect 676239 620610 676244 620666
rect 676300 620610 676350 620666
rect 676239 620605 676350 620610
rect 676290 620490 676350 620605
rect 675130 619866 675136 619930
rect 675200 619928 675206 619930
rect 675200 619868 676320 619928
rect 675200 619866 675206 619868
rect 675514 619422 675520 619486
rect 675584 619484 675590 619486
rect 675584 619424 676320 619484
rect 675584 619422 675590 619424
rect 676047 618966 676113 618969
rect 676047 618964 676320 618966
rect 676047 618908 676052 618964
rect 676108 618908 676320 618964
rect 676047 618906 676320 618908
rect 676047 618903 676113 618906
rect 676239 618596 676305 618599
rect 676239 618594 676350 618596
rect 676239 618538 676244 618594
rect 676300 618538 676350 618594
rect 676239 618533 676350 618538
rect 676290 618418 676350 618533
rect 58959 618004 59025 618007
rect 58959 618002 64638 618004
rect 58959 617946 58964 618002
rect 59020 617946 64638 618002
rect 58959 617944 64638 617946
rect 58959 617941 59025 617944
rect 40378 617646 40384 617710
rect 40448 617708 40454 617710
rect 42831 617708 42897 617711
rect 40448 617706 42897 617708
rect 40448 617650 42836 617706
rect 42892 617650 42897 617706
rect 40448 617648 42897 617650
rect 40448 617646 40454 617648
rect 42831 617645 42897 617648
rect 64578 617416 64638 617944
rect 675898 617942 675904 618006
rect 675968 618004 675974 618006
rect 675968 617944 676320 618004
rect 675968 617942 675974 617944
rect 678159 617708 678225 617711
rect 678159 617706 678270 617708
rect 678159 617650 678164 617706
rect 678220 617650 678270 617706
rect 678159 617645 678270 617650
rect 678210 617456 678270 617645
rect 40762 617202 40768 617266
rect 40832 617264 40838 617266
rect 42735 617264 42801 617267
rect 40832 617262 42801 617264
rect 40832 617206 42740 617262
rect 42796 617206 42801 617262
rect 40832 617204 42801 617206
rect 40832 617202 40838 617204
rect 42735 617201 42801 617204
rect 676239 617116 676305 617119
rect 676239 617114 676350 617116
rect 676239 617058 676244 617114
rect 676300 617058 676350 617114
rect 676239 617053 676350 617058
rect 676290 616938 676350 617053
rect 676047 616524 676113 616527
rect 676047 616522 676320 616524
rect 676047 616466 676052 616522
rect 676108 616466 676320 616522
rect 676047 616464 676320 616466
rect 676047 616461 676113 616464
rect 59631 616228 59697 616231
rect 64578 616228 64638 616234
rect 59631 616226 64638 616228
rect 59631 616170 59636 616226
rect 59692 616170 64638 616226
rect 59631 616168 64638 616170
rect 59631 616165 59697 616168
rect 676047 615932 676113 615935
rect 676047 615930 676320 615932
rect 676047 615874 676052 615930
rect 676108 615874 676320 615930
rect 676047 615872 676320 615874
rect 676047 615869 676113 615872
rect 677050 615722 677056 615786
rect 677120 615722 677126 615786
rect 45903 615636 45969 615639
rect 45903 615634 64638 615636
rect 45903 615578 45908 615634
rect 45964 615578 64638 615634
rect 45903 615576 64638 615578
rect 45903 615573 45969 615576
rect 64578 615052 64638 615576
rect 677058 615458 677118 615722
rect 676239 615192 676305 615195
rect 676239 615190 676350 615192
rect 676239 615134 676244 615190
rect 676300 615134 676350 615190
rect 676239 615129 676350 615134
rect 676290 615014 676350 615129
rect 58959 614452 59025 614455
rect 676047 614452 676113 614455
rect 58959 614450 64638 614452
rect 58959 614394 58964 614450
rect 59020 614394 64638 614450
rect 58959 614392 64638 614394
rect 58959 614389 59025 614392
rect 64578 613870 64638 614392
rect 676047 614450 676320 614452
rect 676047 614394 676052 614450
rect 676108 614394 676320 614450
rect 676047 614392 676320 614394
rect 676047 614389 676113 614392
rect 679938 613715 679998 613904
rect 679938 613710 680049 613715
rect 679938 613654 679988 613710
rect 680044 613654 680049 613710
rect 679938 613652 680049 613654
rect 679983 613649 680049 613652
rect 679746 613271 679806 613534
rect 59631 613268 59697 613271
rect 59631 613266 64638 613268
rect 59631 613210 59636 613266
rect 59692 613210 64638 613266
rect 59631 613208 64638 613210
rect 679746 613266 679857 613271
rect 679983 613268 680049 613271
rect 679746 613210 679796 613266
rect 679852 613210 679857 613266
rect 679746 613208 679857 613210
rect 59631 613205 59697 613208
rect 64578 612688 64638 613208
rect 679791 613205 679857 613208
rect 679938 613266 680049 613268
rect 679938 613210 679988 613266
rect 680044 613210 680049 613266
rect 679938 613205 680049 613210
rect 679938 612942 679998 613205
rect 679791 612824 679857 612827
rect 679746 612822 679857 612824
rect 679746 612766 679796 612822
rect 679852 612766 679857 612822
rect 679746 612761 679857 612766
rect 679746 612424 679806 612761
rect 59535 612084 59601 612087
rect 59535 612082 64638 612084
rect 59535 612026 59540 612082
rect 59596 612026 64638 612082
rect 59535 612024 64638 612026
rect 59535 612021 59601 612024
rect 64578 611506 64638 612024
rect 674170 607730 674176 607794
rect 674240 607792 674246 607794
rect 675183 607792 675249 607795
rect 674240 607790 675249 607792
rect 674240 607734 675188 607790
rect 675244 607734 675249 607790
rect 674240 607732 675249 607734
rect 674240 607730 674246 607732
rect 675183 607729 675249 607732
rect 675183 606018 675249 606019
rect 675130 606016 675136 606018
rect 675092 605956 675136 606016
rect 675200 606014 675249 606018
rect 675244 605958 675249 606014
rect 675130 605954 675136 605956
rect 675200 605954 675249 605958
rect 675183 605953 675249 605954
rect 674554 604770 674560 604834
rect 674624 604832 674630 604834
rect 675279 604832 675345 604835
rect 674624 604830 675345 604832
rect 674624 604774 675284 604830
rect 675340 604774 675345 604830
rect 674624 604772 675345 604774
rect 674624 604770 674630 604772
rect 675279 604769 675345 604772
rect 40335 602168 40401 602171
rect 41722 602168 41728 602170
rect 40335 602166 41728 602168
rect 40335 602110 40340 602166
rect 40396 602110 41728 602166
rect 40335 602108 41728 602110
rect 40335 602105 40401 602108
rect 41722 602106 41728 602108
rect 41792 602168 41798 602170
rect 62319 602168 62385 602171
rect 41792 602166 62385 602168
rect 41792 602110 62324 602166
rect 62380 602110 62385 602166
rect 41792 602108 62385 602110
rect 41792 602106 41798 602108
rect 62319 602105 62385 602108
rect 41775 600540 41841 600543
rect 41568 600538 41841 600540
rect 41568 600482 41780 600538
rect 41836 600482 41841 600538
rect 41568 600480 41841 600482
rect 41775 600477 41841 600480
rect 675471 600246 675537 600247
rect 675471 600242 675520 600246
rect 675584 600244 675590 600246
rect 675471 600186 675476 600242
rect 675471 600182 675520 600186
rect 675584 600184 675628 600244
rect 675584 600182 675590 600184
rect 675471 600181 675537 600182
rect 41538 599803 41598 599918
rect 41538 599798 41649 599803
rect 41538 599742 41588 599798
rect 41644 599742 41649 599798
rect 41538 599740 41649 599742
rect 41583 599737 41649 599740
rect 41775 599430 41841 599433
rect 41568 599428 41841 599430
rect 41568 599372 41780 599428
rect 41836 599372 41841 599428
rect 41568 599370 41841 599372
rect 41775 599367 41841 599370
rect 41775 599060 41841 599063
rect 41568 599058 41841 599060
rect 41568 599002 41780 599058
rect 41836 599002 41841 599058
rect 41568 599000 41841 599002
rect 41775 598997 41841 599000
rect 41538 598323 41598 598438
rect 41538 598318 41649 598323
rect 41538 598262 41588 598318
rect 41644 598262 41649 598318
rect 41538 598260 41649 598262
rect 41583 598257 41649 598260
rect 41914 597950 41920 597952
rect 41568 597890 41920 597950
rect 41914 597888 41920 597890
rect 41984 597888 41990 597952
rect 649986 597876 650046 598336
rect 655215 597876 655281 597879
rect 649986 597874 655281 597876
rect 649986 597818 655220 597874
rect 655276 597818 655281 597874
rect 649986 597816 655281 597818
rect 655215 597813 655281 597816
rect 40335 597728 40401 597731
rect 40335 597726 40446 597728
rect 40335 597670 40340 597726
rect 40396 597670 40446 597726
rect 40335 597665 40446 597670
rect 40386 597550 40446 597665
rect 41722 596988 41728 596990
rect 41568 596928 41728 596988
rect 41722 596926 41728 596928
rect 41792 596926 41798 596990
rect 649986 596692 650046 597154
rect 655407 596692 655473 596695
rect 649986 596690 655473 596692
rect 649986 596634 655412 596690
rect 655468 596634 655473 596690
rect 649986 596632 655473 596634
rect 655407 596629 655473 596632
rect 41538 596251 41598 596366
rect 41538 596246 41649 596251
rect 41538 596190 41588 596246
rect 41644 596190 41649 596246
rect 41538 596188 41649 596190
rect 41583 596185 41649 596188
rect 41538 595807 41598 595996
rect 41487 595802 41598 595807
rect 41487 595746 41492 595802
rect 41548 595746 41598 595802
rect 41487 595744 41598 595746
rect 41487 595741 41553 595744
rect 41775 595508 41841 595511
rect 41568 595506 41841 595508
rect 41568 595450 41780 595506
rect 41836 595450 41841 595506
rect 41568 595448 41841 595450
rect 649986 595508 650046 595972
rect 655599 595508 655665 595511
rect 649986 595506 655665 595508
rect 649986 595450 655604 595506
rect 655660 595450 655665 595506
rect 649986 595448 655665 595450
rect 41775 595445 41841 595448
rect 655599 595445 655665 595448
rect 655119 595360 655185 595363
rect 649986 595358 655185 595360
rect 649986 595302 655124 595358
rect 655180 595302 655185 595358
rect 649986 595300 655185 595302
rect 34434 594771 34494 594886
rect 649986 594790 650046 595300
rect 655119 595297 655185 595300
rect 675759 595360 675825 595363
rect 676282 595360 676288 595362
rect 675759 595358 676288 595360
rect 675759 595302 675764 595358
rect 675820 595302 676288 595358
rect 675759 595300 676288 595302
rect 675759 595297 675825 595300
rect 676282 595298 676288 595300
rect 676352 595298 676358 595362
rect 34383 594766 34494 594771
rect 34383 594710 34388 594766
rect 34444 594710 34494 594766
rect 34383 594708 34494 594710
rect 34383 594705 34449 594708
rect 41538 594324 41598 594516
rect 41679 594324 41745 594327
rect 41538 594322 41745 594324
rect 41538 594266 41684 594322
rect 41740 594266 41745 594322
rect 41538 594264 41745 594266
rect 41679 594261 41745 594264
rect 655791 594176 655857 594179
rect 649986 594174 655857 594176
rect 649986 594118 655796 594174
rect 655852 594118 655857 594174
rect 649986 594116 655857 594118
rect 42159 594028 42225 594031
rect 41568 594026 42225 594028
rect 41568 593970 42164 594026
rect 42220 593970 42225 594026
rect 41568 593968 42225 593970
rect 42159 593965 42225 593968
rect 649986 593608 650046 594116
rect 655791 594113 655857 594116
rect 41775 593436 41841 593439
rect 41568 593434 41841 593436
rect 41568 593378 41780 593434
rect 41836 593378 41841 593434
rect 41568 593376 41841 593378
rect 41775 593373 41841 593376
rect 675759 593436 675825 593439
rect 675898 593436 675904 593438
rect 675759 593434 675904 593436
rect 675759 593378 675764 593434
rect 675820 593378 675904 593434
rect 675759 593376 675904 593378
rect 675759 593373 675825 593376
rect 675898 593374 675904 593376
rect 675968 593374 675974 593438
rect 653775 592992 653841 592995
rect 649986 592990 653841 592992
rect 34434 592847 34494 592962
rect 649986 592934 653780 592990
rect 653836 592934 653841 592990
rect 649986 592932 653841 592934
rect 34434 592842 34545 592847
rect 34434 592786 34484 592842
rect 34540 592786 34545 592842
rect 34434 592784 34545 592786
rect 34479 592781 34545 592784
rect 41967 592548 42033 592551
rect 41568 592546 42033 592548
rect 41568 592490 41972 592546
rect 42028 592490 42033 592546
rect 41568 592488 42033 592490
rect 41967 592485 42033 592488
rect 649986 592426 650046 592932
rect 653775 592929 653841 592932
rect 42063 591956 42129 591959
rect 41568 591954 42129 591956
rect 41568 591898 42068 591954
rect 42124 591898 42129 591954
rect 41568 591896 42129 591898
rect 42063 591893 42129 591896
rect 41538 591367 41598 591482
rect 41538 591362 41649 591367
rect 41538 591306 41588 591362
rect 41644 591306 41649 591362
rect 41538 591304 41649 591306
rect 41583 591301 41649 591304
rect 41871 590994 41937 590997
rect 41568 590992 41937 590994
rect 41568 590936 41876 590992
rect 41932 590936 41937 590992
rect 41568 590934 41937 590936
rect 41871 590931 41937 590934
rect 42351 590476 42417 590479
rect 41568 590474 42417 590476
rect 41568 590418 42356 590474
rect 42412 590418 42417 590474
rect 41568 590416 42417 590418
rect 42351 590413 42417 590416
rect 41538 589887 41598 590002
rect 41538 589882 41649 589887
rect 41538 589826 41588 589882
rect 41644 589826 41649 589882
rect 41538 589824 41649 589826
rect 41583 589821 41649 589824
rect 41538 589295 41598 589484
rect 41538 589290 41649 589295
rect 41538 589234 41588 589290
rect 41644 589234 41649 589290
rect 41538 589232 41649 589234
rect 41583 589229 41649 589232
rect 41568 588936 41790 588996
rect 23106 588259 23166 588522
rect 41730 588404 41790 588936
rect 23055 588254 23166 588259
rect 23055 588198 23060 588254
rect 23116 588198 23166 588254
rect 23055 588196 23166 588198
rect 41538 588344 41790 588404
rect 23055 588193 23121 588196
rect 41538 587815 41598 588344
rect 23055 587812 23121 587815
rect 23055 587810 23166 587812
rect 23055 587754 23060 587810
rect 23116 587754 23166 587810
rect 23055 587749 23166 587754
rect 41538 587810 41649 587815
rect 41538 587754 41588 587810
rect 41644 587754 41649 587810
rect 41538 587752 41649 587754
rect 41583 587749 41649 587752
rect 23106 587486 23166 587749
rect 34383 584852 34449 584855
rect 40570 584852 40576 584854
rect 34383 584850 40576 584852
rect 34383 584794 34388 584850
rect 34444 584794 40576 584850
rect 34383 584792 40576 584794
rect 34383 584789 34449 584792
rect 40570 584790 40576 584792
rect 40640 584790 40646 584854
rect 34479 584704 34545 584707
rect 40378 584704 40384 584706
rect 34479 584702 40384 584704
rect 34479 584646 34484 584702
rect 34540 584646 40384 584702
rect 34479 584644 40384 584646
rect 34479 584641 34545 584644
rect 40378 584642 40384 584644
rect 40448 584642 40454 584706
rect 41967 584704 42033 584707
rect 42106 584704 42112 584706
rect 41967 584702 42112 584704
rect 41967 584646 41972 584702
rect 42028 584646 42112 584702
rect 41967 584644 42112 584646
rect 41967 584641 42033 584644
rect 42106 584642 42112 584644
rect 42176 584642 42182 584706
rect 41487 584558 41553 584559
rect 41487 584556 41536 584558
rect 41444 584554 41536 584556
rect 41444 584498 41492 584554
rect 41444 584496 41536 584498
rect 41487 584494 41536 584496
rect 41600 584494 41606 584558
rect 41679 584556 41745 584559
rect 42298 584556 42304 584558
rect 41679 584554 42304 584556
rect 41679 584498 41684 584554
rect 41740 584498 42304 584554
rect 41679 584496 42304 584498
rect 41487 584493 41553 584494
rect 41679 584493 41745 584496
rect 42298 584494 42304 584496
rect 42368 584494 42374 584558
rect 41338 584198 41344 584262
rect 41408 584260 41414 584262
rect 41871 584260 41937 584263
rect 41408 584258 41937 584260
rect 41408 584202 41876 584258
rect 41932 584202 41937 584258
rect 41408 584200 41937 584202
rect 41408 584198 41414 584200
rect 41871 584197 41937 584200
rect 676290 579823 676350 580086
rect 676290 579818 676401 579823
rect 676290 579762 676340 579818
rect 676396 579762 676401 579818
rect 676290 579760 676401 579762
rect 676335 579757 676401 579760
rect 676143 579376 676209 579379
rect 676290 579376 676350 579494
rect 676143 579374 676350 579376
rect 676143 579318 676148 579374
rect 676204 579318 676350 579374
rect 676143 579316 676350 579318
rect 676143 579313 676209 579316
rect 676239 579228 676305 579231
rect 676239 579226 676350 579228
rect 676239 579170 676244 579226
rect 676300 579170 676350 579226
rect 676239 579165 676350 579170
rect 676290 578976 676350 579165
rect 676239 578784 676305 578787
rect 676239 578782 676350 578784
rect 676239 578726 676244 578782
rect 676300 578726 676350 578782
rect 676239 578721 676350 578726
rect 42298 578574 42304 578638
rect 42368 578636 42374 578638
rect 42831 578636 42897 578639
rect 42368 578634 42897 578636
rect 42368 578578 42836 578634
rect 42892 578578 42897 578634
rect 676290 578606 676350 578721
rect 42368 578576 42897 578578
rect 42368 578574 42374 578576
rect 42831 578573 42897 578576
rect 42063 578194 42129 578195
rect 42063 578192 42112 578194
rect 42020 578190 42112 578192
rect 42020 578134 42068 578190
rect 42020 578132 42112 578134
rect 42063 578130 42112 578132
rect 42176 578130 42182 578194
rect 42063 578129 42129 578130
rect 676290 577899 676350 578014
rect 676239 577894 676350 577899
rect 676239 577838 676244 577894
rect 676300 577838 676350 577894
rect 676239 577836 676350 577838
rect 676239 577833 676305 577836
rect 676047 577526 676113 577529
rect 676047 577524 676320 577526
rect 676047 577468 676052 577524
rect 676108 577468 676320 577524
rect 676047 577466 676320 577468
rect 676047 577463 676113 577466
rect 676047 577156 676113 577159
rect 676047 577154 676320 577156
rect 676047 577098 676052 577154
rect 676108 577098 676320 577154
rect 676047 577096 676320 577098
rect 676047 577093 676113 577096
rect 41530 576798 41536 576862
rect 41600 576860 41606 576862
rect 43023 576860 43089 576863
rect 41600 576858 43089 576860
rect 41600 576802 43028 576858
rect 43084 576802 43089 576858
rect 41600 576800 43089 576802
rect 41600 576798 41606 576800
rect 43023 576797 43089 576800
rect 676047 576564 676113 576567
rect 676047 576562 676320 576564
rect 676047 576506 676052 576562
rect 676108 576506 676320 576562
rect 676047 576504 676320 576506
rect 676047 576501 676113 576504
rect 676047 575972 676113 575975
rect 676047 575970 676320 575972
rect 676047 575914 676052 575970
rect 676108 575914 676320 575970
rect 676047 575912 676320 575914
rect 676047 575909 676113 575912
rect 674746 575762 674752 575826
rect 674816 575824 674822 575826
rect 674816 575764 676350 575824
rect 674816 575762 674822 575764
rect 676290 575572 676350 575764
rect 673978 575022 673984 575086
rect 674048 575084 674054 575086
rect 674048 575024 676320 575084
rect 674048 575022 674054 575024
rect 58959 574788 59025 574791
rect 58959 574786 64638 574788
rect 58959 574730 58964 574786
rect 59020 574730 64638 574786
rect 58959 574728 64638 574730
rect 58959 574725 59025 574728
rect 40570 574430 40576 574494
rect 40640 574492 40646 574494
rect 43119 574492 43185 574495
rect 40640 574490 43185 574492
rect 40640 574434 43124 574490
rect 43180 574434 43185 574490
rect 40640 574432 43185 574434
rect 40640 574430 40646 574432
rect 43119 574429 43185 574432
rect 64578 574194 64638 574728
rect 674938 574430 674944 574494
rect 675008 574492 675014 574494
rect 675008 574432 676320 574492
rect 675008 574430 675014 574432
rect 675322 574282 675328 574346
rect 675392 574344 675398 574346
rect 675392 574284 676350 574344
rect 675392 574282 675398 574284
rect 676290 574092 676350 574284
rect 40378 573986 40384 574050
rect 40448 574048 40454 574050
rect 42927 574048 42993 574051
rect 40448 574046 42993 574048
rect 40448 573990 42932 574046
rect 42988 573990 42993 574046
rect 40448 573988 42993 573990
rect 40448 573986 40454 573988
rect 42927 573985 42993 573988
rect 675706 573542 675712 573606
rect 675776 573604 675782 573606
rect 675776 573544 676320 573604
rect 675776 573542 675782 573544
rect 41338 573394 41344 573458
rect 41408 573456 41414 573458
rect 41775 573456 41841 573459
rect 41408 573454 41841 573456
rect 41408 573398 41780 573454
rect 41836 573398 41841 573454
rect 41408 573396 41841 573398
rect 41408 573394 41414 573396
rect 41775 573393 41841 573396
rect 59631 573012 59697 573015
rect 59631 573010 64638 573012
rect 59631 572954 59636 573010
rect 59692 572954 64638 573010
rect 59631 572952 64638 572954
rect 59631 572949 59697 572952
rect 676090 572802 676096 572866
rect 676160 572864 676166 572866
rect 676290 572864 676350 572982
rect 676160 572804 676350 572864
rect 676160 572802 676166 572804
rect 674362 572506 674368 572570
rect 674432 572568 674438 572570
rect 674432 572508 676320 572568
rect 674432 572506 674438 572508
rect 46191 572420 46257 572423
rect 46191 572418 64638 572420
rect 46191 572362 46196 572418
rect 46252 572362 64638 572418
rect 46191 572360 64638 572362
rect 46191 572357 46257 572360
rect 64578 571830 64638 572360
rect 676239 572272 676305 572275
rect 676239 572270 676350 572272
rect 676239 572214 676244 572270
rect 676300 572214 676350 572270
rect 676239 572209 676350 572214
rect 676290 572094 676350 572209
rect 676047 571532 676113 571535
rect 676047 571530 676320 571532
rect 676047 571474 676052 571530
rect 676108 571474 676320 571530
rect 676047 571472 676320 571474
rect 676047 571469 676113 571472
rect 58959 571236 59025 571239
rect 58959 571234 64638 571236
rect 58959 571178 58964 571234
rect 59020 571178 64638 571234
rect 58959 571176 64638 571178
rect 58959 571173 59025 571176
rect 64578 570648 64638 571176
rect 676047 571088 676113 571091
rect 676047 571086 676320 571088
rect 676047 571030 676052 571086
rect 676108 571030 676320 571086
rect 676047 571028 676320 571030
rect 676047 571025 676113 571028
rect 676047 570570 676113 570573
rect 676047 570568 676320 570570
rect 676047 570512 676052 570568
rect 676108 570512 676320 570568
rect 676047 570510 676320 570512
rect 676047 570507 676113 570510
rect 676239 570200 676305 570203
rect 676239 570198 676350 570200
rect 676239 570142 676244 570198
rect 676300 570142 676350 570198
rect 676239 570137 676350 570142
rect 59343 570052 59409 570055
rect 59343 570050 64638 570052
rect 59343 569994 59348 570050
rect 59404 569994 64638 570050
rect 676290 570022 676350 570137
rect 59343 569992 64638 569994
rect 59343 569989 59409 569992
rect 64578 569466 64638 569992
rect 676047 569608 676113 569611
rect 676047 569606 676320 569608
rect 676047 569550 676052 569606
rect 676108 569550 676320 569606
rect 676047 569548 676320 569550
rect 676047 569545 676113 569548
rect 676047 569090 676113 569093
rect 676047 569088 676320 569090
rect 676047 569032 676052 569088
rect 676108 569032 676320 569088
rect 676047 569030 676320 569032
rect 676047 569027 676113 569030
rect 59535 568868 59601 568871
rect 59535 568866 64638 568868
rect 59535 568810 59540 568866
rect 59596 568810 64638 568866
rect 59535 568808 64638 568810
rect 59535 568805 59601 568808
rect 64578 568284 64638 568808
rect 679983 568720 680049 568723
rect 679938 568718 680049 568720
rect 679938 568662 679988 568718
rect 680044 568662 680049 568718
rect 679938 568657 680049 568662
rect 679938 568542 679998 568657
rect 679746 567835 679806 568098
rect 679746 567830 679857 567835
rect 679983 567832 680049 567835
rect 679746 567774 679796 567830
rect 679852 567774 679857 567830
rect 679746 567772 679857 567774
rect 679791 567769 679857 567772
rect 679938 567830 680049 567832
rect 679938 567774 679988 567830
rect 680044 567774 680049 567830
rect 679938 567769 680049 567774
rect 679938 567506 679998 567769
rect 679791 567388 679857 567391
rect 679746 567386 679857 567388
rect 679746 567330 679796 567386
rect 679852 567330 679857 567386
rect 679746 567325 679857 567330
rect 679746 567062 679806 567325
rect 674938 562886 674944 562950
rect 675008 562948 675014 562950
rect 675183 562948 675249 562951
rect 675008 562946 675249 562948
rect 675008 562890 675188 562946
rect 675244 562890 675249 562946
rect 675008 562888 675249 562890
rect 675008 562886 675014 562888
rect 675183 562885 675249 562888
rect 675322 561702 675328 561766
rect 675392 561764 675398 561766
rect 675471 561764 675537 561767
rect 675392 561762 675537 561764
rect 675392 561706 675476 561762
rect 675532 561706 675537 561762
rect 675392 561704 675537 561706
rect 675392 561702 675398 561704
rect 675471 561701 675537 561704
rect 674362 561406 674368 561470
rect 674432 561468 674438 561470
rect 675375 561468 675441 561471
rect 674432 561466 675441 561468
rect 674432 561410 675380 561466
rect 675436 561410 675441 561466
rect 674432 561408 675441 561410
rect 674432 561406 674438 561408
rect 675375 561405 675441 561408
rect 674746 558890 674752 558954
rect 674816 558952 674822 558954
rect 675471 558952 675537 558955
rect 674816 558950 675537 558952
rect 674816 558894 675476 558950
rect 675532 558894 675537 558950
rect 674816 558892 675537 558894
rect 674816 558890 674822 558892
rect 675471 558889 675537 558892
rect 649986 553328 650046 553914
rect 655119 553328 655185 553331
rect 649986 553326 655185 553328
rect 649986 553270 655124 553326
rect 655180 553270 655185 553326
rect 649986 553268 655185 553270
rect 655119 553265 655185 553268
rect 649986 552144 650046 552732
rect 655311 552144 655377 552147
rect 649986 552142 655377 552144
rect 649986 552086 655316 552142
rect 655372 552086 655377 552142
rect 649986 552084 655377 552086
rect 655311 552081 655377 552084
rect 649986 551108 650046 551550
rect 655503 551108 655569 551111
rect 649986 551106 655569 551108
rect 649986 551050 655508 551106
rect 655564 551050 655569 551106
rect 649986 551048 655569 551050
rect 655503 551045 655569 551048
rect 655695 550960 655761 550963
rect 649986 550958 655761 550960
rect 649986 550902 655700 550958
rect 655756 550902 655761 550958
rect 649986 550900 655761 550902
rect 649986 550368 650046 550900
rect 655695 550897 655761 550900
rect 656559 549776 656625 549779
rect 649986 549774 656625 549776
rect 649986 549718 656564 549774
rect 656620 549718 656625 549774
rect 649986 549716 656625 549718
rect 649986 549186 650046 549716
rect 656559 549713 656625 549716
rect 654159 548592 654225 548595
rect 649986 548590 654225 548592
rect 649986 548534 654164 548590
rect 654220 548534 654225 548590
rect 649986 548532 654225 548534
rect 649986 548004 650046 548532
rect 654159 548529 654225 548532
rect 41914 547198 41920 547262
rect 41984 547260 41990 547262
rect 62511 547260 62577 547263
rect 41984 547258 62577 547260
rect 41984 547202 62516 547258
rect 62572 547202 62577 547258
rect 41984 547200 62577 547202
rect 41984 547198 41990 547200
rect 62511 547197 62577 547200
rect 41722 544386 41728 544450
rect 41792 544448 41798 544450
rect 43023 544448 43089 544451
rect 62703 544448 62769 544451
rect 41792 544446 62769 544448
rect 41792 544390 43028 544446
rect 43084 544390 62708 544446
rect 62764 544390 62769 544446
rect 41792 544388 62769 544390
rect 41792 544386 41798 544388
rect 43023 544385 43089 544388
rect 62703 544385 62769 544388
rect 41538 543119 41598 543234
rect 41538 543114 41649 543119
rect 41538 543058 41588 543114
rect 41644 543058 41649 543114
rect 41538 543056 41649 543058
rect 41583 543053 41649 543056
rect 41775 542746 41841 542749
rect 41568 542744 41841 542746
rect 41568 542688 41780 542744
rect 41836 542688 41841 542744
rect 41568 542686 41841 542688
rect 41775 542683 41841 542686
rect 41775 542228 41841 542231
rect 41568 542226 41841 542228
rect 41568 542170 41780 542226
rect 41836 542170 41841 542226
rect 41568 542168 41841 542170
rect 41775 542165 41841 542168
rect 41775 541784 41841 541787
rect 41568 541782 41841 541784
rect 41568 541726 41780 541782
rect 41836 541726 41841 541782
rect 41568 541724 41841 541726
rect 41775 541721 41841 541724
rect 41538 541192 41598 541236
rect 43503 541192 43569 541195
rect 41538 541190 43569 541192
rect 41538 541134 43508 541190
rect 43564 541134 43569 541190
rect 41538 541132 43569 541134
rect 43503 541129 43569 541132
rect 43407 540748 43473 540751
rect 41568 540746 43473 540748
rect 41568 540690 43412 540746
rect 43468 540690 43473 540746
rect 41568 540688 43473 540690
rect 43407 540685 43473 540688
rect 41914 540304 41920 540306
rect 41568 540244 41920 540304
rect 41914 540242 41920 540244
rect 41984 540242 41990 540306
rect 40578 539566 40638 539682
rect 40570 539502 40576 539566
rect 40640 539502 40646 539566
rect 43023 539268 43089 539271
rect 41568 539266 43089 539268
rect 41568 539210 43028 539266
rect 43084 539210 43089 539266
rect 41568 539208 43089 539210
rect 43023 539205 43089 539208
rect 43119 538824 43185 538827
rect 41568 538822 43185 538824
rect 41568 538766 43124 538822
rect 43180 538766 43185 538822
rect 41568 538764 43185 538766
rect 43119 538761 43185 538764
rect 41775 538232 41841 538235
rect 41568 538230 41841 538232
rect 41568 538174 41780 538230
rect 41836 538174 41841 538230
rect 41568 538172 41841 538174
rect 41775 538169 41841 538172
rect 41538 537640 41598 537684
rect 42298 537640 42304 537642
rect 41538 537580 42304 537640
rect 42298 537578 42304 537580
rect 42368 537578 42374 537642
rect 43023 537344 43089 537347
rect 41568 537342 43089 537344
rect 41568 537286 43028 537342
rect 43084 537286 43089 537342
rect 41568 537284 43089 537286
rect 43023 537281 43089 537284
rect 42735 536752 42801 536755
rect 41568 536750 42801 536752
rect 41568 536694 42740 536750
rect 42796 536694 42801 536750
rect 41568 536692 42801 536694
rect 42735 536689 42801 536692
rect 42927 536604 42993 536607
rect 41538 536602 42993 536604
rect 41538 536546 42932 536602
rect 42988 536546 42993 536602
rect 41538 536544 42993 536546
rect 41538 536204 41598 536544
rect 42927 536541 42993 536544
rect 41775 536310 41841 536311
rect 41722 536246 41728 536310
rect 41792 536308 41841 536310
rect 41792 536306 41884 536308
rect 41836 536250 41884 536306
rect 41792 536248 41884 536250
rect 41792 536246 41841 536248
rect 41775 536245 41841 536246
rect 42106 535864 42112 535866
rect 41568 535804 42112 535864
rect 42106 535802 42112 535804
rect 42176 535802 42182 535866
rect 41538 534978 41598 535242
rect 41967 534978 42033 534979
rect 41530 534914 41536 534978
rect 41600 534914 41606 534978
rect 41914 534976 41920 534978
rect 41876 534916 41920 534976
rect 41984 534974 42033 534978
rect 42028 534918 42033 534974
rect 41914 534914 41920 534916
rect 41984 534914 42033 534918
rect 41967 534913 42033 534914
rect 676143 534976 676209 534979
rect 676290 534976 676350 535242
rect 676143 534974 676350 534976
rect 676143 534918 676148 534974
rect 676204 534918 676350 534974
rect 676143 534916 676350 534918
rect 676143 534913 676209 534916
rect 42831 534680 42897 534683
rect 41568 534678 42897 534680
rect 41568 534622 42836 534678
rect 42892 534622 42897 534678
rect 41568 534620 42897 534622
rect 42831 534617 42897 534620
rect 676290 534387 676350 534724
rect 41722 534384 41728 534386
rect 41538 534324 41728 534384
rect 41538 534280 41598 534324
rect 41722 534322 41728 534324
rect 41792 534322 41798 534386
rect 676239 534382 676350 534387
rect 676239 534326 676244 534382
rect 676300 534326 676350 534382
rect 676239 534324 676350 534326
rect 676239 534321 676305 534324
rect 41775 534234 41841 534239
rect 41775 534178 41780 534234
rect 41836 534178 41841 534234
rect 41775 534173 41841 534178
rect 676047 534236 676113 534239
rect 676047 534234 676320 534236
rect 676047 534178 676052 534234
rect 676108 534178 676320 534234
rect 676047 534176 676320 534178
rect 676047 534173 676113 534176
rect 41778 534088 41838 534173
rect 41538 534028 41838 534088
rect 41538 533762 41598 534028
rect 41775 533942 41841 533943
rect 41722 533940 41728 533942
rect 41684 533880 41728 533940
rect 41792 533938 41841 533942
rect 41836 533882 41841 533938
rect 41722 533878 41728 533880
rect 41792 533878 41841 533882
rect 41775 533877 41841 533878
rect 675951 533792 676017 533795
rect 675951 533790 676320 533792
rect 675951 533734 675956 533790
rect 676012 533734 676320 533790
rect 675951 533732 676320 533734
rect 675951 533729 676017 533732
rect 42735 533200 42801 533203
rect 41568 533198 42801 533200
rect 41568 533142 42740 533198
rect 42796 533142 42801 533198
rect 41568 533140 42801 533142
rect 42735 533137 42801 533140
rect 676674 533055 676734 533170
rect 676674 533050 676785 533055
rect 676674 532994 676724 533050
rect 676780 532994 676785 533050
rect 676674 532992 676785 532994
rect 676719 532989 676785 532992
rect 41722 532830 41728 532832
rect 41568 532770 41728 532830
rect 41722 532768 41728 532770
rect 41792 532768 41798 532832
rect 42298 532694 42304 532758
rect 42368 532756 42374 532758
rect 42927 532756 42993 532759
rect 42368 532754 42993 532756
rect 42368 532698 42932 532754
rect 42988 532698 42993 532754
rect 42368 532696 42993 532698
rect 42368 532694 42374 532696
rect 42927 532693 42993 532696
rect 676047 532756 676113 532759
rect 676047 532754 676320 532756
rect 676047 532698 676052 532754
rect 676108 532698 676320 532754
rect 676047 532696 676320 532698
rect 676047 532693 676113 532696
rect 41914 532312 41920 532314
rect 41568 532252 41920 532312
rect 41914 532250 41920 532252
rect 41984 532250 41990 532314
rect 676674 532019 676734 532282
rect 676623 532014 676734 532019
rect 676623 531958 676628 532014
rect 676684 531958 676734 532014
rect 676623 531956 676734 531958
rect 676623 531953 676689 531956
rect 57711 531720 57777 531723
rect 57711 531718 64638 531720
rect 41346 531537 41406 531690
rect 57711 531662 57716 531718
rect 57772 531662 64638 531718
rect 57711 531660 64638 531662
rect 57711 531657 57777 531660
rect 41338 531473 41344 531537
rect 41408 531473 41414 531537
rect 41538 530980 41598 531246
rect 64578 531172 64638 531660
rect 676290 531575 676350 531690
rect 676239 531570 676350 531575
rect 676239 531514 676244 531570
rect 676300 531514 676350 531570
rect 676239 531512 676350 531514
rect 676239 531509 676305 531512
rect 676482 530983 676542 531246
rect 41538 530920 41790 530980
rect 676482 530978 676593 530983
rect 676482 530922 676532 530978
rect 676588 530922 676593 530978
rect 676482 530920 676593 530922
rect 41346 530433 41406 530802
rect 41730 530536 41790 530920
rect 676527 530917 676593 530920
rect 675130 530770 675136 530834
rect 675200 530832 675206 530834
rect 675200 530772 676320 530832
rect 675200 530770 675206 530772
rect 42106 530622 42112 530686
rect 42176 530684 42182 530686
rect 42831 530684 42897 530687
rect 42176 530682 42897 530684
rect 42176 530626 42836 530682
rect 42892 530626 42897 530682
rect 42176 530624 42897 530626
rect 42176 530622 42182 530624
rect 42831 530621 42897 530624
rect 41538 530476 41790 530536
rect 57615 530536 57681 530539
rect 57615 530534 64638 530536
rect 57615 530478 57620 530534
rect 57676 530478 64638 530534
rect 57615 530476 64638 530478
rect 41338 530369 41344 530433
rect 41408 530369 41414 530433
rect 41538 530210 41598 530476
rect 57615 530473 57681 530476
rect 64578 529990 64638 530476
rect 676282 530474 676288 530538
rect 676352 530474 676358 530538
rect 676290 530210 676350 530474
rect 674170 529882 674176 529946
rect 674240 529944 674246 529946
rect 674240 529884 676350 529944
rect 674240 529882 674246 529884
rect 676290 529692 676350 529884
rect 41530 529586 41536 529650
rect 41600 529648 41606 529650
rect 41775 529648 41841 529651
rect 41600 529646 41841 529648
rect 41600 529590 41780 529646
rect 41836 529590 41841 529646
rect 41600 529588 41841 529590
rect 41600 529586 41606 529588
rect 41775 529585 41841 529588
rect 46671 529352 46737 529355
rect 46671 529350 64638 529352
rect 46671 529294 46676 529350
rect 46732 529294 64638 529350
rect 46671 529292 64638 529294
rect 46671 529289 46737 529292
rect 64578 528808 64638 529292
rect 674554 529290 674560 529354
rect 674624 529352 674630 529354
rect 674624 529292 676320 529352
rect 674624 529290 674630 529292
rect 675514 528698 675520 528762
rect 675584 528760 675590 528762
rect 675584 528700 676320 528760
rect 675584 528698 675590 528700
rect 675898 528106 675904 528170
rect 675968 528168 675974 528170
rect 675968 528108 676320 528168
rect 675968 528106 675974 528108
rect 676239 528020 676305 528023
rect 676239 528018 676350 528020
rect 676239 527962 676244 528018
rect 676300 527962 676350 528018
rect 676239 527957 676350 527962
rect 676290 527842 676350 527957
rect 59631 527576 59697 527579
rect 64578 527576 64638 527626
rect 59631 527574 64638 527576
rect 59631 527518 59636 527574
rect 59692 527518 64638 527574
rect 59631 527516 64638 527518
rect 59631 527513 59697 527516
rect 676239 527428 676305 527431
rect 676239 527426 676350 527428
rect 676239 527370 676244 527426
rect 676300 527370 676350 527426
rect 676239 527365 676350 527370
rect 676290 527250 676350 527365
rect 676047 526688 676113 526691
rect 676047 526686 676320 526688
rect 676047 526630 676052 526686
rect 676108 526630 676320 526686
rect 676047 526628 676320 526630
rect 676047 526625 676113 526628
rect 59343 525948 59409 525951
rect 64578 525948 64638 526444
rect 676047 526318 676113 526321
rect 676047 526316 676320 526318
rect 676047 526260 676052 526316
rect 676108 526260 676320 526316
rect 676047 526258 676320 526260
rect 676047 526255 676113 526258
rect 59343 525946 64638 525948
rect 59343 525890 59348 525946
rect 59404 525890 64638 525946
rect 59343 525888 64638 525890
rect 676239 525948 676305 525951
rect 676239 525946 676350 525948
rect 676239 525890 676244 525946
rect 676300 525890 676350 525946
rect 59343 525885 59409 525888
rect 676239 525885 676350 525890
rect 676290 525770 676350 525885
rect 41338 524998 41344 525062
rect 41408 525060 41414 525062
rect 41679 525060 41745 525063
rect 41408 525058 41745 525060
rect 41408 525002 41684 525058
rect 41740 525002 41745 525058
rect 41408 525000 41745 525002
rect 41408 524998 41414 525000
rect 41679 524997 41745 525000
rect 59631 525060 59697 525063
rect 64578 525060 64638 525262
rect 676047 525208 676113 525211
rect 676047 525206 676320 525208
rect 676047 525150 676052 525206
rect 676108 525150 676320 525206
rect 676047 525148 676320 525150
rect 676047 525145 676113 525148
rect 59631 525058 64638 525060
rect 59631 525002 59636 525058
rect 59692 525002 64638 525058
rect 59631 525000 64638 525002
rect 59631 524997 59697 525000
rect 676047 524838 676113 524841
rect 676047 524836 676320 524838
rect 676047 524780 676052 524836
rect 676108 524780 676320 524836
rect 676047 524778 676320 524780
rect 676047 524775 676113 524778
rect 676239 524468 676305 524471
rect 676239 524466 676350 524468
rect 676239 524410 676244 524466
rect 676300 524410 676350 524466
rect 676239 524405 676350 524410
rect 676290 524290 676350 524405
rect 679746 523583 679806 523698
rect 679746 523578 679857 523583
rect 679746 523522 679796 523578
rect 679852 523522 679857 523578
rect 679746 523520 679857 523522
rect 679791 523517 679857 523520
rect 685506 522991 685566 523254
rect 679791 522988 679857 522991
rect 679746 522986 679857 522988
rect 679746 522930 679796 522986
rect 679852 522930 679857 522986
rect 679746 522925 679857 522930
rect 685455 522986 685566 522991
rect 685455 522930 685460 522986
rect 685516 522930 685566 522986
rect 685455 522928 685566 522930
rect 685455 522925 685521 522928
rect 679746 522810 679806 522925
rect 685455 522544 685521 522547
rect 685455 522542 685566 522544
rect 685455 522486 685460 522542
rect 685516 522486 685566 522542
rect 685455 522481 685566 522486
rect 685506 522218 685566 522481
rect 676143 490576 676209 490579
rect 676290 490576 676350 490842
rect 676143 490574 676350 490576
rect 676143 490518 676148 490574
rect 676204 490518 676350 490574
rect 676143 490516 676350 490518
rect 676143 490513 676209 490516
rect 676290 490135 676350 490324
rect 676290 490130 676401 490135
rect 676290 490074 676340 490130
rect 676396 490074 676401 490130
rect 676290 490072 676401 490074
rect 676335 490069 676401 490072
rect 676239 489984 676305 489987
rect 676239 489982 676350 489984
rect 676239 489926 676244 489982
rect 676300 489926 676350 489982
rect 676239 489921 676350 489926
rect 676290 489806 676350 489921
rect 676674 489247 676734 489362
rect 676674 489242 676785 489247
rect 676674 489186 676724 489242
rect 676780 489186 676785 489242
rect 676674 489184 676785 489186
rect 676719 489181 676785 489184
rect 676674 488655 676734 488770
rect 676674 488650 676785 488655
rect 676674 488594 676724 488650
rect 676780 488594 676785 488650
rect 676674 488592 676785 488594
rect 676719 488589 676785 488592
rect 676047 488356 676113 488359
rect 676047 488354 676320 488356
rect 676047 488298 676052 488354
rect 676108 488298 676320 488354
rect 676047 488296 676320 488298
rect 676047 488293 676113 488296
rect 675279 487912 675345 487915
rect 675279 487910 676320 487912
rect 675279 487854 675284 487910
rect 675340 487854 676320 487910
rect 675279 487852 676320 487854
rect 675279 487849 675345 487852
rect 676290 487175 676350 487290
rect 676239 487170 676350 487175
rect 676239 487114 676244 487170
rect 676300 487114 676350 487170
rect 676239 487112 676350 487114
rect 676239 487109 676305 487112
rect 679746 486583 679806 486846
rect 679695 486578 679806 486583
rect 679695 486522 679700 486578
rect 679756 486522 679806 486578
rect 679695 486520 679806 486522
rect 679695 486517 679761 486520
rect 674362 486370 674368 486434
rect 674432 486432 674438 486434
rect 674432 486372 676320 486432
rect 674432 486370 674438 486372
rect 675951 485840 676017 485843
rect 675951 485838 676320 485840
rect 675951 485782 675956 485838
rect 676012 485782 676320 485838
rect 675951 485780 676320 485782
rect 675951 485777 676017 485780
rect 674938 485630 674944 485694
rect 675008 485692 675014 485694
rect 675008 485632 676350 485692
rect 675008 485630 675014 485632
rect 676290 485292 676350 485632
rect 676239 485100 676305 485103
rect 676239 485098 676350 485100
rect 676239 485042 676244 485098
rect 676300 485042 676350 485098
rect 676239 485037 676350 485042
rect 676290 484922 676350 485037
rect 676047 484360 676113 484363
rect 676047 484358 676320 484360
rect 676047 484302 676052 484358
rect 676108 484302 676320 484358
rect 676047 484300 676320 484302
rect 676047 484297 676113 484300
rect 675951 483768 676017 483771
rect 675951 483766 676320 483768
rect 675951 483710 675956 483766
rect 676012 483710 676320 483766
rect 675951 483708 676320 483710
rect 675951 483705 676017 483708
rect 675322 483410 675328 483474
rect 675392 483472 675398 483474
rect 675392 483412 676320 483472
rect 675392 483410 675398 483412
rect 674746 482818 674752 482882
rect 674816 482880 674822 482882
rect 674816 482820 676320 482880
rect 674816 482818 674822 482820
rect 676047 482288 676113 482291
rect 676047 482286 676320 482288
rect 676047 482230 676052 482286
rect 676108 482230 676320 482286
rect 676047 482228 676320 482230
rect 676047 482225 676113 482228
rect 676047 481918 676113 481921
rect 676047 481916 676320 481918
rect 676047 481860 676052 481916
rect 676108 481860 676320 481916
rect 676047 481858 676320 481860
rect 676047 481855 676113 481858
rect 676239 481548 676305 481551
rect 676239 481546 676350 481548
rect 676239 481490 676244 481546
rect 676300 481490 676350 481546
rect 676239 481485 676350 481490
rect 676290 481370 676350 481485
rect 676047 480808 676113 480811
rect 676047 480806 676320 480808
rect 676047 480750 676052 480806
rect 676108 480750 676320 480806
rect 676047 480748 676320 480750
rect 676047 480745 676113 480748
rect 676047 480438 676113 480441
rect 676047 480436 676320 480438
rect 676047 480380 676052 480436
rect 676108 480380 676320 480436
rect 676047 480378 676320 480380
rect 676047 480375 676113 480378
rect 676239 480068 676305 480071
rect 676239 480066 676350 480068
rect 676239 480010 676244 480066
rect 676300 480010 676350 480066
rect 676239 480005 676350 480010
rect 676290 479890 676350 480005
rect 679938 479183 679998 479298
rect 679887 479178 679998 479183
rect 679887 479122 679892 479178
rect 679948 479122 679998 479178
rect 679887 479120 679998 479122
rect 679887 479117 679953 479120
rect 679746 478591 679806 478854
rect 679695 478586 679806 478591
rect 679695 478530 679700 478586
rect 679756 478530 679806 478586
rect 679695 478528 679806 478530
rect 679887 478588 679953 478591
rect 679887 478586 679998 478588
rect 679887 478530 679892 478586
rect 679948 478530 679998 478586
rect 679695 478525 679761 478528
rect 679887 478525 679998 478530
rect 679938 478410 679998 478525
rect 679695 478144 679761 478147
rect 679695 478142 679806 478144
rect 679695 478086 679700 478142
rect 679756 478086 679806 478142
rect 679695 478081 679806 478086
rect 679746 477818 679806 478081
rect 41538 429307 41598 429422
rect 41538 429302 41649 429307
rect 41538 429246 41588 429302
rect 41644 429246 41649 429302
rect 41538 429244 41649 429246
rect 41583 429241 41649 429244
rect 41775 429008 41841 429011
rect 41568 429006 41841 429008
rect 41568 428950 41780 429006
rect 41836 428950 41841 429006
rect 41568 428948 41841 428950
rect 41775 428945 41841 428948
rect 41775 428416 41841 428419
rect 41568 428414 41841 428416
rect 41568 428358 41780 428414
rect 41836 428358 41841 428414
rect 41568 428356 41841 428358
rect 41775 428353 41841 428356
rect 41775 427972 41841 427975
rect 41568 427970 41841 427972
rect 41568 427914 41780 427970
rect 41836 427914 41841 427970
rect 41568 427912 41841 427914
rect 41775 427909 41841 427912
rect 41775 427454 41841 427457
rect 41568 427452 41841 427454
rect 41568 427396 41780 427452
rect 41836 427396 41841 427452
rect 41568 427394 41841 427396
rect 41775 427391 41841 427394
rect 41775 426936 41841 426939
rect 41568 426934 41841 426936
rect 41568 426878 41780 426934
rect 41836 426878 41841 426934
rect 41568 426876 41841 426878
rect 41775 426873 41841 426876
rect 43503 426492 43569 426495
rect 45231 426492 45297 426495
rect 41568 426490 45297 426492
rect 41568 426434 43508 426490
rect 43564 426434 45236 426490
rect 45292 426434 45297 426490
rect 41568 426432 45297 426434
rect 43503 426429 43569 426432
rect 45231 426429 45297 426432
rect 25794 425607 25854 425944
rect 25794 425602 25905 425607
rect 25794 425546 25844 425602
rect 25900 425546 25905 425602
rect 25794 425544 25905 425546
rect 25839 425541 25905 425544
rect 40378 425542 40384 425606
rect 40448 425542 40454 425606
rect 40386 425456 40446 425542
rect 41775 425456 41841 425459
rect 40386 425454 41841 425456
rect 40386 425426 41780 425454
rect 40416 425398 41780 425426
rect 41836 425398 41841 425454
rect 40416 425396 41841 425398
rect 41775 425393 41841 425396
rect 40578 424718 40638 424982
rect 40570 424654 40576 424718
rect 40640 424654 40646 424718
rect 41722 424420 41728 424422
rect 41568 424360 41728 424420
rect 41722 424358 41728 424360
rect 41792 424358 41798 424422
rect 40770 423682 40830 423946
rect 40762 423618 40768 423682
rect 40832 423618 40838 423682
rect 41346 423238 41406 423502
rect 41338 423174 41344 423238
rect 41408 423174 41414 423238
rect 41914 422940 41920 422942
rect 41568 422880 41920 422940
rect 41914 422878 41920 422880
rect 41984 422878 41990 422942
rect 41538 422200 41598 422392
rect 41679 422200 41745 422203
rect 41538 422198 41745 422200
rect 41538 422142 41684 422198
rect 41740 422142 41745 422198
rect 41538 422140 41745 422142
rect 41679 422137 41745 422140
rect 40962 421758 41022 422022
rect 40954 421694 40960 421758
rect 41024 421694 41030 421758
rect 41538 421166 41598 421430
rect 41530 421102 41536 421166
rect 41600 421102 41606 421166
rect 41154 420722 41214 420912
rect 41146 420658 41152 420722
rect 41216 420658 41222 420722
rect 41538 420279 41598 420542
rect 41538 420274 41649 420279
rect 41538 420218 41588 420274
rect 41644 420218 41649 420274
rect 41538 420216 41649 420218
rect 41583 420213 41649 420216
rect 41775 419980 41841 419983
rect 41568 419978 41841 419980
rect 41568 419922 41780 419978
rect 41836 419922 41841 419978
rect 41568 419920 41841 419922
rect 41775 419917 41841 419920
rect 42106 419388 42112 419390
rect 41568 419328 42112 419388
rect 42106 419326 42112 419328
rect 42176 419326 42182 419390
rect 41775 419018 41841 419021
rect 41568 419016 41841 419018
rect 41568 418960 41780 419016
rect 41836 418960 41841 419016
rect 41568 418958 41841 418960
rect 41775 418955 41841 418958
rect 25839 418796 25905 418799
rect 40378 418796 40384 418798
rect 25839 418794 40384 418796
rect 25839 418738 25844 418794
rect 25900 418738 40384 418794
rect 25839 418736 40384 418738
rect 25839 418733 25905 418736
rect 40378 418734 40384 418736
rect 40448 418734 40454 418798
rect 41775 418500 41841 418503
rect 41568 418498 41841 418500
rect 41568 418442 41780 418498
rect 41836 418442 41841 418498
rect 41568 418440 41841 418442
rect 41775 418437 41841 418440
rect 41538 417760 41598 417878
rect 41538 417700 41790 417760
rect 28866 417171 28926 417508
rect 41730 417316 41790 417700
rect 28815 417166 28926 417171
rect 28815 417110 28820 417166
rect 28876 417110 28926 417166
rect 28815 417108 28926 417110
rect 41538 417256 41790 417316
rect 28815 417105 28881 417108
rect 41538 417020 41598 417256
rect 41775 417020 41841 417023
rect 41538 417018 41841 417020
rect 41538 416990 41780 417018
rect 41568 416962 41780 416990
rect 41836 416962 41841 417018
rect 41568 416960 41841 416962
rect 41775 416957 41841 416960
rect 28815 416724 28881 416727
rect 28815 416722 28926 416724
rect 28815 416666 28820 416722
rect 28876 416666 28926 416722
rect 28815 416661 28926 416666
rect 28866 416398 28926 416661
rect 41722 411186 41728 411250
rect 41792 411248 41798 411250
rect 41871 411248 41937 411251
rect 41792 411246 41937 411248
rect 41792 411190 41876 411246
rect 41932 411190 41937 411246
rect 41792 411188 41937 411190
rect 41792 411186 41798 411188
rect 41871 411185 41937 411188
rect 41871 406070 41937 406071
rect 41871 406066 41920 406070
rect 41984 406068 41990 406070
rect 41871 406010 41876 406066
rect 41871 406006 41920 406010
rect 41984 406008 42028 406068
rect 41984 406006 41990 406008
rect 41871 406005 41937 406006
rect 58479 404144 58545 404147
rect 58479 404142 64638 404144
rect 58479 404086 58484 404142
rect 58540 404086 64638 404142
rect 58479 404084 64638 404086
rect 58479 404081 58545 404084
rect 42063 403850 42129 403851
rect 42063 403846 42112 403850
rect 42176 403848 42182 403850
rect 42063 403790 42068 403846
rect 42063 403786 42112 403790
rect 42176 403788 42220 403848
rect 42176 403786 42182 403788
rect 42063 403785 42129 403786
rect 64578 403550 64638 404084
rect 41146 403046 41152 403110
rect 41216 403108 41222 403110
rect 41775 403108 41841 403111
rect 41216 403106 41841 403108
rect 41216 403050 41780 403106
rect 41836 403050 41841 403106
rect 41216 403048 41841 403050
rect 41216 403046 41222 403048
rect 41775 403045 41841 403048
rect 41530 402602 41536 402666
rect 41600 402664 41606 402666
rect 41775 402664 41841 402667
rect 41600 402662 41841 402664
rect 41600 402606 41780 402662
rect 41836 402606 41841 402662
rect 41600 402604 41841 402606
rect 41600 402602 41606 402604
rect 41775 402601 41841 402604
rect 59343 402368 59409 402371
rect 676143 402368 676209 402371
rect 676290 402368 676350 402634
rect 59343 402366 64638 402368
rect 59343 402310 59348 402366
rect 59404 402310 64638 402366
rect 59343 402308 64638 402310
rect 676143 402366 676350 402368
rect 676143 402310 676148 402366
rect 676204 402310 676350 402366
rect 676143 402308 676350 402310
rect 59343 402305 59409 402308
rect 676143 402305 676209 402308
rect 41338 401862 41344 401926
rect 41408 401924 41414 401926
rect 41775 401924 41841 401927
rect 41408 401922 41841 401924
rect 41408 401866 41780 401922
rect 41836 401866 41841 401922
rect 41408 401864 41841 401866
rect 41408 401862 41414 401864
rect 41775 401861 41841 401864
rect 676290 401779 676350 402116
rect 676239 401774 676350 401779
rect 676239 401718 676244 401774
rect 676300 401718 676350 401774
rect 676239 401716 676350 401718
rect 676239 401713 676305 401716
rect 676047 401628 676113 401631
rect 676047 401626 676320 401628
rect 676047 401570 676052 401626
rect 676108 401570 676320 401626
rect 676047 401568 676320 401570
rect 676047 401565 676113 401568
rect 57711 400592 57777 400595
rect 64578 400592 64638 401186
rect 676674 401039 676734 401154
rect 676674 401034 676785 401039
rect 676674 400978 676724 401034
rect 676780 400978 676785 401034
rect 676674 400976 676785 400978
rect 676719 400973 676785 400976
rect 57711 400590 64638 400592
rect 57711 400534 57716 400590
rect 57772 400534 64638 400590
rect 57711 400532 64638 400534
rect 57711 400529 57777 400532
rect 676290 400447 676350 400636
rect 676239 400442 676350 400447
rect 676239 400386 676244 400442
rect 676300 400386 676350 400442
rect 676239 400384 676350 400386
rect 676239 400381 676305 400384
rect 40570 400086 40576 400150
rect 40640 400148 40646 400150
rect 41775 400148 41841 400151
rect 40640 400146 41841 400148
rect 40640 400090 41780 400146
rect 41836 400090 41841 400146
rect 40640 400088 41841 400090
rect 40640 400086 40646 400088
rect 41775 400085 41841 400088
rect 676047 400148 676113 400151
rect 676047 400146 676320 400148
rect 676047 400090 676052 400146
rect 676108 400090 676320 400146
rect 676047 400088 676320 400090
rect 676047 400085 676113 400088
rect 59631 400000 59697 400003
rect 64578 400000 64638 400004
rect 59631 399998 64638 400000
rect 59631 399942 59636 399998
rect 59692 399942 64638 399998
rect 59631 399940 64638 399942
rect 59631 399937 59697 399940
rect 676047 399704 676113 399707
rect 676047 399702 676320 399704
rect 676047 399646 676052 399702
rect 676108 399646 676320 399702
rect 676047 399644 676320 399646
rect 676047 399641 676113 399644
rect 40954 399494 40960 399558
rect 41024 399556 41030 399558
rect 41775 399556 41841 399559
rect 41024 399554 41841 399556
rect 41024 399498 41780 399554
rect 41836 399498 41841 399554
rect 41024 399496 41841 399498
rect 41024 399494 41030 399496
rect 41775 399493 41841 399496
rect 59727 399408 59793 399411
rect 676623 399408 676689 399411
rect 59727 399406 64638 399408
rect 59727 399350 59732 399406
rect 59788 399350 64638 399406
rect 59727 399348 64638 399350
rect 59727 399345 59793 399348
rect 64578 398822 64638 399348
rect 676623 399406 676734 399408
rect 676623 399350 676628 399406
rect 676684 399350 676734 399406
rect 676623 399345 676734 399350
rect 676674 399082 676734 399345
rect 40762 398754 40768 398818
rect 40832 398816 40838 398818
rect 41775 398816 41841 398819
rect 40832 398814 41841 398816
rect 40832 398758 41780 398814
rect 41836 398758 41841 398814
rect 40832 398756 41841 398758
rect 40832 398754 40838 398756
rect 41775 398753 41841 398756
rect 675951 398668 676017 398671
rect 675951 398666 676320 398668
rect 675951 398610 675956 398666
rect 676012 398610 676320 398666
rect 675951 398608 676320 398610
rect 675951 398605 676017 398608
rect 59535 398224 59601 398227
rect 59535 398222 64638 398224
rect 59535 398166 59540 398222
rect 59596 398166 64638 398222
rect 59535 398164 64638 398166
rect 59535 398161 59601 398164
rect 64578 397640 64638 398164
rect 675898 398162 675904 398226
rect 675968 398224 675974 398226
rect 675968 398164 676320 398224
rect 675968 398162 675974 398164
rect 673978 397570 673984 397634
rect 674048 397632 674054 397634
rect 674048 397572 676320 397632
rect 674048 397570 674054 397572
rect 675130 396830 675136 396894
rect 675200 396892 675206 396894
rect 676290 396892 676350 397084
rect 675200 396832 676350 396892
rect 675200 396830 675206 396832
rect 676674 396450 676734 396714
rect 676666 396386 676672 396450
rect 676736 396386 676742 396450
rect 674938 396090 674944 396154
rect 675008 396152 675014 396154
rect 675008 396092 676320 396152
rect 675008 396090 675014 396092
rect 676047 395634 676113 395637
rect 676047 395632 676320 395634
rect 676047 395576 676052 395632
rect 676108 395576 676320 395632
rect 676047 395574 676320 395576
rect 676047 395571 676113 395574
rect 675706 395202 675712 395266
rect 675776 395264 675782 395266
rect 675776 395204 676320 395264
rect 675776 395202 675782 395204
rect 675322 394610 675328 394674
rect 675392 394672 675398 394674
rect 675392 394612 676320 394672
rect 675392 394610 675398 394612
rect 676482 393934 676542 394050
rect 676474 393870 676480 393934
rect 676544 393870 676550 393934
rect 676290 393342 676350 393680
rect 676282 393278 676288 393342
rect 676352 393278 676358 393342
rect 674362 393130 674368 393194
rect 674432 393192 674438 393194
rect 674432 393132 676320 393192
rect 674432 393130 674438 393132
rect 675514 392538 675520 392602
rect 675584 392600 675590 392602
rect 675584 392540 676320 392600
rect 675584 392538 675590 392540
rect 676090 391798 676096 391862
rect 676160 391860 676166 391862
rect 676290 391860 676350 392200
rect 676160 391800 676350 391860
rect 676160 391798 676166 391800
rect 674170 391650 674176 391714
rect 674240 391712 674246 391714
rect 674240 391652 676320 391712
rect 674240 391650 674246 391652
rect 679746 390975 679806 391090
rect 679746 390970 679857 390975
rect 679746 390914 679796 390970
rect 679852 390914 679857 390970
rect 679746 390912 679857 390914
rect 679791 390909 679857 390912
rect 685506 390383 685566 390646
rect 679791 390380 679857 390383
rect 679746 390378 679857 390380
rect 679746 390322 679796 390378
rect 679852 390322 679857 390378
rect 679746 390317 679857 390322
rect 685455 390378 685566 390383
rect 685455 390322 685460 390378
rect 685516 390322 685566 390378
rect 685455 390320 685566 390322
rect 685455 390317 685521 390320
rect 679746 390202 679806 390317
rect 685455 389936 685521 389939
rect 685455 389934 685566 389936
rect 685455 389878 685460 389934
rect 685516 389878 685566 389934
rect 685455 389873 685566 389878
rect 685506 389610 685566 389873
rect 41775 386532 41841 386535
rect 41568 386530 41841 386532
rect 41568 386474 41780 386530
rect 41836 386474 41841 386530
rect 41568 386472 41841 386474
rect 41775 386469 41841 386472
rect 675183 385942 675249 385943
rect 41538 385795 41598 385910
rect 675130 385878 675136 385942
rect 675200 385940 675249 385942
rect 675200 385938 675292 385940
rect 675244 385882 675292 385938
rect 675200 385880 675292 385882
rect 675200 385878 675249 385880
rect 675183 385877 675249 385878
rect 41538 385790 41649 385795
rect 41538 385734 41588 385790
rect 41644 385734 41649 385790
rect 41538 385732 41649 385734
rect 41583 385729 41649 385732
rect 675759 385646 675825 385647
rect 675706 385582 675712 385646
rect 675776 385644 675825 385646
rect 675776 385642 675868 385644
rect 675820 385586 675868 385642
rect 675776 385584 675868 385586
rect 675776 385582 675825 385584
rect 675759 385581 675825 385582
rect 41775 385422 41841 385425
rect 41568 385420 41841 385422
rect 41568 385364 41780 385420
rect 41836 385364 41841 385420
rect 41568 385362 41841 385364
rect 41775 385359 41841 385362
rect 41583 385200 41649 385203
rect 41538 385198 41649 385200
rect 41538 385142 41588 385198
rect 41644 385142 41649 385198
rect 41538 385137 41649 385142
rect 41538 385022 41598 385137
rect 675759 384904 675825 384907
rect 675898 384904 675904 384906
rect 675759 384902 675904 384904
rect 675759 384846 675764 384902
rect 675820 384846 675904 384902
rect 675759 384844 675904 384846
rect 675759 384841 675825 384844
rect 675898 384842 675904 384844
rect 675968 384842 675974 384906
rect 41775 384460 41841 384463
rect 41568 384458 41841 384460
rect 41568 384402 41780 384458
rect 41836 384402 41841 384458
rect 41568 384400 41841 384402
rect 41775 384397 41841 384400
rect 34434 383723 34494 383838
rect 34434 383718 34545 383723
rect 34434 383662 34484 383718
rect 34540 383662 34545 383718
rect 34434 383660 34545 383662
rect 34479 383657 34545 383660
rect 41775 383498 41841 383501
rect 41568 383496 41841 383498
rect 41568 383440 41780 383496
rect 41836 383440 41841 383496
rect 41568 383438 41841 383440
rect 41775 383435 41841 383438
rect 675759 382980 675825 382983
rect 676666 382980 676672 382982
rect 675759 382978 676672 382980
rect 40194 382687 40254 382950
rect 675759 382922 675764 382978
rect 675820 382922 676672 382978
rect 675759 382920 676672 382922
rect 675759 382917 675825 382920
rect 676666 382918 676672 382920
rect 676736 382918 676742 382982
rect 40194 382682 40305 382687
rect 40194 382626 40244 382682
rect 40300 382626 40305 382682
rect 40194 382624 40305 382626
rect 40239 382621 40305 382624
rect 40378 382622 40384 382686
rect 40448 382622 40454 382686
rect 40386 382388 40446 382622
rect 41722 382388 41728 382390
rect 40386 382358 41728 382388
rect 40416 382328 41728 382358
rect 41722 382326 41728 382328
rect 41792 382326 41798 382390
rect 675322 382326 675328 382390
rect 675392 382388 675398 382390
rect 675471 382388 675537 382391
rect 675392 382386 675537 382388
rect 675392 382330 675476 382386
rect 675532 382330 675537 382386
rect 675392 382328 675537 382330
rect 675392 382326 675398 382328
rect 675471 382325 675537 382328
rect 28674 381651 28734 381988
rect 675759 381796 675825 381799
rect 676474 381796 676480 381798
rect 675759 381794 676480 381796
rect 675759 381738 675764 381794
rect 675820 381738 676480 381794
rect 675759 381736 676480 381738
rect 675759 381733 675825 381736
rect 676474 381734 676480 381736
rect 676544 381734 676550 381798
rect 28674 381646 28785 381651
rect 28674 381590 28724 381646
rect 28780 381590 28785 381646
rect 28674 381588 28785 381590
rect 28719 381585 28785 381588
rect 39810 381206 39870 381470
rect 675567 381206 675633 381207
rect 39802 381142 39808 381206
rect 39872 381142 39878 381206
rect 675514 381142 675520 381206
rect 675584 381204 675633 381206
rect 675584 381202 675676 381204
rect 675628 381146 675676 381202
rect 675584 381144 675676 381146
rect 675584 381142 675633 381144
rect 675567 381141 675633 381142
rect 39426 380763 39486 380878
rect 39375 380758 39486 380763
rect 39375 380702 39380 380758
rect 39436 380702 39486 380758
rect 39375 380700 39486 380702
rect 39375 380697 39441 380700
rect 40002 380318 40062 380434
rect 39994 380254 40000 380318
rect 40064 380254 40070 380318
rect 39810 379727 39870 379990
rect 39279 379724 39345 379727
rect 39234 379722 39345 379724
rect 39234 379666 39284 379722
rect 39340 379666 39345 379722
rect 39234 379661 39345 379666
rect 39810 379722 39921 379727
rect 39810 379666 39860 379722
rect 39916 379666 39921 379722
rect 39810 379664 39921 379666
rect 39855 379661 39921 379664
rect 39234 379398 39294 379661
rect 39810 378839 39870 378954
rect 39759 378834 39870 378839
rect 39759 378778 39764 378834
rect 39820 378778 39870 378834
rect 39759 378776 39870 378778
rect 39759 378773 39825 378776
rect 674938 378774 674944 378838
rect 675008 378836 675014 378838
rect 675471 378836 675537 378839
rect 675008 378834 675537 378836
rect 675008 378778 675476 378834
rect 675532 378778 675537 378834
rect 675008 378776 675537 378778
rect 675008 378774 675014 378776
rect 675471 378773 675537 378776
rect 39426 378247 39486 378436
rect 39426 378242 39537 378247
rect 39426 378186 39476 378242
rect 39532 378186 39537 378242
rect 39426 378184 39537 378186
rect 39471 378181 39537 378184
rect 40570 378034 40576 378098
rect 40640 378034 40646 378098
rect 675759 378096 675825 378099
rect 676090 378096 676096 378098
rect 675759 378094 676096 378096
rect 675759 378038 675764 378094
rect 675820 378038 676096 378094
rect 675759 378036 676096 378038
rect 40578 377918 40638 378034
rect 675759 378033 675825 378036
rect 676090 378034 676096 378036
rect 676160 378034 676166 378098
rect 39618 377211 39678 377474
rect 39618 377206 39729 377211
rect 39618 377150 39668 377206
rect 39724 377150 39729 377206
rect 39618 377148 39729 377150
rect 39663 377145 39729 377148
rect 674362 377146 674368 377210
rect 674432 377208 674438 377210
rect 675375 377208 675441 377211
rect 674432 377206 675441 377208
rect 674432 377150 675380 377206
rect 675436 377150 675441 377206
rect 674432 377148 675441 377150
rect 674432 377146 674438 377148
rect 675375 377145 675441 377148
rect 41775 376986 41841 376989
rect 41568 376984 41841 376986
rect 41568 376928 41780 376984
rect 41836 376928 41841 376984
rect 41568 376926 41841 376928
rect 41775 376923 41841 376926
rect 674170 376702 674176 376766
rect 674240 376764 674246 376766
rect 675471 376764 675537 376767
rect 674240 376762 675537 376764
rect 674240 376706 675476 376762
rect 675532 376706 675537 376762
rect 674240 376704 675537 376706
rect 674240 376702 674246 376704
rect 675471 376701 675537 376704
rect 41914 376468 41920 376470
rect 41568 376408 41920 376468
rect 41914 376406 41920 376408
rect 41984 376406 41990 376470
rect 41775 376024 41841 376027
rect 41568 376022 41841 376024
rect 41568 375966 41780 376022
rect 41836 375966 41841 376022
rect 41568 375964 41841 375966
rect 41775 375961 41841 375964
rect 675759 375728 675825 375731
rect 676282 375728 676288 375730
rect 675759 375726 676288 375728
rect 675759 375670 675764 375726
rect 675820 375670 676288 375726
rect 675759 375668 676288 375670
rect 675759 375665 675825 375668
rect 676282 375666 676288 375668
rect 676352 375666 676358 375730
rect 41538 375287 41598 375402
rect 41538 375282 41649 375287
rect 41538 375226 41588 375282
rect 41644 375226 41649 375282
rect 41538 375224 41649 375226
rect 41583 375221 41649 375224
rect 41538 374692 41598 374958
rect 41538 374632 41790 374692
rect 23106 374251 23166 374514
rect 23055 374246 23166 374251
rect 23055 374190 23060 374246
rect 23116 374190 23166 374246
rect 23055 374188 23166 374190
rect 39759 374248 39825 374251
rect 40762 374248 40768 374250
rect 39759 374246 40768 374248
rect 39759 374190 39764 374246
rect 39820 374190 40768 374246
rect 39759 374188 40768 374190
rect 23055 374185 23121 374188
rect 39759 374185 39825 374188
rect 40762 374186 40768 374188
rect 40832 374186 40838 374250
rect 41730 374248 41790 374632
rect 655503 374396 655569 374399
rect 41538 374188 41790 374248
rect 649986 374394 655569 374396
rect 649986 374338 655508 374394
rect 655564 374338 655569 374394
rect 649986 374336 655569 374338
rect 41538 373952 41598 374188
rect 41871 373952 41937 373955
rect 41538 373950 41937 373952
rect 41538 373922 41876 373950
rect 41568 373894 41876 373922
rect 41932 373894 41937 373950
rect 41568 373892 41937 373894
rect 649986 373892 650046 374336
rect 655503 374333 655569 374336
rect 41871 373889 41937 373892
rect 673978 373890 673984 373954
rect 674048 373952 674054 373954
rect 675471 373952 675537 373955
rect 674048 373950 675537 373952
rect 674048 373894 675476 373950
rect 675532 373894 675537 373950
rect 674048 373892 675537 373894
rect 674048 373890 674054 373892
rect 675471 373889 675537 373892
rect 23055 373804 23121 373807
rect 39855 373804 39921 373807
rect 41530 373804 41536 373806
rect 23055 373802 23166 373804
rect 23055 373746 23060 373802
rect 23116 373746 23166 373802
rect 23055 373741 23166 373746
rect 39855 373802 41536 373804
rect 39855 373746 39860 373802
rect 39916 373746 41536 373802
rect 39855 373744 41536 373746
rect 39855 373741 39921 373744
rect 41530 373742 41536 373744
rect 41600 373742 41606 373806
rect 23106 373404 23166 373741
rect 39994 373594 40000 373658
rect 40064 373656 40070 373658
rect 41338 373656 41344 373658
rect 40064 373596 41344 373656
rect 40064 373594 40070 373596
rect 41338 373594 41344 373596
rect 41408 373594 41414 373658
rect 655119 373360 655185 373363
rect 649986 373358 655185 373360
rect 649986 373302 655124 373358
rect 655180 373302 655185 373358
rect 649986 373300 655185 373302
rect 39471 373212 39537 373215
rect 42106 373212 42112 373214
rect 39471 373210 42112 373212
rect 39471 373154 39476 373210
rect 39532 373154 42112 373210
rect 39471 373152 42112 373154
rect 39471 373149 39537 373152
rect 42106 373150 42112 373152
rect 42176 373150 42182 373214
rect 39375 372768 39441 372771
rect 42298 372768 42304 372770
rect 39375 372766 42304 372768
rect 39375 372710 39380 372766
rect 39436 372710 42304 372766
rect 39375 372708 42304 372710
rect 39375 372705 39441 372708
rect 42298 372706 42304 372708
rect 42368 372706 42374 372770
rect 649986 372710 650046 373300
rect 655119 373297 655185 373300
rect 28719 372472 28785 372475
rect 40954 372472 40960 372474
rect 28719 372470 40960 372472
rect 28719 372414 28724 372470
rect 28780 372414 40960 372470
rect 28719 372412 40960 372414
rect 28719 372409 28785 372412
rect 40954 372410 40960 372412
rect 41024 372410 41030 372474
rect 655311 372176 655377 372179
rect 649986 372174 655377 372176
rect 649986 372118 655316 372174
rect 655372 372118 655377 372174
rect 649986 372116 655377 372118
rect 649986 371528 650046 372116
rect 655311 372113 655377 372116
rect 653775 370992 653841 370995
rect 649986 370990 653841 370992
rect 649986 370934 653780 370990
rect 653836 370934 653841 370990
rect 649986 370932 653841 370934
rect 649986 370346 650046 370932
rect 653775 370929 653841 370932
rect 40378 368118 40384 368182
rect 40448 368180 40454 368182
rect 41775 368180 41841 368183
rect 40448 368178 41841 368180
rect 40448 368122 41780 368178
rect 41836 368122 41841 368178
rect 40448 368120 41841 368122
rect 40448 368118 40454 368120
rect 41775 368117 41841 368120
rect 41530 362790 41536 362854
rect 41600 362852 41606 362854
rect 41775 362852 41841 362855
rect 41600 362850 41841 362852
rect 41600 362794 41780 362850
rect 41836 362794 41841 362850
rect 41600 362792 41841 362794
rect 41600 362790 41606 362792
rect 41775 362789 41841 362792
rect 58479 360928 58545 360931
rect 58479 360926 64638 360928
rect 58479 360870 58484 360926
rect 58540 360870 64638 360926
rect 58479 360868 64638 360870
rect 58479 360865 58545 360868
rect 41967 360634 42033 360635
rect 41914 360632 41920 360634
rect 41876 360572 41920 360632
rect 41984 360630 42033 360634
rect 42028 360574 42033 360630
rect 41914 360570 41920 360572
rect 41984 360570 42033 360574
rect 41967 360569 42033 360570
rect 64578 360328 64638 360868
rect 40570 359830 40576 359894
rect 40640 359892 40646 359894
rect 41775 359892 41841 359895
rect 40640 359890 41841 359892
rect 40640 359834 41780 359890
rect 41836 359834 41841 359890
rect 40640 359832 41841 359834
rect 40640 359830 40646 359832
rect 41775 359829 41841 359832
rect 59151 359744 59217 359747
rect 59151 359742 64638 359744
rect 59151 359686 59156 359742
rect 59212 359686 64638 359742
rect 59151 359684 64638 359686
rect 59151 359681 59217 359684
rect 42063 359302 42129 359303
rect 42063 359298 42112 359302
rect 42176 359300 42182 359302
rect 42063 359242 42068 359298
rect 42063 359238 42112 359242
rect 42176 359240 42220 359300
rect 42176 359238 42182 359240
rect 42063 359237 42129 359238
rect 64578 359146 64638 359684
rect 41338 358794 41344 358858
rect 41408 358856 41414 358858
rect 41775 358856 41841 358859
rect 41408 358854 41841 358856
rect 41408 358798 41780 358854
rect 41836 358798 41841 358854
rect 41408 358796 41841 358798
rect 41408 358794 41414 358796
rect 41775 358793 41841 358796
rect 57711 357524 57777 357527
rect 64578 357524 64638 357964
rect 57711 357522 64638 357524
rect 57711 357466 57716 357522
rect 57772 357466 64638 357522
rect 57711 357464 64638 357466
rect 57711 357461 57777 357464
rect 676290 357231 676350 357494
rect 676239 357226 676350 357231
rect 676239 357170 676244 357226
rect 676300 357170 676350 357226
rect 676239 357168 676350 357170
rect 676239 357165 676305 357168
rect 40954 356870 40960 356934
rect 41024 356932 41030 356934
rect 41871 356932 41937 356935
rect 41024 356930 41937 356932
rect 41024 356874 41876 356930
rect 41932 356874 41937 356930
rect 41024 356872 41937 356874
rect 41024 356870 41030 356872
rect 41871 356869 41937 356872
rect 59631 356784 59697 356787
rect 676143 356784 676209 356787
rect 676290 356784 676350 356902
rect 59631 356782 64638 356784
rect 59631 356726 59636 356782
rect 59692 356726 64638 356782
rect 59631 356724 64638 356726
rect 676143 356782 676350 356784
rect 676143 356726 676148 356782
rect 676204 356726 676350 356782
rect 676143 356724 676350 356726
rect 59631 356721 59697 356724
rect 676143 356721 676209 356724
rect 676047 356414 676113 356417
rect 676047 356412 676320 356414
rect 676047 356356 676052 356412
rect 676108 356356 676320 356412
rect 676047 356354 676320 356356
rect 676047 356351 676113 356354
rect 40762 356130 40768 356194
rect 40832 356192 40838 356194
rect 41775 356192 41841 356195
rect 40832 356190 41841 356192
rect 40832 356134 41780 356190
rect 41836 356134 41841 356190
rect 40832 356132 41841 356134
rect 40832 356130 40838 356132
rect 41775 356129 41841 356132
rect 58383 356192 58449 356195
rect 676239 356192 676305 356195
rect 58383 356190 64638 356192
rect 58383 356134 58388 356190
rect 58444 356134 64638 356190
rect 58383 356132 64638 356134
rect 58383 356129 58449 356132
rect 42159 355748 42225 355751
rect 42298 355748 42304 355750
rect 42159 355746 42304 355748
rect 42159 355690 42164 355746
rect 42220 355690 42304 355746
rect 42159 355688 42304 355690
rect 42159 355685 42225 355688
rect 42298 355686 42304 355688
rect 42368 355686 42374 355750
rect 64578 355600 64638 356132
rect 676239 356190 676350 356192
rect 676239 356134 676244 356190
rect 676300 356134 676350 356190
rect 676239 356129 676350 356134
rect 676290 356014 676350 356129
rect 673978 355390 673984 355454
rect 674048 355452 674054 355454
rect 674048 355392 676320 355452
rect 674048 355390 674054 355392
rect 58479 355008 58545 355011
rect 58479 355006 64638 355008
rect 58479 354950 58484 355006
rect 58540 354950 64638 355006
rect 58479 354948 64638 354950
rect 58479 354945 58545 354948
rect 64578 354418 64638 354948
rect 675951 354860 676017 354863
rect 675951 354858 676320 354860
rect 675951 354802 675956 354858
rect 676012 354802 676320 354858
rect 675951 354800 676320 354802
rect 675951 354797 676017 354800
rect 674170 354502 674176 354566
rect 674240 354564 674246 354566
rect 674240 354504 676320 354564
rect 674240 354502 674246 354504
rect 676047 353972 676113 353975
rect 676047 353970 676320 353972
rect 676047 353914 676052 353970
rect 676108 353914 676320 353970
rect 676047 353912 676320 353914
rect 676047 353909 676113 353912
rect 674362 353318 674368 353382
rect 674432 353380 674438 353382
rect 674432 353320 676320 353380
rect 674432 353318 674438 353320
rect 675706 352948 675712 353012
rect 675776 353010 675782 353012
rect 675776 352950 676320 353010
rect 675776 352948 675782 352950
rect 676866 352199 676926 352462
rect 676866 352194 676977 352199
rect 676866 352138 676916 352194
rect 676972 352138 676977 352194
rect 676866 352136 676977 352138
rect 676911 352133 676977 352136
rect 675567 351900 675633 351903
rect 675567 351898 676320 351900
rect 675567 351842 675572 351898
rect 675628 351842 676320 351898
rect 675567 351840 676320 351842
rect 675567 351837 675633 351840
rect 675898 351394 675904 351458
rect 675968 351456 675974 351458
rect 675968 351396 676320 351456
rect 675968 351394 675974 351396
rect 674554 350950 674560 351014
rect 674624 351012 674630 351014
rect 674624 350952 676320 351012
rect 674624 350950 674630 350952
rect 676866 350275 676926 350390
rect 676815 350270 676926 350275
rect 676815 350214 676820 350270
rect 676876 350214 676926 350270
rect 676815 350212 676926 350214
rect 676815 350209 676881 350212
rect 676290 349831 676350 349946
rect 676239 349826 676350 349831
rect 676239 349770 676244 349826
rect 676300 349770 676350 349826
rect 676239 349768 676350 349770
rect 676239 349765 676305 349768
rect 676047 349532 676113 349535
rect 676047 349530 676320 349532
rect 676047 349474 676052 349530
rect 676108 349474 676320 349530
rect 676047 349472 676320 349474
rect 676047 349469 676113 349472
rect 675951 348940 676017 348943
rect 675951 348938 676320 348940
rect 675951 348882 675956 348938
rect 676012 348882 676320 348938
rect 675951 348880 676320 348882
rect 675951 348877 676017 348880
rect 675514 348434 675520 348498
rect 675584 348496 675590 348498
rect 675584 348436 676320 348496
rect 675584 348434 675590 348436
rect 676047 347978 676113 347981
rect 676047 347976 676320 347978
rect 676047 347920 676052 347976
rect 676108 347920 676320 347976
rect 676047 347918 676320 347920
rect 676047 347915 676113 347918
rect 676047 347460 676113 347463
rect 676047 347458 676320 347460
rect 676047 347402 676052 347458
rect 676108 347402 676320 347458
rect 676047 347400 676320 347402
rect 676047 347397 676113 347400
rect 676290 346871 676350 346986
rect 676239 346866 676350 346871
rect 676239 346810 676244 346866
rect 676300 346810 676350 346866
rect 676239 346808 676350 346810
rect 676239 346805 676305 346808
rect 676143 346276 676209 346279
rect 676290 346276 676350 346394
rect 676143 346274 676350 346276
rect 676143 346218 676148 346274
rect 676204 346218 676350 346274
rect 676143 346216 676350 346218
rect 676143 346213 676209 346216
rect 679746 345687 679806 345950
rect 679695 345682 679806 345687
rect 679695 345626 679700 345682
rect 679756 345626 679806 345682
rect 679695 345624 679806 345626
rect 679695 345621 679761 345624
rect 685506 345243 685566 345506
rect 679695 345240 679761 345243
rect 679695 345238 679806 345240
rect 679695 345182 679700 345238
rect 679756 345182 679806 345238
rect 679695 345177 679806 345182
rect 685455 345238 685566 345243
rect 685455 345182 685460 345238
rect 685516 345182 685566 345238
rect 685455 345180 685566 345182
rect 685455 345177 685521 345180
rect 679746 344914 679806 345177
rect 685455 344796 685521 344799
rect 685455 344794 685566 344796
rect 685455 344738 685460 344794
rect 685516 344738 685566 344794
rect 685455 344733 685566 344738
rect 685506 344470 685566 344733
rect 41538 343319 41598 343434
rect 41538 343314 41649 343319
rect 41538 343258 41588 343314
rect 41644 343258 41649 343314
rect 41538 343256 41649 343258
rect 41583 343253 41649 343256
rect 676474 342958 676480 343022
rect 676544 343020 676550 343022
rect 676815 343020 676881 343023
rect 676544 343018 676881 343020
rect 676544 342962 676820 343018
rect 676876 342962 676881 343018
rect 676544 342960 676881 342962
rect 676544 342958 676550 342960
rect 676815 342957 676881 342960
rect 41775 342946 41841 342949
rect 41568 342944 41841 342946
rect 41568 342888 41780 342944
rect 41836 342888 41841 342944
rect 41568 342886 41841 342888
rect 41775 342883 41841 342886
rect 676666 342810 676672 342874
rect 676736 342872 676742 342874
rect 676911 342872 676977 342875
rect 676736 342870 676977 342872
rect 676736 342814 676916 342870
rect 676972 342814 676977 342870
rect 676736 342812 676977 342814
rect 676736 342810 676742 342812
rect 676911 342809 676977 342812
rect 41775 342428 41841 342431
rect 41568 342426 41841 342428
rect 41568 342370 41780 342426
rect 41836 342370 41841 342426
rect 41568 342368 41841 342370
rect 41775 342365 41841 342368
rect 41775 341984 41841 341987
rect 41568 341982 41841 341984
rect 41568 341926 41780 341982
rect 41836 341926 41841 341982
rect 41568 341924 41841 341926
rect 41775 341921 41841 341924
rect 41775 341466 41841 341469
rect 41568 341464 41841 341466
rect 41568 341408 41780 341464
rect 41836 341408 41841 341464
rect 41568 341406 41841 341408
rect 41775 341403 41841 341406
rect 41775 340948 41841 340951
rect 41568 340946 41841 340948
rect 41568 340890 41780 340946
rect 41836 340890 41841 340946
rect 41568 340888 41841 340890
rect 41775 340885 41841 340888
rect 41775 340504 41841 340507
rect 41568 340502 41841 340504
rect 41568 340446 41780 340502
rect 41836 340446 41841 340502
rect 41568 340444 41841 340446
rect 41775 340441 41841 340444
rect 41775 339912 41841 339915
rect 41568 339910 41841 339912
rect 41568 339854 41780 339910
rect 41836 339854 41841 339910
rect 41568 339852 41841 339854
rect 41775 339849 41841 339852
rect 41583 339764 41649 339767
rect 41538 339762 41649 339764
rect 41538 339706 41588 339762
rect 41644 339706 41649 339762
rect 41538 339701 41649 339706
rect 41538 339438 41598 339701
rect 675759 339618 675825 339619
rect 675706 339616 675712 339618
rect 675668 339556 675712 339616
rect 675776 339614 675825 339618
rect 675820 339558 675825 339614
rect 675706 339554 675712 339556
rect 675776 339554 675825 339558
rect 675759 339553 675825 339554
rect 28674 338731 28734 338994
rect 28674 338726 28785 338731
rect 28674 338670 28724 338726
rect 28780 338670 28785 338726
rect 28674 338668 28785 338670
rect 28719 338665 28785 338668
rect 39810 338286 39870 338402
rect 39802 338222 39808 338286
rect 39872 338222 39878 338286
rect 39234 337695 39294 337884
rect 675759 337840 675825 337843
rect 675898 337840 675904 337842
rect 675759 337838 675904 337840
rect 675759 337782 675764 337838
rect 675820 337782 675904 337838
rect 675759 337780 675904 337782
rect 675759 337777 675825 337780
rect 675898 337778 675904 337780
rect 675968 337778 675974 337842
rect 39234 337690 39345 337695
rect 39234 337634 39284 337690
rect 39340 337634 39345 337690
rect 39234 337632 39345 337634
rect 39279 337629 39345 337632
rect 40386 337250 40446 337514
rect 40378 337186 40384 337250
rect 40448 337186 40454 337250
rect 40578 336806 40638 336922
rect 40570 336742 40576 336806
rect 40640 336742 40646 336806
rect 41538 336212 41598 336404
rect 41679 336212 41745 336215
rect 41538 336210 41745 336212
rect 41538 336154 41684 336210
rect 41740 336154 41745 336210
rect 41538 336152 41745 336154
rect 41679 336149 41745 336152
rect 40962 335770 41022 336034
rect 40954 335706 40960 335770
rect 41024 335706 41030 335770
rect 41154 335178 41214 335442
rect 41146 335114 41152 335178
rect 41216 335114 41222 335178
rect 41914 334880 41920 334882
rect 41568 334820 41920 334880
rect 41914 334818 41920 334820
rect 41984 334818 41990 334882
rect 41538 334143 41598 334480
rect 41538 334138 41649 334143
rect 41538 334082 41588 334138
rect 41644 334082 41649 334138
rect 41538 334080 41649 334082
rect 41583 334077 41649 334080
rect 41775 333992 41841 333995
rect 41568 333990 41841 333992
rect 41568 333934 41780 333990
rect 41836 333934 41841 333990
rect 41568 333932 41841 333934
rect 41775 333929 41841 333932
rect 674554 333486 674560 333550
rect 674624 333548 674630 333550
rect 675375 333548 675441 333551
rect 674624 333546 675441 333548
rect 674624 333490 675380 333546
rect 675436 333490 675441 333546
rect 674624 333488 675441 333490
rect 674624 333486 674630 333488
rect 675375 333485 675441 333488
rect 42106 333400 42112 333402
rect 41568 333340 42112 333400
rect 42106 333338 42112 333340
rect 42176 333338 42182 333402
rect 41538 332660 41598 333000
rect 42490 332660 42496 332662
rect 41538 332600 42496 332660
rect 42490 332598 42496 332600
rect 42560 332598 42566 332662
rect 41775 332512 41841 332515
rect 41568 332510 41841 332512
rect 41568 332454 41780 332510
rect 41836 332454 41841 332510
rect 41568 332452 41841 332454
rect 41775 332449 41841 332452
rect 41538 331772 41598 331890
rect 41538 331712 41790 331772
rect 23106 331183 23166 331446
rect 41730 331328 41790 331712
rect 41538 331268 41790 331328
rect 23055 331178 23166 331183
rect 23055 331122 23060 331178
rect 23116 331122 23166 331178
rect 23055 331120 23166 331122
rect 39279 331180 39345 331183
rect 40762 331180 40768 331182
rect 39279 331178 40768 331180
rect 39279 331122 39284 331178
rect 39340 331122 40768 331178
rect 39279 331120 40768 331122
rect 23055 331117 23121 331120
rect 39279 331117 39345 331120
rect 40762 331118 40768 331120
rect 40832 331118 40838 331182
rect 41538 331032 41598 331268
rect 41871 331032 41937 331035
rect 41538 331030 41937 331032
rect 41538 331002 41876 331030
rect 41568 330974 41876 331002
rect 41932 330974 41937 331030
rect 41568 330972 41937 330974
rect 41871 330969 41937 330972
rect 23055 330736 23121 330739
rect 23055 330734 23166 330736
rect 23055 330678 23060 330734
rect 23116 330678 23166 330734
rect 23055 330673 23166 330678
rect 39802 330674 39808 330738
rect 39872 330736 39878 330738
rect 41530 330736 41536 330738
rect 39872 330676 41536 330736
rect 39872 330674 39878 330676
rect 41530 330674 41536 330676
rect 41600 330674 41606 330738
rect 23106 330410 23166 330673
rect 675567 330590 675633 330591
rect 675514 330526 675520 330590
rect 675584 330588 675633 330590
rect 675584 330586 675676 330588
rect 675628 330530 675676 330586
rect 675584 330528 675676 330530
rect 675584 330526 675633 330528
rect 675567 330525 675633 330526
rect 655215 329848 655281 329851
rect 649986 329846 655281 329848
rect 649986 329790 655220 329846
rect 655276 329790 655281 329846
rect 649986 329788 655281 329790
rect 28719 329256 28785 329259
rect 42298 329256 42304 329258
rect 28719 329254 42304 329256
rect 28719 329198 28724 329254
rect 28780 329198 42304 329254
rect 28719 329196 42304 329198
rect 28719 329193 28785 329196
rect 42298 329194 42304 329196
rect 42368 329194 42374 329258
rect 649986 329234 650046 329788
rect 655215 329785 655281 329788
rect 40378 328306 40384 328370
rect 40448 328368 40454 328370
rect 41338 328368 41344 328370
rect 40448 328308 41344 328368
rect 40448 328306 40454 328308
rect 41338 328306 41344 328308
rect 41408 328306 41414 328370
rect 655119 328072 655185 328075
rect 649986 328070 655185 328072
rect 649986 328014 655124 328070
rect 655180 328014 655185 328070
rect 649986 328012 655185 328014
rect 655119 328009 655185 328012
rect 675759 328072 675825 328075
rect 676666 328072 676672 328074
rect 675759 328070 676672 328072
rect 675759 328014 675764 328070
rect 675820 328014 676672 328070
rect 675759 328012 676672 328014
rect 675759 328009 675825 328012
rect 676666 328010 676672 328012
rect 676736 328010 676742 328074
rect 655311 327480 655377 327483
rect 649986 327478 655377 327480
rect 649986 327422 655316 327478
rect 655372 327422 655377 327478
rect 649986 327420 655377 327422
rect 649986 326870 650046 327420
rect 655311 327417 655377 327420
rect 675759 326888 675825 326891
rect 676474 326888 676480 326890
rect 675759 326886 676480 326888
rect 675759 326830 675764 326886
rect 675820 326830 676480 326886
rect 675759 326828 676480 326830
rect 675759 326825 675825 326828
rect 676474 326826 676480 326828
rect 676544 326826 676550 326890
rect 654159 326296 654225 326299
rect 649986 326294 654225 326296
rect 649986 326238 654164 326294
rect 654220 326238 654225 326294
rect 649986 326236 654225 326238
rect 649986 325688 650046 326236
rect 654159 326233 654225 326236
rect 41530 324902 41536 324966
rect 41600 324964 41606 324966
rect 41775 324964 41841 324967
rect 41600 324962 41841 324964
rect 41600 324906 41780 324962
rect 41836 324906 41841 324962
rect 41600 324904 41841 324906
rect 41600 324902 41606 324904
rect 41775 324901 41841 324904
rect 42159 320524 42225 320527
rect 42490 320524 42496 320526
rect 42159 320522 42496 320524
rect 42159 320466 42164 320522
rect 42220 320466 42496 320522
rect 42159 320464 42496 320466
rect 42159 320461 42225 320464
rect 42490 320462 42496 320464
rect 42560 320462 42566 320526
rect 40570 319722 40576 319786
rect 40640 319784 40646 319786
rect 41775 319784 41841 319787
rect 40640 319782 41841 319784
rect 40640 319726 41780 319782
rect 41836 319726 41841 319782
rect 40640 319724 41841 319726
rect 40640 319722 40646 319724
rect 41775 319721 41841 319724
rect 58479 317712 58545 317715
rect 58479 317710 64638 317712
rect 58479 317654 58484 317710
rect 58540 317654 64638 317710
rect 58479 317652 64638 317654
rect 58479 317649 58545 317652
rect 42159 317418 42225 317419
rect 42106 317416 42112 317418
rect 42068 317356 42112 317416
rect 42176 317414 42225 317418
rect 42220 317358 42225 317414
rect 42106 317354 42112 317356
rect 42176 317354 42225 317358
rect 42159 317353 42225 317354
rect 64578 317106 64638 317652
rect 41871 316826 41937 316827
rect 41871 316822 41920 316826
rect 41984 316824 41990 316826
rect 41871 316766 41876 316822
rect 41871 316762 41920 316766
rect 41984 316764 42028 316824
rect 41984 316762 41990 316764
rect 41871 316761 41937 316762
rect 59151 316528 59217 316531
rect 59151 316526 64638 316528
rect 59151 316470 59156 316526
rect 59212 316470 64638 316526
rect 59151 316468 64638 316470
rect 59151 316465 59217 316468
rect 41146 316022 41152 316086
rect 41216 316084 41222 316086
rect 41775 316084 41841 316087
rect 41216 316082 41841 316084
rect 41216 316026 41780 316082
rect 41836 316026 41841 316082
rect 41216 316024 41841 316026
rect 41216 316022 41222 316024
rect 41775 316021 41841 316024
rect 64578 315924 64638 316468
rect 41338 315578 41344 315642
rect 41408 315640 41414 315642
rect 41775 315640 41841 315643
rect 41408 315638 41841 315640
rect 41408 315582 41780 315638
rect 41836 315582 41841 315638
rect 41408 315580 41841 315582
rect 41408 315578 41414 315580
rect 41775 315577 41841 315580
rect 59055 314160 59121 314163
rect 64578 314160 64638 314742
rect 59055 314158 64638 314160
rect 59055 314102 59060 314158
rect 59116 314102 64638 314158
rect 59055 314100 64638 314102
rect 59055 314097 59121 314100
rect 42063 313716 42129 313719
rect 42298 313716 42304 313718
rect 42063 313714 42304 313716
rect 42063 313658 42068 313714
rect 42124 313658 42304 313714
rect 42063 313656 42304 313658
rect 42063 313653 42129 313656
rect 42298 313654 42304 313656
rect 42368 313654 42374 313718
rect 59631 313568 59697 313571
rect 59631 313566 64638 313568
rect 59631 313510 59636 313566
rect 59692 313510 64638 313566
rect 59631 313508 64638 313510
rect 59631 313505 59697 313508
rect 40954 313062 40960 313126
rect 41024 313124 41030 313126
rect 41775 313124 41841 313127
rect 41024 313122 41841 313124
rect 41024 313066 41780 313122
rect 41836 313066 41841 313122
rect 41024 313064 41841 313066
rect 41024 313062 41030 313064
rect 41775 313061 41841 313064
rect 59727 312976 59793 312979
rect 59727 312974 64638 312976
rect 59727 312918 59732 312974
rect 59788 312918 64638 312974
rect 59727 312916 64638 312918
rect 59727 312913 59793 312916
rect 40762 312322 40768 312386
rect 40832 312384 40838 312386
rect 41775 312384 41841 312387
rect 40832 312382 41841 312384
rect 40832 312326 41780 312382
rect 41836 312326 41841 312382
rect 64578 312378 64638 312916
rect 40832 312324 41841 312326
rect 40832 312322 40838 312324
rect 41775 312321 41841 312324
rect 676290 312239 676350 312502
rect 676290 312234 676401 312239
rect 676290 312178 676340 312234
rect 676396 312178 676401 312234
rect 676290 312176 676401 312178
rect 676335 312173 676401 312176
rect 59535 311792 59601 311795
rect 59535 311790 64638 311792
rect 59535 311734 59540 311790
rect 59596 311734 64638 311790
rect 59535 311732 64638 311734
rect 59535 311729 59601 311732
rect 64578 311196 64638 311732
rect 676143 311644 676209 311647
rect 676290 311644 676350 311910
rect 676143 311642 676350 311644
rect 676143 311586 676148 311642
rect 676204 311586 676350 311642
rect 676143 311584 676350 311586
rect 676143 311581 676209 311584
rect 676290 311203 676350 311392
rect 676239 311198 676350 311203
rect 676239 311142 676244 311198
rect 676300 311142 676350 311198
rect 676239 311140 676350 311142
rect 676239 311137 676305 311140
rect 673978 310990 673984 311054
rect 674048 311052 674054 311054
rect 674048 310992 676320 311052
rect 674048 310990 674054 310992
rect 675322 310398 675328 310462
rect 675392 310460 675398 310462
rect 675392 310400 676320 310460
rect 675392 310398 675398 310400
rect 674170 309806 674176 309870
rect 674240 309868 674246 309870
rect 674240 309808 676320 309868
rect 674240 309806 674246 309808
rect 675130 309066 675136 309130
rect 675200 309128 675206 309130
rect 676290 309128 676350 309468
rect 675200 309068 676350 309128
rect 675200 309066 675206 309068
rect 670479 308980 670545 308983
rect 674362 308980 674368 308982
rect 670479 308978 674368 308980
rect 670479 308922 670484 308978
rect 670540 308922 674368 308978
rect 670479 308920 674368 308922
rect 670479 308917 670545 308920
rect 674362 308918 674368 308920
rect 674432 308980 674438 308982
rect 674432 308920 676320 308980
rect 674432 308918 674438 308920
rect 675514 308326 675520 308390
rect 675584 308388 675590 308390
rect 675584 308328 676320 308388
rect 675584 308326 675590 308328
rect 676047 308018 676113 308021
rect 676047 308016 676320 308018
rect 676047 307960 676052 308016
rect 676108 307960 676320 308016
rect 676047 307958 676320 307960
rect 676047 307955 676113 307958
rect 674554 307438 674560 307502
rect 674624 307500 674630 307502
rect 674624 307440 676320 307500
rect 674624 307438 674630 307440
rect 676290 306763 676350 306878
rect 676239 306758 676350 306763
rect 676239 306702 676244 306758
rect 676300 306702 676350 306758
rect 676239 306700 676350 306702
rect 676239 306697 676305 306700
rect 673978 306402 673984 306466
rect 674048 306464 674054 306466
rect 674048 306404 676320 306464
rect 674048 306402 674054 306404
rect 674746 305958 674752 306022
rect 674816 306020 674822 306022
rect 674816 305960 676320 306020
rect 674816 305958 674822 305960
rect 676911 305724 676977 305727
rect 676866 305722 676977 305724
rect 676866 305666 676916 305722
rect 676972 305666 676977 305722
rect 676866 305661 676977 305666
rect 676866 305398 676926 305661
rect 676290 304839 676350 304954
rect 676239 304834 676350 304839
rect 676239 304778 676244 304834
rect 676300 304778 676350 304834
rect 676239 304776 676350 304778
rect 676239 304773 676305 304776
rect 676047 304466 676113 304469
rect 676047 304464 676320 304466
rect 676047 304408 676052 304464
rect 676108 304408 676320 304464
rect 676047 304406 676320 304408
rect 676047 304403 676113 304406
rect 675951 303948 676017 303951
rect 675951 303946 676320 303948
rect 675951 303890 675956 303946
rect 676012 303890 676320 303946
rect 675951 303888 676320 303890
rect 675951 303885 676017 303888
rect 676866 303359 676926 303474
rect 654159 303356 654225 303359
rect 649986 303354 654225 303356
rect 649986 303298 654164 303354
rect 654220 303298 654225 303354
rect 649986 303296 654225 303298
rect 649986 302776 650046 303296
rect 654159 303293 654225 303296
rect 676815 303354 676926 303359
rect 676815 303298 676820 303354
rect 676876 303298 676926 303354
rect 676815 303296 676926 303298
rect 676815 303293 676881 303296
rect 674938 302554 674944 302618
rect 675008 302616 675014 302618
rect 676290 302616 676350 302956
rect 675008 302556 676350 302616
rect 675008 302554 675014 302556
rect 676047 302468 676113 302471
rect 676047 302466 676320 302468
rect 676047 302410 676052 302466
rect 676108 302410 676320 302466
rect 676047 302408 676320 302410
rect 676047 302405 676113 302408
rect 654063 302172 654129 302175
rect 649986 302170 654129 302172
rect 649986 302114 654068 302170
rect 654124 302114 654129 302170
rect 649986 302112 654129 302114
rect 649986 301594 650046 302112
rect 654063 302109 654129 302112
rect 676047 302024 676113 302027
rect 676047 302022 676320 302024
rect 676047 301966 676052 302022
rect 676108 301966 676320 302022
rect 676047 301964 676320 301966
rect 676047 301961 676113 301964
rect 676290 301287 676350 301402
rect 676239 301282 676350 301287
rect 676239 301226 676244 301282
rect 676300 301226 676350 301282
rect 676239 301224 676350 301226
rect 676239 301221 676305 301224
rect 654255 300988 654321 300991
rect 649986 300986 654321 300988
rect 649986 300930 654260 300986
rect 654316 300930 654321 300986
rect 649986 300928 654321 300930
rect 649986 300412 650046 300928
rect 654255 300925 654321 300928
rect 679938 300695 679998 300958
rect 679938 300690 680049 300695
rect 679938 300634 679988 300690
rect 680044 300634 680049 300690
rect 679938 300632 680049 300634
rect 679983 300629 680049 300632
rect 679746 300251 679806 300514
rect 679746 300246 679857 300251
rect 679983 300248 680049 300251
rect 41538 299955 41598 300218
rect 679746 300190 679796 300246
rect 679852 300190 679857 300246
rect 679746 300188 679857 300190
rect 679791 300185 679857 300188
rect 679938 300246 680049 300248
rect 679938 300190 679988 300246
rect 680044 300190 680049 300246
rect 679938 300185 680049 300190
rect 41538 299950 41649 299955
rect 41538 299894 41588 299950
rect 41644 299894 41649 299950
rect 679938 299922 679998 300185
rect 41538 299892 41649 299894
rect 41583 299889 41649 299892
rect 41775 299804 41841 299807
rect 679791 299804 679857 299807
rect 41568 299802 41841 299804
rect 41568 299746 41780 299802
rect 41836 299746 41841 299802
rect 41568 299744 41841 299746
rect 41775 299741 41841 299744
rect 679746 299802 679857 299804
rect 679746 299746 679796 299802
rect 679852 299746 679857 299802
rect 679746 299741 679857 299746
rect 39663 299508 39729 299511
rect 39618 299506 39729 299508
rect 39618 299450 39668 299506
rect 39724 299450 39729 299506
rect 39618 299445 39729 299450
rect 39618 299182 39678 299445
rect 679746 299404 679806 299741
rect 41775 298768 41841 298771
rect 41568 298766 41841 298768
rect 41568 298710 41780 298766
rect 41836 298710 41841 298766
rect 41568 298708 41841 298710
rect 649986 298768 650046 299230
rect 675706 299150 675712 299214
rect 675776 299212 675782 299214
rect 676815 299212 676881 299215
rect 675776 299210 676881 299212
rect 675776 299154 676820 299210
rect 676876 299154 676881 299210
rect 675776 299152 676881 299154
rect 675776 299150 675782 299152
rect 676815 299149 676881 299152
rect 654159 298768 654225 298771
rect 649986 298766 654225 298768
rect 649986 298710 654164 298766
rect 654220 298710 654225 298766
rect 649986 298708 654225 298710
rect 41775 298705 41841 298708
rect 654159 298705 654225 298708
rect 676666 298706 676672 298770
rect 676736 298768 676742 298770
rect 676911 298768 676977 298771
rect 676736 298766 676977 298768
rect 676736 298710 676916 298766
rect 676972 298710 676977 298766
rect 676736 298708 676977 298710
rect 676736 298706 676742 298708
rect 676911 298705 676977 298708
rect 41775 298250 41841 298253
rect 41568 298248 41841 298250
rect 41568 298192 41780 298248
rect 41836 298192 41841 298248
rect 41568 298190 41841 298192
rect 41775 298187 41841 298190
rect 41775 297732 41841 297735
rect 41568 297730 41841 297732
rect 41568 297674 41780 297730
rect 41836 297674 41841 297730
rect 41568 297672 41841 297674
rect 41775 297669 41841 297672
rect 649986 297584 650046 298048
rect 656463 297584 656529 297587
rect 649986 297582 656529 297584
rect 649986 297526 656468 297582
rect 656524 297526 656529 297582
rect 649986 297524 656529 297526
rect 656463 297521 656529 297524
rect 41871 297288 41937 297291
rect 41568 297286 41937 297288
rect 41568 297230 41876 297286
rect 41932 297230 41937 297286
rect 41568 297228 41937 297230
rect 41871 297225 41937 297228
rect 649986 296844 650046 296866
rect 656079 296844 656145 296847
rect 649986 296842 656145 296844
rect 649986 296786 656084 296842
rect 656140 296786 656145 296842
rect 649986 296784 656145 296786
rect 656079 296781 656145 296784
rect 41775 296770 41841 296773
rect 41568 296768 41841 296770
rect 41568 296712 41780 296768
rect 41836 296712 41841 296768
rect 41568 296710 41841 296712
rect 41775 296707 41841 296710
rect 654159 296696 654225 296699
rect 675375 296696 675441 296699
rect 654159 296694 675441 296696
rect 654159 296638 654164 296694
rect 654220 296638 675380 296694
rect 675436 296638 675441 296694
rect 654159 296636 675441 296638
rect 654159 296633 654225 296636
rect 675375 296633 675441 296636
rect 39855 296548 39921 296551
rect 39810 296546 39921 296548
rect 39810 296490 39860 296546
rect 39916 296490 39921 296546
rect 39810 296485 39921 296490
rect 39810 296222 39870 296485
rect 28674 295515 28734 295778
rect 28674 295510 28785 295515
rect 28674 295454 28724 295510
rect 28780 295454 28785 295510
rect 28674 295452 28785 295454
rect 28719 295449 28785 295452
rect 59247 295216 59313 295219
rect 64578 295216 64638 295684
rect 59247 295214 64638 295216
rect 41538 294922 41598 295186
rect 59247 295158 59252 295214
rect 59308 295158 64638 295214
rect 59247 295156 64638 295158
rect 649986 295216 650046 295684
rect 656559 295216 656625 295219
rect 649986 295214 656625 295216
rect 649986 295158 656564 295214
rect 656620 295158 656625 295214
rect 649986 295156 656625 295158
rect 59247 295153 59313 295156
rect 656559 295153 656625 295156
rect 41530 294858 41536 294922
rect 41600 294858 41606 294922
rect 42298 294772 42304 294774
rect 41568 294712 42304 294772
rect 42298 294710 42304 294712
rect 42368 294710 42374 294774
rect 40386 294034 40446 294298
rect 40378 293970 40384 294034
rect 40448 293970 40454 294034
rect 60303 294032 60369 294035
rect 64578 294032 64638 294502
rect 60303 294030 64638 294032
rect 60303 293974 60308 294030
rect 60364 293974 64638 294030
rect 60303 293972 64638 293974
rect 649986 294032 650046 294502
rect 655887 294032 655953 294035
rect 649986 294030 655953 294032
rect 649986 293974 655892 294030
rect 655948 293974 655953 294030
rect 649986 293972 655953 293974
rect 60303 293969 60369 293972
rect 655887 293969 655953 293972
rect 41914 293736 41920 293738
rect 41568 293676 41920 293736
rect 41914 293674 41920 293676
rect 41984 293674 41990 293738
rect 41538 292996 41598 293188
rect 41679 292996 41745 292999
rect 41538 292994 41745 292996
rect 41538 292938 41684 292994
rect 41740 292938 41745 292994
rect 41538 292936 41745 292938
rect 41679 292933 41745 292936
rect 59631 292848 59697 292851
rect 64578 292848 64638 293320
rect 59631 292846 64638 292848
rect 40962 292554 41022 292818
rect 59631 292790 59636 292846
rect 59692 292790 64638 292846
rect 59631 292788 64638 292790
rect 649986 292848 650046 293320
rect 655983 292848 656049 292851
rect 649986 292846 656049 292848
rect 649986 292790 655988 292846
rect 656044 292790 656049 292846
rect 649986 292788 656049 292790
rect 59631 292785 59697 292788
rect 655983 292785 656049 292788
rect 673978 292786 673984 292850
rect 674048 292848 674054 292850
rect 675375 292848 675441 292851
rect 674048 292846 675441 292848
rect 674048 292790 675380 292846
rect 675436 292790 675441 292846
rect 674048 292788 675441 292790
rect 674048 292786 674054 292788
rect 675375 292785 675441 292788
rect 58191 292700 58257 292703
rect 58191 292698 64638 292700
rect 58191 292642 58196 292698
rect 58252 292642 64638 292698
rect 58191 292640 64638 292642
rect 58191 292637 58257 292640
rect 40954 292490 40960 292554
rect 41024 292490 41030 292554
rect 41154 292110 41214 292226
rect 64578 292138 64638 292640
rect 41146 292046 41152 292110
rect 41216 292046 41222 292110
rect 41346 291518 41406 291708
rect 649986 291664 650046 292138
rect 656175 291664 656241 291667
rect 649986 291662 656241 291664
rect 649986 291606 656180 291662
rect 656236 291606 656241 291662
rect 649986 291604 656241 291606
rect 656175 291601 656241 291604
rect 41338 291454 41344 291518
rect 41408 291454 41414 291518
rect 60207 291516 60273 291519
rect 60207 291514 64638 291516
rect 60207 291458 60212 291514
rect 60268 291458 64638 291514
rect 60207 291456 64638 291458
rect 60207 291453 60273 291456
rect 41538 291075 41598 291338
rect 41538 291070 41649 291075
rect 41538 291014 41588 291070
rect 41644 291014 41649 291070
rect 41538 291012 41649 291014
rect 41583 291009 41649 291012
rect 64578 290956 64638 291456
rect 649986 290924 650046 290956
rect 655791 290924 655857 290927
rect 649986 290922 655857 290924
rect 649986 290866 655796 290922
rect 655852 290866 655857 290922
rect 649986 290864 655857 290866
rect 655791 290861 655857 290864
rect 42447 290776 42513 290779
rect 41568 290774 42513 290776
rect 41568 290718 42452 290774
rect 42508 290718 42513 290774
rect 41568 290716 42513 290718
rect 42447 290713 42513 290716
rect 40578 290038 40638 290154
rect 40570 289974 40576 290038
rect 40640 289974 40646 290038
rect 41775 289814 41841 289817
rect 41568 289812 41841 289814
rect 41568 289756 41780 289812
rect 41836 289756 41841 289812
rect 41568 289754 41841 289756
rect 41775 289751 41841 289754
rect 41775 289296 41841 289299
rect 41568 289294 41841 289296
rect 41568 289238 41780 289294
rect 41836 289238 41841 289294
rect 41568 289236 41841 289238
rect 41775 289233 41841 289236
rect 59535 289296 59601 289299
rect 64578 289296 64638 289774
rect 59535 289294 64638 289296
rect 59535 289238 59540 289294
rect 59596 289238 64638 289294
rect 59535 289236 64638 289238
rect 649986 289296 650046 289774
rect 655599 289296 655665 289299
rect 649986 289294 655665 289296
rect 649986 289238 655604 289294
rect 655660 289238 655665 289294
rect 649986 289236 655665 289238
rect 59535 289233 59601 289236
rect 655599 289233 655665 289236
rect 41538 288556 41598 288674
rect 41538 288496 41790 288556
rect 23106 287967 23166 288304
rect 41730 288112 41790 288496
rect 23055 287962 23166 287967
rect 23055 287906 23060 287962
rect 23116 287906 23166 287962
rect 23055 287904 23166 287906
rect 41538 288052 41790 288112
rect 59151 288112 59217 288115
rect 64578 288112 64638 288592
rect 59151 288110 64638 288112
rect 59151 288054 59156 288110
rect 59212 288054 64638 288110
rect 59151 288052 64638 288054
rect 649986 288112 650046 288592
rect 674746 288494 674752 288558
rect 674816 288556 674822 288558
rect 675471 288556 675537 288559
rect 674816 288554 675537 288556
rect 674816 288498 675476 288554
rect 675532 288498 675537 288554
rect 674816 288496 675537 288498
rect 674816 288494 674822 288496
rect 675471 288493 675537 288496
rect 655407 288112 655473 288115
rect 649986 288110 655473 288112
rect 649986 288054 655412 288110
rect 655468 288054 655473 288110
rect 649986 288052 655473 288054
rect 23055 287901 23121 287904
rect 41538 287816 41598 288052
rect 59151 288049 59217 288052
rect 655407 288049 655473 288052
rect 41914 287902 41920 287966
rect 41984 287964 41990 287966
rect 42490 287964 42496 287966
rect 41984 287904 42496 287964
rect 41984 287902 41990 287904
rect 42490 287902 42496 287904
rect 42560 287902 42566 287966
rect 41871 287816 41937 287819
rect 41538 287814 41937 287816
rect 41538 287786 41876 287814
rect 41568 287758 41876 287786
rect 41932 287758 41937 287814
rect 41568 287756 41937 287758
rect 41871 287753 41937 287756
rect 23055 287520 23121 287523
rect 23055 287518 23166 287520
rect 23055 287462 23060 287518
rect 23116 287462 23166 287518
rect 23055 287457 23166 287462
rect 23106 287194 23166 287457
rect 59247 286928 59313 286931
rect 64578 286928 64638 287410
rect 59247 286926 64638 286928
rect 59247 286870 59252 286926
rect 59308 286870 64638 286926
rect 59247 286868 64638 286870
rect 649986 286928 650046 287410
rect 674938 287310 674944 287374
rect 675008 287372 675014 287374
rect 675471 287372 675537 287375
rect 675008 287370 675537 287372
rect 675008 287314 675476 287370
rect 675532 287314 675537 287370
rect 675008 287312 675537 287314
rect 675008 287310 675014 287312
rect 675471 287309 675537 287312
rect 655695 286928 655761 286931
rect 649986 286926 655761 286928
rect 649986 286870 655700 286926
rect 655756 286870 655761 286926
rect 649986 286868 655761 286870
rect 59247 286865 59313 286868
rect 655695 286865 655761 286868
rect 58959 285744 59025 285747
rect 64578 285744 64638 286228
rect 58959 285742 64638 285744
rect 58959 285686 58964 285742
rect 59020 285686 64638 285742
rect 58959 285684 64638 285686
rect 649986 285744 650046 286228
rect 655503 285744 655569 285747
rect 649986 285742 655569 285744
rect 649986 285686 655508 285742
rect 655564 285686 655569 285742
rect 649986 285684 655569 285686
rect 58959 285681 59025 285684
rect 655503 285681 655569 285684
rect 675663 285302 675729 285303
rect 675663 285298 675712 285302
rect 675776 285300 675782 285302
rect 675663 285242 675668 285298
rect 675663 285238 675712 285242
rect 675776 285240 675820 285300
rect 675776 285238 675782 285240
rect 675663 285237 675729 285238
rect 28719 285152 28785 285155
rect 41722 285152 41728 285154
rect 28719 285150 41728 285152
rect 28719 285094 28724 285150
rect 28780 285094 41728 285150
rect 28719 285092 41728 285094
rect 28719 285089 28785 285092
rect 41722 285090 41728 285092
rect 41792 285090 41798 285154
rect 57615 284560 57681 284563
rect 64578 284560 64638 285046
rect 57615 284558 64638 284560
rect 57615 284502 57620 284558
rect 57676 284502 64638 284558
rect 57615 284500 64638 284502
rect 649986 284560 650046 285046
rect 653775 284560 653841 284563
rect 649986 284558 653841 284560
rect 649986 284502 653780 284558
rect 653836 284502 653841 284558
rect 649986 284500 653841 284502
rect 57615 284497 57681 284500
rect 653775 284497 653841 284500
rect 58575 283376 58641 283379
rect 64578 283376 64638 283864
rect 58575 283374 64638 283376
rect 58575 283318 58580 283374
rect 58636 283318 64638 283374
rect 58575 283316 64638 283318
rect 649986 283376 650046 283864
rect 674554 283610 674560 283674
rect 674624 283672 674630 283674
rect 675375 283672 675441 283675
rect 674624 283670 675441 283672
rect 674624 283614 675380 283670
rect 675436 283614 675441 283670
rect 674624 283612 675441 283614
rect 674624 283610 674630 283612
rect 675375 283609 675441 283612
rect 655119 283376 655185 283379
rect 649986 283374 655185 283376
rect 649986 283318 655124 283374
rect 655180 283318 655185 283374
rect 649986 283316 655185 283318
rect 58575 283313 58641 283316
rect 655119 283313 655185 283316
rect 59631 282488 59697 282491
rect 64578 282488 64638 282682
rect 59631 282486 64638 282488
rect 59631 282430 59636 282486
rect 59692 282430 64638 282486
rect 59631 282428 64638 282430
rect 59631 282425 59697 282428
rect 649986 282340 650046 282682
rect 655311 282340 655377 282343
rect 649986 282338 655377 282340
rect 649986 282282 655316 282338
rect 655372 282282 655377 282338
rect 649986 282280 655377 282282
rect 655311 282277 655377 282280
rect 675759 281896 675825 281899
rect 676666 281896 676672 281898
rect 675759 281894 676672 281896
rect 675759 281838 675764 281894
rect 675820 281838 676672 281894
rect 675759 281836 676672 281838
rect 675759 281833 675825 281836
rect 676666 281834 676672 281836
rect 676736 281834 676742 281898
rect 41530 281686 41536 281750
rect 41600 281748 41606 281750
rect 41871 281748 41937 281751
rect 41600 281746 41937 281748
rect 41600 281690 41876 281746
rect 41932 281690 41937 281746
rect 41600 281688 41937 281690
rect 41600 281686 41606 281688
rect 41871 281685 41937 281688
rect 41914 281538 41920 281602
rect 41984 281600 41990 281602
rect 42447 281600 42513 281603
rect 41984 281598 42513 281600
rect 41984 281542 42452 281598
rect 42508 281542 42513 281598
rect 41984 281540 42513 281542
rect 41984 281538 41990 281540
rect 42447 281537 42513 281540
rect 58383 281008 58449 281011
rect 64578 281008 64638 281500
rect 58383 281006 64638 281008
rect 58383 280950 58388 281006
rect 58444 280950 64638 281006
rect 58383 280948 64638 280950
rect 649986 281008 650046 281500
rect 655215 281008 655281 281011
rect 649986 281006 655281 281008
rect 649986 280950 655220 281006
rect 655276 280950 655281 281006
rect 649986 280948 655281 280950
rect 58383 280945 58449 280948
rect 655215 280945 655281 280948
rect 58575 279824 58641 279827
rect 64578 279824 64638 280318
rect 58575 279822 64638 279824
rect 58575 279766 58580 279822
rect 58636 279766 64638 279822
rect 58575 279764 64638 279766
rect 649986 279824 650046 280318
rect 654255 279824 654321 279827
rect 649986 279822 654321 279824
rect 649986 279766 654260 279822
rect 654316 279766 654321 279822
rect 649986 279764 654321 279766
rect 58575 279761 58641 279764
rect 654255 279761 654321 279764
rect 45039 278640 45105 278643
rect 670479 278640 670545 278643
rect 45039 278638 670545 278640
rect 45039 278582 45044 278638
rect 45100 278582 670484 278638
rect 670540 278582 670545 278638
rect 45039 278580 670545 278582
rect 45039 278577 45105 278580
rect 670479 278577 670545 278580
rect 61935 278492 62001 278495
rect 675130 278492 675136 278494
rect 61935 278490 675136 278492
rect 61935 278434 61940 278490
rect 61996 278434 675136 278490
rect 61935 278432 675136 278434
rect 61935 278429 62001 278432
rect 675130 278430 675136 278432
rect 675200 278492 675206 278494
rect 675279 278492 675345 278495
rect 675200 278490 675345 278492
rect 675200 278434 675284 278490
rect 675340 278434 675345 278490
rect 675200 278432 675345 278434
rect 675200 278430 675206 278432
rect 675279 278429 675345 278432
rect 62127 278344 62193 278347
rect 675514 278344 675520 278346
rect 62127 278342 675520 278344
rect 62127 278286 62132 278342
rect 62188 278286 675520 278342
rect 62127 278284 675520 278286
rect 62127 278281 62193 278284
rect 675514 278282 675520 278284
rect 675584 278344 675590 278346
rect 675759 278344 675825 278347
rect 675584 278342 675825 278344
rect 675584 278286 675764 278342
rect 675820 278286 675825 278342
rect 675584 278284 675825 278286
rect 675584 278282 675590 278284
rect 675759 278281 675825 278284
rect 62319 278196 62385 278199
rect 674170 278196 674176 278198
rect 62319 278194 674176 278196
rect 62319 278138 62324 278194
rect 62380 278138 674176 278194
rect 62319 278136 674176 278138
rect 62319 278133 62385 278136
rect 674170 278134 674176 278136
rect 674240 278134 674246 278198
rect 41967 278050 42033 278051
rect 41914 277986 41920 278050
rect 41984 278048 42033 278050
rect 62607 278048 62673 278051
rect 670287 278048 670353 278051
rect 41984 278046 42076 278048
rect 42028 277990 42076 278046
rect 41984 277988 42076 277990
rect 62607 278046 670353 278048
rect 62607 277990 62612 278046
rect 62668 277990 670292 278046
rect 670348 277990 670353 278046
rect 62607 277988 670353 277990
rect 41984 277986 42033 277988
rect 41967 277985 42033 277986
rect 62607 277985 62673 277988
rect 670287 277985 670353 277988
rect 62895 277900 62961 277903
rect 670095 277900 670161 277903
rect 62895 277898 670161 277900
rect 62895 277842 62900 277898
rect 62956 277842 670100 277898
rect 670156 277842 670161 277898
rect 62895 277840 670161 277842
rect 62895 277837 62961 277840
rect 670095 277837 670161 277840
rect 62991 277752 63057 277755
rect 669903 277752 669969 277755
rect 62991 277750 669969 277752
rect 62991 277694 62996 277750
rect 63052 277694 669908 277750
rect 669964 277694 669969 277750
rect 62991 277692 669969 277694
rect 62991 277689 63057 277692
rect 669903 277689 669969 277692
rect 402543 276864 402609 276867
rect 526959 276864 527025 276867
rect 402543 276862 527025 276864
rect 402543 276806 402548 276862
rect 402604 276806 526964 276862
rect 527020 276806 527025 276862
rect 402543 276804 527025 276806
rect 402543 276801 402609 276804
rect 526959 276801 527025 276804
rect 393903 276716 393969 276719
rect 603663 276716 603729 276719
rect 393903 276714 603729 276716
rect 393903 276658 393908 276714
rect 393964 276658 603668 276714
rect 603724 276658 603729 276714
rect 393903 276656 603729 276658
rect 393903 276653 393969 276656
rect 603663 276653 603729 276656
rect 42159 276568 42225 276571
rect 42490 276568 42496 276570
rect 42159 276566 42496 276568
rect 42159 276510 42164 276566
rect 42220 276510 42496 276566
rect 42159 276508 42496 276510
rect 42159 276505 42225 276508
rect 42490 276506 42496 276508
rect 42560 276506 42566 276570
rect 396687 276568 396753 276571
rect 610767 276568 610833 276571
rect 396687 276566 610833 276568
rect 396687 276510 396692 276566
rect 396748 276510 610772 276566
rect 610828 276510 610833 276566
rect 396687 276508 610833 276510
rect 396687 276505 396753 276508
rect 610767 276505 610833 276508
rect 45711 276272 45777 276275
rect 672399 276272 672465 276275
rect 45711 276270 672465 276272
rect 45711 276214 45716 276270
rect 45772 276214 672404 276270
rect 672460 276214 672465 276270
rect 45711 276212 672465 276214
rect 45711 276209 45777 276212
rect 672399 276209 672465 276212
rect 379023 276124 379089 276127
rect 566991 276124 567057 276127
rect 379023 276122 567057 276124
rect 379023 276066 379028 276122
rect 379084 276066 566996 276122
rect 567052 276066 567057 276122
rect 379023 276064 567057 276066
rect 379023 276061 379089 276064
rect 566991 276061 567057 276064
rect 383439 275976 383505 275979
rect 577647 275976 577713 275979
rect 383439 275974 577713 275976
rect 383439 275918 383444 275974
rect 383500 275918 577652 275974
rect 577708 275918 577713 275974
rect 383439 275916 577713 275918
rect 383439 275913 383505 275916
rect 577647 275913 577713 275916
rect 390351 275828 390417 275831
rect 595407 275828 595473 275831
rect 390351 275826 595473 275828
rect 390351 275770 390356 275826
rect 390412 275770 595412 275826
rect 595468 275770 595473 275826
rect 390351 275768 595473 275770
rect 390351 275765 390417 275768
rect 595407 275765 595473 275768
rect 398895 275680 398961 275683
rect 616623 275680 616689 275683
rect 398895 275678 616689 275680
rect 398895 275622 398900 275678
rect 398956 275622 616628 275678
rect 616684 275622 616689 275678
rect 398895 275620 616689 275622
rect 398895 275617 398961 275620
rect 616623 275617 616689 275620
rect 407823 275532 407889 275535
rect 637935 275532 638001 275535
rect 407823 275530 638001 275532
rect 407823 275474 407828 275530
rect 407884 275474 637940 275530
rect 637996 275474 638001 275530
rect 407823 275472 638001 275474
rect 407823 275469 407889 275472
rect 637935 275469 638001 275472
rect 44751 275384 44817 275387
rect 646479 275384 646545 275387
rect 44751 275382 646545 275384
rect 44751 275326 44756 275382
rect 44812 275326 646484 275382
rect 646540 275326 646545 275382
rect 44751 275324 646545 275326
rect 44751 275321 44817 275324
rect 646479 275321 646545 275324
rect 50607 275236 50673 275239
rect 669711 275236 669777 275239
rect 50607 275234 669777 275236
rect 50607 275178 50612 275234
rect 50668 275178 669716 275234
rect 669772 275178 669777 275234
rect 50607 275176 669777 275178
rect 50607 275173 50673 275176
rect 669711 275173 669777 275176
rect 50415 275088 50481 275091
rect 669519 275088 669585 275091
rect 50415 275086 669585 275088
rect 50415 275030 50420 275086
rect 50476 275030 669524 275086
rect 669580 275030 669585 275086
rect 50415 275028 669585 275030
rect 50415 275025 50481 275028
rect 669519 275025 669585 275028
rect 353391 274940 353457 274943
rect 503151 274940 503217 274943
rect 353391 274938 503217 274940
rect 353391 274882 353396 274938
rect 353452 274882 503156 274938
rect 503212 274882 503217 274938
rect 353391 274880 503217 274882
rect 353391 274877 353457 274880
rect 503151 274877 503217 274880
rect 350223 274792 350289 274795
rect 496047 274792 496113 274795
rect 350223 274790 496113 274792
rect 350223 274734 350228 274790
rect 350284 274734 496052 274790
rect 496108 274734 496113 274790
rect 350223 274732 496113 274734
rect 350223 274729 350289 274732
rect 496047 274729 496113 274732
rect 347631 274644 347697 274647
rect 489039 274644 489105 274647
rect 347631 274642 489105 274644
rect 347631 274586 347636 274642
rect 347692 274586 489044 274642
rect 489100 274586 489105 274642
rect 347631 274584 489105 274586
rect 347631 274581 347697 274584
rect 489039 274581 489105 274584
rect 341679 274496 341745 274499
rect 474831 274496 474897 274499
rect 341679 274494 474897 274496
rect 341679 274438 341684 274494
rect 341740 274438 474836 274494
rect 474892 274438 474897 274494
rect 341679 274436 474897 274438
rect 341679 274433 341745 274436
rect 474831 274433 474897 274436
rect 42106 274286 42112 274350
rect 42176 274348 42182 274350
rect 670191 274348 670257 274351
rect 42176 274346 670257 274348
rect 42176 274290 670196 274346
rect 670252 274290 670257 274346
rect 42176 274288 670257 274290
rect 42176 274286 42182 274288
rect 670191 274285 670257 274288
rect 40570 274138 40576 274202
rect 40640 274200 40646 274202
rect 41775 274200 41841 274203
rect 40640 274198 41841 274200
rect 40640 274142 41780 274198
rect 41836 274142 41841 274198
rect 40640 274140 41841 274142
rect 40640 274138 40646 274140
rect 41775 274137 41841 274140
rect 41338 273546 41344 273610
rect 41408 273608 41414 273610
rect 41775 273608 41841 273611
rect 41408 273606 41841 273608
rect 41408 273550 41780 273606
rect 41836 273550 41841 273606
rect 41408 273548 41841 273550
rect 41408 273546 41414 273548
rect 41775 273545 41841 273548
rect 62703 273608 62769 273611
rect 672783 273608 672849 273611
rect 62703 273606 672849 273608
rect 62703 273550 62708 273606
rect 62764 273550 672788 273606
rect 672844 273550 672849 273606
rect 62703 273548 672849 273550
rect 62703 273545 62769 273548
rect 672783 273545 672849 273548
rect 62511 273460 62577 273463
rect 672591 273460 672657 273463
rect 62511 273458 672657 273460
rect 62511 273402 62516 273458
rect 62572 273402 672596 273458
rect 672652 273402 672657 273458
rect 62511 273400 672657 273402
rect 62511 273397 62577 273400
rect 672591 273397 672657 273400
rect 45231 273312 45297 273315
rect 408879 273312 408945 273315
rect 45231 273310 408945 273312
rect 45231 273254 45236 273310
rect 45292 273254 408884 273310
rect 408940 273254 408945 273310
rect 45231 273252 408945 273254
rect 45231 273249 45297 273252
rect 408879 273249 408945 273252
rect 382959 273164 383025 273167
rect 576495 273164 576561 273167
rect 382959 273162 576561 273164
rect 382959 273106 382964 273162
rect 383020 273106 576500 273162
rect 576556 273106 576561 273162
rect 382959 273104 576561 273106
rect 382959 273101 383025 273104
rect 576495 273101 576561 273104
rect 390159 273016 390225 273019
rect 594159 273016 594225 273019
rect 390159 273014 594225 273016
rect 390159 272958 390164 273014
rect 390220 272958 594164 273014
rect 594220 272958 594225 273014
rect 390159 272956 594225 272958
rect 390159 272953 390225 272956
rect 594159 272953 594225 272956
rect 41146 272806 41152 272870
rect 41216 272868 41222 272870
rect 41775 272868 41841 272871
rect 41216 272866 41841 272868
rect 41216 272810 41780 272866
rect 41836 272810 41841 272866
rect 41216 272808 41841 272810
rect 41216 272806 41222 272808
rect 41775 272805 41841 272808
rect 392751 272868 392817 272871
rect 601263 272868 601329 272871
rect 392751 272866 601329 272868
rect 392751 272810 392756 272866
rect 392812 272810 601268 272866
rect 601324 272810 601329 272866
rect 392751 272808 601329 272810
rect 392751 272805 392817 272808
rect 601263 272805 601329 272808
rect 91887 272720 91953 272723
rect 200463 272720 200529 272723
rect 91887 272718 200529 272720
rect 91887 272662 91892 272718
rect 91948 272662 200468 272718
rect 200524 272662 200529 272718
rect 91887 272660 200529 272662
rect 91887 272657 91953 272660
rect 200463 272657 200529 272660
rect 398703 272720 398769 272723
rect 615471 272720 615537 272723
rect 398703 272718 615537 272720
rect 398703 272662 398708 272718
rect 398764 272662 615476 272718
rect 615532 272662 615537 272718
rect 398703 272660 615537 272662
rect 398703 272657 398769 272660
rect 615471 272657 615537 272660
rect 88335 272572 88401 272575
rect 199215 272572 199281 272575
rect 88335 272570 199281 272572
rect 88335 272514 88340 272570
rect 88396 272514 199220 272570
rect 199276 272514 199281 272570
rect 88335 272512 199281 272514
rect 88335 272509 88401 272512
rect 199215 272509 199281 272512
rect 404175 272572 404241 272575
rect 629679 272572 629745 272575
rect 404175 272570 629745 272572
rect 404175 272514 404180 272570
rect 404236 272514 629684 272570
rect 629740 272514 629745 272570
rect 404175 272512 629745 272514
rect 404175 272509 404241 272512
rect 629679 272509 629745 272512
rect 78831 272424 78897 272427
rect 196623 272424 196689 272427
rect 78831 272422 196689 272424
rect 78831 272366 78836 272422
rect 78892 272366 196628 272422
rect 196684 272366 196689 272422
rect 78831 272364 196689 272366
rect 78831 272361 78897 272364
rect 196623 272361 196689 272364
rect 407247 272424 407313 272427
rect 636783 272424 636849 272427
rect 407247 272422 636849 272424
rect 407247 272366 407252 272422
rect 407308 272366 636788 272422
rect 636844 272366 636849 272422
rect 407247 272364 636849 272366
rect 407247 272361 407313 272364
rect 636783 272361 636849 272364
rect 40378 272214 40384 272278
rect 40448 272276 40454 272278
rect 41775 272276 41841 272279
rect 40448 272274 41841 272276
rect 40448 272218 41780 272274
rect 41836 272218 41841 272274
rect 40448 272216 41841 272218
rect 40448 272214 40454 272216
rect 41775 272213 41841 272216
rect 72975 272276 73041 272279
rect 194415 272276 194481 272279
rect 72975 272274 194481 272276
rect 72975 272218 72980 272274
rect 73036 272218 194420 272274
rect 194476 272218 194481 272274
rect 72975 272216 194481 272218
rect 72975 272213 73041 272216
rect 194415 272213 194481 272216
rect 410895 272276 410961 272279
rect 646191 272276 646257 272279
rect 410895 272274 646257 272276
rect 410895 272218 410900 272274
rect 410956 272218 646196 272274
rect 646252 272218 646257 272274
rect 410895 272216 646257 272218
rect 410895 272213 410961 272216
rect 646191 272213 646257 272216
rect 70575 272128 70641 272131
rect 193743 272128 193809 272131
rect 70575 272126 193809 272128
rect 70575 272070 70580 272126
rect 70636 272070 193748 272126
rect 193804 272070 193809 272126
rect 70575 272068 193809 272070
rect 70575 272065 70641 272068
rect 193743 272065 193809 272068
rect 411759 272128 411825 272131
rect 648591 272128 648657 272131
rect 411759 272126 648657 272128
rect 411759 272070 411764 272126
rect 411820 272070 648596 272126
rect 648652 272070 648657 272126
rect 411759 272068 648657 272070
rect 411759 272065 411825 272068
rect 648591 272065 648657 272068
rect 378639 271980 378705 271983
rect 565839 271980 565905 271983
rect 378639 271978 565905 271980
rect 378639 271922 378644 271978
rect 378700 271922 565844 271978
rect 565900 271922 565905 271978
rect 378639 271920 565905 271922
rect 378639 271917 378705 271920
rect 565839 271917 565905 271920
rect 375567 271832 375633 271835
rect 558735 271832 558801 271835
rect 375567 271830 558801 271832
rect 375567 271774 375572 271830
rect 375628 271774 558740 271830
rect 558796 271774 558801 271830
rect 375567 271772 558801 271774
rect 375567 271769 375633 271772
rect 558735 271769 558801 271772
rect 370095 271684 370161 271687
rect 544527 271684 544593 271687
rect 370095 271682 544593 271684
rect 370095 271626 370100 271682
rect 370156 271626 544532 271682
rect 544588 271626 544593 271682
rect 370095 271624 544593 271626
rect 370095 271621 370161 271624
rect 544527 271621 544593 271624
rect 369615 271536 369681 271539
rect 543375 271536 543441 271539
rect 369615 271534 543441 271536
rect 369615 271478 369620 271534
rect 369676 271478 543380 271534
rect 543436 271478 543441 271534
rect 369615 271476 543441 271478
rect 369615 271473 369681 271476
rect 543375 271473 543441 271476
rect 382383 270796 382449 270799
rect 388719 270796 388785 270799
rect 382383 270794 388785 270796
rect 382383 270738 382388 270794
rect 382444 270738 388724 270794
rect 388780 270738 388785 270794
rect 382383 270736 388785 270738
rect 382383 270733 382449 270736
rect 388719 270733 388785 270736
rect 41775 270650 41841 270651
rect 41722 270648 41728 270650
rect 41684 270588 41728 270648
rect 41792 270646 41841 270650
rect 41836 270590 41841 270646
rect 41722 270586 41728 270588
rect 41792 270586 41841 270590
rect 41775 270585 41841 270586
rect 45423 270648 45489 270651
rect 669999 270648 670065 270651
rect 45423 270646 670065 270648
rect 45423 270590 45428 270646
rect 45484 270590 670004 270646
rect 670060 270590 670065 270646
rect 45423 270588 670065 270590
rect 45423 270585 45489 270588
rect 669999 270585 670065 270588
rect 367887 270500 367953 270503
rect 539823 270500 539889 270503
rect 367887 270498 539889 270500
rect 367887 270442 367892 270498
rect 367948 270442 539828 270498
rect 539884 270442 539889 270498
rect 367887 270440 539889 270442
rect 367887 270437 367953 270440
rect 539823 270437 539889 270440
rect 377007 270352 377073 270355
rect 562287 270352 562353 270355
rect 377007 270350 562353 270352
rect 377007 270294 377012 270350
rect 377068 270294 562292 270350
rect 562348 270294 562353 270350
rect 377007 270292 562353 270294
rect 377007 270289 377073 270292
rect 562287 270289 562353 270292
rect 385551 270204 385617 270207
rect 583599 270204 583665 270207
rect 385551 270202 583665 270204
rect 385551 270146 385556 270202
rect 385612 270146 583604 270202
rect 583660 270146 583665 270202
rect 385551 270144 583665 270146
rect 385551 270141 385617 270144
rect 583599 270141 583665 270144
rect 40954 269994 40960 270058
rect 41024 270056 41030 270058
rect 41775 270056 41841 270059
rect 41024 270054 41841 270056
rect 41024 269998 41780 270054
rect 41836 269998 41841 270054
rect 41024 269996 41841 269998
rect 41024 269994 41030 269996
rect 41775 269993 41841 269996
rect 388431 270056 388497 270059
rect 590607 270056 590673 270059
rect 388431 270054 590673 270056
rect 388431 269998 388436 270054
rect 388492 269998 590612 270054
rect 590668 269998 590673 270054
rect 388431 269996 590673 269998
rect 388431 269993 388497 269996
rect 590607 269993 590673 269996
rect 139119 269908 139185 269911
rect 213327 269908 213393 269911
rect 139119 269906 213393 269908
rect 139119 269850 139124 269906
rect 139180 269850 213332 269906
rect 213388 269850 213393 269906
rect 139119 269848 213393 269850
rect 139119 269845 139185 269848
rect 213327 269845 213393 269848
rect 391503 269908 391569 269911
rect 597711 269908 597777 269911
rect 391503 269906 597777 269908
rect 391503 269850 391508 269906
rect 391564 269850 597716 269906
rect 597772 269850 597777 269906
rect 391503 269848 597777 269850
rect 391503 269845 391569 269848
rect 597711 269845 597777 269848
rect 77583 269760 77649 269763
rect 196143 269760 196209 269763
rect 77583 269758 196209 269760
rect 77583 269702 77588 269758
rect 77644 269702 196148 269758
rect 196204 269702 196209 269758
rect 77583 269700 196209 269702
rect 77583 269697 77649 269700
rect 196143 269697 196209 269700
rect 403023 269760 403089 269763
rect 626127 269760 626193 269763
rect 403023 269758 626193 269760
rect 403023 269702 403028 269758
rect 403084 269702 626132 269758
rect 626188 269702 626193 269758
rect 403023 269700 626193 269702
rect 403023 269697 403089 269700
rect 626127 269697 626193 269700
rect 69423 269612 69489 269615
rect 193071 269612 193137 269615
rect 69423 269610 193137 269612
rect 69423 269554 69428 269610
rect 69484 269554 193076 269610
rect 193132 269554 193137 269610
rect 69423 269552 193137 269554
rect 69423 269549 69489 269552
rect 193071 269549 193137 269552
rect 405615 269612 405681 269615
rect 633231 269612 633297 269615
rect 405615 269610 633297 269612
rect 405615 269554 405620 269610
rect 405676 269554 633236 269610
rect 633292 269554 633297 269610
rect 405615 269552 633297 269554
rect 405615 269549 405681 269552
rect 633231 269549 633297 269552
rect 67023 269464 67089 269467
rect 192591 269464 192657 269467
rect 67023 269462 192657 269464
rect 67023 269406 67028 269462
rect 67084 269406 192596 269462
rect 192652 269406 192657 269462
rect 67023 269404 192657 269406
rect 67023 269401 67089 269404
rect 192591 269401 192657 269404
rect 410415 269464 410481 269467
rect 645039 269464 645105 269467
rect 410415 269462 645105 269464
rect 410415 269406 410420 269462
rect 410476 269406 645044 269462
rect 645100 269406 645105 269462
rect 410415 269404 645105 269406
rect 410415 269401 410481 269404
rect 645039 269401 645105 269404
rect 42159 269316 42225 269319
rect 42298 269316 42304 269318
rect 42159 269314 42304 269316
rect 42159 269258 42164 269314
rect 42220 269258 42304 269314
rect 42159 269256 42304 269258
rect 42159 269253 42225 269256
rect 42298 269254 42304 269256
rect 42368 269254 42374 269318
rect 71727 269316 71793 269319
rect 194223 269316 194289 269319
rect 71727 269314 194289 269316
rect 71727 269258 71732 269314
rect 71788 269258 194228 269314
rect 194284 269258 194289 269314
rect 71727 269256 194289 269258
rect 71727 269253 71793 269256
rect 194223 269253 194289 269256
rect 411567 269316 411633 269319
rect 647343 269316 647409 269319
rect 411567 269314 647409 269316
rect 411567 269258 411572 269314
rect 411628 269258 647348 269314
rect 647404 269258 647409 269314
rect 411567 269256 647409 269258
rect 411567 269253 411633 269256
rect 647343 269253 647409 269256
rect 368367 269168 368433 269171
rect 540975 269168 541041 269171
rect 368367 269166 541041 269168
rect 368367 269110 368372 269166
rect 368428 269110 540980 269166
rect 541036 269110 541041 269166
rect 368367 269108 541041 269110
rect 368367 269105 368433 269108
rect 540975 269105 541041 269108
rect 397071 269020 397137 269023
rect 532815 269020 532881 269023
rect 397071 269018 532881 269020
rect 397071 268962 397076 269018
rect 397132 268962 532820 269018
rect 532876 268962 532881 269018
rect 397071 268960 532881 268962
rect 397071 268957 397137 268960
rect 532815 268957 532881 268960
rect 374319 268872 374385 268875
rect 508239 268872 508305 268875
rect 374319 268870 508305 268872
rect 374319 268814 374324 268870
rect 374380 268814 508244 268870
rect 508300 268814 508305 268870
rect 374319 268812 508305 268814
rect 374319 268809 374385 268812
rect 508239 268809 508305 268812
rect 208143 268132 208209 268135
rect 214287 268132 214353 268135
rect 208143 268130 214353 268132
rect 208143 268074 208148 268130
rect 208204 268074 214292 268130
rect 214348 268074 214353 268130
rect 208143 268072 214353 268074
rect 208143 268069 208209 268072
rect 214287 268069 214353 268072
rect 44655 267392 44721 267395
rect 646575 267392 646641 267395
rect 44655 267390 646641 267392
rect 44655 267334 44660 267390
rect 44716 267334 646580 267390
rect 646636 267334 646641 267390
rect 44655 267332 646641 267334
rect 44655 267329 44721 267332
rect 646575 267329 646641 267332
rect 676290 267247 676350 267510
rect 43503 267244 43569 267247
rect 652239 267244 652305 267247
rect 43503 267242 652305 267244
rect 43503 267186 43508 267242
rect 43564 267186 652244 267242
rect 652300 267186 652305 267242
rect 43503 267184 652305 267186
rect 676290 267242 676401 267247
rect 676290 267186 676340 267242
rect 676396 267186 676401 267242
rect 676290 267184 676401 267186
rect 43503 267181 43569 267184
rect 652239 267181 652305 267184
rect 676335 267181 676401 267184
rect 62415 267096 62481 267099
rect 672783 267096 672849 267099
rect 62415 267094 672849 267096
rect 62415 267038 62420 267094
rect 62476 267038 672788 267094
rect 672844 267038 672849 267094
rect 62415 267036 672849 267038
rect 62415 267033 62481 267036
rect 672783 267033 672849 267036
rect 62031 266948 62097 266951
rect 672591 266948 672657 266951
rect 62031 266946 672657 266948
rect 62031 266890 62036 266946
rect 62092 266890 672596 266946
rect 672652 266890 672657 266946
rect 62031 266888 672657 266890
rect 62031 266885 62097 266888
rect 672591 266885 672657 266888
rect 61839 266800 61905 266803
rect 672399 266800 672465 266803
rect 61839 266798 672465 266800
rect 61839 266742 61844 266798
rect 61900 266742 672404 266798
rect 672460 266742 672465 266798
rect 61839 266740 672465 266742
rect 61839 266737 61905 266740
rect 672399 266737 672465 266740
rect 62223 266652 62289 266655
rect 672975 266652 673041 266655
rect 62223 266650 673041 266652
rect 62223 266594 62228 266650
rect 62284 266594 672980 266650
rect 673036 266594 673041 266650
rect 62223 266592 673041 266594
rect 62223 266589 62289 266592
rect 672975 266589 673041 266592
rect 676143 266652 676209 266655
rect 676290 266652 676350 266918
rect 676143 266650 676350 266652
rect 676143 266594 676148 266650
rect 676204 266594 676350 266650
rect 676143 266592 676350 266594
rect 676143 266589 676209 266592
rect 44943 266504 45009 266507
rect 671823 266504 671889 266507
rect 44943 266502 671889 266504
rect 44943 266446 44948 266502
rect 45004 266446 671828 266502
rect 671884 266446 671889 266502
rect 44943 266444 671889 266446
rect 44943 266441 45009 266444
rect 671823 266441 671889 266444
rect 45135 266356 45201 266359
rect 673455 266356 673521 266359
rect 45135 266354 673521 266356
rect 45135 266298 45140 266354
rect 45196 266298 673460 266354
rect 673516 266298 673521 266354
rect 45135 266296 673521 266298
rect 45135 266293 45201 266296
rect 673455 266293 673521 266296
rect 676290 266211 676350 266326
rect 676239 266206 676350 266211
rect 676239 266150 676244 266206
rect 676300 266150 676350 266206
rect 676239 266148 676350 266150
rect 676239 266145 676305 266148
rect 675322 265998 675328 266062
rect 675392 266060 675398 266062
rect 675392 266000 676320 266060
rect 675392 265998 675398 266000
rect 673978 265406 673984 265470
rect 674048 265468 674054 265470
rect 674048 265408 676320 265468
rect 674048 265406 674054 265408
rect 679695 265172 679761 265175
rect 679695 265170 679806 265172
rect 679695 265114 679700 265170
rect 679756 265114 679806 265170
rect 679695 265109 679806 265114
rect 679746 264846 679806 265109
rect 676239 264728 676305 264731
rect 676239 264726 676350 264728
rect 676239 264670 676244 264726
rect 676300 264670 676350 264726
rect 676239 264665 676350 264670
rect 676290 264476 676350 264665
rect 679791 264284 679857 264287
rect 679746 264282 679857 264284
rect 679746 264226 679796 264282
rect 679852 264226 679857 264282
rect 679746 264221 679857 264226
rect 679746 263958 679806 264221
rect 47823 263544 47889 263547
rect 668175 263544 668241 263547
rect 47823 263542 668241 263544
rect 47823 263486 47828 263542
rect 47884 263486 668180 263542
rect 668236 263486 668241 263542
rect 47823 263484 668241 263486
rect 47823 263481 47889 263484
rect 668175 263481 668241 263484
rect 43311 263396 43377 263399
rect 649743 263396 649809 263399
rect 43311 263394 649809 263396
rect 43311 263338 43316 263394
rect 43372 263338 649748 263394
rect 649804 263338 649809 263394
rect 43311 263336 649809 263338
rect 43311 263333 43377 263336
rect 649743 263333 649809 263336
rect 673455 263396 673521 263399
rect 673455 263394 676320 263396
rect 673455 263338 673460 263394
rect 673516 263338 676320 263394
rect 673455 263336 676320 263338
rect 673455 263333 673521 263336
rect 676290 262807 676350 262922
rect 676239 262802 676350 262807
rect 676239 262746 676244 262802
rect 676300 262746 676350 262802
rect 676239 262744 676350 262746
rect 676239 262741 676305 262744
rect 676866 262215 676926 262478
rect 420399 262212 420465 262215
rect 412512 262210 420465 262212
rect 412512 262154 420404 262210
rect 420460 262154 420465 262210
rect 412512 262152 420465 262154
rect 676866 262210 676977 262215
rect 676866 262154 676916 262210
rect 676972 262154 676977 262210
rect 676866 262152 676977 262154
rect 420399 262149 420465 262152
rect 676911 262149 676977 262152
rect 676290 261770 676350 261886
rect 676282 261706 676288 261770
rect 676352 261706 676358 261770
rect 676290 261327 676350 261442
rect 676239 261322 676350 261327
rect 676239 261266 676244 261322
rect 676300 261266 676350 261322
rect 676239 261264 676350 261266
rect 676239 261261 676305 261264
rect 675706 260966 675712 261030
rect 675776 261028 675782 261030
rect 675776 260968 676320 261028
rect 675776 260966 675782 260968
rect 676815 260584 676881 260587
rect 676815 260582 676926 260584
rect 676815 260526 676820 260582
rect 676876 260526 676926 260582
rect 676815 260521 676926 260526
rect 676866 260406 676926 260521
rect 676290 259847 676350 259962
rect 420399 259844 420465 259847
rect 412512 259842 420465 259844
rect 412512 259786 420404 259842
rect 420460 259786 420465 259842
rect 412512 259784 420465 259786
rect 420399 259781 420465 259784
rect 676239 259842 676350 259847
rect 676239 259786 676244 259842
rect 676300 259786 676350 259842
rect 676239 259784 676350 259786
rect 676239 259781 676305 259784
rect 676047 259474 676113 259477
rect 676047 259472 676320 259474
rect 676047 259416 676052 259472
rect 676108 259416 676320 259472
rect 676047 259414 676320 259416
rect 676047 259411 676113 259414
rect 191535 259400 191601 259403
rect 191535 259398 191904 259400
rect 191535 259342 191540 259398
rect 191596 259342 191904 259398
rect 191535 259340 191904 259342
rect 191535 259337 191601 259340
rect 675514 258894 675520 258958
rect 675584 258956 675590 258958
rect 675584 258896 676320 258956
rect 675584 258894 675590 258896
rect 674938 258450 674944 258514
rect 675008 258512 675014 258514
rect 675008 258452 676320 258512
rect 675008 258450 675014 258452
rect 674554 257858 674560 257922
rect 674624 257920 674630 257922
rect 674624 257860 676320 257920
rect 674624 257858 674630 257860
rect 41538 256887 41598 257076
rect 412482 257032 412542 257520
rect 676047 257476 676113 257479
rect 676047 257474 676320 257476
rect 676047 257418 676052 257474
rect 676108 257418 676320 257474
rect 676047 257416 676320 257418
rect 676047 257413 676113 257416
rect 420399 257032 420465 257035
rect 412482 257030 420465 257032
rect 412482 256974 420404 257030
rect 420460 256974 420465 257030
rect 412482 256972 420465 256974
rect 420399 256969 420465 256972
rect 675951 257032 676017 257035
rect 675951 257030 676320 257032
rect 675951 256974 675956 257030
rect 676012 256974 676320 257030
rect 675951 256972 676320 256974
rect 675951 256969 676017 256972
rect 41538 256882 41649 256887
rect 41538 256826 41588 256882
rect 41644 256826 41649 256882
rect 41538 256824 41649 256826
rect 41583 256821 41649 256824
rect 41775 256588 41841 256591
rect 41568 256586 41841 256588
rect 41568 256530 41780 256586
rect 41836 256530 41841 256586
rect 41568 256528 41841 256530
rect 41775 256525 41841 256528
rect 674746 256378 674752 256442
rect 674816 256440 674822 256442
rect 674816 256380 676320 256440
rect 674816 256378 674822 256380
rect 41775 255996 41841 255999
rect 41568 255994 41841 255996
rect 41568 255938 41780 255994
rect 41836 255938 41841 255994
rect 41568 255936 41841 255938
rect 41775 255933 41841 255936
rect 679746 255703 679806 255966
rect 679746 255698 679857 255703
rect 679746 255642 679796 255698
rect 679852 255642 679857 255698
rect 679746 255640 679857 255642
rect 679791 255637 679857 255640
rect 41775 255552 41841 255555
rect 41568 255550 41841 255552
rect 41568 255494 41780 255550
rect 41836 255494 41841 255550
rect 41568 255492 41841 255494
rect 41775 255489 41841 255492
rect 685506 255259 685566 255522
rect 420399 255256 420465 255259
rect 679791 255256 679857 255259
rect 412512 255254 420465 255256
rect 412512 255198 420404 255254
rect 420460 255198 420465 255254
rect 412512 255196 420465 255198
rect 420399 255193 420465 255196
rect 679746 255254 679857 255256
rect 679746 255198 679796 255254
rect 679852 255198 679857 255254
rect 679746 255193 679857 255198
rect 685506 255254 685617 255259
rect 685506 255198 685556 255254
rect 685612 255198 685617 255254
rect 685506 255196 685617 255198
rect 685551 255193 685617 255196
rect 41775 255108 41841 255111
rect 41568 255106 41841 255108
rect 41568 255050 41780 255106
rect 41836 255050 41841 255106
rect 41568 255048 41841 255050
rect 41775 255045 41841 255048
rect 679746 254930 679806 255193
rect 23343 254812 23409 254815
rect 685551 254812 685617 254815
rect 23298 254810 23409 254812
rect 23298 254754 23348 254810
rect 23404 254754 23409 254810
rect 23298 254749 23409 254754
rect 685506 254810 685617 254812
rect 685506 254754 685556 254810
rect 685612 254754 685617 254810
rect 685506 254749 685617 254754
rect 23298 254486 23358 254749
rect 685506 254412 685566 254749
rect 23490 253927 23550 254042
rect 23151 253924 23217 253927
rect 23106 253922 23217 253924
rect 23106 253866 23156 253922
rect 23212 253866 23217 253922
rect 23106 253861 23217 253866
rect 23490 253922 23601 253927
rect 23490 253866 23540 253922
rect 23596 253866 23601 253922
rect 23490 253864 23601 253866
rect 23535 253861 23601 253864
rect 23106 253524 23166 253861
rect 23055 253332 23121 253335
rect 23055 253330 23166 253332
rect 23055 253274 23060 253330
rect 23116 253274 23166 253330
rect 23055 253269 23166 253274
rect 675898 253270 675904 253334
rect 675968 253332 675974 253334
rect 676815 253332 676881 253335
rect 675968 253330 676881 253332
rect 675968 253274 676820 253330
rect 676876 253274 676881 253330
rect 675968 253272 676881 253274
rect 675968 253270 675974 253272
rect 676815 253269 676881 253272
rect 23106 253006 23166 253269
rect 676090 253122 676096 253186
rect 676160 253184 676166 253186
rect 676911 253184 676977 253187
rect 676160 253182 676977 253184
rect 676160 253126 676916 253182
rect 676972 253126 676977 253182
rect 676160 253124 676977 253126
rect 676160 253122 676166 253124
rect 676911 253121 676977 253124
rect 420399 252888 420465 252891
rect 412512 252886 420465 252888
rect 412512 252830 420404 252886
rect 420460 252830 420465 252886
rect 412512 252828 420465 252830
rect 420399 252825 420465 252828
rect 40770 252298 40830 252562
rect 40762 252234 40768 252298
rect 40832 252234 40838 252298
rect 41722 252074 41728 252076
rect 41568 252014 41728 252074
rect 41722 252012 41728 252014
rect 41792 252012 41798 252076
rect 40570 251642 40576 251706
rect 40640 251642 40646 251706
rect 190191 251704 190257 251707
rect 190191 251702 191904 251704
rect 190191 251646 190196 251702
rect 190252 251646 191904 251702
rect 190191 251644 191904 251646
rect 40578 251526 40638 251642
rect 190191 251641 190257 251644
rect 40962 250818 41022 251082
rect 40954 250754 40960 250818
rect 41024 250754 41030 250818
rect 675759 250816 675825 250819
rect 676282 250816 676288 250818
rect 675759 250814 676288 250816
rect 675759 250758 675764 250814
rect 675820 250758 676288 250814
rect 675759 250756 676288 250758
rect 675759 250753 675825 250756
rect 676282 250754 676288 250756
rect 676352 250754 676358 250818
rect 420303 250520 420369 250523
rect 412512 250518 420369 250520
rect 41538 250374 41598 250490
rect 412512 250462 420308 250518
rect 420364 250462 420369 250518
rect 412512 250460 420369 250462
rect 420303 250457 420369 250460
rect 41530 250310 41536 250374
rect 41600 250310 41606 250374
rect 41775 250076 41841 250079
rect 41568 250074 41841 250076
rect 41568 250018 41780 250074
rect 41836 250018 41841 250074
rect 41568 250016 41841 250018
rect 41775 250013 41841 250016
rect 41914 249632 41920 249634
rect 41568 249572 41920 249632
rect 41914 249570 41920 249572
rect 41984 249570 41990 249634
rect 41154 248894 41214 249010
rect 41146 248830 41152 248894
rect 41216 248830 41222 248894
rect 41346 248302 41406 248492
rect 41338 248238 41344 248302
rect 41408 248238 41414 248302
rect 420399 248152 420465 248155
rect 412512 248150 420465 248152
rect 41538 247859 41598 248122
rect 412512 248094 420404 248150
rect 420460 248094 420465 248150
rect 412512 248092 420465 248094
rect 420399 248089 420465 248092
rect 41487 247854 41598 247859
rect 41487 247798 41492 247854
rect 41548 247798 41598 247854
rect 41487 247796 41598 247798
rect 41487 247793 41553 247796
rect 41538 247415 41598 247530
rect 41538 247410 41649 247415
rect 41538 247354 41588 247410
rect 41644 247354 41649 247410
rect 41538 247352 41649 247354
rect 41583 247349 41649 247352
rect 40386 246822 40446 247012
rect 40378 246758 40384 246822
rect 40448 246758 40454 246822
rect 41871 246672 41937 246675
rect 675567 246674 675633 246675
rect 41568 246670 41937 246672
rect 41568 246614 41876 246670
rect 41932 246614 41937 246670
rect 41568 246612 41937 246614
rect 41871 246609 41937 246612
rect 675514 246610 675520 246674
rect 675584 246672 675633 246674
rect 675584 246670 675676 246672
rect 675628 246614 675676 246670
rect 675584 246612 675676 246614
rect 675584 246610 675633 246612
rect 675567 246609 675633 246610
rect 41538 245932 41598 246050
rect 41679 245932 41745 245935
rect 41538 245930 41745 245932
rect 41538 245874 41684 245930
rect 41740 245874 41745 245930
rect 41538 245872 41745 245874
rect 41679 245869 41745 245872
rect 41538 245340 41598 245458
rect 41679 245340 41745 245343
rect 41538 245338 41745 245340
rect 41538 245282 41684 245338
rect 41740 245282 41745 245338
rect 41538 245280 41745 245282
rect 412482 245340 412542 245828
rect 420399 245340 420465 245343
rect 412482 245338 420465 245340
rect 412482 245282 420404 245338
rect 420460 245282 420465 245338
rect 412482 245280 420465 245282
rect 41679 245277 41745 245280
rect 420399 245277 420465 245280
rect 41538 244899 41598 245088
rect 41538 244894 41649 244899
rect 41538 244838 41588 244894
rect 41644 244838 41649 244894
rect 41538 244836 41649 244838
rect 41583 244833 41649 244836
rect 148335 244600 148401 244603
rect 143904 244598 148401 244600
rect 41538 244307 41598 244570
rect 143904 244542 148340 244598
rect 148396 244542 148401 244598
rect 143904 244540 148401 244542
rect 148335 244537 148401 244540
rect 41538 244302 41649 244307
rect 41538 244246 41588 244302
rect 41644 244246 41649 244302
rect 41538 244244 41649 244246
rect 41583 244241 41649 244244
rect 148527 243416 148593 243419
rect 143904 243414 148593 243416
rect 143904 243358 148532 243414
rect 148588 243358 148593 243414
rect 143904 243356 148593 243358
rect 148527 243353 148593 243356
rect 187119 243416 187185 243419
rect 191874 243416 191934 243904
rect 420303 243564 420369 243567
rect 412512 243562 420369 243564
rect 412512 243506 420308 243562
rect 420364 243506 420369 243562
rect 412512 243504 420369 243506
rect 420303 243501 420369 243504
rect 675663 243566 675729 243567
rect 675663 243562 675712 243566
rect 675776 243564 675782 243566
rect 675663 243506 675668 243562
rect 675663 243502 675712 243506
rect 675776 243504 675820 243564
rect 675776 243502 675782 243504
rect 675663 243501 675729 243502
rect 187119 243414 191934 243416
rect 187119 243358 187124 243414
rect 187180 243358 191934 243414
rect 187119 243356 191934 243358
rect 187119 243353 187185 243356
rect 143874 242084 143934 242128
rect 148719 242084 148785 242087
rect 143874 242082 148785 242084
rect 143874 242026 148724 242082
rect 148780 242026 148785 242082
rect 143874 242024 148785 242026
rect 148719 242021 148785 242024
rect 674554 242022 674560 242086
rect 674624 242084 674630 242086
rect 675375 242084 675441 242087
rect 674624 242082 675441 242084
rect 674624 242026 675380 242082
rect 675436 242026 675441 242082
rect 674624 242024 675441 242026
rect 674624 242022 674630 242024
rect 675375 242021 675441 242024
rect 674746 241726 674752 241790
rect 674816 241788 674822 241790
rect 675471 241788 675537 241791
rect 674816 241786 675537 241788
rect 674816 241730 675476 241786
rect 675532 241730 675537 241786
rect 674816 241728 675537 241730
rect 674816 241726 674822 241728
rect 675471 241725 675537 241728
rect 412431 241492 412497 241495
rect 567375 241492 567441 241495
rect 412431 241490 567441 241492
rect 412431 241434 412436 241490
rect 412492 241434 567380 241490
rect 567436 241434 567441 241490
rect 412431 241432 567441 241434
rect 412431 241429 412497 241432
rect 567375 241429 567441 241432
rect 420303 241196 420369 241199
rect 412512 241194 420369 241196
rect 412512 241138 420308 241194
rect 420364 241138 420369 241194
rect 412512 241136 420369 241138
rect 420303 241133 420369 241136
rect 149007 240900 149073 240903
rect 143904 240898 149073 240900
rect 143904 240842 149012 240898
rect 149068 240842 149073 240898
rect 143904 240840 149073 240842
rect 149007 240837 149073 240840
rect 412719 240900 412785 240903
rect 581775 240900 581841 240903
rect 412719 240898 581841 240900
rect 412719 240842 412724 240898
rect 412780 240842 581780 240898
rect 581836 240842 581841 240898
rect 412719 240840 581841 240842
rect 412719 240837 412785 240840
rect 581775 240837 581841 240840
rect 412239 240752 412305 240755
rect 566703 240752 566769 240755
rect 412239 240750 566769 240752
rect 412239 240694 412244 240750
rect 412300 240694 566708 240750
rect 566764 240694 566769 240750
rect 412239 240692 566769 240694
rect 412239 240689 412305 240692
rect 566703 240689 566769 240692
rect 412623 240604 412689 240607
rect 610479 240604 610545 240607
rect 412623 240602 610545 240604
rect 412623 240546 412628 240602
rect 412684 240546 610484 240602
rect 610540 240546 610545 240602
rect 412623 240544 610545 240546
rect 412623 240541 412689 240544
rect 610479 240541 610545 240544
rect 674938 240542 674944 240606
rect 675008 240604 675014 240606
rect 675471 240604 675537 240607
rect 675008 240602 675537 240604
rect 675008 240546 675476 240602
rect 675532 240546 675537 240602
rect 675008 240544 675537 240546
rect 675008 240542 675014 240544
rect 675471 240541 675537 240544
rect 412143 240456 412209 240459
rect 627183 240456 627249 240459
rect 412143 240454 627249 240456
rect 412143 240398 412148 240454
rect 412204 240398 627188 240454
rect 627244 240398 627249 240454
rect 412143 240396 627249 240398
rect 412143 240393 412209 240396
rect 627183 240393 627249 240396
rect 412047 240308 412113 240311
rect 544815 240308 544881 240311
rect 412047 240306 544881 240308
rect 412047 240250 412052 240306
rect 412108 240250 544820 240306
rect 544876 240250 544881 240306
rect 412047 240248 544881 240250
rect 412047 240245 412113 240248
rect 544815 240245 544881 240248
rect 412527 240160 412593 240163
rect 541455 240160 541521 240163
rect 412527 240158 541521 240160
rect 412527 240102 412532 240158
rect 412588 240102 541460 240158
rect 541516 240102 541521 240158
rect 412527 240100 541521 240102
rect 412527 240097 412593 240100
rect 541455 240097 541521 240100
rect 412335 240012 412401 240015
rect 550863 240012 550929 240015
rect 412335 240010 550929 240012
rect 412335 239954 412340 240010
rect 412396 239954 550868 240010
rect 550924 239954 550929 240010
rect 412335 239952 550929 239954
rect 412335 239949 412401 239952
rect 550863 239949 550929 239952
rect 148239 239716 148305 239719
rect 143904 239714 148305 239716
rect 143904 239658 148244 239714
rect 148300 239658 148305 239714
rect 143904 239656 148305 239658
rect 148239 239653 148305 239656
rect 413391 238976 413457 238979
rect 553935 238976 554001 238979
rect 413391 238974 554001 238976
rect 413391 238918 413396 238974
rect 413452 238918 553940 238974
rect 553996 238918 554001 238974
rect 413391 238916 554001 238918
rect 413391 238913 413457 238916
rect 553935 238913 554001 238916
rect 413679 238680 413745 238683
rect 550191 238680 550257 238683
rect 413679 238678 550257 238680
rect 413679 238622 413684 238678
rect 413740 238622 550196 238678
rect 550252 238622 550257 238678
rect 413679 238620 550257 238622
rect 413679 238617 413745 238620
rect 550191 238617 550257 238620
rect 675759 238680 675825 238683
rect 676090 238680 676096 238682
rect 675759 238678 676096 238680
rect 675759 238622 675764 238678
rect 675820 238622 676096 238678
rect 675759 238620 676096 238622
rect 675759 238617 675825 238620
rect 676090 238618 676096 238620
rect 676160 238618 676166 238682
rect 148815 238532 148881 238535
rect 143904 238530 148881 238532
rect 143904 238474 148820 238530
rect 148876 238474 148881 238530
rect 143904 238472 148881 238474
rect 148815 238469 148881 238472
rect 413967 238384 414033 238387
rect 544335 238384 544401 238387
rect 413967 238382 544401 238384
rect 413967 238326 413972 238382
rect 414028 238326 544340 238382
rect 544396 238326 544401 238382
rect 413967 238324 544401 238326
rect 413967 238321 414033 238324
rect 544335 238321 544401 238324
rect 414255 238236 414321 238239
rect 559887 238236 559953 238239
rect 414255 238234 559953 238236
rect 414255 238178 414260 238234
rect 414316 238178 559892 238234
rect 559948 238178 559953 238234
rect 414255 238176 559953 238178
rect 414255 238173 414321 238176
rect 559887 238173 559953 238176
rect 414447 238088 414513 238091
rect 537999 238088 538065 238091
rect 414447 238086 538065 238088
rect 414447 238030 414452 238086
rect 414508 238030 538004 238086
rect 538060 238030 538065 238086
rect 414447 238028 538065 238030
rect 414447 238025 414513 238028
rect 537999 238025 538065 238028
rect 41775 237942 41841 237943
rect 41722 237940 41728 237942
rect 41684 237880 41728 237940
rect 41792 237938 41841 237942
rect 41836 237882 41841 237938
rect 41722 237878 41728 237880
rect 41792 237878 41841 237882
rect 41775 237877 41841 237878
rect 40762 237138 40768 237202
rect 40832 237200 40838 237202
rect 41530 237200 41536 237202
rect 40832 237140 41536 237200
rect 40832 237138 40838 237140
rect 41530 237138 41536 237140
rect 41600 237138 41606 237202
rect 143874 236756 143934 237244
rect 372207 237052 372273 237055
rect 388719 237052 388785 237055
rect 398991 237052 399057 237055
rect 408687 237052 408753 237055
rect 372207 237050 388542 237052
rect 372207 236994 372212 237050
rect 372268 236994 388542 237050
rect 372207 236992 388542 236994
rect 372207 236989 372273 236992
rect 373455 236904 373521 236907
rect 387951 236904 388017 236907
rect 373455 236902 388017 236904
rect 373455 236846 373460 236902
rect 373516 236846 387956 236902
rect 388012 236846 388017 236902
rect 373455 236844 388017 236846
rect 373455 236841 373521 236844
rect 387951 236841 388017 236844
rect 148623 236756 148689 236759
rect 143874 236754 148689 236756
rect 143874 236698 148628 236754
rect 148684 236698 148689 236754
rect 143874 236696 148689 236698
rect 148623 236693 148689 236696
rect 370383 236756 370449 236759
rect 382575 236756 382641 236759
rect 370383 236754 382641 236756
rect 370383 236698 370388 236754
rect 370444 236698 382580 236754
rect 382636 236698 382641 236754
rect 370383 236696 382641 236698
rect 370383 236693 370449 236696
rect 382575 236693 382641 236696
rect 382767 236756 382833 236759
rect 388335 236756 388401 236759
rect 382767 236754 388401 236756
rect 382767 236698 382772 236754
rect 382828 236698 388340 236754
rect 388396 236698 388401 236754
rect 382767 236696 388401 236698
rect 388482 236756 388542 236992
rect 388719 237050 398910 237052
rect 388719 236994 388724 237050
rect 388780 236994 398910 237050
rect 388719 236992 398910 236994
rect 388719 236989 388785 236992
rect 388719 236904 388785 236907
rect 398703 236904 398769 236907
rect 388719 236902 398769 236904
rect 388719 236846 388724 236902
rect 388780 236846 398708 236902
rect 398764 236846 398769 236902
rect 388719 236844 398769 236846
rect 398850 236904 398910 236992
rect 398991 237050 408753 237052
rect 398991 236994 398996 237050
rect 399052 236994 408692 237050
rect 408748 236994 408753 237050
rect 398991 236992 408753 236994
rect 398991 236989 399057 236992
rect 408687 236989 408753 236992
rect 408879 237052 408945 237055
rect 573135 237052 573201 237055
rect 408879 237050 573201 237052
rect 408879 236994 408884 237050
rect 408940 236994 573140 237050
rect 573196 236994 573201 237050
rect 408879 236992 573201 236994
rect 408879 236989 408945 236992
rect 573135 236989 573201 236992
rect 408975 236904 409041 236907
rect 398850 236902 409041 236904
rect 398850 236846 408980 236902
rect 409036 236846 409041 236902
rect 398850 236844 409041 236846
rect 388719 236841 388785 236844
rect 398703 236841 398769 236844
rect 408975 236841 409041 236844
rect 409359 236904 409425 236907
rect 566031 236904 566097 236907
rect 409359 236902 566097 236904
rect 409359 236846 409364 236902
rect 409420 236846 566036 236902
rect 566092 236846 566097 236902
rect 409359 236844 566097 236846
rect 409359 236841 409425 236844
rect 566031 236841 566097 236844
rect 675759 236904 675825 236907
rect 675898 236904 675904 236906
rect 675759 236902 675904 236904
rect 675759 236846 675764 236902
rect 675820 236846 675904 236902
rect 675759 236844 675904 236846
rect 675759 236841 675825 236844
rect 675898 236842 675904 236844
rect 675968 236842 675974 236906
rect 408783 236756 408849 236759
rect 388482 236754 408849 236756
rect 388482 236698 408788 236754
rect 408844 236698 408849 236754
rect 388482 236696 408849 236698
rect 382767 236693 382833 236696
rect 388335 236693 388401 236696
rect 408783 236693 408849 236696
rect 409018 236694 409024 236758
rect 409088 236756 409094 236758
rect 562191 236756 562257 236759
rect 409088 236754 562257 236756
rect 409088 236698 562196 236754
rect 562252 236698 562257 236754
rect 409088 236696 562257 236698
rect 409088 236694 409094 236696
rect 562191 236693 562257 236696
rect 374895 236608 374961 236611
rect 559215 236608 559281 236611
rect 374895 236606 559281 236608
rect 374895 236550 374900 236606
rect 374956 236550 559220 236606
rect 559276 236550 559281 236606
rect 374895 236548 559281 236550
rect 374895 236545 374961 236548
rect 559215 236545 559281 236548
rect 376719 236460 376785 236463
rect 388623 236460 388689 236463
rect 557679 236460 557745 236463
rect 376719 236458 388542 236460
rect 376719 236402 376724 236458
rect 376780 236402 388542 236458
rect 376719 236400 388542 236402
rect 376719 236397 376785 236400
rect 368943 236312 369009 236315
rect 377775 236312 377841 236315
rect 368943 236310 377841 236312
rect 368943 236254 368948 236310
rect 369004 236254 377780 236310
rect 377836 236254 377841 236310
rect 368943 236252 377841 236254
rect 368943 236249 369009 236252
rect 377775 236249 377841 236252
rect 377967 236312 378033 236315
rect 388482 236312 388542 236400
rect 388623 236458 557745 236460
rect 388623 236402 388628 236458
rect 388684 236402 557684 236458
rect 557740 236402 557745 236458
rect 388623 236400 557745 236402
rect 388623 236397 388689 236400
rect 557679 236397 557745 236400
rect 388815 236312 388881 236315
rect 377967 236310 388350 236312
rect 377967 236254 377972 236310
rect 378028 236254 388350 236310
rect 377967 236252 388350 236254
rect 388482 236310 388881 236312
rect 388482 236254 388820 236310
rect 388876 236254 388881 236310
rect 388482 236252 388881 236254
rect 377967 236249 378033 236252
rect 388290 236164 388350 236252
rect 388815 236249 388881 236252
rect 389007 236312 389073 236315
rect 408687 236312 408753 236315
rect 389007 236310 408753 236312
rect 389007 236254 389012 236310
rect 389068 236254 408692 236310
rect 408748 236254 408753 236310
rect 389007 236252 408753 236254
rect 389007 236249 389073 236252
rect 408687 236249 408753 236252
rect 409167 236312 409233 236315
rect 414447 236312 414513 236315
rect 409167 236310 414513 236312
rect 409167 236254 409172 236310
rect 409228 236254 414452 236310
rect 414508 236254 414513 236310
rect 409167 236252 414513 236254
rect 409167 236249 409233 236252
rect 414447 236249 414513 236252
rect 414639 236312 414705 236315
rect 621135 236312 621201 236315
rect 414639 236310 621201 236312
rect 414639 236254 414644 236310
rect 414700 236254 621140 236310
rect 621196 236254 621201 236310
rect 414639 236252 621201 236254
rect 414639 236249 414705 236252
rect 621135 236249 621201 236252
rect 389007 236164 389073 236167
rect 408634 236164 408640 236166
rect 388290 236104 388926 236164
rect 149103 236016 149169 236019
rect 143904 236014 149169 236016
rect 143904 235958 149108 236014
rect 149164 235958 149169 236014
rect 143904 235956 149169 235958
rect 149103 235953 149169 235956
rect 342543 236016 342609 236019
rect 385935 236016 386001 236019
rect 342543 236014 386001 236016
rect 342543 235958 342548 236014
rect 342604 235958 385940 236014
rect 385996 235958 386001 236014
rect 342543 235956 386001 235958
rect 388866 236016 388926 236104
rect 389007 236162 408640 236164
rect 389007 236106 389012 236162
rect 389068 236106 408640 236162
rect 389007 236104 408640 236106
rect 389007 236101 389073 236104
rect 408634 236102 408640 236104
rect 408704 236102 408710 236166
rect 408783 236164 408849 236167
rect 593007 236164 593073 236167
rect 408783 236162 593073 236164
rect 408783 236106 408788 236162
rect 408844 236106 593012 236162
rect 593068 236106 593073 236162
rect 408783 236104 593073 236106
rect 408783 236101 408849 236104
rect 593007 236101 593073 236104
rect 389391 236016 389457 236019
rect 388866 236014 389457 236016
rect 388866 235958 389396 236014
rect 389452 235958 389457 236014
rect 388866 235956 389457 235958
rect 342543 235953 342609 235956
rect 385935 235953 386001 235956
rect 389391 235953 389457 235956
rect 403119 236016 403185 236019
rect 595887 236016 595953 236019
rect 403119 236014 595953 236016
rect 403119 235958 403124 236014
rect 403180 235958 595892 236014
rect 595948 235958 595953 236014
rect 403119 235956 595953 235958
rect 403119 235953 403185 235956
rect 595887 235953 595953 235956
rect 392559 235868 392625 235871
rect 393135 235868 393201 235871
rect 392559 235866 393201 235868
rect 392559 235810 392564 235866
rect 392620 235810 393140 235866
rect 393196 235810 393201 235866
rect 392559 235808 393201 235810
rect 392559 235805 392625 235808
rect 393135 235805 393201 235808
rect 401391 235868 401457 235871
rect 408783 235868 408849 235871
rect 401391 235866 408849 235868
rect 401391 235810 401396 235866
rect 401452 235810 408788 235866
rect 408844 235810 408849 235866
rect 401391 235808 408849 235810
rect 401391 235805 401457 235808
rect 408783 235805 408849 235808
rect 409018 235806 409024 235870
rect 409088 235868 409094 235870
rect 591471 235868 591537 235871
rect 409088 235866 591537 235868
rect 409088 235810 591476 235866
rect 591532 235810 591537 235866
rect 409088 235808 591537 235810
rect 409088 235806 409094 235808
rect 591471 235805 591537 235808
rect 354927 235720 354993 235723
rect 403311 235720 403377 235723
rect 354927 235718 403377 235720
rect 354927 235662 354932 235718
rect 354988 235662 403316 235718
rect 403372 235662 403377 235718
rect 354927 235660 403377 235662
rect 354927 235657 354993 235660
rect 403311 235657 403377 235660
rect 405519 235720 405585 235723
rect 597423 235720 597489 235723
rect 405519 235718 597489 235720
rect 405519 235662 405524 235718
rect 405580 235662 597428 235718
rect 597484 235662 597489 235718
rect 405519 235660 597489 235662
rect 405519 235657 405585 235660
rect 597423 235657 597489 235660
rect 385839 235572 385905 235575
rect 580335 235572 580401 235575
rect 385839 235570 580401 235572
rect 385839 235514 385844 235570
rect 385900 235514 580340 235570
rect 580396 235514 580401 235570
rect 385839 235512 580401 235514
rect 385839 235509 385905 235512
rect 580335 235509 580401 235512
rect 403983 235424 404049 235427
rect 596175 235424 596241 235427
rect 403983 235422 596241 235424
rect 403983 235366 403988 235422
rect 404044 235366 596180 235422
rect 596236 235366 596241 235422
rect 403983 235364 596241 235366
rect 403983 235361 404049 235364
rect 596175 235361 596241 235364
rect 387663 235276 387729 235279
rect 583407 235276 583473 235279
rect 387663 235274 583473 235276
rect 387663 235218 387668 235274
rect 387724 235218 583412 235274
rect 583468 235218 583473 235274
rect 387663 235216 583473 235218
rect 387663 235213 387729 235216
rect 583407 235213 583473 235216
rect 301647 235128 301713 235131
rect 344175 235128 344241 235131
rect 301647 235126 344241 235128
rect 301647 235070 301652 235126
rect 301708 235070 344180 235126
rect 344236 235070 344241 235126
rect 301647 235068 344241 235070
rect 301647 235065 301713 235068
rect 344175 235065 344241 235068
rect 344367 235128 344433 235131
rect 391791 235128 391857 235131
rect 344367 235126 391857 235128
rect 344367 235070 344372 235126
rect 344428 235070 391796 235126
rect 391852 235070 391857 235126
rect 344367 235068 391857 235070
rect 344367 235065 344433 235068
rect 391791 235065 391857 235068
rect 399855 235128 399921 235131
rect 408442 235128 408448 235130
rect 399855 235126 408448 235128
rect 399855 235070 399860 235126
rect 399916 235070 408448 235126
rect 399855 235068 408448 235070
rect 399855 235065 399921 235068
rect 408442 235066 408448 235068
rect 408512 235066 408518 235130
rect 595407 235128 595473 235131
rect 408642 235126 595473 235128
rect 408642 235070 595412 235126
rect 595468 235070 595473 235126
rect 408642 235068 595473 235070
rect 299343 234980 299409 234983
rect 349743 234980 349809 234983
rect 299343 234978 349809 234980
rect 299343 234922 299348 234978
rect 299404 234922 349748 234978
rect 349804 234922 349809 234978
rect 299343 234920 349809 234922
rect 299343 234917 299409 234920
rect 349743 234917 349809 234920
rect 393423 234980 393489 234983
rect 408642 234980 408702 235068
rect 595407 235065 595473 235068
rect 393423 234978 408702 234980
rect 393423 234922 393428 234978
rect 393484 234922 408702 234978
rect 393423 234920 408702 234922
rect 408783 234980 408849 234983
rect 594639 234980 594705 234983
rect 408783 234978 594705 234980
rect 408783 234922 408788 234978
rect 408844 234922 594644 234978
rect 594700 234922 594705 234978
rect 408783 234920 594705 234922
rect 393423 234917 393489 234920
rect 408783 234917 408849 234920
rect 594639 234917 594705 234920
rect 148431 234832 148497 234835
rect 143904 234830 148497 234832
rect 143904 234774 148436 234830
rect 148492 234774 148497 234830
rect 143904 234772 148497 234774
rect 148431 234769 148497 234772
rect 299439 234832 299505 234835
rect 354351 234832 354417 234835
rect 299439 234830 354417 234832
rect 299439 234774 299444 234830
rect 299500 234774 354356 234830
rect 354412 234774 354417 234830
rect 299439 234772 354417 234774
rect 299439 234769 299505 234772
rect 354351 234769 354417 234772
rect 356751 234832 356817 234835
rect 400431 234832 400497 234835
rect 356751 234830 400497 234832
rect 356751 234774 356756 234830
rect 356812 234774 400436 234830
rect 400492 234774 400497 234830
rect 356751 234772 400497 234774
rect 356751 234769 356817 234772
rect 400431 234769 400497 234772
rect 405423 234832 405489 234835
rect 618831 234832 618897 234835
rect 405423 234830 618897 234832
rect 405423 234774 405428 234830
rect 405484 234774 618836 234830
rect 618892 234774 618897 234830
rect 405423 234772 618897 234774
rect 405423 234769 405489 234772
rect 618831 234769 618897 234772
rect 298959 234684 299025 234687
rect 354255 234684 354321 234687
rect 298959 234682 354321 234684
rect 298959 234626 298964 234682
rect 299020 234626 354260 234682
rect 354316 234626 354321 234682
rect 298959 234624 354321 234626
rect 298959 234621 299025 234624
rect 354255 234621 354321 234624
rect 356847 234684 356913 234687
rect 392847 234684 392913 234687
rect 356847 234682 392913 234684
rect 356847 234626 356852 234682
rect 356908 234626 392852 234682
rect 392908 234626 392913 234682
rect 356847 234624 392913 234626
rect 356847 234621 356913 234624
rect 392847 234621 392913 234624
rect 393039 234684 393105 234687
rect 407919 234684 407985 234687
rect 393039 234682 407985 234684
rect 393039 234626 393044 234682
rect 393100 234626 407924 234682
rect 407980 234626 407985 234682
rect 393039 234624 407985 234626
rect 393039 234621 393105 234624
rect 407919 234621 407985 234624
rect 408111 234684 408177 234687
rect 624879 234684 624945 234687
rect 408111 234682 624945 234684
rect 408111 234626 408116 234682
rect 408172 234626 624884 234682
rect 624940 234626 624945 234682
rect 408111 234624 624945 234626
rect 408111 234621 408177 234624
rect 624879 234621 624945 234624
rect 341583 234536 341649 234539
rect 490479 234536 490545 234539
rect 341583 234534 490545 234536
rect 341583 234478 341588 234534
rect 341644 234478 490484 234534
rect 490540 234478 490545 234534
rect 341583 234476 490545 234478
rect 341583 234473 341649 234476
rect 490479 234473 490545 234476
rect 379119 234388 379185 234391
rect 392559 234388 392625 234391
rect 379119 234386 392625 234388
rect 379119 234330 379124 234386
rect 379180 234330 392564 234386
rect 392620 234330 392625 234386
rect 379119 234328 392625 234330
rect 379119 234325 379185 234328
rect 392559 234325 392625 234328
rect 392847 234388 392913 234391
rect 405711 234388 405777 234391
rect 392847 234386 405777 234388
rect 392847 234330 392852 234386
rect 392908 234330 405716 234386
rect 405772 234330 405777 234386
rect 392847 234328 405777 234330
rect 392847 234325 392913 234328
rect 405711 234325 405777 234328
rect 408495 234388 408561 234391
rect 512175 234388 512241 234391
rect 408495 234386 512241 234388
rect 408495 234330 408500 234386
rect 408556 234330 512180 234386
rect 512236 234330 512241 234386
rect 408495 234328 512241 234330
rect 408495 234325 408561 234328
rect 512175 234325 512241 234328
rect 367215 234240 367281 234243
rect 405903 234240 405969 234243
rect 367215 234238 405969 234240
rect 367215 234182 367220 234238
rect 367276 234182 405908 234238
rect 405964 234182 405969 234238
rect 367215 234180 405969 234182
rect 367215 234177 367281 234180
rect 405903 234177 405969 234180
rect 407247 234240 407313 234243
rect 495375 234240 495441 234243
rect 407247 234238 495441 234240
rect 407247 234182 407252 234238
rect 407308 234182 495380 234238
rect 495436 234182 495441 234238
rect 407247 234180 495441 234182
rect 407247 234177 407313 234180
rect 495375 234177 495441 234180
rect 370287 234092 370353 234095
rect 428271 234092 428337 234095
rect 370287 234090 428337 234092
rect 370287 234034 370292 234090
rect 370348 234034 428276 234090
rect 428332 234034 428337 234090
rect 370287 234032 428337 234034
rect 370287 234029 370353 234032
rect 428271 234029 428337 234032
rect 376335 233944 376401 233947
rect 414255 233944 414321 233947
rect 376335 233942 414321 233944
rect 376335 233886 376340 233942
rect 376396 233886 414260 233942
rect 414316 233886 414321 233942
rect 376335 233884 414321 233886
rect 376335 233881 376401 233884
rect 414255 233881 414321 233884
rect 347631 233796 347697 233799
rect 411567 233796 411633 233799
rect 347631 233794 411633 233796
rect 347631 233738 347636 233794
rect 347692 233738 411572 233794
rect 411628 233738 411633 233794
rect 347631 233736 411633 233738
rect 347631 233733 347697 233736
rect 411567 233733 411633 233736
rect 148911 233648 148977 233651
rect 143904 233646 148977 233648
rect 143904 233590 148916 233646
rect 148972 233590 148977 233646
rect 143904 233588 148977 233590
rect 148911 233585 148977 233588
rect 392559 233648 392625 233651
rect 406959 233648 407025 233651
rect 392559 233646 407025 233648
rect 392559 233590 392564 233646
rect 392620 233590 406964 233646
rect 407020 233590 407025 233646
rect 392559 233588 407025 233590
rect 392559 233585 392625 233588
rect 406959 233585 407025 233588
rect 41775 233354 41841 233355
rect 41722 233352 41728 233354
rect 41684 233292 41728 233352
rect 41792 233350 41841 233354
rect 41836 233294 41841 233350
rect 41722 233290 41728 233292
rect 41792 233290 41841 233294
rect 41775 233289 41841 233290
rect 330255 233204 330321 233207
rect 470127 233204 470193 233207
rect 330255 233202 470193 233204
rect 330255 233146 330260 233202
rect 330316 233146 470132 233202
rect 470188 233146 470193 233202
rect 330255 233144 470193 233146
rect 330255 233141 330321 233144
rect 470127 233141 470193 233144
rect 334863 233056 334929 233059
rect 479151 233056 479217 233059
rect 334863 233054 479217 233056
rect 334863 232998 334868 233054
rect 334924 232998 479156 233054
rect 479212 232998 479217 233054
rect 334863 232996 479217 232998
rect 334863 232993 334929 232996
rect 479151 232993 479217 232996
rect 359055 232908 359121 232911
rect 525231 232908 525297 232911
rect 359055 232906 525297 232908
rect 359055 232850 359060 232906
rect 359116 232850 525236 232906
rect 525292 232850 525297 232906
rect 359055 232848 525297 232850
rect 359055 232845 359121 232848
rect 525231 232845 525297 232848
rect 370767 232760 370833 232763
rect 551631 232760 551697 232763
rect 370767 232758 551697 232760
rect 370767 232702 370772 232758
rect 370828 232702 551636 232758
rect 551692 232702 551697 232758
rect 370767 232700 551697 232702
rect 370767 232697 370833 232700
rect 551631 232697 551697 232700
rect 375375 232612 375441 232615
rect 560751 232612 560817 232615
rect 375375 232610 560817 232612
rect 375375 232554 375380 232610
rect 375436 232554 560756 232610
rect 560812 232554 560817 232610
rect 375375 232552 560817 232554
rect 375375 232549 375441 232552
rect 560751 232549 560817 232552
rect 378927 232464 378993 232467
rect 564495 232464 564561 232467
rect 378927 232462 564561 232464
rect 378927 232406 378932 232462
rect 378988 232406 564500 232462
rect 564556 232406 564561 232462
rect 378927 232404 564561 232406
rect 378927 232401 378993 232404
rect 564495 232401 564561 232404
rect 147663 232316 147729 232319
rect 143904 232314 147729 232316
rect 143904 232258 147668 232314
rect 147724 232258 147729 232314
rect 143904 232256 147729 232258
rect 147663 232253 147729 232256
rect 381711 232316 381777 232319
rect 570447 232316 570513 232319
rect 381711 232314 570513 232316
rect 381711 232258 381716 232314
rect 381772 232258 570452 232314
rect 570508 232258 570513 232314
rect 381711 232256 570513 232258
rect 381711 232253 381777 232256
rect 570447 232253 570513 232256
rect 384975 232168 385041 232171
rect 576591 232168 576657 232171
rect 384975 232166 576657 232168
rect 384975 232110 384980 232166
rect 385036 232110 576596 232166
rect 576652 232110 576657 232166
rect 384975 232108 576657 232110
rect 384975 232105 385041 232108
rect 576591 232105 576657 232108
rect 385359 232020 385425 232023
rect 578031 232020 578097 232023
rect 385359 232018 578097 232020
rect 385359 231962 385364 232018
rect 385420 231962 578036 232018
rect 578092 231962 578097 232018
rect 385359 231960 578097 231962
rect 385359 231957 385425 231960
rect 578031 231957 578097 231960
rect 382959 231872 383025 231875
rect 575823 231872 575889 231875
rect 382959 231870 575889 231872
rect 382959 231814 382964 231870
rect 383020 231814 575828 231870
rect 575884 231814 575889 231870
rect 382959 231812 575889 231814
rect 382959 231809 383025 231812
rect 575823 231809 575889 231812
rect 322479 231724 322545 231727
rect 455151 231724 455217 231727
rect 322479 231722 455217 231724
rect 322479 231666 322484 231722
rect 322540 231666 455156 231722
rect 455212 231666 455217 231722
rect 322479 231664 455217 231666
rect 322479 231661 322545 231664
rect 455151 231661 455217 231664
rect 319503 231576 319569 231579
rect 448911 231576 448977 231579
rect 319503 231574 448977 231576
rect 319503 231518 319508 231574
rect 319564 231518 448916 231574
rect 448972 231518 448977 231574
rect 319503 231516 448977 231518
rect 319503 231513 319569 231516
rect 448911 231513 448977 231516
rect 316719 231428 316785 231431
rect 442863 231428 442929 231431
rect 316719 231426 442929 231428
rect 316719 231370 316724 231426
rect 316780 231370 442868 231426
rect 442924 231370 442929 231426
rect 316719 231368 442929 231370
rect 316719 231365 316785 231368
rect 442863 231365 442929 231368
rect 307599 231280 307665 231283
rect 424719 231280 424785 231283
rect 307599 231278 424785 231280
rect 307599 231222 307604 231278
rect 307660 231222 424724 231278
rect 424780 231222 424785 231278
rect 307599 231220 424785 231222
rect 307599 231217 307665 231220
rect 424719 231217 424785 231220
rect 40378 231070 40384 231134
rect 40448 231132 40454 231134
rect 41775 231132 41841 231135
rect 149391 231132 149457 231135
rect 40448 231130 41841 231132
rect 40448 231074 41780 231130
rect 41836 231074 41841 231130
rect 40448 231072 41841 231074
rect 143904 231130 149457 231132
rect 143904 231074 149396 231130
rect 149452 231074 149457 231130
rect 143904 231072 149457 231074
rect 40448 231070 40454 231072
rect 41775 231069 41841 231072
rect 149391 231069 149457 231072
rect 302895 231132 302961 231135
rect 415695 231132 415761 231135
rect 302895 231130 415761 231132
rect 302895 231074 302900 231130
rect 302956 231074 415700 231130
rect 415756 231074 415761 231130
rect 302895 231072 415761 231074
rect 302895 231069 302961 231072
rect 415695 231069 415761 231072
rect 41338 230330 41344 230394
rect 41408 230392 41414 230394
rect 41775 230392 41841 230395
rect 41408 230390 41841 230392
rect 41408 230334 41780 230390
rect 41836 230334 41841 230390
rect 41408 230332 41841 230334
rect 41408 230330 41414 230332
rect 41775 230329 41841 230332
rect 342159 230392 342225 230395
rect 494223 230392 494289 230395
rect 342159 230390 494289 230392
rect 342159 230334 342164 230390
rect 342220 230334 494228 230390
rect 494284 230334 494289 230390
rect 342159 230332 494289 230334
rect 342159 230329 342225 230332
rect 494223 230329 494289 230332
rect 345519 230244 345585 230247
rect 497967 230244 498033 230247
rect 345519 230242 498033 230244
rect 345519 230186 345524 230242
rect 345580 230186 497972 230242
rect 498028 230186 498033 230242
rect 345519 230184 498033 230186
rect 345519 230181 345585 230184
rect 497967 230181 498033 230184
rect 363567 230096 363633 230099
rect 534255 230096 534321 230099
rect 363567 230094 534321 230096
rect 363567 230038 363572 230094
rect 363628 230038 534260 230094
rect 534316 230038 534321 230094
rect 363567 230036 534321 230038
rect 363567 230033 363633 230036
rect 534255 230033 534321 230036
rect 146895 229948 146961 229951
rect 143904 229946 146961 229948
rect 143904 229890 146900 229946
rect 146956 229890 146961 229946
rect 143904 229888 146961 229890
rect 146895 229885 146961 229888
rect 358959 229948 359025 229951
rect 527535 229948 527601 229951
rect 358959 229946 527601 229948
rect 358959 229890 358964 229946
rect 359020 229890 527540 229946
rect 527596 229890 527601 229946
rect 358959 229888 527601 229890
rect 358959 229885 359025 229888
rect 527535 229885 527601 229888
rect 365775 229800 365841 229803
rect 538863 229800 538929 229803
rect 365775 229798 538929 229800
rect 365775 229742 365780 229798
rect 365836 229742 538868 229798
rect 538924 229742 538929 229798
rect 365775 229740 538929 229742
rect 365775 229737 365841 229740
rect 538863 229737 538929 229740
rect 41146 229590 41152 229654
rect 41216 229652 41222 229654
rect 41775 229652 41841 229655
rect 41216 229650 41841 229652
rect 41216 229594 41780 229650
rect 41836 229594 41841 229650
rect 41216 229592 41841 229594
rect 41216 229590 41222 229592
rect 41775 229589 41841 229592
rect 373071 229652 373137 229655
rect 553935 229652 554001 229655
rect 373071 229650 554001 229652
rect 373071 229594 373076 229650
rect 373132 229594 553940 229650
rect 553996 229594 554001 229650
rect 373071 229592 554001 229594
rect 373071 229589 373137 229592
rect 553935 229589 554001 229592
rect 383535 229504 383601 229507
rect 573519 229504 573585 229507
rect 383535 229502 573585 229504
rect 383535 229446 383540 229502
rect 383596 229446 573524 229502
rect 573580 229446 573585 229502
rect 383535 229444 573585 229446
rect 383535 229441 383601 229444
rect 573519 229441 573585 229444
rect 381327 229356 381393 229359
rect 572751 229356 572817 229359
rect 381327 229354 572817 229356
rect 381327 229298 381332 229354
rect 381388 229298 572756 229354
rect 572812 229298 572817 229354
rect 381327 229296 572817 229298
rect 381327 229293 381393 229296
rect 572751 229293 572817 229296
rect 384399 229208 384465 229211
rect 578895 229208 578961 229211
rect 384399 229206 578961 229208
rect 384399 229150 384404 229206
rect 384460 229150 578900 229206
rect 578956 229150 578961 229206
rect 384399 229148 578961 229150
rect 384399 229145 384465 229148
rect 578895 229145 578961 229148
rect 40954 228998 40960 229062
rect 41024 229060 41030 229062
rect 41775 229060 41841 229063
rect 41024 229058 41841 229060
rect 41024 229002 41780 229058
rect 41836 229002 41841 229058
rect 41024 229000 41841 229002
rect 41024 228998 41030 229000
rect 41775 228997 41841 229000
rect 403119 229060 403185 229063
rect 599919 229060 599985 229063
rect 403119 229058 599985 229060
rect 403119 229002 403124 229058
rect 403180 229002 599924 229058
rect 599980 229002 599985 229058
rect 403119 229000 599985 229002
rect 403119 228997 403185 229000
rect 599919 228997 599985 229000
rect 292143 228912 292209 228915
rect 359823 228912 359889 228915
rect 292143 228910 359889 228912
rect 292143 228854 292148 228910
rect 292204 228854 359828 228910
rect 359884 228854 359889 228910
rect 292143 228852 359889 228854
rect 292143 228849 292209 228852
rect 359823 228849 359889 228852
rect 399471 228912 399537 228915
rect 607503 228912 607569 228915
rect 399471 228910 607569 228912
rect 399471 228854 399476 228910
rect 399532 228854 607508 228910
rect 607564 228854 607569 228910
rect 399471 228852 607569 228854
rect 399471 228849 399537 228852
rect 607503 228849 607569 228852
rect 339375 228764 339441 228767
rect 488271 228764 488337 228767
rect 339375 228762 488337 228764
rect 339375 228706 339380 228762
rect 339436 228706 488276 228762
rect 488332 228706 488337 228762
rect 339375 228704 488337 228706
rect 339375 228701 339441 228704
rect 488271 228701 488337 228704
rect 143874 228172 143934 228660
rect 333039 228616 333105 228619
rect 476175 228616 476241 228619
rect 333039 228614 476241 228616
rect 333039 228558 333044 228614
rect 333100 228558 476180 228614
rect 476236 228558 476241 228614
rect 333039 228556 476241 228558
rect 333039 228553 333105 228556
rect 476175 228553 476241 228556
rect 313455 228468 313521 228471
rect 436911 228468 436977 228471
rect 313455 228466 436977 228468
rect 313455 228410 313460 228466
rect 313516 228410 436916 228466
rect 436972 228410 436977 228466
rect 313455 228408 436977 228410
rect 313455 228405 313521 228408
rect 436911 228405 436977 228408
rect 310671 228320 310737 228323
rect 430863 228320 430929 228323
rect 310671 228318 430929 228320
rect 310671 228262 310676 228318
rect 310732 228262 430868 228318
rect 430924 228262 430929 228318
rect 310671 228260 430929 228262
rect 310671 228257 310737 228260
rect 430863 228257 430929 228260
rect 149391 228172 149457 228175
rect 143874 228170 149457 228172
rect 143874 228114 149396 228170
rect 149452 228114 149457 228170
rect 143874 228112 149457 228114
rect 149391 228109 149457 228112
rect 41530 227370 41536 227434
rect 41600 227432 41606 227434
rect 41775 227432 41841 227435
rect 149295 227432 149361 227435
rect 41600 227430 41841 227432
rect 41600 227374 41780 227430
rect 41836 227374 41841 227430
rect 41600 227372 41841 227374
rect 143904 227430 149361 227432
rect 143904 227374 149300 227430
rect 149356 227374 149361 227430
rect 143904 227372 149361 227374
rect 41600 227370 41606 227372
rect 41775 227369 41841 227372
rect 149295 227369 149361 227372
rect 330831 227432 330897 227435
rect 469359 227432 469425 227435
rect 330831 227430 469425 227432
rect 330831 227374 330836 227430
rect 330892 227374 469364 227430
rect 469420 227374 469425 227430
rect 330831 227372 469425 227374
rect 330831 227369 330897 227372
rect 469359 227369 469425 227372
rect 333807 227284 333873 227287
rect 475311 227284 475377 227287
rect 333807 227282 475377 227284
rect 333807 227226 333812 227282
rect 333868 227226 475316 227282
rect 475372 227226 475377 227282
rect 333807 227224 475377 227226
rect 333807 227221 333873 227224
rect 475311 227221 475377 227224
rect 336879 227136 336945 227139
rect 481455 227136 481521 227139
rect 336879 227134 481521 227136
rect 336879 227078 336884 227134
rect 336940 227078 481460 227134
rect 481516 227078 481521 227134
rect 336879 227076 481521 227078
rect 336879 227073 336945 227076
rect 481455 227073 481521 227076
rect 343023 226988 343089 226991
rect 493455 226988 493521 226991
rect 343023 226986 493521 226988
rect 343023 226930 343028 226986
rect 343084 226930 493460 226986
rect 493516 226930 493521 226986
rect 343023 226928 493521 226930
rect 343023 226925 343089 226928
rect 493455 226925 493521 226928
rect 41871 226842 41937 226843
rect 41871 226838 41920 226842
rect 41984 226840 41990 226842
rect 344751 226840 344817 226843
rect 498831 226840 498897 226843
rect 41871 226782 41876 226838
rect 41871 226778 41920 226782
rect 41984 226780 42028 226840
rect 344751 226838 498897 226840
rect 344751 226782 344756 226838
rect 344812 226782 498836 226838
rect 498892 226782 498897 226838
rect 344751 226780 498897 226782
rect 41984 226778 41990 226780
rect 41871 226777 41937 226778
rect 344751 226777 344817 226780
rect 498831 226777 498897 226780
rect 391599 226692 391665 226695
rect 591663 226692 591729 226695
rect 391599 226690 591729 226692
rect 391599 226634 391604 226690
rect 391660 226634 591668 226690
rect 591724 226634 591729 226690
rect 391599 226632 591729 226634
rect 391599 226629 391665 226632
rect 591663 226629 591729 226632
rect 394479 226544 394545 226547
rect 596943 226544 597009 226547
rect 394479 226542 597009 226544
rect 394479 226486 394484 226542
rect 394540 226486 596948 226542
rect 597004 226486 597009 226542
rect 394479 226484 597009 226486
rect 394479 226481 394545 226484
rect 596943 226481 597009 226484
rect 149391 226396 149457 226399
rect 143904 226394 149457 226396
rect 143904 226338 149396 226394
rect 149452 226338 149457 226394
rect 143904 226336 149457 226338
rect 149391 226333 149457 226336
rect 394095 226396 394161 226399
rect 596175 226396 596241 226399
rect 394095 226394 596241 226396
rect 394095 226338 394100 226394
rect 394156 226338 596180 226394
rect 596236 226338 596241 226394
rect 394095 226336 596241 226338
rect 394095 226333 394161 226336
rect 596175 226333 596241 226336
rect 405807 226248 405873 226251
rect 620367 226248 620433 226251
rect 405807 226246 620433 226248
rect 405807 226190 405812 226246
rect 405868 226190 620372 226246
rect 620428 226190 620433 226246
rect 405807 226188 620433 226190
rect 405807 226185 405873 226188
rect 620367 226185 620433 226188
rect 407631 226100 407697 226103
rect 623343 226100 623409 226103
rect 407631 226098 623409 226100
rect 407631 226042 407636 226098
rect 407692 226042 623348 226098
rect 623404 226042 623409 226098
rect 407631 226040 623409 226042
rect 407631 226037 407697 226040
rect 623343 226037 623409 226040
rect 40570 225890 40576 225954
rect 40640 225952 40646 225954
rect 41775 225952 41841 225955
rect 40640 225950 41841 225952
rect 40640 225894 41780 225950
rect 41836 225894 41841 225950
rect 40640 225892 41841 225894
rect 40640 225890 40646 225892
rect 41775 225889 41841 225892
rect 351375 225952 351441 225955
rect 487503 225952 487569 225955
rect 351375 225950 487569 225952
rect 351375 225894 351380 225950
rect 351436 225894 487508 225950
rect 487564 225894 487569 225950
rect 351375 225892 487569 225894
rect 351375 225889 351441 225892
rect 487503 225889 487569 225892
rect 328047 225804 328113 225807
rect 463311 225804 463377 225807
rect 328047 225802 463377 225804
rect 328047 225746 328052 225802
rect 328108 225746 463316 225802
rect 463372 225746 463377 225802
rect 328047 225744 463377 225746
rect 328047 225741 328113 225744
rect 463311 225741 463377 225744
rect 321711 225656 321777 225659
rect 451215 225656 451281 225659
rect 321711 225654 451281 225656
rect 321711 225598 321716 225654
rect 321772 225598 451220 225654
rect 451276 225598 451281 225654
rect 321711 225596 451281 225598
rect 321711 225593 321777 225596
rect 451215 225593 451281 225596
rect 318927 225508 318993 225511
rect 445167 225508 445233 225511
rect 318927 225506 445233 225508
rect 318927 225450 318932 225506
rect 318988 225450 445172 225506
rect 445228 225450 445233 225506
rect 318927 225448 445233 225450
rect 318927 225445 318993 225448
rect 445167 225445 445233 225448
rect 342639 225360 342705 225363
rect 457263 225360 457329 225363
rect 342639 225358 457329 225360
rect 342639 225302 342644 225358
rect 342700 225302 457268 225358
rect 457324 225302 457329 225358
rect 342639 225300 457329 225302
rect 342639 225297 342705 225300
rect 457263 225297 457329 225300
rect 149487 225212 149553 225215
rect 143904 225210 149553 225212
rect 143904 225154 149492 225210
rect 149548 225154 149553 225210
rect 143904 225152 149553 225154
rect 149487 225149 149553 225152
rect 354159 224620 354225 224623
rect 518415 224620 518481 224623
rect 354159 224618 518481 224620
rect 354159 224562 354164 224618
rect 354220 224562 518420 224618
rect 518476 224562 518481 224618
rect 354159 224560 518481 224562
rect 354159 224557 354225 224560
rect 518415 224557 518481 224560
rect 357519 224472 357585 224475
rect 524463 224472 524529 224475
rect 357519 224470 524529 224472
rect 357519 224414 357524 224470
rect 357580 224414 524468 224470
rect 524524 224414 524529 224470
rect 357519 224412 524529 224414
rect 357519 224409 357585 224412
rect 524463 224409 524529 224412
rect 359727 224324 359793 224327
rect 528975 224324 529041 224327
rect 359727 224322 529041 224324
rect 359727 224266 359732 224322
rect 359788 224266 528980 224322
rect 529036 224266 529041 224322
rect 359727 224264 529041 224266
rect 359727 224261 359793 224264
rect 528975 224261 529041 224264
rect 361455 224176 361521 224179
rect 532047 224176 532113 224179
rect 361455 224174 532113 224176
rect 361455 224118 361460 224174
rect 361516 224118 532052 224174
rect 532108 224118 532113 224174
rect 361455 224116 532113 224118
rect 361455 224113 361521 224116
rect 532047 224113 532113 224116
rect 360303 224028 360369 224031
rect 530511 224028 530577 224031
rect 360303 224026 530577 224028
rect 360303 223970 360308 224026
rect 360364 223970 530516 224026
rect 530572 223970 530577 224026
rect 360303 223968 530577 223970
rect 360303 223965 360369 223968
rect 530511 223965 530577 223968
rect 149487 223880 149553 223883
rect 143904 223878 149553 223880
rect 143904 223822 149492 223878
rect 149548 223822 149553 223878
rect 143904 223820 149553 223822
rect 149487 223817 149553 223820
rect 363471 223880 363537 223883
rect 536559 223880 536625 223883
rect 363471 223878 536625 223880
rect 363471 223822 363476 223878
rect 363532 223822 536564 223878
rect 536620 223822 536625 223878
rect 363471 223820 536625 223822
rect 363471 223817 363537 223820
rect 536559 223817 536625 223820
rect 367599 223732 367665 223735
rect 544047 223732 544113 223735
rect 367599 223730 544113 223732
rect 367599 223674 367604 223730
rect 367660 223674 544052 223730
rect 544108 223674 544113 223730
rect 367599 223672 544113 223674
rect 367599 223669 367665 223672
rect 544047 223669 544113 223672
rect 377583 223584 377649 223587
rect 562959 223584 563025 223587
rect 377583 223582 563025 223584
rect 377583 223526 377588 223582
rect 377644 223526 562964 223582
rect 563020 223526 563025 223582
rect 377583 223524 563025 223526
rect 377583 223521 377649 223524
rect 562959 223521 563025 223524
rect 381231 223436 381297 223439
rect 571311 223436 571377 223439
rect 381231 223434 571377 223436
rect 381231 223378 381236 223434
rect 381292 223378 571316 223434
rect 571372 223378 571377 223434
rect 381231 223376 571377 223378
rect 381231 223373 381297 223376
rect 571311 223373 571377 223376
rect 379791 223288 379857 223291
rect 568239 223288 568305 223291
rect 379791 223286 568305 223288
rect 379791 223230 379796 223286
rect 379852 223230 568244 223286
rect 568300 223230 568305 223286
rect 379791 223228 568305 223230
rect 379791 223225 379857 223228
rect 568239 223225 568305 223228
rect 384303 223140 384369 223143
rect 577263 223140 577329 223143
rect 384303 223138 577329 223140
rect 384303 223082 384308 223138
rect 384364 223082 577268 223138
rect 577324 223082 577329 223138
rect 384303 223080 577329 223082
rect 384303 223077 384369 223080
rect 577263 223077 577329 223080
rect 359439 222992 359505 222995
rect 526671 222992 526737 222995
rect 359439 222990 526737 222992
rect 359439 222934 359444 222990
rect 359500 222934 526676 222990
rect 526732 222934 526737 222990
rect 359439 222932 526737 222934
rect 359439 222929 359505 222932
rect 526671 222929 526737 222932
rect 382767 222844 382833 222847
rect 541071 222844 541137 222847
rect 382767 222842 541137 222844
rect 382767 222786 382772 222842
rect 382828 222786 541076 222842
rect 541132 222786 541137 222842
rect 382767 222784 541137 222786
rect 382767 222781 382833 222784
rect 541071 222781 541137 222784
rect 149391 222696 149457 222699
rect 143904 222694 149457 222696
rect 143904 222638 149396 222694
rect 149452 222638 149457 222694
rect 143904 222636 149457 222638
rect 149391 222633 149457 222636
rect 405711 222696 405777 222699
rect 522927 222696 522993 222699
rect 405711 222694 522993 222696
rect 405711 222638 405716 222694
rect 405772 222638 522932 222694
rect 522988 222638 522993 222694
rect 405711 222636 522993 222638
rect 405711 222633 405777 222636
rect 522927 222633 522993 222636
rect 676290 222107 676350 222222
rect 676239 222102 676350 222107
rect 676239 222046 676244 222102
rect 676300 222046 676350 222102
rect 676239 222044 676350 222046
rect 676239 222041 676305 222044
rect 676239 221956 676305 221959
rect 676239 221954 676350 221956
rect 676239 221898 676244 221954
rect 676300 221898 676350 221954
rect 676239 221893 676350 221898
rect 676290 221778 676350 221893
rect 149487 221512 149553 221515
rect 143904 221510 149553 221512
rect 143904 221454 149492 221510
rect 149548 221454 149553 221510
rect 143904 221452 149553 221454
rect 149487 221449 149553 221452
rect 676047 221216 676113 221219
rect 676047 221214 676320 221216
rect 676047 221158 676052 221214
rect 676108 221158 676320 221214
rect 676047 221156 676320 221158
rect 676047 221153 676113 221156
rect 186831 221068 186897 221071
rect 186831 221066 190560 221068
rect 186831 221010 186836 221066
rect 186892 221010 190560 221066
rect 186831 221008 190560 221010
rect 186831 221005 186897 221008
rect 673978 220710 673984 220774
rect 674048 220772 674054 220774
rect 674048 220712 676320 220772
rect 674048 220710 674054 220712
rect 187023 220328 187089 220331
rect 187023 220326 190560 220328
rect 187023 220270 187028 220326
rect 187084 220270 190560 220326
rect 187023 220268 190560 220270
rect 187023 220265 187089 220268
rect 143874 219736 143934 220224
rect 149391 219736 149457 219739
rect 143874 219734 149457 219736
rect 143874 219678 149396 219734
rect 149452 219678 149457 219734
rect 143874 219676 149457 219678
rect 149391 219673 149457 219676
rect 184335 219588 184401 219591
rect 184335 219586 190560 219588
rect 184335 219530 184340 219586
rect 184396 219530 190560 219586
rect 184335 219528 190560 219530
rect 184335 219525 184401 219528
rect 147663 218996 147729 218999
rect 143904 218994 147729 218996
rect 143904 218938 147668 218994
rect 147724 218938 147729 218994
rect 143904 218936 147729 218938
rect 147663 218933 147729 218936
rect 184335 218848 184401 218851
rect 184335 218846 190560 218848
rect 184335 218790 184340 218846
rect 184396 218790 190560 218846
rect 184335 218788 190560 218790
rect 184335 218785 184401 218788
rect 639810 218670 639870 220594
rect 674362 219970 674368 220034
rect 674432 220032 674438 220034
rect 676290 220032 676350 220224
rect 674432 219972 676350 220032
rect 674432 219970 674438 219972
rect 676239 219884 676305 219887
rect 676239 219882 676350 219884
rect 676239 219826 676244 219882
rect 676300 219826 676350 219882
rect 676239 219821 676350 219826
rect 676290 219706 676350 219821
rect 672975 219292 673041 219295
rect 673978 219292 673984 219294
rect 672975 219290 673984 219292
rect 672975 219234 672980 219290
rect 673036 219234 673984 219290
rect 672975 219232 673984 219234
rect 672975 219229 673041 219232
rect 673978 219230 673984 219232
rect 674048 219292 674054 219294
rect 674048 219232 676320 219292
rect 674048 219230 674054 219232
rect 676047 218774 676113 218777
rect 676047 218772 676320 218774
rect 676047 218716 676052 218772
rect 676108 218716 676320 218772
rect 676047 218714 676320 218716
rect 676047 218711 676113 218714
rect 672783 218256 672849 218259
rect 674170 218256 674176 218258
rect 672783 218254 674176 218256
rect 672783 218198 672788 218254
rect 672844 218198 674176 218254
rect 672783 218196 674176 218198
rect 672783 218193 672849 218196
rect 674170 218194 674176 218196
rect 674240 218256 674246 218258
rect 674240 218196 676320 218256
rect 674240 218194 674246 218196
rect 186927 218108 186993 218111
rect 186927 218106 190560 218108
rect 186927 218050 186932 218106
rect 186988 218050 190560 218106
rect 186927 218048 190560 218050
rect 186927 218045 186993 218048
rect 147279 217812 147345 217815
rect 143904 217810 147345 217812
rect 143904 217754 147284 217810
rect 147340 217754 147345 217810
rect 143904 217752 147345 217754
rect 147279 217749 147345 217752
rect 190146 217294 190206 218048
rect 675898 217750 675904 217814
rect 675968 217812 675974 217814
rect 675968 217752 676320 217812
rect 675968 217750 675974 217752
rect 190146 217234 190560 217294
rect 677058 217075 677118 217190
rect 677007 217070 677118 217075
rect 677007 217014 677012 217070
rect 677068 217014 677118 217070
rect 677007 217012 677118 217014
rect 677007 217009 677073 217012
rect 675759 216776 675825 216779
rect 675759 216774 676320 216776
rect 149391 216628 149457 216631
rect 143904 216626 149457 216628
rect 143904 216570 149396 216626
rect 149452 216570 149457 216626
rect 143904 216568 149457 216570
rect 149391 216565 149457 216568
rect 186735 216480 186801 216483
rect 186735 216478 190560 216480
rect 186735 216422 186740 216478
rect 186796 216422 190560 216478
rect 186735 216420 190560 216422
rect 186735 216417 186801 216420
rect 190146 215814 190206 216420
rect 190146 215754 190560 215814
rect 143874 214852 143934 215340
rect 186255 215000 186321 215003
rect 186255 214998 190560 215000
rect 186255 214942 186260 214998
rect 186316 214942 190560 214998
rect 186255 214940 190560 214942
rect 186255 214937 186321 214940
rect 147375 214852 147441 214855
rect 143874 214850 147441 214852
rect 143874 214794 147380 214850
rect 147436 214794 147441 214850
rect 143874 214792 147441 214794
rect 147375 214789 147441 214792
rect 190146 214334 190206 214940
rect 640386 214822 640446 216746
rect 675759 216718 675764 216774
rect 675820 216718 676320 216774
rect 675759 216716 676320 216718
rect 675759 216713 675825 216716
rect 675706 216270 675712 216334
rect 675776 216332 675782 216334
rect 675776 216272 676320 216332
rect 675776 216270 675782 216272
rect 675514 215678 675520 215742
rect 675584 215740 675590 215742
rect 675584 215680 676320 215740
rect 675584 215678 675590 215680
rect 676866 215003 676926 215192
rect 676866 214998 676977 215003
rect 676866 214942 676916 214998
rect 676972 214942 676977 214998
rect 676866 214940 676977 214942
rect 676911 214937 676977 214940
rect 675279 214852 675345 214855
rect 675279 214850 676320 214852
rect 675279 214794 675284 214850
rect 675340 214794 676320 214850
rect 675279 214792 676320 214794
rect 675279 214789 675345 214792
rect 190146 214274 190560 214334
rect 676290 214115 676350 214230
rect 147567 214112 147633 214115
rect 143904 214110 147633 214112
rect 143904 214054 147572 214110
rect 147628 214054 147633 214110
rect 143904 214052 147633 214054
rect 147567 214049 147633 214052
rect 676239 214110 676350 214115
rect 676239 214054 676244 214110
rect 676300 214054 676350 214110
rect 676239 214052 676350 214054
rect 676239 214049 676305 214052
rect 676047 213742 676113 213745
rect 676047 213740 676320 213742
rect 676047 213684 676052 213740
rect 676108 213684 676320 213740
rect 676047 213682 676320 213684
rect 676047 213679 676113 213682
rect 41775 213668 41841 213671
rect 41568 213666 41841 213668
rect 41568 213610 41780 213666
rect 41836 213610 41841 213666
rect 41568 213608 41841 213610
rect 41775 213605 41841 213608
rect 186063 213520 186129 213523
rect 186063 213518 190560 213520
rect 186063 213462 186068 213518
rect 186124 213462 190560 213518
rect 186063 213460 190560 213462
rect 186063 213457 186129 213460
rect 41775 213150 41841 213153
rect 41568 213148 41841 213150
rect 41568 213092 41780 213148
rect 41836 213092 41841 213148
rect 41568 213090 41841 213092
rect 41775 213087 41841 213090
rect 146895 212928 146961 212931
rect 143904 212926 146961 212928
rect 143904 212870 146900 212926
rect 146956 212870 146961 212926
rect 143904 212868 146961 212870
rect 146895 212865 146961 212868
rect 41583 212780 41649 212783
rect 41538 212778 41649 212780
rect 41538 212722 41588 212778
rect 41644 212722 41649 212778
rect 41538 212717 41649 212722
rect 41538 212602 41598 212717
rect 190146 212706 190206 213460
rect 676866 213079 676926 213342
rect 676815 213074 676926 213079
rect 676815 213018 676820 213074
rect 676876 213018 676926 213074
rect 676815 213016 676926 213018
rect 676815 213013 676881 213016
rect 190146 212646 190560 212706
rect 640194 212339 640254 212898
rect 676047 212780 676113 212783
rect 676047 212778 676320 212780
rect 676047 212722 676052 212778
rect 676108 212722 676320 212778
rect 676047 212720 676320 212722
rect 676047 212717 676113 212720
rect 640143 212334 640254 212339
rect 640143 212278 640148 212334
rect 640204 212278 640254 212334
rect 640143 212276 640254 212278
rect 640143 212273 640209 212276
rect 41775 212188 41841 212191
rect 41568 212186 41841 212188
rect 41568 212130 41780 212186
rect 41836 212130 41841 212186
rect 41568 212128 41841 212130
rect 41775 212125 41841 212128
rect 676290 212043 676350 212158
rect 187023 212040 187089 212043
rect 187023 212038 190560 212040
rect 187023 211982 187028 212038
rect 187084 211982 190560 212038
rect 187023 211980 190560 211982
rect 676239 212038 676350 212043
rect 676239 211982 676244 212038
rect 676300 211982 676350 212038
rect 676239 211980 676350 211982
rect 187023 211977 187089 211980
rect 147375 211744 147441 211747
rect 143904 211742 147441 211744
rect 143904 211686 147380 211742
rect 147436 211686 147441 211742
rect 143904 211684 147441 211686
rect 147375 211681 147441 211684
rect 41775 211670 41841 211673
rect 41568 211668 41841 211670
rect 41568 211612 41780 211668
rect 41836 211612 41841 211668
rect 41568 211610 41841 211612
rect 41775 211607 41841 211610
rect 41583 211300 41649 211303
rect 41538 211298 41649 211300
rect 41538 211242 41588 211298
rect 41644 211242 41649 211298
rect 41538 211237 41649 211242
rect 41538 211122 41598 211237
rect 190146 211152 190206 211980
rect 676239 211977 676305 211980
rect 676047 211818 676113 211821
rect 676047 211816 676320 211818
rect 676047 211760 676052 211816
rect 676108 211760 676320 211816
rect 676047 211758 676320 211760
rect 676047 211755 676113 211758
rect 640143 211596 640209 211599
rect 640143 211594 640254 211596
rect 640143 211538 640148 211594
rect 640204 211538 640254 211594
rect 640143 211533 640254 211538
rect 190146 211092 190560 211152
rect 640194 210974 640254 211533
rect 675951 211300 676017 211303
rect 675951 211298 676320 211300
rect 675951 211242 675956 211298
rect 676012 211242 676320 211298
rect 675951 211240 676320 211242
rect 675951 211237 676017 211240
rect 41775 210708 41841 210711
rect 41568 210706 41841 210708
rect 41568 210650 41780 210706
rect 41836 210650 41841 210706
rect 41568 210648 41841 210650
rect 41775 210645 41841 210648
rect 679938 210563 679998 210678
rect 186447 210560 186513 210563
rect 186447 210558 190206 210560
rect 186447 210502 186452 210558
rect 186508 210502 190206 210558
rect 186447 210500 190206 210502
rect 679938 210558 680049 210563
rect 679938 210502 679988 210558
rect 680044 210502 680049 210558
rect 679938 210500 680049 210502
rect 186447 210497 186513 210500
rect 190146 210486 190206 210500
rect 679983 210497 680049 210500
rect 190146 210426 190560 210486
rect 147375 210412 147441 210415
rect 143904 210410 147441 210412
rect 143904 210354 147380 210410
rect 147436 210354 147441 210410
rect 143904 210352 147441 210354
rect 147375 210349 147441 210352
rect 41775 210116 41841 210119
rect 41568 210114 41841 210116
rect 41568 210058 41780 210114
rect 41836 210058 41841 210114
rect 41568 210056 41841 210058
rect 41775 210053 41841 210056
rect 41583 209820 41649 209823
rect 41538 209818 41649 209820
rect 41538 209762 41588 209818
rect 41644 209762 41649 209818
rect 41538 209757 41649 209762
rect 41538 209642 41598 209757
rect 190146 209672 190206 210426
rect 679746 209971 679806 210308
rect 679746 209966 679857 209971
rect 679983 209968 680049 209971
rect 679746 209910 679796 209966
rect 679852 209910 679857 209966
rect 679746 209908 679857 209910
rect 679791 209905 679857 209908
rect 679938 209966 680049 209968
rect 679938 209910 679988 209966
rect 680044 209910 680049 209966
rect 679938 209905 680049 209910
rect 679938 209790 679998 209905
rect 190146 209612 190560 209672
rect 679791 209524 679857 209527
rect 679746 209522 679857 209524
rect 679746 209466 679796 209522
rect 679852 209466 679857 209522
rect 679746 209461 679857 209466
rect 146895 209228 146961 209231
rect 143904 209226 146961 209228
rect 25602 208935 25662 209198
rect 143904 209170 146900 209226
rect 146956 209170 146961 209226
rect 679746 209198 679806 209461
rect 143904 209168 146961 209170
rect 146895 209165 146961 209168
rect 186639 209080 186705 209083
rect 186639 209078 190206 209080
rect 186639 209022 186644 209078
rect 186700 209022 190206 209078
rect 186639 209020 190206 209022
rect 186639 209017 186705 209020
rect 190146 209006 190206 209020
rect 190146 208946 190560 209006
rect 25602 208930 25713 208935
rect 25602 208874 25652 208930
rect 25708 208874 25713 208930
rect 25602 208872 25713 208874
rect 25647 208869 25713 208872
rect 25794 208343 25854 208606
rect 25794 208338 25905 208343
rect 25794 208282 25844 208338
rect 25900 208282 25905 208338
rect 25794 208280 25905 208282
rect 25839 208277 25905 208280
rect 190146 208192 190206 208946
rect 190146 208132 190560 208192
rect 25602 207899 25662 208088
rect 146991 208044 147057 208047
rect 143904 208042 147057 208044
rect 143904 207986 146996 208042
rect 147052 207986 147057 208042
rect 143904 207984 147057 207986
rect 146991 207981 147057 207984
rect 25551 207894 25662 207899
rect 25551 207838 25556 207894
rect 25612 207838 25662 207894
rect 25551 207836 25662 207838
rect 25551 207833 25617 207836
rect 34242 207455 34302 207718
rect 34242 207450 34353 207455
rect 34242 207394 34292 207450
rect 34348 207394 34353 207450
rect 34242 207392 34353 207394
rect 34287 207389 34353 207392
rect 190146 207318 190560 207378
rect 186351 207304 186417 207307
rect 190146 207304 190206 207318
rect 186351 207302 190206 207304
rect 186351 207246 186356 207302
rect 186412 207246 190206 207302
rect 639810 207274 639870 209124
rect 676282 207686 676288 207750
rect 676352 207748 676358 207750
rect 677007 207748 677073 207751
rect 676352 207746 677073 207748
rect 676352 207690 677012 207746
rect 677068 207690 677073 207746
rect 676352 207688 677073 207690
rect 676352 207686 676358 207688
rect 677007 207685 677073 207688
rect 676666 207538 676672 207602
rect 676736 207600 676742 207602
rect 676911 207600 676977 207603
rect 676736 207598 676977 207600
rect 676736 207542 676916 207598
rect 676972 207542 676977 207598
rect 676736 207540 676977 207542
rect 676736 207538 676742 207540
rect 676911 207537 676977 207540
rect 676474 207390 676480 207454
rect 676544 207452 676550 207454
rect 676815 207452 676881 207455
rect 676544 207450 676881 207452
rect 676544 207394 676820 207450
rect 676876 207394 676881 207450
rect 676544 207392 676881 207394
rect 676544 207390 676550 207392
rect 676815 207389 676881 207392
rect 186351 207244 190206 207246
rect 186351 207241 186417 207244
rect 25794 206863 25854 207126
rect 25743 206858 25854 206863
rect 25743 206802 25748 206858
rect 25804 206802 25854 206858
rect 25743 206800 25854 206802
rect 25743 206797 25809 206800
rect 41871 206638 41937 206641
rect 41568 206636 41937 206638
rect 41568 206580 41876 206636
rect 41932 206580 41937 206636
rect 41568 206578 41937 206580
rect 41871 206575 41937 206578
rect 143874 206416 143934 206904
rect 190146 206712 190206 207244
rect 190146 206652 190560 206712
rect 147087 206416 147153 206419
rect 143874 206414 147153 206416
rect 143874 206358 147092 206414
rect 147148 206358 147153 206414
rect 143874 206356 147153 206358
rect 147087 206353 147153 206356
rect 41154 205974 41214 206238
rect 41146 205910 41152 205974
rect 41216 205910 41222 205974
rect 190146 205838 190560 205898
rect 149391 205676 149457 205679
rect 143904 205674 149457 205676
rect 41346 205382 41406 205646
rect 143904 205618 149396 205674
rect 149452 205618 149457 205674
rect 143904 205616 149457 205618
rect 149391 205613 149457 205616
rect 41338 205318 41344 205382
rect 41408 205318 41414 205382
rect 186543 205232 186609 205235
rect 190146 205232 190206 205838
rect 186543 205230 190560 205232
rect 186543 205174 186548 205230
rect 186604 205174 190560 205230
rect 186543 205172 190560 205174
rect 186543 205169 186609 205172
rect 40770 204938 40830 205054
rect 40762 204874 40768 204938
rect 40832 204874 40838 204938
rect 41538 204347 41598 204684
rect 147663 204492 147729 204495
rect 143904 204490 147729 204492
rect 143904 204434 147668 204490
rect 147724 204434 147729 204490
rect 143904 204432 147729 204434
rect 147663 204429 147729 204432
rect 41538 204342 41649 204347
rect 41538 204286 41588 204342
rect 41644 204286 41649 204342
rect 41538 204284 41649 204286
rect 41583 204281 41649 204284
rect 186159 204344 186225 204347
rect 186159 204342 190560 204344
rect 186159 204286 186164 204342
rect 186220 204286 190560 204342
rect 186159 204284 190560 204286
rect 186159 204281 186225 204284
rect 41775 204196 41841 204199
rect 41568 204194 41841 204196
rect 41568 204138 41780 204194
rect 41836 204138 41841 204194
rect 41568 204136 41841 204138
rect 41775 204133 41841 204136
rect 41914 203604 41920 203606
rect 41568 203544 41920 203604
rect 41914 203542 41920 203544
rect 41984 203542 41990 203606
rect 190146 203604 190206 204284
rect 190146 203544 190560 203604
rect 639810 203426 639870 205350
rect 675759 204492 675825 204495
rect 675898 204492 675904 204494
rect 675759 204490 675904 204492
rect 675759 204434 675764 204490
rect 675820 204434 675904 204490
rect 675759 204432 675904 204434
rect 675759 204429 675825 204432
rect 675898 204430 675904 204432
rect 675968 204430 675974 204494
rect 149487 203308 149553 203311
rect 143904 203306 149553 203308
rect 143904 203250 149492 203306
rect 149548 203250 149553 203306
rect 143904 203248 149553 203250
rect 149487 203245 149553 203248
rect 41775 203234 41841 203237
rect 41568 203232 41841 203234
rect 41568 203176 41780 203232
rect 41836 203176 41841 203232
rect 41568 203174 41841 203176
rect 41775 203171 41841 203174
rect 185967 202864 186033 202867
rect 185967 202862 190560 202864
rect 185967 202806 185972 202862
rect 186028 202806 190560 202862
rect 185967 202804 190560 202806
rect 185967 202801 186033 202804
rect 41775 202716 41841 202719
rect 41568 202714 41841 202716
rect 41568 202658 41780 202714
rect 41836 202658 41841 202714
rect 41568 202656 41841 202658
rect 41775 202653 41841 202656
rect 41967 202124 42033 202127
rect 41568 202122 42033 202124
rect 41568 202066 41972 202122
rect 42028 202066 42033 202122
rect 41568 202064 42033 202066
rect 190146 202124 190206 202804
rect 675663 202718 675729 202719
rect 675663 202714 675712 202718
rect 675776 202716 675782 202718
rect 675663 202658 675668 202714
rect 675663 202654 675712 202658
rect 675776 202656 675820 202716
rect 675776 202654 675782 202656
rect 675663 202653 675729 202654
rect 190146 202064 190560 202124
rect 41967 202061 42033 202064
rect 41967 201680 42033 201683
rect 41568 201678 42033 201680
rect 41568 201622 41972 201678
rect 42028 201622 42033 201678
rect 41568 201620 42033 201622
rect 143874 201680 143934 202020
rect 149391 201680 149457 201683
rect 143874 201678 149457 201680
rect 143874 201622 149396 201678
rect 149452 201622 149457 201678
rect 143874 201620 149457 201622
rect 41967 201617 42033 201620
rect 149391 201617 149457 201620
rect 34287 201532 34353 201535
rect 40954 201532 40960 201534
rect 34287 201530 40960 201532
rect 34287 201474 34292 201530
rect 34348 201474 40960 201530
rect 34287 201472 40960 201474
rect 34287 201469 34353 201472
rect 40954 201470 40960 201472
rect 41024 201470 41030 201534
rect 190287 201384 190353 201387
rect 190287 201382 190560 201384
rect 190287 201326 190292 201382
rect 190348 201326 190560 201382
rect 190287 201324 190560 201326
rect 190287 201321 190353 201324
rect 41775 201236 41841 201239
rect 41568 201234 41841 201236
rect 41568 201178 41780 201234
rect 41836 201178 41841 201234
rect 41568 201176 41841 201178
rect 41775 201173 41841 201176
rect 640194 200943 640254 201502
rect 25647 200940 25713 200943
rect 25602 200938 25713 200940
rect 25602 200882 25652 200938
rect 25708 200882 25713 200938
rect 25602 200877 25713 200882
rect 25839 200940 25905 200943
rect 41722 200940 41728 200942
rect 25839 200938 41728 200940
rect 25839 200882 25844 200938
rect 25900 200882 41728 200938
rect 25839 200880 41728 200882
rect 25839 200877 25905 200880
rect 41722 200878 41728 200880
rect 41792 200878 41798 200942
rect 640143 200938 640254 200943
rect 640143 200882 640148 200938
rect 640204 200882 640254 200938
rect 640143 200880 640254 200882
rect 640143 200877 640209 200880
rect 25602 200792 25662 200877
rect 42298 200792 42304 200794
rect 25602 200732 42304 200792
rect 42298 200730 42304 200732
rect 42368 200730 42374 200794
rect 149391 200792 149457 200795
rect 143904 200790 149457 200792
rect 143904 200734 149396 200790
rect 149452 200734 149457 200790
rect 143904 200732 149457 200734
rect 149391 200729 149457 200732
rect 190287 200570 190353 200573
rect 190287 200568 190560 200570
rect 190287 200512 190292 200568
rect 190348 200512 190560 200568
rect 190287 200510 190560 200512
rect 190287 200507 190353 200510
rect 640143 200200 640209 200203
rect 640143 200198 640254 200200
rect 640143 200142 640148 200198
rect 640204 200142 640254 200198
rect 640143 200137 640254 200142
rect 25551 200052 25617 200055
rect 42106 200052 42112 200054
rect 25551 200050 42112 200052
rect 25551 199994 25556 200050
rect 25612 199994 42112 200050
rect 25551 199992 42112 199994
rect 25551 199989 25617 199992
rect 42106 199990 42112 199992
rect 42176 199990 42182 200054
rect 25743 199756 25809 199759
rect 41530 199756 41536 199758
rect 25743 199754 41536 199756
rect 25743 199698 25748 199754
rect 25804 199698 41536 199754
rect 25743 199696 41536 199698
rect 25743 199693 25809 199696
rect 41530 199694 41536 199696
rect 41600 199694 41606 199758
rect 184335 199756 184401 199759
rect 184335 199754 190560 199756
rect 184335 199698 184340 199754
rect 184396 199698 190560 199754
rect 184335 199696 190560 199698
rect 184335 199693 184401 199696
rect 147471 199608 147537 199611
rect 143904 199606 147537 199608
rect 143904 199550 147476 199606
rect 147532 199550 147537 199606
rect 640194 199578 640254 200137
rect 143904 199548 147537 199550
rect 147471 199545 147537 199548
rect 187215 199164 187281 199167
rect 187215 199162 190014 199164
rect 187215 199106 187220 199162
rect 187276 199106 190014 199162
rect 187215 199104 190014 199106
rect 187215 199101 187281 199104
rect 189954 199090 190014 199104
rect 189954 199030 190560 199090
rect 149295 198424 149361 198427
rect 675567 198426 675633 198427
rect 143904 198422 149361 198424
rect 143904 198366 149300 198422
rect 149356 198366 149361 198422
rect 143904 198364 149361 198366
rect 149295 198361 149361 198364
rect 675514 198362 675520 198426
rect 675584 198424 675633 198426
rect 675584 198422 675676 198424
rect 675628 198366 675676 198422
rect 675584 198364 675676 198366
rect 675584 198362 675633 198364
rect 675567 198361 675633 198362
rect 185487 198276 185553 198279
rect 185487 198274 190560 198276
rect 185487 198218 185492 198274
rect 185548 198218 190560 198274
rect 185487 198216 190560 198218
rect 185487 198213 185553 198216
rect 184239 197684 184305 197687
rect 184239 197682 190014 197684
rect 184239 197626 184244 197682
rect 184300 197626 190014 197682
rect 184239 197624 190014 197626
rect 184239 197621 184305 197624
rect 189954 197610 190014 197624
rect 189954 197550 190560 197610
rect 149391 197092 149457 197095
rect 143904 197090 149457 197092
rect 143904 197034 149396 197090
rect 149452 197034 149457 197090
rect 143904 197032 149457 197034
rect 149391 197029 149457 197032
rect 184431 196796 184497 196799
rect 184431 196794 190560 196796
rect 184431 196738 184436 196794
rect 184492 196738 190560 196794
rect 184431 196736 190560 196738
rect 184431 196733 184497 196736
rect 184335 196056 184401 196059
rect 184335 196054 190560 196056
rect 184335 195998 184340 196054
rect 184396 195998 190560 196054
rect 184335 195996 190560 195998
rect 184335 195993 184401 195996
rect 147279 195908 147345 195911
rect 143904 195906 147345 195908
rect 143904 195850 147284 195906
rect 147340 195850 147345 195906
rect 143904 195848 147345 195850
rect 147279 195845 147345 195848
rect 639810 195730 639870 197654
rect 41775 195318 41841 195319
rect 41722 195316 41728 195318
rect 41684 195256 41728 195316
rect 41792 195314 41841 195318
rect 41836 195258 41841 195314
rect 41722 195254 41728 195256
rect 41792 195254 41841 195258
rect 41775 195253 41841 195254
rect 184335 195316 184401 195319
rect 675759 195316 675825 195319
rect 676474 195316 676480 195318
rect 184335 195314 190560 195316
rect 184335 195258 184340 195314
rect 184396 195258 190560 195314
rect 184335 195256 190560 195258
rect 675759 195314 676480 195316
rect 675759 195258 675764 195314
rect 675820 195258 676480 195314
rect 675759 195256 676480 195258
rect 184335 195253 184401 195256
rect 675759 195253 675825 195256
rect 676474 195254 676480 195256
rect 676544 195254 676550 195318
rect 149487 194724 149553 194727
rect 143904 194722 149553 194724
rect 143904 194666 149492 194722
rect 149548 194666 149553 194722
rect 143904 194664 149553 194666
rect 149487 194661 149553 194664
rect 184431 194428 184497 194431
rect 184431 194426 190560 194428
rect 184431 194370 184436 194426
rect 184492 194370 190560 194426
rect 184431 194368 190560 194370
rect 184431 194365 184497 194368
rect 184527 193836 184593 193839
rect 184527 193834 190014 193836
rect 184527 193778 184532 193834
rect 184588 193778 190014 193834
rect 184527 193776 190014 193778
rect 184527 193773 184593 193776
rect 189954 193762 190014 193776
rect 189954 193702 190560 193762
rect 143874 193392 143934 193436
rect 149391 193392 149457 193395
rect 143874 193390 149457 193392
rect 143874 193334 149396 193390
rect 149452 193334 149457 193390
rect 143874 193332 149457 193334
rect 149391 193329 149457 193332
rect 184431 192948 184497 192951
rect 184431 192946 190560 192948
rect 184431 192890 184436 192946
rect 184492 192890 190560 192946
rect 184431 192888 190560 192890
rect 184431 192885 184497 192888
rect 184335 192356 184401 192359
rect 184335 192354 190014 192356
rect 184335 192298 184340 192354
rect 184396 192298 190014 192354
rect 184335 192296 190014 192298
rect 184335 192293 184401 192296
rect 189954 192282 190014 192296
rect 189954 192222 190560 192282
rect 149391 192208 149457 192211
rect 143904 192206 149457 192208
rect 143904 192150 149396 192206
rect 149452 192150 149457 192206
rect 143904 192148 149457 192150
rect 149391 192145 149457 192148
rect 639810 192030 639870 193880
rect 675759 193540 675825 193543
rect 676282 193540 676288 193542
rect 675759 193538 676288 193540
rect 675759 193482 675764 193538
rect 675820 193482 676288 193538
rect 675759 193480 676288 193482
rect 675759 193477 675825 193480
rect 676282 193478 676288 193480
rect 676352 193478 676358 193542
rect 675759 191616 675825 191619
rect 676666 191616 676672 191618
rect 675759 191614 676672 191616
rect 675759 191558 675764 191614
rect 675820 191558 676672 191614
rect 675759 191556 676672 191558
rect 675759 191553 675825 191556
rect 676666 191554 676672 191556
rect 676736 191554 676742 191618
rect 184527 191468 184593 191471
rect 184527 191466 190560 191468
rect 184527 191410 184532 191466
rect 184588 191410 190560 191466
rect 184527 191408 190560 191410
rect 184527 191405 184593 191408
rect 147279 191024 147345 191027
rect 143904 191022 147345 191024
rect 143904 190966 147284 191022
rect 147340 190966 147345 191022
rect 143904 190964 147345 190966
rect 147279 190961 147345 190964
rect 184623 190728 184689 190731
rect 184623 190726 190014 190728
rect 184623 190670 184628 190726
rect 184684 190670 190014 190726
rect 184623 190668 190014 190670
rect 184623 190665 184689 190668
rect 189954 190654 190014 190668
rect 189954 190594 190560 190654
rect 41530 190074 41536 190138
rect 41600 190136 41606 190138
rect 41775 190136 41841 190139
rect 41600 190134 41841 190136
rect 41600 190078 41780 190134
rect 41836 190078 41841 190134
rect 41600 190076 41841 190078
rect 41600 190074 41606 190076
rect 41775 190073 41841 190076
rect 184335 189988 184401 189991
rect 184335 189986 190560 189988
rect 184335 189930 184340 189986
rect 184396 189930 190560 189986
rect 184335 189928 190560 189930
rect 184335 189925 184401 189928
rect 149391 189840 149457 189843
rect 143904 189838 149457 189840
rect 143904 189782 149396 189838
rect 149452 189782 149457 189838
rect 143904 189780 149457 189782
rect 149391 189777 149457 189780
rect 41338 189630 41344 189694
rect 41408 189630 41414 189694
rect 41346 189250 41406 189630
rect 41338 189186 41344 189250
rect 41408 189186 41414 189250
rect 184527 189248 184593 189251
rect 184527 189246 190014 189248
rect 184527 189190 184532 189246
rect 184588 189190 190014 189246
rect 184527 189188 190014 189190
rect 184527 189185 184593 189188
rect 189954 189174 190014 189188
rect 189954 189114 190560 189174
rect 143874 188064 143934 188552
rect 184431 188508 184497 188511
rect 184431 188506 190560 188508
rect 184431 188450 184436 188506
rect 184492 188450 190560 188506
rect 184431 188448 190560 188450
rect 184431 188445 184497 188448
rect 639810 188182 639870 190106
rect 149583 188064 149649 188067
rect 143874 188062 149649 188064
rect 143874 188006 149588 188062
rect 149644 188006 149649 188062
rect 143874 188004 149649 188006
rect 149583 188001 149649 188004
rect 41871 187918 41937 187919
rect 41871 187914 41920 187918
rect 41984 187916 41990 187918
rect 41871 187858 41876 187914
rect 41871 187854 41920 187858
rect 41984 187856 42028 187916
rect 41984 187854 41990 187856
rect 41871 187853 41937 187854
rect 184335 187620 184401 187623
rect 184335 187618 190560 187620
rect 184335 187562 184340 187618
rect 184396 187562 190560 187618
rect 184335 187560 190560 187562
rect 184335 187557 184401 187560
rect 149295 187472 149361 187475
rect 143904 187470 149361 187472
rect 143904 187414 149300 187470
rect 149356 187414 149361 187470
rect 143904 187412 149361 187414
rect 149295 187409 149361 187412
rect 40762 187114 40768 187178
rect 40832 187176 40838 187178
rect 41775 187176 41841 187179
rect 40832 187174 41841 187176
rect 40832 187118 41780 187174
rect 41836 187118 41841 187174
rect 40832 187116 41841 187118
rect 40832 187114 40838 187116
rect 41775 187113 41841 187116
rect 184335 186880 184401 186883
rect 184335 186878 190560 186880
rect 184335 186822 184340 186878
rect 184396 186822 190560 186878
rect 184335 186820 190560 186822
rect 184335 186817 184401 186820
rect 41338 186670 41344 186734
rect 41408 186732 41414 186734
rect 41775 186732 41841 186735
rect 41408 186730 41841 186732
rect 41408 186674 41780 186730
rect 41836 186674 41841 186730
rect 41408 186672 41841 186674
rect 41408 186670 41414 186672
rect 41775 186669 41841 186672
rect 149199 186288 149265 186291
rect 143904 186286 149265 186288
rect 143904 186230 149204 186286
rect 149260 186230 149265 186286
rect 143904 186228 149265 186230
rect 149199 186225 149265 186228
rect 184431 186140 184497 186143
rect 184431 186138 190560 186140
rect 184431 186082 184436 186138
rect 184492 186082 190560 186138
rect 184431 186080 190560 186082
rect 184431 186077 184497 186080
rect 40954 185782 40960 185846
rect 41024 185844 41030 185846
rect 41775 185844 41841 185847
rect 41024 185842 41841 185844
rect 41024 185786 41780 185842
rect 41836 185786 41841 185842
rect 41024 185784 41841 185786
rect 41024 185782 41030 185784
rect 41775 185781 41841 185784
rect 640194 185699 640254 186258
rect 640194 185694 640305 185699
rect 640194 185638 640244 185694
rect 640300 185638 640305 185694
rect 640194 185636 640305 185638
rect 640239 185633 640305 185636
rect 184623 185400 184689 185403
rect 184623 185398 190014 185400
rect 184623 185342 184628 185398
rect 184684 185342 190014 185398
rect 184623 185340 190014 185342
rect 184623 185337 184689 185340
rect 189954 185326 190014 185340
rect 189954 185266 190560 185326
rect 143874 184512 143934 185000
rect 640239 184956 640305 184959
rect 640194 184954 640305 184956
rect 640194 184898 640244 184954
rect 640300 184898 640305 184954
rect 640194 184893 640305 184898
rect 184527 184660 184593 184663
rect 184527 184658 190560 184660
rect 184527 184602 184532 184658
rect 184588 184602 190560 184658
rect 184527 184600 190560 184602
rect 184527 184597 184593 184600
rect 149391 184512 149457 184515
rect 143874 184510 149457 184512
rect 143874 184454 149396 184510
rect 149452 184454 149457 184510
rect 143874 184452 149457 184454
rect 149391 184449 149457 184452
rect 640194 184334 640254 184893
rect 42159 184216 42225 184219
rect 42298 184216 42304 184218
rect 42159 184214 42304 184216
rect 42159 184158 42164 184214
rect 42220 184158 42304 184214
rect 42159 184156 42304 184158
rect 42159 184153 42225 184156
rect 42298 184154 42304 184156
rect 42368 184154 42374 184218
rect 184335 183920 184401 183923
rect 184335 183918 190014 183920
rect 184335 183862 184340 183918
rect 184396 183862 190014 183918
rect 184335 183860 190014 183862
rect 184335 183857 184401 183860
rect 189954 183846 190014 183860
rect 189954 183786 190560 183846
rect 149487 183772 149553 183775
rect 143904 183770 149553 183772
rect 143904 183714 149492 183770
rect 149548 183714 149553 183770
rect 143904 183712 149553 183714
rect 149487 183709 149553 183712
rect 41871 183626 41937 183627
rect 41871 183622 41920 183626
rect 41984 183624 41990 183626
rect 41871 183566 41876 183622
rect 41871 183562 41920 183566
rect 41984 183564 42028 183624
rect 41984 183562 41990 183564
rect 41871 183561 41937 183562
rect 184431 183180 184497 183183
rect 184431 183178 190560 183180
rect 184431 183122 184436 183178
rect 184492 183122 190560 183178
rect 184431 183120 190560 183122
rect 184431 183117 184497 183120
rect 645135 183032 645201 183035
rect 640386 183030 645201 183032
rect 640386 182974 645140 183030
rect 645196 182974 645201 183030
rect 640386 182972 645201 182974
rect 42063 182886 42129 182887
rect 42063 182882 42112 182886
rect 42176 182884 42182 182886
rect 42063 182826 42068 182882
rect 42063 182822 42112 182826
rect 42176 182824 42220 182884
rect 42176 182822 42182 182824
rect 42063 182821 42129 182822
rect 149391 182588 149457 182591
rect 143904 182586 149457 182588
rect 143904 182530 149396 182586
rect 149452 182530 149457 182586
rect 143904 182528 149457 182530
rect 149391 182525 149457 182528
rect 185775 182440 185841 182443
rect 640386 182440 640446 182972
rect 645135 182969 645201 182972
rect 185775 182438 190014 182440
rect 185775 182382 185780 182438
rect 185836 182382 190014 182438
rect 640224 182410 640446 182440
rect 185775 182380 190014 182382
rect 185775 182377 185841 182380
rect 189954 182366 190014 182380
rect 640194 182380 640416 182410
rect 189954 182306 190560 182366
rect 184527 181552 184593 181555
rect 184527 181550 190560 181552
rect 184527 181494 184532 181550
rect 184588 181494 190560 181550
rect 184527 181492 190560 181494
rect 184527 181489 184593 181492
rect 149487 181404 149553 181407
rect 143904 181402 149553 181404
rect 143904 181346 149492 181402
rect 149548 181346 149553 181402
rect 143904 181344 149553 181346
rect 149487 181341 149553 181344
rect 184335 180812 184401 180815
rect 184335 180810 190560 180812
rect 184335 180754 184340 180810
rect 184396 180754 190560 180810
rect 184335 180752 190560 180754
rect 184335 180749 184401 180752
rect 640194 180560 640254 182380
rect 143874 179628 143934 180116
rect 184431 180072 184497 180075
rect 184431 180070 190560 180072
rect 184431 180014 184436 180070
rect 184492 180014 190560 180070
rect 184431 180012 190560 180014
rect 184431 180009 184497 180012
rect 149295 179628 149361 179631
rect 143874 179626 149361 179628
rect 143874 179570 149300 179626
rect 149356 179570 149361 179626
rect 143874 179568 149361 179570
rect 149295 179565 149361 179568
rect 184623 179332 184689 179335
rect 645135 179332 645201 179335
rect 184623 179330 190560 179332
rect 184623 179274 184628 179330
rect 184684 179274 190560 179330
rect 184623 179272 190560 179274
rect 640194 179330 645201 179332
rect 640194 179274 645140 179330
rect 645196 179274 645201 179330
rect 640194 179272 645201 179274
rect 184623 179269 184689 179272
rect 149391 178888 149457 178891
rect 143904 178886 149457 178888
rect 143904 178830 149396 178886
rect 149452 178830 149457 178886
rect 143904 178828 149457 178830
rect 149391 178825 149457 178828
rect 184527 178592 184593 178595
rect 184527 178590 190560 178592
rect 184527 178534 184532 178590
rect 184588 178534 190560 178590
rect 184527 178532 190560 178534
rect 184527 178529 184593 178532
rect 149487 177704 149553 177707
rect 143904 177702 149553 177704
rect 143904 177646 149492 177702
rect 149548 177646 149553 177702
rect 143904 177644 149553 177646
rect 149487 177641 149553 177644
rect 186735 177704 186801 177707
rect 186735 177702 190560 177704
rect 186735 177646 186740 177702
rect 186796 177646 190560 177702
rect 186735 177644 190560 177646
rect 186735 177641 186801 177644
rect 184335 177112 184401 177115
rect 184335 177110 190014 177112
rect 184335 177054 184340 177110
rect 184396 177054 190014 177110
rect 184335 177052 190014 177054
rect 184335 177049 184401 177052
rect 189954 177038 190014 177052
rect 189954 176978 190560 177038
rect 640194 176786 640254 179272
rect 645135 179269 645201 179272
rect 676143 177408 676209 177411
rect 676290 177408 676350 177674
rect 676143 177406 676350 177408
rect 676143 177350 676148 177406
rect 676204 177350 676350 177406
rect 676143 177348 676350 177350
rect 676143 177345 676209 177348
rect 676290 176819 676350 177082
rect 676290 176814 676401 176819
rect 676290 176758 676340 176814
rect 676396 176758 676401 176814
rect 676290 176756 676401 176758
rect 676335 176753 676401 176756
rect 149391 176520 149457 176523
rect 143904 176518 149457 176520
rect 143904 176462 149396 176518
rect 149452 176462 149457 176518
rect 143904 176460 149457 176462
rect 149391 176457 149457 176460
rect 676290 176375 676350 176638
rect 676239 176370 676350 176375
rect 676239 176314 676244 176370
rect 676300 176314 676350 176370
rect 676239 176312 676350 176314
rect 676239 176309 676305 176312
rect 184431 176224 184497 176227
rect 184431 176222 190560 176224
rect 184431 176166 184436 176222
rect 184492 176166 190560 176222
rect 184431 176164 190560 176166
rect 184431 176161 184497 176164
rect 674362 176162 674368 176226
rect 674432 176224 674438 176226
rect 674432 176164 676320 176224
rect 674432 176162 674438 176164
rect 184335 175632 184401 175635
rect 184335 175630 190014 175632
rect 184335 175574 184340 175630
rect 184396 175574 190014 175630
rect 184335 175572 190014 175574
rect 184335 175569 184401 175572
rect 189954 175558 190014 175572
rect 674362 175570 674368 175634
rect 674432 175632 674438 175634
rect 674432 175572 676320 175632
rect 674432 175570 674438 175572
rect 189954 175498 190560 175558
rect 673978 175422 673984 175486
rect 674048 175484 674054 175486
rect 674048 175424 676350 175484
rect 674048 175422 674054 175424
rect 147663 175188 147729 175191
rect 143904 175186 147729 175188
rect 143904 175130 147668 175186
rect 147724 175130 147729 175186
rect 143904 175128 147729 175130
rect 147663 175125 147729 175128
rect 676290 175084 676350 175424
rect 645135 174892 645201 174895
rect 640416 174890 645201 174892
rect 640416 174862 645140 174890
rect 640386 174834 645140 174862
rect 645196 174834 645201 174890
rect 640386 174832 645201 174834
rect 186255 174744 186321 174747
rect 186255 174742 190560 174744
rect 186255 174686 186260 174742
rect 186316 174686 190560 174742
rect 186255 174684 190560 174686
rect 186255 174681 186321 174684
rect 148911 174004 148977 174007
rect 143904 174002 148977 174004
rect 143904 173946 148916 174002
rect 148972 173946 148977 174002
rect 143904 173944 148977 173946
rect 148911 173941 148977 173944
rect 184431 174004 184497 174007
rect 184431 174002 190014 174004
rect 184431 173946 184436 174002
rect 184492 173946 190014 174002
rect 184431 173944 190014 173946
rect 184431 173941 184497 173944
rect 189954 173930 190014 173944
rect 189954 173870 190560 173930
rect 185583 173264 185649 173267
rect 185583 173262 190560 173264
rect 185583 173206 185588 173262
rect 185644 173206 190560 173262
rect 185583 173204 190560 173206
rect 185583 173201 185649 173204
rect 640386 172938 640446 174832
rect 645135 174829 645201 174832
rect 672399 174448 672465 174451
rect 676290 174448 676350 174714
rect 672399 174446 676350 174448
rect 672399 174390 672404 174446
rect 672460 174390 676350 174446
rect 672399 174388 676350 174390
rect 672399 174385 672465 174388
rect 673986 174004 674046 174388
rect 674170 174090 674176 174154
rect 674240 174152 674246 174154
rect 674240 174092 676320 174152
rect 674240 174090 674246 174092
rect 674170 174004 674176 174006
rect 673986 173944 674176 174004
rect 674170 173942 674176 173944
rect 674240 173942 674246 174006
rect 672591 173560 672657 173563
rect 673978 173560 673984 173562
rect 672591 173558 673984 173560
rect 672591 173502 672596 173558
rect 672652 173502 673984 173558
rect 672591 173500 673984 173502
rect 672591 173497 672657 173500
rect 673978 173498 673984 173500
rect 674048 173560 674054 173562
rect 674048 173500 676320 173560
rect 674048 173498 674054 173500
rect 675898 173202 675904 173266
rect 675968 173264 675974 173266
rect 675968 173204 676320 173264
rect 675968 173202 675974 173204
rect 149583 172820 149649 172823
rect 143904 172818 149649 172820
rect 143904 172762 149588 172818
rect 149644 172762 149649 172818
rect 143904 172760 149649 172762
rect 149583 172757 149649 172760
rect 184335 172524 184401 172527
rect 184335 172522 190014 172524
rect 184335 172466 184340 172522
rect 184396 172466 190014 172522
rect 184335 172464 190014 172466
rect 184335 172461 184401 172464
rect 189954 172450 190014 172464
rect 189954 172390 190560 172450
rect 676866 172379 676926 172642
rect 676866 172374 676977 172379
rect 676866 172318 676916 172374
rect 676972 172318 676977 172374
rect 676866 172316 676977 172318
rect 676911 172313 676977 172316
rect 675567 172080 675633 172083
rect 675567 172078 676320 172080
rect 675567 172022 675572 172078
rect 675628 172022 676320 172078
rect 675567 172020 676320 172022
rect 675567 172017 675633 172020
rect 184527 171784 184593 171787
rect 184527 171782 190560 171784
rect 184527 171726 184532 171782
rect 184588 171726 190560 171782
rect 184527 171724 190560 171726
rect 184527 171721 184593 171724
rect 676047 171710 676113 171713
rect 676047 171708 676320 171710
rect 676047 171652 676052 171708
rect 676108 171652 676320 171708
rect 676047 171650 676320 171652
rect 676047 171647 676113 171650
rect 143874 171044 143934 171532
rect 675130 171130 675136 171194
rect 675200 171192 675206 171194
rect 675200 171132 676320 171192
rect 675200 171130 675206 171132
rect 149199 171044 149265 171047
rect 645135 171044 645201 171047
rect 143874 171042 149265 171044
rect 143874 170986 149204 171042
rect 149260 170986 149265 171042
rect 640416 171042 645201 171044
rect 640416 171014 645140 171042
rect 143874 170984 149265 170986
rect 149199 170981 149265 170984
rect 640386 170986 645140 171014
rect 645196 170986 645201 171042
rect 640386 170984 645201 170986
rect 184623 170896 184689 170899
rect 184623 170894 190560 170896
rect 184623 170838 184628 170894
rect 184684 170838 190560 170894
rect 184623 170836 190560 170838
rect 184623 170833 184689 170836
rect 148719 170304 148785 170307
rect 143904 170302 148785 170304
rect 143904 170246 148724 170302
rect 148780 170246 148785 170302
rect 143904 170244 148785 170246
rect 148719 170241 148785 170244
rect 184431 170304 184497 170307
rect 184431 170302 190014 170304
rect 184431 170246 184436 170302
rect 184492 170246 190014 170302
rect 184431 170244 190014 170246
rect 184431 170241 184497 170244
rect 189954 170230 190014 170244
rect 189954 170170 190560 170230
rect 184335 169416 184401 169419
rect 184335 169414 190560 169416
rect 184335 169358 184340 169414
rect 184396 169358 190560 169414
rect 184335 169356 190560 169358
rect 184335 169353 184401 169356
rect 149487 169120 149553 169123
rect 143904 169118 149553 169120
rect 143904 169062 149492 169118
rect 149548 169062 149553 169118
rect 640386 169090 640446 170984
rect 645135 170981 645201 170984
rect 676866 170455 676926 170570
rect 676815 170450 676926 170455
rect 676815 170394 676820 170450
rect 676876 170394 676926 170450
rect 676815 170392 676926 170394
rect 676815 170389 676881 170392
rect 676047 170230 676113 170233
rect 676047 170228 676320 170230
rect 676047 170172 676052 170228
rect 676108 170172 676320 170228
rect 676047 170170 676320 170172
rect 676047 170167 676113 170170
rect 676047 169712 676113 169715
rect 676047 169710 676320 169712
rect 676047 169654 676052 169710
rect 676108 169654 676320 169710
rect 676047 169652 676320 169654
rect 676047 169649 676113 169652
rect 143904 169060 149553 169062
rect 149487 169057 149553 169060
rect 676290 168975 676350 169090
rect 676239 168970 676350 168975
rect 676239 168914 676244 168970
rect 676300 168914 676350 168970
rect 676239 168912 676350 168914
rect 676239 168909 676305 168912
rect 184431 168676 184497 168679
rect 184431 168674 190014 168676
rect 184431 168618 184436 168674
rect 184492 168618 190014 168674
rect 184431 168616 190014 168618
rect 184431 168613 184497 168616
rect 189954 168602 190014 168616
rect 674746 168614 674752 168678
rect 674816 168676 674822 168678
rect 674816 168616 676320 168676
rect 674816 168614 674822 168616
rect 189954 168542 190560 168602
rect 674938 168170 674944 168234
rect 675008 168232 675014 168234
rect 675008 168172 676320 168232
rect 675008 168170 675014 168172
rect 149007 168084 149073 168087
rect 143904 168082 149073 168084
rect 143904 168026 149012 168082
rect 149068 168026 149073 168082
rect 143904 168024 149073 168026
rect 149007 168021 149073 168024
rect 184623 167936 184689 167939
rect 184623 167934 190560 167936
rect 184623 167878 184628 167934
rect 184684 167878 190560 167934
rect 184623 167876 190560 167878
rect 184623 167873 184689 167876
rect 645135 167788 645201 167791
rect 640386 167786 645201 167788
rect 640386 167730 645140 167786
rect 645196 167730 645201 167786
rect 640386 167728 645201 167730
rect 184527 167196 184593 167199
rect 184527 167194 190014 167196
rect 184527 167138 184532 167194
rect 184588 167138 190014 167194
rect 184527 167136 190014 167138
rect 184527 167133 184593 167136
rect 189954 167122 190014 167136
rect 189954 167062 190560 167122
rect 143874 166308 143934 166796
rect 184335 166456 184401 166459
rect 184335 166454 190560 166456
rect 184335 166398 184340 166454
rect 184396 166398 190560 166454
rect 184335 166396 190560 166398
rect 184335 166393 184401 166396
rect 148719 166308 148785 166311
rect 143874 166306 148785 166308
rect 143874 166250 148724 166306
rect 148780 166250 148785 166306
rect 143874 166248 148785 166250
rect 148719 166245 148785 166248
rect 640386 166012 640446 167728
rect 645135 167725 645201 167728
rect 676047 167640 676113 167643
rect 676047 167638 676320 167640
rect 676047 167582 676052 167638
rect 676108 167582 676320 167638
rect 676047 167580 676320 167582
rect 676047 167577 676113 167580
rect 674554 167134 674560 167198
rect 674624 167196 674630 167198
rect 674624 167136 676320 167196
rect 674624 167134 674630 167136
rect 676047 166678 676113 166681
rect 676047 166676 676320 166678
rect 676047 166620 676052 166676
rect 676108 166620 676320 166676
rect 676047 166618 676320 166620
rect 676047 166615 676113 166618
rect 676047 166160 676113 166163
rect 676047 166158 676320 166160
rect 676047 166102 676052 166158
rect 676108 166102 676320 166158
rect 676047 166100 676320 166102
rect 676047 166097 676113 166100
rect 640194 165952 640446 166012
rect 184431 165716 184497 165719
rect 184431 165714 190014 165716
rect 184431 165658 184436 165714
rect 184492 165658 190014 165714
rect 184431 165656 190014 165658
rect 184431 165653 184497 165656
rect 189954 165642 190014 165656
rect 189954 165582 190560 165642
rect 148527 165568 148593 165571
rect 143904 165566 148593 165568
rect 143904 165510 148532 165566
rect 148588 165510 148593 165566
rect 143904 165508 148593 165510
rect 148527 165505 148593 165508
rect 640194 165242 640254 165952
rect 676143 165420 676209 165423
rect 676290 165420 676350 165686
rect 676143 165418 676350 165420
rect 676143 165362 676148 165418
rect 676204 165362 676350 165418
rect 676143 165360 676350 165362
rect 676143 165357 676209 165360
rect 676290 164831 676350 165168
rect 184527 164828 184593 164831
rect 184527 164826 190560 164828
rect 184527 164770 184532 164826
rect 184588 164770 190560 164826
rect 184527 164768 190560 164770
rect 676239 164826 676350 164831
rect 676239 164770 676244 164826
rect 676300 164770 676350 164826
rect 676239 164768 676350 164770
rect 184527 164765 184593 164768
rect 676239 164765 676305 164768
rect 148335 164384 148401 164387
rect 143904 164382 148401 164384
rect 143904 164326 148340 164382
rect 148396 164326 148401 164382
rect 143904 164324 148401 164326
rect 148335 164321 148401 164324
rect 184335 164088 184401 164091
rect 184335 164086 190560 164088
rect 184335 164030 184340 164086
rect 184396 164030 190560 164086
rect 184335 164028 190560 164030
rect 184335 164025 184401 164028
rect 184335 163348 184401 163351
rect 645135 163348 645201 163351
rect 184335 163346 190560 163348
rect 184335 163290 184340 163346
rect 184396 163290 190560 163346
rect 640416 163346 645201 163348
rect 640416 163318 645140 163346
rect 184335 163288 190560 163290
rect 640386 163290 645140 163318
rect 645196 163290 645201 163346
rect 640386 163288 645201 163290
rect 184335 163285 184401 163288
rect 148623 163200 148689 163203
rect 143904 163198 148689 163200
rect 143904 163142 148628 163198
rect 148684 163142 148689 163198
rect 143904 163140 148689 163142
rect 148623 163137 148689 163140
rect 185295 162608 185361 162611
rect 185295 162606 190560 162608
rect 185295 162550 185300 162606
rect 185356 162550 190560 162606
rect 185295 162548 190560 162550
rect 185295 162545 185361 162548
rect 148239 161868 148305 161871
rect 143904 161866 148305 161868
rect 143904 161810 148244 161866
rect 148300 161810 148305 161866
rect 143904 161808 148305 161810
rect 148239 161805 148305 161808
rect 184431 161868 184497 161871
rect 184431 161866 190560 161868
rect 184431 161810 184436 161866
rect 184492 161810 190560 161866
rect 184431 161808 190560 161810
rect 184431 161805 184497 161808
rect 640386 161394 640446 163288
rect 645135 163285 645201 163288
rect 675706 161510 675712 161574
rect 675776 161572 675782 161574
rect 676911 161572 676977 161575
rect 675776 161570 676977 161572
rect 675776 161514 676916 161570
rect 676972 161514 676977 161570
rect 675776 161512 676977 161514
rect 675776 161510 675782 161512
rect 676911 161509 676977 161512
rect 676666 161362 676672 161426
rect 676736 161424 676742 161426
rect 676815 161424 676881 161427
rect 676736 161422 676881 161424
rect 676736 161366 676820 161422
rect 676876 161366 676881 161422
rect 676736 161364 676881 161366
rect 676736 161362 676742 161364
rect 676815 161361 676881 161364
rect 184335 160980 184401 160983
rect 184335 160978 190560 160980
rect 184335 160922 184340 160978
rect 184396 160922 190560 160978
rect 184335 160920 190560 160922
rect 184335 160917 184401 160920
rect 148431 160684 148497 160687
rect 143904 160682 148497 160684
rect 143904 160626 148436 160682
rect 148492 160626 148497 160682
rect 143904 160624 148497 160626
rect 148431 160621 148497 160624
rect 184431 160388 184497 160391
rect 184431 160386 190014 160388
rect 184431 160330 184436 160386
rect 184492 160330 190014 160386
rect 184431 160328 190014 160330
rect 184431 160325 184497 160328
rect 189954 160314 190014 160328
rect 189954 160254 190560 160314
rect 146895 159500 146961 159503
rect 143904 159498 146961 159500
rect 143904 159442 146900 159498
rect 146956 159442 146961 159498
rect 143904 159440 146961 159442
rect 146895 159437 146961 159440
rect 184527 159500 184593 159503
rect 645135 159500 645201 159503
rect 184527 159498 190560 159500
rect 184527 159442 184532 159498
rect 184588 159442 190560 159498
rect 640416 159498 645201 159500
rect 640416 159470 645140 159498
rect 184527 159440 190560 159442
rect 640386 159442 645140 159470
rect 645196 159442 645201 159498
rect 640386 159440 645201 159442
rect 184527 159437 184593 159440
rect 184623 158908 184689 158911
rect 184623 158906 190014 158908
rect 184623 158850 184628 158906
rect 184684 158850 190014 158906
rect 184623 158848 190014 158850
rect 184623 158845 184689 158848
rect 189954 158834 190014 158848
rect 189954 158774 190560 158834
rect 143874 157724 143934 158212
rect 184527 158020 184593 158023
rect 184527 158018 190560 158020
rect 184527 157962 184532 158018
rect 184588 157962 190560 158018
rect 184527 157960 190560 157962
rect 184527 157957 184593 157960
rect 149295 157724 149361 157727
rect 143874 157722 149361 157724
rect 143874 157666 149300 157722
rect 149356 157666 149361 157722
rect 143874 157664 149361 157666
rect 149295 157661 149361 157664
rect 640386 157546 640446 159440
rect 645135 159437 645201 159440
rect 675759 159352 675825 159355
rect 675898 159352 675904 159354
rect 675759 159350 675904 159352
rect 675759 159294 675764 159350
rect 675820 159294 675904 159350
rect 675759 159292 675904 159294
rect 675759 159289 675825 159292
rect 675898 159290 675904 159292
rect 675968 159290 675974 159354
rect 184623 157428 184689 157431
rect 184623 157426 190014 157428
rect 184623 157370 184628 157426
rect 184684 157370 190014 157426
rect 184623 157368 190014 157370
rect 184623 157365 184689 157368
rect 189954 157354 190014 157368
rect 189954 157294 190560 157354
rect 149679 156984 149745 156987
rect 143904 156982 149745 156984
rect 143904 156926 149684 156982
rect 149740 156926 149745 156982
rect 143904 156924 149745 156926
rect 149679 156921 149745 156924
rect 184335 156540 184401 156543
rect 184335 156538 190560 156540
rect 184335 156482 184340 156538
rect 184396 156482 190560 156538
rect 184335 156480 190560 156482
rect 184335 156477 184401 156480
rect 148815 155800 148881 155803
rect 143904 155798 148881 155800
rect 143904 155742 148820 155798
rect 148876 155742 148881 155798
rect 143904 155740 148881 155742
rect 148815 155737 148881 155740
rect 184431 155652 184497 155655
rect 184431 155650 190560 155652
rect 184431 155594 184436 155650
rect 184492 155594 190560 155650
rect 184431 155592 190560 155594
rect 184431 155589 184497 155592
rect 640194 155504 640254 155622
rect 645135 155504 645201 155507
rect 640194 155502 645201 155504
rect 640194 155446 645140 155502
rect 645196 155446 645201 155502
rect 640194 155444 645201 155446
rect 184335 155060 184401 155063
rect 184335 155058 190560 155060
rect 184335 155002 184340 155058
rect 184396 155002 190560 155058
rect 184335 155000 190560 155002
rect 184335 154997 184401 155000
rect 149679 154616 149745 154619
rect 143904 154614 149745 154616
rect 143904 154558 149684 154614
rect 149740 154558 149745 154614
rect 143904 154556 149745 154558
rect 149679 154553 149745 154556
rect 184431 154172 184497 154175
rect 184431 154170 190560 154172
rect 184431 154114 184436 154170
rect 184492 154114 190560 154170
rect 184431 154112 190560 154114
rect 184431 154109 184497 154112
rect 640386 153772 640446 155444
rect 645135 155441 645201 155444
rect 184527 153580 184593 153583
rect 184527 153578 190014 153580
rect 184527 153522 184532 153578
rect 184588 153522 190014 153578
rect 184527 153520 190014 153522
rect 184527 153517 184593 153520
rect 189954 153506 190014 153520
rect 189954 153446 190560 153506
rect 675130 153370 675136 153434
rect 675200 153432 675206 153434
rect 675471 153432 675537 153435
rect 675200 153430 675537 153432
rect 675200 153374 675476 153430
rect 675532 153374 675537 153430
rect 675200 153372 675537 153374
rect 675200 153370 675206 153372
rect 675471 153369 675537 153372
rect 143874 153136 143934 153328
rect 149199 153136 149265 153139
rect 143874 153134 149265 153136
rect 143874 153078 149204 153134
rect 149260 153078 149265 153134
rect 143874 153076 149265 153078
rect 149199 153073 149265 153076
rect 184623 152692 184689 152695
rect 184623 152690 190560 152692
rect 184623 152634 184628 152690
rect 184684 152634 190560 152690
rect 184623 152632 190560 152634
rect 184623 152629 184689 152632
rect 645135 152544 645201 152547
rect 640194 152542 645201 152544
rect 640194 152486 645140 152542
rect 645196 152486 645201 152542
rect 640194 152484 645201 152486
rect 149199 152100 149265 152103
rect 143904 152098 149265 152100
rect 143904 152042 149204 152098
rect 149260 152042 149265 152098
rect 143904 152040 149265 152042
rect 149199 152037 149265 152040
rect 184335 151952 184401 151955
rect 184335 151950 190014 151952
rect 184335 151894 184340 151950
rect 184396 151894 190014 151950
rect 184335 151892 190014 151894
rect 184335 151889 184401 151892
rect 189954 151878 190014 151892
rect 189954 151818 190560 151878
rect 184527 151212 184593 151215
rect 184527 151210 190560 151212
rect 184527 151154 184532 151210
rect 184588 151154 190560 151210
rect 184527 151152 190560 151154
rect 184527 151149 184593 151152
rect 149679 150916 149745 150919
rect 143904 150914 149745 150916
rect 143904 150858 149684 150914
rect 149740 150858 149745 150914
rect 143904 150856 149745 150858
rect 149679 150853 149745 150856
rect 184431 150472 184497 150475
rect 184431 150470 190014 150472
rect 184431 150414 184436 150470
rect 184492 150414 190014 150470
rect 184431 150412 190014 150414
rect 184431 150409 184497 150412
rect 189954 150398 190014 150412
rect 189954 150338 190560 150398
rect 640194 149998 640254 152484
rect 645135 152481 645201 152484
rect 674554 152482 674560 152546
rect 674624 152544 674630 152546
rect 675375 152544 675441 152547
rect 674624 152542 675441 152544
rect 674624 152486 675380 152542
rect 675436 152486 675441 152542
rect 674624 152484 675441 152486
rect 674624 152482 674630 152484
rect 675375 152481 675441 152484
rect 674938 152186 674944 152250
rect 675008 152248 675014 152250
rect 675471 152248 675537 152251
rect 675008 152246 675537 152248
rect 675008 152190 675476 152246
rect 675532 152190 675537 152246
rect 675008 152188 675537 152190
rect 675008 152186 675014 152188
rect 675471 152185 675537 152188
rect 674746 150262 674752 150326
rect 674816 150324 674822 150326
rect 675471 150324 675537 150327
rect 674816 150322 675537 150324
rect 674816 150266 675476 150322
rect 675532 150266 675537 150322
rect 674816 150264 675537 150266
rect 674816 150262 674822 150264
rect 675471 150261 675537 150264
rect 149199 149880 149265 149883
rect 143874 149878 149265 149880
rect 143874 149822 149204 149878
rect 149260 149822 149265 149878
rect 143874 149820 149265 149822
rect 143874 149776 143934 149820
rect 149199 149817 149265 149820
rect 184335 149732 184401 149735
rect 184335 149730 190560 149732
rect 184335 149674 184340 149730
rect 184396 149674 190560 149730
rect 184335 149672 190560 149674
rect 184335 149669 184401 149672
rect 184431 148992 184497 148995
rect 184431 148990 190014 148992
rect 184431 148934 184436 148990
rect 184492 148934 190014 148990
rect 184431 148932 190014 148934
rect 184431 148929 184497 148932
rect 189954 148918 190014 148932
rect 189954 148858 190560 148918
rect 149679 148548 149745 148551
rect 675759 148550 675825 148551
rect 143904 148546 149745 148548
rect 143904 148490 149684 148546
rect 149740 148490 149745 148546
rect 143904 148488 149745 148490
rect 149679 148485 149745 148488
rect 675706 148486 675712 148550
rect 675776 148548 675825 148550
rect 675776 148546 675868 148548
rect 675820 148490 675868 148546
rect 675776 148488 675868 148490
rect 675776 148486 675825 148488
rect 675759 148485 675825 148486
rect 184335 148104 184401 148107
rect 645135 148104 645201 148107
rect 184335 148102 190560 148104
rect 184335 148046 184340 148102
rect 184396 148046 190560 148102
rect 640416 148102 645201 148104
rect 640416 148074 645140 148102
rect 184335 148044 190560 148046
rect 640386 148046 645140 148074
rect 645196 148046 645201 148102
rect 640386 148044 645201 148046
rect 184335 148041 184401 148044
rect 149199 147364 149265 147367
rect 143904 147362 149265 147364
rect 143904 147306 149204 147362
rect 149260 147306 149265 147362
rect 143904 147304 149265 147306
rect 149199 147301 149265 147304
rect 184527 147364 184593 147367
rect 184527 147362 190560 147364
rect 184527 147306 184532 147362
rect 184588 147306 190560 147362
rect 184527 147304 190560 147306
rect 184527 147301 184593 147304
rect 185391 146624 185457 146627
rect 185391 146622 190560 146624
rect 185391 146566 185396 146622
rect 185452 146566 190560 146622
rect 185391 146564 190560 146566
rect 185391 146561 185457 146564
rect 149679 146180 149745 146183
rect 143904 146178 149745 146180
rect 143904 146122 149684 146178
rect 149740 146122 149745 146178
rect 640386 146150 640446 148044
rect 645135 148041 645201 148044
rect 675759 146624 675825 146627
rect 676666 146624 676672 146626
rect 675759 146622 676672 146624
rect 675759 146566 675764 146622
rect 675820 146566 676672 146622
rect 675759 146564 676672 146566
rect 675759 146561 675825 146564
rect 676666 146562 676672 146564
rect 676736 146562 676742 146626
rect 143904 146120 149745 146122
rect 149679 146117 149745 146120
rect 186735 145884 186801 145887
rect 186735 145882 190560 145884
rect 186735 145826 186740 145882
rect 186796 145826 190560 145882
rect 186735 145824 190560 145826
rect 186735 145821 186801 145824
rect 184335 145144 184401 145147
rect 184335 145142 190014 145144
rect 184335 145086 184340 145142
rect 184396 145086 190014 145142
rect 184335 145084 190014 145086
rect 184335 145081 184401 145084
rect 189954 145070 190014 145084
rect 189954 145010 190560 145070
rect 143874 144552 143934 144892
rect 149199 144552 149265 144555
rect 143874 144550 149265 144552
rect 143874 144494 149204 144550
rect 149260 144494 149265 144550
rect 143874 144492 149265 144494
rect 149199 144489 149265 144492
rect 184431 144404 184497 144407
rect 184431 144402 190560 144404
rect 184431 144346 184436 144402
rect 184492 144346 190560 144402
rect 184431 144344 190560 144346
rect 184431 144341 184497 144344
rect 646671 144256 646737 144259
rect 640416 144254 646737 144256
rect 640416 144226 646676 144254
rect 640386 144198 646676 144226
rect 646732 144198 646737 144254
rect 640386 144196 646737 144198
rect 149679 143664 149745 143667
rect 143904 143662 149745 143664
rect 143904 143606 149684 143662
rect 149740 143606 149745 143662
rect 143904 143604 149745 143606
rect 149679 143601 149745 143604
rect 184623 143664 184689 143667
rect 184623 143662 190014 143664
rect 184623 143606 184628 143662
rect 184684 143606 190014 143662
rect 184623 143604 190014 143606
rect 184623 143601 184689 143604
rect 189954 143590 190014 143604
rect 189954 143530 190560 143590
rect 184335 142776 184401 142779
rect 184335 142774 190560 142776
rect 184335 142718 184340 142774
rect 184396 142718 190560 142774
rect 184335 142716 190560 142718
rect 184335 142713 184401 142716
rect 149199 142480 149265 142483
rect 143904 142478 149265 142480
rect 143904 142422 149204 142478
rect 149260 142422 149265 142478
rect 143904 142420 149265 142422
rect 149199 142417 149265 142420
rect 640386 142302 640446 144196
rect 646671 144193 646737 144196
rect 184431 142184 184497 142187
rect 184431 142182 190014 142184
rect 184431 142126 184436 142182
rect 184492 142126 190014 142182
rect 184431 142124 190014 142126
rect 184431 142121 184497 142124
rect 189954 142110 190014 142124
rect 189954 142050 190560 142110
rect 148815 141296 148881 141299
rect 143904 141294 148881 141296
rect 143904 141238 148820 141294
rect 148876 141238 148881 141294
rect 143904 141236 148881 141238
rect 148815 141233 148881 141236
rect 184527 141296 184593 141299
rect 184527 141294 190560 141296
rect 184527 141238 184532 141294
rect 184588 141238 190560 141294
rect 184527 141236 190560 141238
rect 184527 141233 184593 141236
rect 646767 141000 646833 141003
rect 640386 140998 646833 141000
rect 640386 140942 646772 140998
rect 646828 140942 646833 140998
rect 640386 140940 646833 140942
rect 184335 140556 184401 140559
rect 184335 140554 190560 140556
rect 184335 140498 184340 140554
rect 184396 140498 190560 140554
rect 184335 140496 190560 140498
rect 184335 140493 184401 140496
rect 640386 140408 640446 140940
rect 646767 140937 646833 140940
rect 640224 140378 640446 140408
rect 640194 140348 640416 140378
rect 147087 139964 147153 139967
rect 143904 139962 147153 139964
rect 143904 139906 147092 139962
rect 147148 139906 147153 139962
rect 143904 139904 147153 139906
rect 147087 139901 147153 139904
rect 184431 139816 184497 139819
rect 184431 139814 190560 139816
rect 184431 139758 184436 139814
rect 184492 139758 190560 139814
rect 184431 139756 190560 139758
rect 184431 139753 184497 139756
rect 184527 138928 184593 138931
rect 184527 138926 190560 138928
rect 184527 138870 184532 138926
rect 184588 138870 190560 138926
rect 184527 138868 190560 138870
rect 184527 138865 184593 138868
rect 149199 138780 149265 138783
rect 143904 138778 149265 138780
rect 143904 138722 149204 138778
rect 149260 138722 149265 138778
rect 143904 138720 149265 138722
rect 149199 138717 149265 138720
rect 640194 138528 640254 140348
rect 186063 138336 186129 138339
rect 186063 138334 190560 138336
rect 186063 138278 186068 138334
rect 186124 138278 190560 138334
rect 186063 138276 190560 138278
rect 186063 138273 186129 138276
rect 149679 137596 149745 137599
rect 143904 137594 149745 137596
rect 143904 137538 149684 137594
rect 149740 137538 149745 137594
rect 143904 137536 149745 137538
rect 149679 137533 149745 137536
rect 186159 137448 186225 137451
rect 186159 137446 190560 137448
rect 186159 137390 186164 137446
rect 186220 137390 190560 137446
rect 186159 137388 190560 137390
rect 186159 137385 186225 137388
rect 185967 136856 186033 136859
rect 185967 136854 190014 136856
rect 185967 136798 185972 136854
rect 186028 136798 190014 136854
rect 185967 136796 190014 136798
rect 185967 136793 186033 136796
rect 189954 136782 190014 136796
rect 189954 136722 190560 136782
rect 143874 135968 143934 136308
rect 149199 135968 149265 135971
rect 143874 135966 149265 135968
rect 143874 135910 149204 135966
rect 149260 135910 149265 135966
rect 143874 135908 149265 135910
rect 149199 135905 149265 135908
rect 185487 135968 185553 135971
rect 185487 135966 190560 135968
rect 185487 135910 185492 135966
rect 185548 135910 190560 135966
rect 185487 135908 190560 135910
rect 185487 135905 185553 135908
rect 186255 135228 186321 135231
rect 186255 135226 190014 135228
rect 186255 135170 186260 135226
rect 186316 135170 190014 135226
rect 186255 135168 190014 135170
rect 186255 135165 186321 135168
rect 189954 135154 190014 135168
rect 189954 135094 190560 135154
rect 149487 135080 149553 135083
rect 143904 135078 149553 135080
rect 143904 135022 149492 135078
rect 149548 135022 149553 135078
rect 143904 135020 149553 135022
rect 149487 135017 149553 135020
rect 647055 134784 647121 134787
rect 640416 134782 647121 134784
rect 640416 134726 647060 134782
rect 647116 134726 647121 134782
rect 640416 134724 647121 134726
rect 647055 134721 647121 134724
rect 184335 134488 184401 134491
rect 184335 134486 190560 134488
rect 184335 134430 184340 134486
rect 184396 134430 190560 134486
rect 184335 134428 190560 134430
rect 184335 134425 184401 134428
rect 149391 133896 149457 133899
rect 143904 133894 149457 133896
rect 143904 133838 149396 133894
rect 149452 133838 149457 133894
rect 143904 133836 149457 133838
rect 149391 133833 149457 133836
rect 184431 133748 184497 133751
rect 184431 133746 190014 133748
rect 184431 133690 184436 133746
rect 184492 133690 190014 133746
rect 184431 133688 190014 133690
rect 184431 133685 184497 133688
rect 189954 133674 190014 133688
rect 189954 133614 190560 133674
rect 184527 133008 184593 133011
rect 184527 133006 190560 133008
rect 184527 132950 184532 133006
rect 184588 132950 190560 133006
rect 184527 132948 190560 132950
rect 184527 132945 184593 132948
rect 148815 132712 148881 132715
rect 143904 132710 148881 132712
rect 143904 132654 148820 132710
rect 148876 132654 148881 132710
rect 143904 132652 148881 132654
rect 148815 132649 148881 132652
rect 184623 132268 184689 132271
rect 184623 132266 190014 132268
rect 184623 132210 184628 132266
rect 184684 132210 190014 132266
rect 184623 132208 190014 132210
rect 184623 132205 184689 132208
rect 189954 132194 190014 132208
rect 189954 132134 190560 132194
rect 676143 131824 676209 131827
rect 676290 131824 676350 132090
rect 676143 131822 676350 131824
rect 676143 131766 676148 131822
rect 676204 131766 676350 131822
rect 676143 131764 676350 131766
rect 676143 131761 676209 131764
rect 184335 131528 184401 131531
rect 184335 131526 190560 131528
rect 184335 131470 184340 131526
rect 184396 131470 190560 131526
rect 184335 131468 190560 131470
rect 184335 131465 184401 131468
rect 143874 130936 143934 131424
rect 676290 131235 676350 131498
rect 676290 131230 676401 131235
rect 676290 131174 676340 131230
rect 676396 131174 676401 131230
rect 676290 131172 676401 131174
rect 676335 131169 676401 131172
rect 148911 130936 148977 130939
rect 647823 130936 647889 130939
rect 143874 130934 148977 130936
rect 143874 130878 148916 130934
rect 148972 130878 148977 130934
rect 143874 130876 148977 130878
rect 640416 130934 647889 130936
rect 640416 130878 647828 130934
rect 647884 130878 647889 130934
rect 640416 130876 647889 130878
rect 148911 130873 148977 130876
rect 647823 130873 647889 130876
rect 676290 130791 676350 130980
rect 676239 130786 676350 130791
rect 676239 130730 676244 130786
rect 676300 130730 676350 130786
rect 676239 130728 676350 130730
rect 676239 130725 676305 130728
rect 184527 130640 184593 130643
rect 184527 130638 190560 130640
rect 184527 130582 184532 130638
rect 184588 130582 190560 130638
rect 184527 130580 190560 130582
rect 184527 130577 184593 130580
rect 674362 130578 674368 130642
rect 674432 130640 674438 130642
rect 674432 130580 676320 130640
rect 674432 130578 674438 130580
rect 147183 130344 147249 130347
rect 143904 130342 147249 130344
rect 143904 130286 147188 130342
rect 147244 130286 147249 130342
rect 143904 130284 147249 130286
rect 147183 130281 147249 130284
rect 184431 129900 184497 129903
rect 184431 129898 190560 129900
rect 184431 129842 184436 129898
rect 184492 129842 190560 129898
rect 184431 129840 190560 129842
rect 184431 129837 184497 129840
rect 676290 129755 676350 130018
rect 676239 129750 676350 129755
rect 676239 129694 676244 129750
rect 676300 129694 676350 129750
rect 676239 129692 676350 129694
rect 676239 129689 676305 129692
rect 674170 129394 674176 129458
rect 674240 129456 674246 129458
rect 674240 129396 676320 129456
rect 674240 129394 674246 129396
rect 148527 129160 148593 129163
rect 143904 129158 148593 129160
rect 143904 129102 148532 129158
rect 148588 129102 148593 129158
rect 143904 129100 148593 129102
rect 148527 129097 148593 129100
rect 184335 129160 184401 129163
rect 184335 129158 190560 129160
rect 184335 129102 184340 129158
rect 184396 129102 190560 129158
rect 184335 129100 190560 129102
rect 184335 129097 184401 129100
rect 645711 129012 645777 129015
rect 640416 129010 645777 129012
rect 640416 128954 645716 129010
rect 645772 128954 645777 129010
rect 640416 128952 645777 128954
rect 645711 128949 645777 128952
rect 676143 128864 676209 128867
rect 676290 128864 676350 129130
rect 676143 128862 676350 128864
rect 676143 128806 676148 128862
rect 676204 128806 676350 128862
rect 676143 128804 676350 128806
rect 676143 128801 676209 128804
rect 673978 128506 673984 128570
rect 674048 128568 674054 128570
rect 674048 128508 676320 128568
rect 674048 128506 674054 128508
rect 184431 128420 184497 128423
rect 184431 128418 190014 128420
rect 184431 128362 184436 128418
rect 184492 128362 190014 128418
rect 184431 128360 190014 128362
rect 184431 128357 184497 128360
rect 189954 128346 190014 128360
rect 189954 128286 190560 128346
rect 149103 127976 149169 127979
rect 143904 127974 149169 127976
rect 143904 127918 149108 127974
rect 149164 127918 149169 127974
rect 143904 127916 149169 127918
rect 149103 127913 149169 127916
rect 676290 127831 676350 127946
rect 676239 127826 676350 127831
rect 676239 127770 676244 127826
rect 676300 127770 676350 127826
rect 676239 127768 676350 127770
rect 676239 127765 676305 127768
rect 184527 127680 184593 127683
rect 646959 127680 647025 127683
rect 184527 127678 190560 127680
rect 184527 127622 184532 127678
rect 184588 127622 190560 127678
rect 184527 127620 190560 127622
rect 640386 127678 647025 127680
rect 640386 127622 646964 127678
rect 647020 127622 647025 127678
rect 640386 127620 647025 127622
rect 184527 127617 184593 127620
rect 640386 127058 640446 127620
rect 646959 127617 647025 127620
rect 676047 127606 676113 127609
rect 676047 127604 676320 127606
rect 676047 127548 676052 127604
rect 676108 127548 676320 127604
rect 676047 127546 676320 127548
rect 676047 127543 676113 127546
rect 184623 126940 184689 126943
rect 184623 126938 190014 126940
rect 184623 126882 184628 126938
rect 184684 126882 190014 126938
rect 184623 126880 190014 126882
rect 184623 126877 184689 126880
rect 189954 126866 190014 126880
rect 189954 126806 190560 126866
rect 676866 126795 676926 127058
rect 676866 126790 676977 126795
rect 676866 126734 676916 126790
rect 676972 126734 676977 126790
rect 676866 126732 676977 126734
rect 676911 126729 676977 126732
rect 149583 126644 149649 126647
rect 143904 126642 149649 126644
rect 143904 126586 149588 126642
rect 149644 126586 149649 126642
rect 143904 126584 149649 126586
rect 149583 126581 149649 126584
rect 676290 126351 676350 126466
rect 676239 126346 676350 126351
rect 676239 126290 676244 126346
rect 676300 126290 676350 126346
rect 676239 126288 676350 126290
rect 676239 126285 676305 126288
rect 676047 126126 676113 126129
rect 676047 126124 676320 126126
rect 676047 126068 676052 126124
rect 676108 126068 676320 126124
rect 676047 126066 676320 126068
rect 676047 126063 676113 126066
rect 184431 126052 184497 126055
rect 184431 126050 190560 126052
rect 184431 125994 184436 126050
rect 184492 125994 190560 126050
rect 184431 125992 190560 125994
rect 184431 125989 184497 125992
rect 646863 125756 646929 125759
rect 640386 125754 646929 125756
rect 640386 125698 646868 125754
rect 646924 125698 646929 125754
rect 640386 125696 646929 125698
rect 148143 125460 148209 125463
rect 143904 125458 148209 125460
rect 143904 125402 148148 125458
rect 148204 125402 148209 125458
rect 143904 125400 148209 125402
rect 148143 125397 148209 125400
rect 184335 125460 184401 125463
rect 184335 125458 190014 125460
rect 184335 125402 184340 125458
rect 184396 125402 190014 125458
rect 184335 125400 190014 125402
rect 184335 125397 184401 125400
rect 189954 125386 190014 125400
rect 189954 125326 190560 125386
rect 640386 125208 640446 125696
rect 646863 125693 646929 125696
rect 674362 125546 674368 125610
rect 674432 125608 674438 125610
rect 674432 125548 676320 125608
rect 674432 125546 674438 125548
rect 676866 124871 676926 124986
rect 676815 124866 676926 124871
rect 676815 124810 676820 124866
rect 676876 124810 676926 124866
rect 676815 124808 676926 124810
rect 676815 124805 676881 124808
rect 184527 124572 184593 124575
rect 676047 124572 676113 124575
rect 184527 124570 190560 124572
rect 184527 124514 184532 124570
rect 184588 124514 190560 124570
rect 184527 124512 190560 124514
rect 676047 124570 676320 124572
rect 676047 124514 676052 124570
rect 676108 124514 676320 124570
rect 676047 124512 676320 124514
rect 184527 124509 184593 124512
rect 676047 124509 676113 124512
rect 149295 124276 149361 124279
rect 143904 124274 149361 124276
rect 143904 124218 149300 124274
rect 149356 124218 149361 124274
rect 143904 124216 149361 124218
rect 149295 124213 149361 124216
rect 675951 124128 676017 124131
rect 675951 124126 676320 124128
rect 675951 124070 675956 124126
rect 676012 124070 676320 124126
rect 675951 124068 676320 124070
rect 675951 124065 676017 124068
rect 184335 123832 184401 123835
rect 646575 123832 646641 123835
rect 184335 123830 190560 123832
rect 184335 123774 184340 123830
rect 184396 123774 190560 123830
rect 184335 123772 190560 123774
rect 640194 123830 646641 123832
rect 640194 123774 646580 123830
rect 646636 123774 646641 123830
rect 640194 123772 646641 123774
rect 184335 123769 184401 123772
rect 640194 123358 640254 123772
rect 646575 123769 646641 123772
rect 676047 123536 676113 123539
rect 676047 123534 676320 123536
rect 676047 123478 676052 123534
rect 676108 123478 676320 123534
rect 676047 123476 676320 123478
rect 676047 123473 676113 123476
rect 184431 123092 184497 123095
rect 184431 123090 190560 123092
rect 184431 123034 184436 123090
rect 184492 123034 190560 123090
rect 184431 123032 190560 123034
rect 184431 123029 184497 123032
rect 674554 123030 674560 123094
rect 674624 123092 674630 123094
rect 674624 123032 676320 123092
rect 674624 123030 674630 123032
rect 143874 122500 143934 122988
rect 149007 122500 149073 122503
rect 143874 122498 149073 122500
rect 143874 122442 149012 122498
rect 149068 122442 149073 122498
rect 143874 122440 149073 122442
rect 149007 122437 149073 122440
rect 184335 122204 184401 122207
rect 184335 122202 190560 122204
rect 184335 122146 184340 122202
rect 184396 122146 190560 122202
rect 184335 122144 190560 122146
rect 184335 122141 184401 122144
rect 673978 122142 673984 122206
rect 674048 122204 674054 122206
rect 676290 122204 676350 122544
rect 674048 122144 676350 122204
rect 674048 122142 674054 122144
rect 646479 122056 646545 122059
rect 640194 122054 646545 122056
rect 640194 121998 646484 122054
rect 646540 121998 646545 122054
rect 640194 121996 646545 121998
rect 149199 121760 149265 121763
rect 143904 121758 149265 121760
rect 143904 121702 149204 121758
rect 149260 121702 149265 121758
rect 143904 121700 149265 121702
rect 149199 121697 149265 121700
rect 184527 121612 184593 121615
rect 184527 121610 190560 121612
rect 184527 121554 184532 121610
rect 184588 121554 190560 121610
rect 184527 121552 190560 121554
rect 184527 121549 184593 121552
rect 640194 121434 640254 121996
rect 646479 121993 646545 121996
rect 676047 122056 676113 122059
rect 676047 122054 676320 122056
rect 676047 121998 676052 122054
rect 676108 121998 676320 122054
rect 676047 121996 676320 121998
rect 676047 121993 676113 121996
rect 676290 121467 676350 121582
rect 676239 121462 676350 121467
rect 676239 121406 676244 121462
rect 676300 121406 676350 121462
rect 676239 121404 676350 121406
rect 676239 121401 676305 121404
rect 676047 121094 676113 121097
rect 676047 121092 676320 121094
rect 676047 121036 676052 121092
rect 676108 121036 676320 121092
rect 676047 121034 676320 121036
rect 676047 121031 676113 121034
rect 184431 120724 184497 120727
rect 184431 120722 190560 120724
rect 184431 120666 184436 120722
rect 184492 120666 190560 120722
rect 184431 120664 190560 120666
rect 184431 120661 184497 120664
rect 149391 120576 149457 120579
rect 143904 120574 149457 120576
rect 143904 120518 149396 120574
rect 149452 120518 149457 120574
rect 143904 120516 149457 120518
rect 149391 120513 149457 120516
rect 676047 120576 676113 120579
rect 676047 120574 676320 120576
rect 676047 120518 676052 120574
rect 676108 120518 676320 120574
rect 676047 120516 676320 120518
rect 676047 120513 676113 120516
rect 184527 120132 184593 120135
rect 184527 120130 190014 120132
rect 184527 120074 184532 120130
rect 184588 120074 190014 120130
rect 184527 120072 190014 120074
rect 184527 120069 184593 120072
rect 189954 120058 190014 120072
rect 189954 119998 190560 120058
rect 676143 119836 676209 119839
rect 676290 119836 676350 120102
rect 676143 119834 676350 119836
rect 676143 119778 676148 119834
rect 676204 119778 676350 119834
rect 676143 119776 676350 119778
rect 676143 119773 676209 119776
rect 647919 119540 647985 119543
rect 640416 119538 647985 119540
rect 640416 119482 647924 119538
rect 647980 119482 647985 119538
rect 640416 119480 647985 119482
rect 647919 119477 647985 119480
rect 149487 119392 149553 119395
rect 143904 119390 149553 119392
rect 143904 119334 149492 119390
rect 149548 119334 149553 119390
rect 143904 119332 149553 119334
rect 149487 119329 149553 119332
rect 676290 119247 676350 119510
rect 184335 119244 184401 119247
rect 184335 119242 190560 119244
rect 184335 119186 184340 119242
rect 184396 119186 190560 119242
rect 184335 119184 190560 119186
rect 676239 119242 676350 119247
rect 676239 119186 676244 119242
rect 676300 119186 676350 119242
rect 676239 119184 676350 119186
rect 184335 119181 184401 119184
rect 676239 119181 676305 119184
rect 184623 118652 184689 118655
rect 184623 118650 190014 118652
rect 184623 118594 184628 118650
rect 184684 118594 190014 118650
rect 184623 118592 190014 118594
rect 184623 118589 184689 118592
rect 189954 118578 190014 118592
rect 189954 118518 190560 118578
rect 149391 118208 149457 118211
rect 143874 118206 149457 118208
rect 143874 118150 149396 118206
rect 149452 118150 149457 118206
rect 143874 118148 149457 118150
rect 143874 118104 143934 118148
rect 149391 118145 149457 118148
rect 676474 117998 676480 118062
rect 676544 118060 676550 118062
rect 676815 118060 676881 118063
rect 676544 118058 676881 118060
rect 676544 118002 676820 118058
rect 676876 118002 676881 118058
rect 676544 118000 676881 118002
rect 676544 117998 676550 118000
rect 676815 117997 676881 118000
rect 675898 117850 675904 117914
rect 675968 117912 675974 117914
rect 676911 117912 676977 117915
rect 675968 117910 676977 117912
rect 675968 117854 676916 117910
rect 676972 117854 676977 117910
rect 675968 117852 676977 117854
rect 675968 117850 675974 117852
rect 676911 117849 676977 117852
rect 184335 117764 184401 117767
rect 184335 117762 190560 117764
rect 184335 117706 184340 117762
rect 184396 117706 190560 117762
rect 184335 117704 190560 117706
rect 184335 117701 184401 117704
rect 645231 117616 645297 117619
rect 640416 117614 645297 117616
rect 640416 117558 645236 117614
rect 645292 117558 645297 117614
rect 640416 117556 645297 117558
rect 645231 117553 645297 117556
rect 184431 117024 184497 117027
rect 184431 117022 190014 117024
rect 184431 116966 184436 117022
rect 184492 116966 190014 117022
rect 184431 116964 190014 116966
rect 184431 116961 184497 116964
rect 189954 116950 190014 116964
rect 189954 116890 190560 116950
rect 149391 116876 149457 116879
rect 143904 116874 149457 116876
rect 143904 116818 149396 116874
rect 149452 116818 149457 116874
rect 143904 116816 149457 116818
rect 149391 116813 149457 116816
rect 184527 116284 184593 116287
rect 184527 116282 190560 116284
rect 184527 116226 184532 116282
rect 184588 116226 190560 116282
rect 184527 116224 190560 116226
rect 184527 116221 184593 116224
rect 149487 115692 149553 115695
rect 647919 115692 647985 115695
rect 143904 115690 149553 115692
rect 143904 115634 149492 115690
rect 149548 115634 149553 115690
rect 143904 115632 149553 115634
rect 640416 115690 647985 115692
rect 640416 115634 647924 115690
rect 647980 115634 647985 115690
rect 640416 115632 647985 115634
rect 149487 115629 149553 115632
rect 647919 115629 647985 115632
rect 184623 115396 184689 115399
rect 184623 115394 190560 115396
rect 184623 115338 184628 115394
rect 184684 115338 190560 115394
rect 184623 115336 190560 115338
rect 184623 115333 184689 115336
rect 148527 115248 148593 115251
rect 149391 115248 149457 115251
rect 148527 115246 149457 115248
rect 148527 115190 148532 115246
rect 148588 115190 149396 115246
rect 149452 115190 149457 115246
rect 148527 115188 149457 115190
rect 148527 115185 148593 115188
rect 149391 115185 149457 115188
rect 184335 114804 184401 114807
rect 184335 114802 190560 114804
rect 184335 114746 184340 114802
rect 184396 114746 190560 114802
rect 184335 114744 190560 114746
rect 184335 114741 184401 114744
rect 149487 114508 149553 114511
rect 143904 114506 149553 114508
rect 143904 114450 149492 114506
rect 149548 114450 149553 114506
rect 143904 114448 149553 114450
rect 149487 114445 149553 114448
rect 184431 113916 184497 113919
rect 184431 113914 190560 113916
rect 184431 113858 184436 113914
rect 184492 113858 190560 113914
rect 184431 113856 190560 113858
rect 184431 113853 184497 113856
rect 149391 113176 149457 113179
rect 143904 113174 149457 113176
rect 143904 113118 149396 113174
rect 149452 113118 149457 113174
rect 143904 113116 149457 113118
rect 149391 113113 149457 113116
rect 184527 113176 184593 113179
rect 640194 113176 640254 113738
rect 646575 113176 646641 113179
rect 184527 113174 190560 113176
rect 184527 113118 184532 113174
rect 184588 113118 190560 113174
rect 184527 113116 190560 113118
rect 640194 113174 646641 113176
rect 640194 113118 646580 113174
rect 646636 113118 646641 113174
rect 640194 113116 646641 113118
rect 184527 113113 184593 113116
rect 646575 113113 646641 113116
rect 185679 112436 185745 112439
rect 185679 112434 190560 112436
rect 185679 112378 185684 112434
rect 185740 112378 190560 112434
rect 185679 112376 190560 112378
rect 185679 112373 185745 112376
rect 148239 111992 148305 111995
rect 143904 111990 148305 111992
rect 143904 111934 148244 111990
rect 148300 111934 148305 111990
rect 143904 111932 148305 111934
rect 148239 111929 148305 111932
rect 184335 111696 184401 111699
rect 184335 111694 190014 111696
rect 184335 111638 184340 111694
rect 184396 111638 190014 111694
rect 184335 111636 190014 111638
rect 184335 111633 184401 111636
rect 189954 111622 190014 111636
rect 189954 111562 190560 111622
rect 640386 111400 640446 111888
rect 647055 111400 647121 111403
rect 640386 111398 647121 111400
rect 640386 111342 647060 111398
rect 647116 111342 647121 111398
rect 640386 111340 647121 111342
rect 647055 111337 647121 111340
rect 148431 110956 148497 110959
rect 143904 110954 148497 110956
rect 143904 110898 148436 110954
rect 148492 110898 148497 110954
rect 143904 110896 148497 110898
rect 148431 110893 148497 110896
rect 184431 110956 184497 110959
rect 184431 110954 190560 110956
rect 184431 110898 184436 110954
rect 184492 110898 190560 110954
rect 184431 110896 190560 110898
rect 184431 110893 184497 110896
rect 184527 110216 184593 110219
rect 184527 110214 190014 110216
rect 184527 110158 184532 110214
rect 184588 110158 190014 110214
rect 184527 110156 190014 110158
rect 184527 110153 184593 110156
rect 189954 110142 190014 110156
rect 189954 110082 190560 110142
rect 143874 109624 143934 109668
rect 149391 109624 149457 109627
rect 143874 109622 149457 109624
rect 143874 109566 149396 109622
rect 149452 109566 149457 109622
rect 143874 109564 149457 109566
rect 149391 109561 149457 109564
rect 640386 109476 640446 109890
rect 646671 109476 646737 109479
rect 640386 109474 646737 109476
rect 640386 109418 646676 109474
rect 646732 109418 646737 109474
rect 640386 109416 646737 109418
rect 646671 109413 646737 109416
rect 184431 109328 184497 109331
rect 184431 109326 190560 109328
rect 184431 109270 184436 109326
rect 184492 109270 190560 109326
rect 184431 109268 190560 109270
rect 184431 109265 184497 109268
rect 185583 108736 185649 108739
rect 185583 108734 190014 108736
rect 185583 108678 185588 108734
rect 185644 108678 190014 108734
rect 185583 108676 190014 108678
rect 185583 108673 185649 108676
rect 189954 108662 190014 108676
rect 189954 108602 190560 108662
rect 147663 108440 147729 108443
rect 143904 108438 147729 108440
rect 143904 108382 147668 108438
rect 147724 108382 147729 108438
rect 143904 108380 147729 108382
rect 147663 108377 147729 108380
rect 674362 108082 674368 108146
rect 674432 108144 674438 108146
rect 675375 108144 675441 108147
rect 674432 108142 675441 108144
rect 674432 108086 675380 108142
rect 675436 108086 675441 108142
rect 674432 108084 675441 108086
rect 674432 108082 674438 108084
rect 675375 108081 675441 108084
rect 646767 107996 646833 107999
rect 640416 107994 646833 107996
rect 640416 107938 646772 107994
rect 646828 107938 646833 107994
rect 640416 107936 646833 107938
rect 646767 107933 646833 107936
rect 186159 107848 186225 107851
rect 186159 107846 190560 107848
rect 186159 107790 186164 107846
rect 186220 107790 190560 107846
rect 186159 107788 190560 107790
rect 186159 107785 186225 107788
rect 146991 107256 147057 107259
rect 143904 107254 147057 107256
rect 143904 107198 146996 107254
rect 147052 107198 147057 107254
rect 143904 107196 147057 107198
rect 146991 107193 147057 107196
rect 184335 107108 184401 107111
rect 184335 107106 190560 107108
rect 184335 107050 184340 107106
rect 184396 107050 190560 107106
rect 184335 107048 190560 107050
rect 184335 107045 184401 107048
rect 673978 106602 673984 106666
rect 674048 106664 674054 106666
rect 675471 106664 675537 106667
rect 674048 106662 675537 106664
rect 674048 106606 675476 106662
rect 675532 106606 675537 106662
rect 674048 106604 675537 106606
rect 674048 106602 674054 106604
rect 675471 106601 675537 106604
rect 184335 106368 184401 106371
rect 668175 106368 668241 106371
rect 184335 106366 190560 106368
rect 184335 106310 184340 106366
rect 184396 106310 190560 106366
rect 184335 106308 190560 106310
rect 665346 106366 668241 106368
rect 665346 106310 668180 106366
rect 668236 106310 668241 106366
rect 665346 106308 668241 106310
rect 184335 106305 184401 106308
rect 665346 106082 665406 106308
rect 668175 106305 668241 106308
rect 148527 106072 148593 106075
rect 645711 106072 645777 106075
rect 143904 106070 148593 106072
rect 143904 106014 148532 106070
rect 148588 106014 148593 106070
rect 143904 106012 148593 106014
rect 640416 106070 645777 106072
rect 640416 106014 645716 106070
rect 645772 106014 645777 106070
rect 640416 106012 645777 106014
rect 148527 106009 148593 106012
rect 645711 106009 645777 106012
rect 184527 105628 184593 105631
rect 184527 105626 190560 105628
rect 184527 105570 184532 105626
rect 184588 105570 190560 105626
rect 184527 105568 190560 105570
rect 184527 105565 184593 105568
rect 665346 105184 665406 105361
rect 668367 105184 668433 105187
rect 665346 105182 668433 105184
rect 665346 105126 668372 105182
rect 668428 105126 668433 105182
rect 665346 105124 668433 105126
rect 668367 105121 668433 105124
rect 674554 105122 674560 105186
rect 674624 105184 674630 105186
rect 675375 105184 675441 105187
rect 674624 105182 675441 105184
rect 674624 105126 675380 105182
rect 675436 105126 675441 105182
rect 674624 105124 675441 105126
rect 674624 105122 674630 105124
rect 675375 105121 675441 105124
rect 665346 104891 665406 104996
rect 184431 104888 184497 104891
rect 184431 104886 190014 104888
rect 184431 104830 184436 104886
rect 184492 104830 190014 104886
rect 184431 104828 190014 104830
rect 184431 104825 184497 104828
rect 189954 104814 190014 104828
rect 665295 104886 665406 104891
rect 665295 104830 665300 104886
rect 665356 104830 665406 104886
rect 665295 104828 665406 104830
rect 665295 104825 665361 104828
rect 189954 104754 190560 104814
rect 148335 104740 148401 104743
rect 143904 104738 148401 104740
rect 143904 104682 148340 104738
rect 148396 104682 148401 104738
rect 143904 104680 148401 104682
rect 148335 104677 148401 104680
rect 647919 104148 647985 104151
rect 640416 104146 647985 104148
rect 640416 104090 647924 104146
rect 647980 104090 647985 104146
rect 640416 104088 647985 104090
rect 647919 104085 647985 104088
rect 184623 104000 184689 104003
rect 184623 103998 190560 104000
rect 184623 103942 184628 103998
rect 184684 103942 190560 103998
rect 184623 103940 190560 103942
rect 184623 103937 184689 103940
rect 149583 103556 149649 103559
rect 143904 103554 149649 103556
rect 143904 103498 149588 103554
rect 149644 103498 149649 103554
rect 143904 103496 149649 103498
rect 149583 103493 149649 103496
rect 184335 103408 184401 103411
rect 184335 103406 190014 103408
rect 184335 103350 184340 103406
rect 184396 103350 190014 103406
rect 184335 103348 190014 103350
rect 184335 103345 184401 103348
rect 189954 103334 190014 103348
rect 189954 103274 190560 103334
rect 675759 103260 675825 103263
rect 675898 103260 675904 103262
rect 675759 103258 675904 103260
rect 675759 103202 675764 103258
rect 675820 103202 675904 103258
rect 675759 103200 675904 103202
rect 675759 103197 675825 103200
rect 675898 103198 675904 103200
rect 675968 103198 675974 103262
rect 184431 102520 184497 102523
rect 184431 102518 190560 102520
rect 184431 102462 184436 102518
rect 184492 102462 190560 102518
rect 184431 102460 190560 102462
rect 184431 102457 184497 102460
rect 148623 102372 148689 102375
rect 143904 102370 148689 102372
rect 143904 102314 148628 102370
rect 148684 102314 148689 102370
rect 143904 102312 148689 102314
rect 148623 102309 148689 102312
rect 645135 102224 645201 102227
rect 640416 102222 645201 102224
rect 640416 102166 645140 102222
rect 645196 102166 645201 102222
rect 640416 102164 645201 102166
rect 645135 102161 645201 102164
rect 184719 101928 184785 101931
rect 184719 101926 190014 101928
rect 184719 101870 184724 101926
rect 184780 101870 190014 101926
rect 184719 101868 190014 101870
rect 184719 101865 184785 101868
rect 189954 101854 190014 101868
rect 189954 101794 190560 101854
rect 675759 101484 675825 101487
rect 676474 101484 676480 101486
rect 675759 101482 676480 101484
rect 675759 101426 675764 101482
rect 675820 101426 676480 101482
rect 675759 101424 676480 101426
rect 675759 101421 675825 101424
rect 676474 101422 676480 101424
rect 676544 101422 676550 101486
rect 143874 100892 143934 101084
rect 184527 101040 184593 101043
rect 184527 101038 190560 101040
rect 184527 100982 184532 101038
rect 184588 100982 190560 101038
rect 184527 100980 190560 100982
rect 184527 100977 184593 100980
rect 149391 100892 149457 100895
rect 143874 100890 149457 100892
rect 143874 100834 149396 100890
rect 149452 100834 149457 100890
rect 143874 100832 149457 100834
rect 149391 100829 149457 100832
rect 184335 100300 184401 100303
rect 184335 100298 190014 100300
rect 184335 100242 184340 100298
rect 184396 100242 190014 100298
rect 184335 100240 190014 100242
rect 184335 100237 184401 100240
rect 189954 100226 190014 100240
rect 189954 100166 190560 100226
rect 149487 99856 149553 99859
rect 143904 99854 149553 99856
rect 143904 99798 149492 99854
rect 149548 99798 149553 99854
rect 143904 99796 149553 99798
rect 149487 99793 149553 99796
rect 640194 99708 640254 100270
rect 647919 99708 647985 99711
rect 640194 99706 647985 99708
rect 640194 99650 647924 99706
rect 647980 99650 647985 99706
rect 640194 99648 647985 99650
rect 647919 99645 647985 99648
rect 184431 99560 184497 99563
rect 184431 99558 190560 99560
rect 184431 99502 184436 99558
rect 184492 99502 190560 99558
rect 184431 99500 190560 99502
rect 184431 99497 184497 99500
rect 149391 98672 149457 98675
rect 143904 98670 149457 98672
rect 143904 98614 149396 98670
rect 149452 98614 149457 98670
rect 143904 98612 149457 98614
rect 149391 98609 149457 98612
rect 184527 98672 184593 98675
rect 184527 98670 190560 98672
rect 184527 98614 184532 98670
rect 184588 98614 190560 98670
rect 184527 98612 190560 98614
rect 184527 98609 184593 98612
rect 184623 98080 184689 98083
rect 640386 98080 640446 98420
rect 646959 98080 647025 98083
rect 184623 98078 190560 98080
rect 184623 98022 184628 98078
rect 184684 98022 190560 98078
rect 184623 98020 190560 98022
rect 640386 98078 647025 98080
rect 640386 98022 646964 98078
rect 647020 98022 647025 98078
rect 640386 98020 647025 98022
rect 184623 98017 184689 98020
rect 646959 98017 647025 98020
rect 149487 97488 149553 97491
rect 143904 97486 149553 97488
rect 143904 97430 149492 97486
rect 149548 97430 149553 97486
rect 143904 97428 149553 97430
rect 149487 97425 149553 97428
rect 184335 97192 184401 97195
rect 184335 97190 190560 97192
rect 184335 97134 184340 97190
rect 184396 97134 190560 97190
rect 184335 97132 190560 97134
rect 184335 97129 184401 97132
rect 184431 96452 184497 96455
rect 184431 96450 190560 96452
rect 184431 96394 184436 96450
rect 184492 96394 190560 96450
rect 184431 96392 190560 96394
rect 184431 96389 184497 96392
rect 143874 95712 143934 96200
rect 640386 96008 640446 96570
rect 645423 96008 645489 96011
rect 640386 96006 645489 96008
rect 640386 95950 645428 96006
rect 645484 95950 645489 96006
rect 640386 95948 645489 95950
rect 645423 95945 645489 95948
rect 149391 95712 149457 95715
rect 143874 95710 149457 95712
rect 143874 95654 149396 95710
rect 149452 95654 149457 95710
rect 143874 95652 149457 95654
rect 149391 95649 149457 95652
rect 184527 95712 184593 95715
rect 184527 95710 190560 95712
rect 184527 95654 184532 95710
rect 184588 95654 190560 95710
rect 184527 95652 190560 95654
rect 184527 95649 184593 95652
rect 149679 94972 149745 94975
rect 143904 94970 149745 94972
rect 143904 94914 149684 94970
rect 149740 94914 149745 94970
rect 143904 94912 149745 94914
rect 149679 94909 149745 94912
rect 184335 94972 184401 94975
rect 184335 94970 190014 94972
rect 184335 94914 184340 94970
rect 184396 94914 190014 94970
rect 184335 94912 190014 94914
rect 184335 94909 184401 94912
rect 189954 94898 190014 94912
rect 189954 94838 190560 94898
rect 186255 94232 186321 94235
rect 186255 94230 190560 94232
rect 186255 94174 186260 94230
rect 186316 94174 190560 94230
rect 186255 94172 190560 94174
rect 186255 94169 186321 94172
rect 640386 94084 640446 94646
rect 647727 94084 647793 94087
rect 640386 94082 647793 94084
rect 640386 94026 647732 94082
rect 647788 94026 647793 94082
rect 640386 94024 647793 94026
rect 647727 94021 647793 94024
rect 149487 93788 149553 93791
rect 143904 93786 149553 93788
rect 143904 93730 149492 93786
rect 149548 93730 149553 93786
rect 143904 93728 149553 93730
rect 149487 93725 149553 93728
rect 184335 93492 184401 93495
rect 184335 93490 190014 93492
rect 184335 93434 184340 93490
rect 184396 93434 190014 93490
rect 184335 93432 190014 93434
rect 184335 93429 184401 93432
rect 189954 93418 190014 93432
rect 189954 93358 190560 93418
rect 184623 92752 184689 92755
rect 647823 92752 647889 92755
rect 184623 92750 190560 92752
rect 184623 92694 184628 92750
rect 184684 92694 190560 92750
rect 184623 92692 190560 92694
rect 640416 92750 647889 92752
rect 640416 92694 647828 92750
rect 647884 92694 647889 92750
rect 640416 92692 647889 92694
rect 184623 92689 184689 92692
rect 647823 92689 647889 92692
rect 149391 92604 149457 92607
rect 143904 92602 149457 92604
rect 143904 92546 149396 92602
rect 149452 92546 149457 92602
rect 143904 92544 149457 92546
rect 149391 92541 149457 92544
rect 189954 91878 190560 91938
rect 184335 91864 184401 91867
rect 189954 91864 190014 91878
rect 184335 91862 190014 91864
rect 184335 91806 184340 91862
rect 184396 91806 190014 91862
rect 184335 91804 190014 91806
rect 184335 91801 184401 91804
rect 149199 91420 149265 91423
rect 143904 91418 149265 91420
rect 143904 91362 149204 91418
rect 149260 91362 149265 91418
rect 143904 91360 149265 91362
rect 149199 91357 149265 91360
rect 184431 91124 184497 91127
rect 184431 91122 190560 91124
rect 184431 91066 184436 91122
rect 184492 91066 190560 91122
rect 184431 91064 190560 91066
rect 184431 91061 184497 91064
rect 659343 90828 659409 90831
rect 640416 90826 659409 90828
rect 640416 90770 659348 90826
rect 659404 90770 659409 90826
rect 640416 90768 659409 90770
rect 659343 90765 659409 90768
rect 184527 90384 184593 90387
rect 184527 90382 190560 90384
rect 184527 90326 184532 90382
rect 184588 90326 190560 90382
rect 184527 90324 190560 90326
rect 184527 90321 184593 90324
rect 149295 90236 149361 90239
rect 143904 90234 149361 90236
rect 143904 90178 149300 90234
rect 149356 90178 149361 90234
rect 143904 90176 149361 90178
rect 149295 90173 149361 90176
rect 184623 89644 184689 89647
rect 184623 89642 190560 89644
rect 184623 89586 184628 89642
rect 184684 89586 190560 89642
rect 184623 89584 190560 89586
rect 184623 89581 184689 89584
rect 149391 89052 149457 89055
rect 143904 89050 149457 89052
rect 143904 88994 149396 89050
rect 149452 88994 149457 89050
rect 143904 88992 149457 88994
rect 149391 88989 149457 88992
rect 184335 88904 184401 88907
rect 645903 88904 645969 88907
rect 184335 88902 190560 88904
rect 184335 88846 184340 88902
rect 184396 88846 190560 88902
rect 184335 88844 190560 88846
rect 640416 88902 645969 88904
rect 640416 88846 645908 88902
rect 645964 88846 645969 88902
rect 640416 88844 645969 88846
rect 184335 88841 184401 88844
rect 645903 88841 645969 88844
rect 184431 88164 184497 88167
rect 184431 88162 190014 88164
rect 184431 88106 184436 88162
rect 184492 88106 190014 88162
rect 184431 88104 190014 88106
rect 184431 88101 184497 88104
rect 189954 88090 190014 88104
rect 189954 88030 190560 88090
rect 143874 87424 143934 87764
rect 149487 87424 149553 87427
rect 143874 87422 149553 87424
rect 143874 87366 149492 87422
rect 149548 87366 149553 87422
rect 143874 87364 149553 87366
rect 149487 87361 149553 87364
rect 184527 87276 184593 87279
rect 184527 87274 190560 87276
rect 184527 87218 184532 87274
rect 184588 87218 190560 87274
rect 184527 87216 190560 87218
rect 184527 87213 184593 87216
rect 647919 87128 647985 87131
rect 640386 87126 647985 87128
rect 640386 87070 647924 87126
rect 647980 87070 647985 87126
rect 640386 87068 647985 87070
rect 640386 86950 640446 87068
rect 647919 87065 647985 87068
rect 653679 86980 653745 86983
rect 653679 86978 656736 86980
rect 653679 86922 653684 86978
rect 653740 86922 656736 86978
rect 653679 86920 656736 86922
rect 653679 86917 653745 86920
rect 184623 86684 184689 86687
rect 184623 86682 190014 86684
rect 184623 86626 184628 86682
rect 184684 86626 190014 86682
rect 184623 86624 190014 86626
rect 184623 86621 184689 86624
rect 189954 86610 190014 86624
rect 189954 86550 190560 86610
rect 148719 86536 148785 86539
rect 143904 86534 148785 86536
rect 143904 86478 148724 86534
rect 148780 86478 148785 86534
rect 143904 86476 148785 86478
rect 148719 86473 148785 86476
rect 663279 86388 663345 86391
rect 663234 86386 663345 86388
rect 663234 86330 663284 86386
rect 663340 86330 663345 86386
rect 663234 86325 663345 86330
rect 650895 86240 650961 86243
rect 650895 86238 656736 86240
rect 650895 86182 650900 86238
rect 650956 86182 656736 86238
rect 663234 86210 663294 86325
rect 650895 86180 656736 86182
rect 650895 86177 650961 86180
rect 184431 85796 184497 85799
rect 184431 85794 190560 85796
rect 184431 85738 184436 85794
rect 184492 85738 190560 85794
rect 184431 85736 190560 85738
rect 184431 85733 184497 85736
rect 148431 85352 148497 85355
rect 143904 85350 148497 85352
rect 143904 85294 148436 85350
rect 148492 85294 148497 85350
rect 143904 85292 148497 85294
rect 148431 85289 148497 85292
rect 652335 85352 652401 85355
rect 652335 85350 656736 85352
rect 652335 85294 652340 85350
rect 652396 85294 656736 85350
rect 652335 85292 656736 85294
rect 652335 85289 652401 85292
rect 184335 85204 184401 85207
rect 184335 85202 190014 85204
rect 184335 85146 184340 85202
rect 184396 85146 190014 85202
rect 184335 85144 190014 85146
rect 184335 85141 184401 85144
rect 189954 85130 190014 85144
rect 189954 85070 190560 85130
rect 640194 84464 640254 85026
rect 663234 84763 663294 85322
rect 663234 84758 663345 84763
rect 663234 84702 663284 84758
rect 663340 84702 663345 84758
rect 663234 84700 663345 84702
rect 663279 84697 663345 84700
rect 645903 84464 645969 84467
rect 640194 84462 645969 84464
rect 640194 84406 645908 84462
rect 645964 84406 645969 84462
rect 640194 84404 645969 84406
rect 645903 84401 645969 84404
rect 184527 84316 184593 84319
rect 651759 84316 651825 84319
rect 184527 84314 190560 84316
rect 184527 84258 184532 84314
rect 184588 84258 190560 84314
rect 184527 84256 190560 84258
rect 651759 84314 656736 84316
rect 651759 84258 651764 84314
rect 651820 84258 656736 84314
rect 651759 84256 656736 84258
rect 184527 84253 184593 84256
rect 651759 84253 651825 84256
rect 147087 84168 147153 84171
rect 143904 84166 147153 84168
rect 143904 84110 147092 84166
rect 147148 84110 147153 84166
rect 143904 84108 147153 84110
rect 147087 84105 147153 84108
rect 663426 84023 663486 84582
rect 663426 84018 663537 84023
rect 663426 83962 663476 84018
rect 663532 83962 663537 84018
rect 663426 83960 663537 83962
rect 663471 83957 663537 83960
rect 189954 83442 190560 83502
rect 184335 83428 184401 83431
rect 189954 83428 190014 83442
rect 184335 83426 190014 83428
rect 184335 83370 184340 83426
rect 184396 83370 190014 83426
rect 184335 83368 190014 83370
rect 652239 83428 652305 83431
rect 652239 83426 656736 83428
rect 652239 83370 652244 83426
rect 652300 83370 656736 83426
rect 652239 83368 656736 83370
rect 184335 83365 184401 83368
rect 652239 83365 652305 83368
rect 143874 82392 143934 82880
rect 186159 82836 186225 82839
rect 186159 82834 190560 82836
rect 186159 82778 186164 82834
rect 186220 82778 190560 82834
rect 186159 82776 190560 82778
rect 186159 82773 186225 82776
rect 640386 82688 640446 83176
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 647919 82688 647985 82691
rect 640386 82686 647985 82688
rect 640386 82630 647924 82686
rect 647980 82630 647985 82686
rect 640386 82628 647985 82630
rect 647919 82625 647985 82628
rect 652431 82688 652497 82691
rect 652431 82686 656736 82688
rect 652431 82630 652436 82686
rect 652492 82630 656736 82686
rect 652431 82628 656736 82630
rect 652431 82625 652497 82628
rect 149103 82392 149169 82395
rect 143874 82390 149169 82392
rect 143874 82334 149108 82390
rect 149164 82334 149169 82390
rect 143874 82332 149169 82334
rect 149103 82329 149169 82332
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 184239 81948 184305 81951
rect 184239 81946 190560 81948
rect 184239 81890 184244 81946
rect 184300 81890 190560 81946
rect 184239 81888 190560 81890
rect 184239 81885 184305 81888
rect 148239 81652 148305 81655
rect 143904 81650 148305 81652
rect 143904 81594 148244 81650
rect 148300 81594 148305 81650
rect 143904 81592 148305 81594
rect 148239 81589 148305 81592
rect 662415 81652 662481 81655
rect 663042 81652 663102 81770
rect 662415 81650 663102 81652
rect 662415 81594 662420 81650
rect 662476 81594 663102 81650
rect 662415 81592 663102 81594
rect 662415 81589 662481 81592
rect 184431 81356 184497 81359
rect 184431 81354 190560 81356
rect 184431 81298 184436 81354
rect 184492 81298 190560 81354
rect 184431 81296 190560 81298
rect 184431 81293 184497 81296
rect 640386 81060 640446 81326
rect 647919 81060 647985 81063
rect 640386 81058 647985 81060
rect 640386 81002 647924 81058
rect 647980 81002 647985 81058
rect 640386 81000 647985 81002
rect 647919 80997 647985 81000
rect 149583 80468 149649 80471
rect 143904 80466 149649 80468
rect 143904 80410 149588 80466
rect 149644 80410 149649 80466
rect 143904 80408 149649 80410
rect 149583 80405 149649 80408
rect 184623 80468 184689 80471
rect 184623 80466 190560 80468
rect 184623 80410 184628 80466
rect 184684 80410 190560 80466
rect 184623 80408 190560 80410
rect 184623 80405 184689 80408
rect 184431 79876 184497 79879
rect 184431 79874 190014 79876
rect 184431 79818 184436 79874
rect 184492 79818 190014 79874
rect 184431 79816 190014 79818
rect 184431 79813 184497 79816
rect 189954 79802 190014 79816
rect 189954 79742 190560 79802
rect 645519 79432 645585 79435
rect 640416 79430 645585 79432
rect 640416 79374 645524 79430
rect 645580 79374 645585 79430
rect 640416 79372 645585 79374
rect 645519 79369 645585 79372
rect 149679 79284 149745 79287
rect 143904 79282 149745 79284
rect 143904 79226 149684 79282
rect 149740 79226 149745 79282
rect 143904 79224 149745 79226
rect 149679 79221 149745 79224
rect 184335 78988 184401 78991
rect 184335 78986 190560 78988
rect 184335 78930 184340 78986
rect 184396 78930 190560 78986
rect 184335 78928 190560 78930
rect 184335 78925 184401 78928
rect 184527 78248 184593 78251
rect 184527 78246 190014 78248
rect 184527 78190 184532 78246
rect 184588 78190 190014 78246
rect 184527 78188 190014 78190
rect 184527 78185 184593 78188
rect 189954 78174 190014 78188
rect 189954 78114 190560 78174
rect 148815 77952 148881 77955
rect 143904 77950 148881 77952
rect 143904 77894 148820 77950
rect 148876 77894 148881 77950
rect 143904 77892 148881 77894
rect 148815 77889 148881 77892
rect 184335 77508 184401 77511
rect 647919 77508 647985 77511
rect 184335 77506 190560 77508
rect 184335 77450 184340 77506
rect 184396 77450 190560 77506
rect 184335 77448 190560 77450
rect 640416 77506 647985 77508
rect 640416 77450 647924 77506
rect 647980 77450 647985 77506
rect 640416 77448 647985 77450
rect 184335 77445 184401 77448
rect 647919 77445 647985 77448
rect 149199 76768 149265 76771
rect 143904 76766 149265 76768
rect 143904 76710 149204 76766
rect 149260 76710 149265 76766
rect 143904 76708 149265 76710
rect 149199 76705 149265 76708
rect 184431 76768 184497 76771
rect 184431 76766 190014 76768
rect 184431 76710 184436 76766
rect 184492 76710 190014 76766
rect 184431 76708 190014 76710
rect 184431 76705 184497 76708
rect 189954 76694 190014 76708
rect 189954 76634 190560 76694
rect 184527 76028 184593 76031
rect 184527 76026 190560 76028
rect 184527 75970 184532 76026
rect 184588 75970 190560 76026
rect 184527 75968 190560 75970
rect 184527 75965 184593 75968
rect 149391 75584 149457 75587
rect 645999 75584 646065 75587
rect 143904 75582 149457 75584
rect 143904 75526 149396 75582
rect 149452 75526 149457 75582
rect 143904 75524 149457 75526
rect 640416 75582 646065 75584
rect 640416 75526 646004 75582
rect 646060 75526 646065 75582
rect 640416 75524 646065 75526
rect 149391 75521 149457 75524
rect 645999 75521 646065 75524
rect 184623 75140 184689 75143
rect 184623 75138 190560 75140
rect 184623 75082 184628 75138
rect 184684 75082 190560 75138
rect 184623 75080 190560 75082
rect 184623 75077 184689 75080
rect 184335 74400 184401 74403
rect 184335 74398 190560 74400
rect 184335 74342 184340 74398
rect 184396 74342 190560 74398
rect 184335 74340 190560 74342
rect 184335 74337 184401 74340
rect 143874 73808 143934 74296
rect 149295 73808 149361 73811
rect 143874 73806 149361 73808
rect 143874 73750 149300 73806
rect 149356 73750 149361 73806
rect 143874 73748 149361 73750
rect 149295 73745 149361 73748
rect 184527 73660 184593 73663
rect 647919 73660 647985 73663
rect 184527 73658 190560 73660
rect 184527 73602 184532 73658
rect 184588 73602 190560 73658
rect 184527 73600 190560 73602
rect 640416 73658 647985 73660
rect 640416 73602 647924 73658
rect 647980 73602 647985 73658
rect 640416 73600 647985 73602
rect 184527 73597 184593 73600
rect 647919 73597 647985 73600
rect 149007 73068 149073 73071
rect 143904 73066 149073 73068
rect 143904 73010 149012 73066
rect 149068 73010 149073 73066
rect 143904 73008 149073 73010
rect 149007 73005 149073 73008
rect 184431 72920 184497 72923
rect 184431 72918 190560 72920
rect 184431 72862 184436 72918
rect 184492 72862 190560 72918
rect 184431 72860 190560 72862
rect 184431 72857 184497 72860
rect 184623 72180 184689 72183
rect 184623 72178 190560 72180
rect 184623 72122 184628 72178
rect 184684 72122 190560 72178
rect 184623 72120 190560 72122
rect 184623 72117 184689 72120
rect 149103 72032 149169 72035
rect 143904 72030 149169 72032
rect 143904 71974 149108 72030
rect 149164 71974 149169 72030
rect 143904 71972 149169 71974
rect 149103 71969 149169 71972
rect 647151 71884 647217 71887
rect 640386 71882 647217 71884
rect 640386 71826 647156 71882
rect 647212 71826 647217 71882
rect 640386 71824 647217 71826
rect 640386 71706 640446 71824
rect 647151 71821 647217 71824
rect 184431 71440 184497 71443
rect 184431 71438 190014 71440
rect 184431 71382 184436 71438
rect 184492 71382 190014 71438
rect 184431 71380 190014 71382
rect 184431 71377 184497 71380
rect 189954 71366 190014 71380
rect 189954 71306 190560 71366
rect 149487 70848 149553 70851
rect 143904 70846 149553 70848
rect 143904 70790 149492 70846
rect 149548 70790 149553 70846
rect 143904 70788 149553 70790
rect 149487 70785 149553 70788
rect 184335 70552 184401 70555
rect 184335 70550 190560 70552
rect 184335 70494 184340 70550
rect 184396 70494 190560 70550
rect 184335 70492 190560 70494
rect 184335 70489 184401 70492
rect 184527 69960 184593 69963
rect 184527 69958 190014 69960
rect 184527 69902 184532 69958
rect 184588 69902 190014 69958
rect 184527 69900 190014 69902
rect 184527 69897 184593 69900
rect 189954 69886 190014 69900
rect 189954 69826 190560 69886
rect 640386 69664 640446 69856
rect 647919 69664 647985 69667
rect 640386 69662 647985 69664
rect 640386 69606 647924 69662
rect 647980 69606 647985 69662
rect 640386 69604 647985 69606
rect 647919 69601 647985 69604
rect 149391 69516 149457 69519
rect 143904 69514 149457 69516
rect 143904 69458 149396 69514
rect 149452 69458 149457 69514
rect 143904 69456 149457 69458
rect 149391 69453 149457 69456
rect 184335 69072 184401 69075
rect 184335 69070 190560 69072
rect 184335 69014 184340 69070
rect 184396 69014 190560 69070
rect 184335 69012 190560 69014
rect 184335 69009 184401 69012
rect 646863 68628 646929 68631
rect 640194 68626 646929 68628
rect 640194 68570 646868 68626
rect 646924 68570 646929 68626
rect 640194 68568 646929 68570
rect 184431 68480 184497 68483
rect 184431 68478 190014 68480
rect 184431 68422 184436 68478
rect 184492 68422 190014 68478
rect 184431 68420 190014 68422
rect 184431 68417 184497 68420
rect 189954 68406 190014 68420
rect 189954 68346 190560 68406
rect 149199 68332 149265 68335
rect 143904 68330 149265 68332
rect 143904 68274 149204 68330
rect 149260 68274 149265 68330
rect 143904 68272 149265 68274
rect 149199 68269 149265 68272
rect 640194 68006 640254 68568
rect 646863 68565 646929 68568
rect 184335 67592 184401 67595
rect 184335 67590 190560 67592
rect 184335 67534 184340 67590
rect 184396 67534 190560 67590
rect 184335 67532 190560 67534
rect 184335 67529 184401 67532
rect 149583 67148 149649 67151
rect 143904 67146 149649 67148
rect 143904 67090 149588 67146
rect 149644 67090 149649 67146
rect 143904 67088 149649 67090
rect 149583 67085 149649 67088
rect 184527 66852 184593 66855
rect 184527 66850 190560 66852
rect 184527 66794 184532 66850
rect 184588 66794 190560 66850
rect 184527 66792 190560 66794
rect 184527 66789 184593 66792
rect 645999 66260 646065 66263
rect 640194 66258 646065 66260
rect 640194 66202 646004 66258
rect 646060 66202 646065 66258
rect 640194 66200 646065 66202
rect 184335 66112 184401 66115
rect 184335 66110 190560 66112
rect 184335 66054 184340 66110
rect 184396 66054 190560 66110
rect 640194 66082 640254 66200
rect 645999 66197 646065 66200
rect 184335 66052 190560 66054
rect 184335 66049 184401 66052
rect 143874 65372 143934 65860
rect 149295 65372 149361 65375
rect 143874 65370 149361 65372
rect 143874 65314 149300 65370
rect 149356 65314 149361 65370
rect 143874 65312 149361 65314
rect 149295 65309 149361 65312
rect 184527 65224 184593 65227
rect 184527 65222 190560 65224
rect 184527 65166 184532 65222
rect 184588 65166 190560 65222
rect 184527 65164 190560 65166
rect 184527 65161 184593 65164
rect 149391 64632 149457 64635
rect 143904 64630 149457 64632
rect 143904 64574 149396 64630
rect 149452 64574 149457 64630
rect 143904 64572 149457 64574
rect 149391 64569 149457 64572
rect 184431 64632 184497 64635
rect 184431 64630 190014 64632
rect 184431 64574 184436 64630
rect 184492 64574 190014 64630
rect 184431 64572 190014 64574
rect 184431 64569 184497 64572
rect 189954 64558 190014 64572
rect 189954 64498 190560 64558
rect 647919 64188 647985 64191
rect 640416 64186 647985 64188
rect 640416 64130 647924 64186
rect 647980 64130 647985 64186
rect 640416 64128 647985 64130
rect 647919 64125 647985 64128
rect 184623 63744 184689 63747
rect 184623 63742 190560 63744
rect 184623 63686 184628 63742
rect 184684 63686 190560 63742
rect 184623 63684 190560 63686
rect 184623 63681 184689 63684
rect 149487 63448 149553 63451
rect 143904 63446 149553 63448
rect 143904 63390 149492 63446
rect 149548 63390 149553 63446
rect 143904 63388 149553 63390
rect 149487 63385 149553 63388
rect 184335 63152 184401 63155
rect 184335 63150 190014 63152
rect 184335 63094 184340 63150
rect 184396 63094 190014 63150
rect 184335 63092 190014 63094
rect 184335 63089 184401 63092
rect 189954 63078 190014 63092
rect 189954 63018 190560 63078
rect 149391 62264 149457 62267
rect 143904 62262 149457 62264
rect 143904 62206 149396 62262
rect 149452 62206 149457 62262
rect 143904 62204 149457 62206
rect 149391 62201 149457 62204
rect 184527 62264 184593 62267
rect 647919 62264 647985 62267
rect 184527 62262 190560 62264
rect 184527 62206 184532 62262
rect 184588 62206 190560 62262
rect 184527 62204 190560 62206
rect 640416 62262 647985 62264
rect 640416 62206 647924 62262
rect 647980 62206 647985 62262
rect 640416 62204 647985 62206
rect 184527 62201 184593 62204
rect 647919 62201 647985 62204
rect 184431 61524 184497 61527
rect 184431 61522 190014 61524
rect 184431 61466 184436 61522
rect 184492 61466 190014 61522
rect 184431 61464 190014 61466
rect 184431 61461 184497 61464
rect 189954 61450 190014 61464
rect 189954 61390 190560 61450
rect 143874 60636 143934 60976
rect 184623 60784 184689 60787
rect 184623 60782 190560 60784
rect 184623 60726 184628 60782
rect 184684 60726 190560 60782
rect 184623 60724 190560 60726
rect 184623 60721 184689 60724
rect 149295 60636 149361 60639
rect 143874 60634 149361 60636
rect 143874 60578 149300 60634
rect 149356 60578 149361 60634
rect 143874 60576 149361 60578
rect 149295 60573 149361 60576
rect 647055 60340 647121 60343
rect 640416 60338 647121 60340
rect 640416 60282 647060 60338
rect 647116 60282 647121 60338
rect 640416 60280 647121 60282
rect 647055 60277 647121 60280
rect 184335 60044 184401 60047
rect 184335 60042 190014 60044
rect 184335 59986 184340 60042
rect 184396 59986 190014 60042
rect 184335 59984 190014 59986
rect 184335 59981 184401 59984
rect 189954 59970 190014 59984
rect 189954 59910 190560 59970
rect 149391 59748 149457 59751
rect 143904 59746 149457 59748
rect 143904 59690 149396 59746
rect 149452 59690 149457 59746
rect 143904 59688 149457 59690
rect 149391 59685 149457 59688
rect 184431 59304 184497 59307
rect 184431 59302 190560 59304
rect 184431 59246 184436 59302
rect 184492 59246 190560 59302
rect 184431 59244 190560 59246
rect 184431 59241 184497 59244
rect 645999 59008 646065 59011
rect 640386 59006 646065 59008
rect 640386 58950 646004 59006
rect 646060 58950 646065 59006
rect 640386 58948 646065 58950
rect 149391 58564 149457 58567
rect 143904 58562 149457 58564
rect 143904 58506 149396 58562
rect 149452 58506 149457 58562
rect 143904 58504 149457 58506
rect 149391 58501 149457 58504
rect 184527 58416 184593 58419
rect 184527 58414 190560 58416
rect 184527 58358 184532 58414
rect 184588 58358 190560 58414
rect 640386 58386 640446 58948
rect 645999 58945 646065 58948
rect 184527 58356 190560 58358
rect 184527 58353 184593 58356
rect 184335 57676 184401 57679
rect 184335 57674 190560 57676
rect 184335 57618 184340 57674
rect 184396 57618 190560 57674
rect 184335 57616 190560 57618
rect 184335 57613 184401 57616
rect 149487 57380 149553 57383
rect 143904 57378 149553 57380
rect 143904 57322 149492 57378
rect 149548 57322 149553 57378
rect 143904 57320 149553 57322
rect 149487 57317 149553 57320
rect 646767 57084 646833 57087
rect 640386 57082 646833 57084
rect 640386 57026 646772 57082
rect 646828 57026 646833 57082
rect 640386 57024 646833 57026
rect 184335 56936 184401 56939
rect 184335 56934 190560 56936
rect 184335 56878 184340 56934
rect 184396 56878 190560 56934
rect 184335 56876 190560 56878
rect 184335 56873 184401 56876
rect 640386 56536 640446 57024
rect 646767 57021 646833 57024
rect 149391 56196 149457 56199
rect 143874 56194 149457 56196
rect 143874 56138 149396 56194
rect 149452 56138 149457 56194
rect 143874 56136 149457 56138
rect 143874 56092 143934 56136
rect 149391 56133 149457 56136
rect 184335 56196 184401 56199
rect 184335 56194 190560 56196
rect 184335 56138 184340 56194
rect 184396 56138 190560 56194
rect 184335 56136 190560 56138
rect 184335 56133 184401 56136
rect 184431 55456 184497 55459
rect 184431 55454 190560 55456
rect 184431 55398 184436 55454
rect 184492 55398 190560 55454
rect 184431 55396 190560 55398
rect 184431 55393 184497 55396
rect 149679 54864 149745 54867
rect 143904 54862 149745 54864
rect 143904 54806 149684 54862
rect 149740 54806 149745 54862
rect 143904 54804 149745 54806
rect 149679 54801 149745 54804
rect 184335 54716 184401 54719
rect 646479 54716 646545 54719
rect 184335 54714 190014 54716
rect 184335 54658 184340 54714
rect 184396 54658 190014 54714
rect 184335 54656 190014 54658
rect 184335 54653 184401 54656
rect 189954 54642 190014 54656
rect 640386 54714 646545 54716
rect 640386 54658 646484 54714
rect 646540 54658 646545 54714
rect 640386 54656 646545 54658
rect 189954 54582 190560 54642
rect 640386 54612 640446 54656
rect 646479 54653 646545 54656
rect 184335 53976 184401 53979
rect 184335 53974 190560 53976
rect 184335 53918 184340 53974
rect 184396 53918 190560 53974
rect 184335 53916 190560 53918
rect 184335 53913 184401 53916
rect 149391 53828 149457 53831
rect 143904 53826 149457 53828
rect 143904 53770 149396 53826
rect 149452 53770 149457 53826
rect 143904 53768 149457 53770
rect 149391 53765 149457 53768
rect 426159 44948 426225 44951
rect 472239 44948 472305 44951
rect 419394 44946 426225 44948
rect 419394 44890 426164 44946
rect 426220 44890 426225 44946
rect 419394 44888 426225 44890
rect 419394 44404 419454 44888
rect 426159 44885 426225 44888
rect 472194 44946 472305 44948
rect 472194 44890 472244 44946
rect 472300 44890 472305 44946
rect 472194 44885 472305 44890
rect 472194 44404 472254 44885
rect 517359 42136 517425 42139
rect 520335 42136 520401 42139
rect 517359 42134 520401 42136
rect 517359 42078 517364 42134
rect 517420 42078 520340 42134
rect 520396 42078 520401 42134
rect 517359 42076 520401 42078
rect 517359 42073 517425 42076
rect 520335 42073 520401 42076
rect 187599 41988 187665 41991
rect 216399 41988 216465 41991
rect 187599 41986 216465 41988
rect 187599 41930 187604 41986
rect 187660 41930 216404 41986
rect 216460 41930 216465 41986
rect 187599 41928 216465 41930
rect 187599 41925 187665 41928
rect 216399 41925 216465 41928
rect 415215 41988 415281 41991
rect 434895 41988 434961 41991
rect 415215 41986 434961 41988
rect 415215 41930 415220 41986
rect 415276 41930 434900 41986
rect 434956 41930 434961 41986
rect 415215 41928 434961 41930
rect 415215 41925 415281 41928
rect 434895 41925 434961 41928
rect 194319 41840 194385 41843
rect 302895 41840 302961 41843
rect 357711 41840 357777 41843
rect 394575 41840 394641 41843
rect 194319 41838 195870 41840
rect 194319 41782 194324 41838
rect 194380 41782 195870 41838
rect 194319 41780 195870 41782
rect 194319 41777 194385 41780
rect 195810 40508 195870 41780
rect 302895 41838 316830 41840
rect 302895 41782 302900 41838
rect 302956 41782 316830 41838
rect 302895 41780 316830 41782
rect 302895 41777 302961 41780
rect 224559 40508 224625 40511
rect 195810 40506 224625 40508
rect 195810 40450 224564 40506
rect 224620 40450 224625 40506
rect 195810 40448 224625 40450
rect 316770 40508 316830 41780
rect 357711 41838 394641 41840
rect 357711 41782 357716 41838
rect 357772 41782 394580 41838
rect 394636 41782 394641 41838
rect 357711 41780 394641 41782
rect 357711 41777 357777 41780
rect 394575 41777 394641 41780
rect 416847 41840 416913 41843
rect 470319 41840 470385 41843
rect 471663 41840 471729 41843
rect 416847 41838 417630 41840
rect 416847 41782 416852 41838
rect 416908 41782 417630 41838
rect 416847 41780 417630 41782
rect 416847 41777 416913 41780
rect 345615 40508 345681 40511
rect 316770 40506 345681 40508
rect 316770 40450 345620 40506
rect 345676 40450 345681 40506
rect 316770 40448 345681 40450
rect 417570 40508 417630 41780
rect 470319 41838 471102 41840
rect 470319 41782 470324 41838
rect 470380 41782 471102 41838
rect 470319 41780 471102 41782
rect 470319 41777 470385 41780
rect 458607 40508 458673 40511
rect 417570 40506 458673 40508
rect 417570 40450 458612 40506
rect 458668 40450 458673 40506
rect 417570 40448 458673 40450
rect 471042 40508 471102 41780
rect 471663 41838 478110 41840
rect 471663 41782 471668 41838
rect 471724 41782 478110 41838
rect 471663 41780 478110 41782
rect 471663 41777 471729 41780
rect 478050 40656 478110 41780
rect 505359 40656 505425 40659
rect 478050 40654 505425 40656
rect 478050 40598 505364 40654
rect 505420 40598 505425 40654
rect 478050 40596 505425 40598
rect 505359 40593 505425 40596
rect 545199 40508 545265 40511
rect 471042 40506 545265 40508
rect 471042 40450 545204 40506
rect 545260 40450 545265 40506
rect 471042 40448 545265 40450
rect 224559 40445 224625 40448
rect 345615 40445 345681 40448
rect 458607 40445 458673 40448
rect 545199 40445 545265 40448
rect 142095 40212 142161 40215
rect 141762 40210 142161 40212
rect 141762 40154 142100 40210
rect 142156 40154 142161 40210
rect 141762 40152 142161 40154
rect 141762 39886 141822 40152
rect 142095 40149 142161 40152
rect 311055 37252 311121 37255
rect 324303 37252 324369 37255
rect 311055 37250 324369 37252
rect 311055 37194 311060 37250
rect 311116 37194 324308 37250
rect 324364 37194 324369 37250
rect 311055 37192 324369 37194
rect 311055 37189 311121 37192
rect 324303 37189 324369 37192
<< via3 >>
rect 40384 813894 40448 813958
rect 40576 812710 40640 812774
rect 41536 808862 41600 808926
rect 41152 801314 41216 801378
rect 41728 800486 41792 800490
rect 41728 800430 41740 800486
rect 41740 800430 41792 800486
rect 41728 800426 41792 800430
rect 41920 800338 41984 800342
rect 41920 800282 41972 800338
rect 41972 800282 41984 800338
rect 41920 800278 41984 800282
rect 42304 800278 42368 800342
rect 41920 798118 41984 798122
rect 41920 798062 41972 798118
rect 41972 798062 41984 798118
rect 41920 798058 41984 798062
rect 42304 795394 42368 795458
rect 41728 792938 41792 792942
rect 41728 792882 41780 792938
rect 41780 792882 41792 792938
rect 41728 792878 41792 792882
rect 41536 791842 41600 791906
rect 41152 791694 41216 791758
rect 675136 787994 675200 788058
rect 675712 787166 675776 787170
rect 675712 787110 675724 787166
rect 675724 787110 675776 787166
rect 675712 787106 675776 787110
rect 674176 786662 674240 786726
rect 675328 784798 675392 784802
rect 675328 784742 675380 784798
rect 675380 784742 675392 784798
rect 675328 784738 675392 784742
rect 676096 784146 676160 784210
rect 673984 783406 674048 783470
rect 675520 780654 675584 780658
rect 675520 780598 675532 780654
rect 675532 780598 675584 780654
rect 675520 780594 675584 780598
rect 676288 779854 676352 779918
rect 676480 779114 676544 779178
rect 676672 777634 676736 777698
rect 675904 775414 675968 775478
rect 40384 774526 40448 774590
rect 40576 773934 40640 773998
rect 675712 771862 675776 771926
rect 40384 770678 40448 770742
rect 40576 769642 40640 769706
rect 40768 758838 40832 758902
rect 43072 758010 43136 758014
rect 43072 757954 43084 758010
rect 43084 757954 43136 758010
rect 43072 757950 43136 757954
rect 40960 757506 41024 757570
rect 42880 757210 42944 757274
rect 42112 757062 42176 757126
rect 42112 754694 42176 754758
rect 42880 751586 42944 751650
rect 43072 750402 43136 750466
rect 40768 747146 40832 747210
rect 40960 746850 41024 746914
rect 676288 745814 676352 745878
rect 677440 745814 677504 745878
rect 674368 741078 674432 741142
rect 674944 740338 675008 740402
rect 674560 739598 674624 739662
rect 676864 737970 676928 738034
rect 675712 735514 675776 735518
rect 675712 735458 675724 735514
rect 675724 735458 675776 735514
rect 675712 735454 675776 735458
rect 676480 732938 676544 733002
rect 677056 732938 677120 733002
rect 676864 732494 676928 732558
rect 676864 732050 676928 732114
rect 674752 731606 674816 731670
rect 40384 731458 40448 731522
rect 40576 731310 40640 731374
rect 676288 728498 676352 728562
rect 676672 728054 676736 728118
rect 42688 715830 42752 715834
rect 42688 715774 42740 715830
rect 42740 715774 42752 715830
rect 42688 715770 42752 715774
rect 40384 715622 40448 715686
rect 41344 714882 41408 714946
rect 42880 714498 42944 714502
rect 42880 714442 42892 714498
rect 42892 714442 42944 714498
rect 42880 714438 42944 714442
rect 42112 714202 42176 714206
rect 42112 714146 42164 714202
rect 42164 714146 42176 714202
rect 42112 714142 42176 714146
rect 42496 713994 42560 714058
rect 42304 713846 42368 713910
rect 674176 711182 674240 711246
rect 42304 711034 42368 711098
rect 42496 710738 42560 710802
rect 675904 710590 675968 710654
rect 675136 710442 675200 710506
rect 675328 709702 675392 709766
rect 675520 709110 675584 709174
rect 42880 708222 42944 708286
rect 42112 707986 42176 707990
rect 42112 707930 42164 707986
rect 42164 707930 42176 707986
rect 42112 707926 42176 707930
rect 676096 707926 676160 707990
rect 42688 707186 42752 707250
rect 673984 707038 674048 707102
rect 677248 706446 677312 706510
rect 677440 705410 677504 705474
rect 41344 705114 41408 705178
rect 40384 704078 40448 704142
rect 675136 697862 675200 697926
rect 675904 697122 675968 697186
rect 674176 696974 674240 697038
rect 675520 694814 675584 694818
rect 675520 694758 675572 694814
rect 675572 694758 675584 694814
rect 675520 694754 675584 694758
rect 676672 694162 676736 694226
rect 677056 686466 677120 686530
rect 40576 684098 40640 684162
rect 40384 682914 40448 682978
rect 41536 673590 41600 673654
rect 41344 671074 41408 671138
rect 41728 670986 41792 670990
rect 41728 670930 41740 670986
rect 41740 670930 41792 670986
rect 41728 670926 41792 670930
rect 41920 670838 41984 670842
rect 41920 670782 41932 670838
rect 41932 670782 41984 670838
rect 41920 670778 41984 670782
rect 42112 670690 42176 670694
rect 42112 670634 42124 670690
rect 42124 670634 42176 670690
rect 42112 670630 42176 670634
rect 41920 666694 41984 666698
rect 41920 666638 41932 666694
rect 41932 666638 41984 666694
rect 41920 666634 41984 666638
rect 42112 664770 42176 664774
rect 42112 664714 42164 664770
rect 42164 664714 42176 664770
rect 42112 664710 42176 664714
rect 674368 664562 674432 664626
rect 676288 663822 676352 663886
rect 674944 663082 675008 663146
rect 675712 662490 675776 662554
rect 674752 661602 674816 661666
rect 41728 660922 41792 660926
rect 41728 660866 41780 660922
rect 41780 660866 41792 660922
rect 41728 660862 41792 660866
rect 674560 661010 674624 661074
rect 41344 660270 41408 660334
rect 41536 659678 41600 659742
rect 676864 659234 676928 659298
rect 674944 652574 675008 652638
rect 674368 652130 674432 652194
rect 674752 651390 674816 651454
rect 675328 649674 675392 649678
rect 675328 649618 675380 649674
rect 675380 649618 675392 649674
rect 675328 649614 675392 649618
rect 675712 645382 675776 645386
rect 675712 645326 675724 645382
rect 675724 645326 675776 645382
rect 675712 645322 675776 645326
rect 40576 645026 40640 645090
rect 40384 644878 40448 644942
rect 41728 641030 41792 641094
rect 673984 639994 674048 640058
rect 676096 638514 676160 638578
rect 41536 638218 41600 638282
rect 676672 636590 676736 636654
rect 40384 628006 40448 628070
rect 40768 627858 40832 627922
rect 42304 627414 42368 627478
rect 41536 625194 41600 625258
rect 42304 624750 42368 624814
rect 674176 620902 674240 620966
rect 675136 619866 675200 619930
rect 675520 619422 675584 619486
rect 40384 617646 40448 617710
rect 675904 617942 675968 618006
rect 40768 617202 40832 617266
rect 677056 615722 677120 615786
rect 674176 607730 674240 607794
rect 675136 606014 675200 606018
rect 675136 605958 675188 606014
rect 675188 605958 675200 606014
rect 675136 605954 675200 605958
rect 674560 604770 674624 604834
rect 41728 602106 41792 602170
rect 675520 600242 675584 600246
rect 675520 600186 675532 600242
rect 675532 600186 675584 600242
rect 675520 600182 675584 600186
rect 41920 597888 41984 597952
rect 41728 596926 41792 596990
rect 676288 595298 676352 595362
rect 675904 593374 675968 593438
rect 40576 584790 40640 584854
rect 40384 584642 40448 584706
rect 42112 584642 42176 584706
rect 41536 584554 41600 584558
rect 41536 584498 41548 584554
rect 41548 584498 41600 584554
rect 41536 584494 41600 584498
rect 42304 584494 42368 584558
rect 41344 584198 41408 584262
rect 42304 578574 42368 578638
rect 42112 578190 42176 578194
rect 42112 578134 42124 578190
rect 42124 578134 42176 578190
rect 42112 578130 42176 578134
rect 41536 576798 41600 576862
rect 674752 575762 674816 575826
rect 673984 575022 674048 575086
rect 40576 574430 40640 574494
rect 674944 574430 675008 574494
rect 675328 574282 675392 574346
rect 40384 573986 40448 574050
rect 675712 573542 675776 573606
rect 41344 573394 41408 573458
rect 676096 572802 676160 572866
rect 674368 572506 674432 572570
rect 674944 562886 675008 562950
rect 675328 561702 675392 561766
rect 674368 561406 674432 561470
rect 674752 558890 674816 558954
rect 41920 547198 41984 547262
rect 41728 544386 41792 544450
rect 41920 540242 41984 540306
rect 40576 539502 40640 539566
rect 42304 537578 42368 537642
rect 41728 536306 41792 536310
rect 41728 536250 41780 536306
rect 41780 536250 41792 536306
rect 41728 536246 41792 536250
rect 42112 535802 42176 535866
rect 41536 534914 41600 534978
rect 41920 534974 41984 534978
rect 41920 534918 41972 534974
rect 41972 534918 41984 534974
rect 41920 534914 41984 534918
rect 41728 534322 41792 534386
rect 41728 533938 41792 533942
rect 41728 533882 41780 533938
rect 41780 533882 41792 533938
rect 41728 533878 41792 533882
rect 41728 532768 41792 532832
rect 42304 532694 42368 532758
rect 41920 532250 41984 532314
rect 41344 531473 41408 531537
rect 675136 530770 675200 530834
rect 42112 530622 42176 530686
rect 41344 530369 41408 530433
rect 676288 530474 676352 530538
rect 674176 529882 674240 529946
rect 41536 529586 41600 529650
rect 674560 529290 674624 529354
rect 675520 528698 675584 528762
rect 675904 528106 675968 528170
rect 41344 524998 41408 525062
rect 674368 486370 674432 486434
rect 674944 485630 675008 485694
rect 675328 483410 675392 483474
rect 674752 482818 674816 482882
rect 40384 425542 40448 425606
rect 40576 424654 40640 424718
rect 41728 424358 41792 424422
rect 40768 423618 40832 423682
rect 41344 423174 41408 423238
rect 41920 422878 41984 422942
rect 40960 421694 41024 421758
rect 41536 421102 41600 421166
rect 41152 420658 41216 420722
rect 42112 419326 42176 419390
rect 40384 418734 40448 418798
rect 41728 411186 41792 411250
rect 41920 406066 41984 406070
rect 41920 406010 41932 406066
rect 41932 406010 41984 406066
rect 41920 406006 41984 406010
rect 42112 403846 42176 403850
rect 42112 403790 42124 403846
rect 42124 403790 42176 403846
rect 42112 403786 42176 403790
rect 41152 403046 41216 403110
rect 41536 402602 41600 402666
rect 41344 401862 41408 401926
rect 40576 400086 40640 400150
rect 40960 399494 41024 399558
rect 40768 398754 40832 398818
rect 675904 398162 675968 398226
rect 673984 397570 674048 397634
rect 675136 396830 675200 396894
rect 676672 396386 676736 396450
rect 674944 396090 675008 396154
rect 675712 395202 675776 395266
rect 675328 394610 675392 394674
rect 676480 393870 676544 393934
rect 676288 393278 676352 393342
rect 674368 393130 674432 393194
rect 675520 392538 675584 392602
rect 676096 391798 676160 391862
rect 674176 391650 674240 391714
rect 675136 385938 675200 385942
rect 675136 385882 675188 385938
rect 675188 385882 675200 385938
rect 675136 385878 675200 385882
rect 675712 385642 675776 385646
rect 675712 385586 675764 385642
rect 675764 385586 675776 385642
rect 675712 385582 675776 385586
rect 675904 384842 675968 384906
rect 676672 382918 676736 382982
rect 40384 382622 40448 382686
rect 41728 382326 41792 382390
rect 675328 382326 675392 382390
rect 676480 381734 676544 381798
rect 39808 381142 39872 381206
rect 675520 381202 675584 381206
rect 675520 381146 675572 381202
rect 675572 381146 675584 381202
rect 675520 381142 675584 381146
rect 40000 380254 40064 380318
rect 674944 378774 675008 378838
rect 40576 378034 40640 378098
rect 676096 378034 676160 378098
rect 674368 377146 674432 377210
rect 674176 376702 674240 376766
rect 41920 376406 41984 376470
rect 676288 375666 676352 375730
rect 40768 374186 40832 374250
rect 673984 373890 674048 373954
rect 41536 373742 41600 373806
rect 40000 373594 40064 373658
rect 41344 373594 41408 373658
rect 42112 373150 42176 373214
rect 42304 372706 42368 372770
rect 40960 372410 41024 372474
rect 40384 368118 40448 368182
rect 41536 362790 41600 362854
rect 41920 360630 41984 360634
rect 41920 360574 41972 360630
rect 41972 360574 41984 360630
rect 41920 360570 41984 360574
rect 40576 359830 40640 359894
rect 42112 359298 42176 359302
rect 42112 359242 42124 359298
rect 42124 359242 42176 359298
rect 42112 359238 42176 359242
rect 41344 358794 41408 358858
rect 40960 356870 41024 356934
rect 40768 356130 40832 356194
rect 42304 355686 42368 355750
rect 673984 355390 674048 355454
rect 674176 354502 674240 354566
rect 674368 353318 674432 353382
rect 675712 352948 675776 353012
rect 675904 351394 675968 351458
rect 674560 350950 674624 351014
rect 675520 348434 675584 348498
rect 676480 342958 676544 343022
rect 676672 342810 676736 342874
rect 675712 339614 675776 339618
rect 675712 339558 675764 339614
rect 675764 339558 675776 339614
rect 675712 339554 675776 339558
rect 39808 338222 39872 338286
rect 675904 337778 675968 337842
rect 40384 337186 40448 337250
rect 40576 336742 40640 336806
rect 40960 335706 41024 335770
rect 41152 335114 41216 335178
rect 41920 334818 41984 334882
rect 674560 333486 674624 333550
rect 42112 333338 42176 333402
rect 42496 332598 42560 332662
rect 40768 331118 40832 331182
rect 39808 330674 39872 330738
rect 41536 330674 41600 330738
rect 675520 330586 675584 330590
rect 675520 330530 675572 330586
rect 675572 330530 675584 330586
rect 675520 330526 675584 330530
rect 42304 329194 42368 329258
rect 40384 328306 40448 328370
rect 41344 328306 41408 328370
rect 676672 328010 676736 328074
rect 676480 326826 676544 326890
rect 41536 324902 41600 324966
rect 42496 320462 42560 320526
rect 40576 319722 40640 319786
rect 42112 317414 42176 317418
rect 42112 317358 42164 317414
rect 42164 317358 42176 317414
rect 42112 317354 42176 317358
rect 41920 316822 41984 316826
rect 41920 316766 41932 316822
rect 41932 316766 41984 316822
rect 41920 316762 41984 316766
rect 41152 316022 41216 316086
rect 41344 315578 41408 315642
rect 42304 313654 42368 313718
rect 40960 313062 41024 313126
rect 40768 312322 40832 312386
rect 673984 310990 674048 311054
rect 675328 310398 675392 310462
rect 674176 309806 674240 309870
rect 675136 309066 675200 309130
rect 674368 308918 674432 308982
rect 675520 308326 675584 308390
rect 674560 307438 674624 307502
rect 673984 306402 674048 306466
rect 674752 305958 674816 306022
rect 674944 302554 675008 302618
rect 675712 299150 675776 299214
rect 676672 298706 676736 298770
rect 41536 294858 41600 294922
rect 42304 294710 42368 294774
rect 40384 293970 40448 294034
rect 41920 293674 41984 293738
rect 673984 292786 674048 292850
rect 40960 292490 41024 292554
rect 41152 292046 41216 292110
rect 41344 291454 41408 291518
rect 40576 289974 40640 290038
rect 674752 288494 674816 288558
rect 41920 287902 41984 287966
rect 42496 287902 42560 287966
rect 674944 287310 675008 287374
rect 675712 285298 675776 285302
rect 675712 285242 675724 285298
rect 675724 285242 675776 285298
rect 675712 285238 675776 285242
rect 41728 285090 41792 285154
rect 674560 283610 674624 283674
rect 676672 281834 676736 281898
rect 41536 281686 41600 281750
rect 41920 281538 41984 281602
rect 675136 278430 675200 278494
rect 675520 278282 675584 278346
rect 674176 278134 674240 278198
rect 41920 278046 41984 278050
rect 41920 277990 41972 278046
rect 41972 277990 41984 278046
rect 41920 277986 41984 277990
rect 42496 276506 42560 276570
rect 42112 274286 42176 274350
rect 40576 274138 40640 274202
rect 41344 273546 41408 273610
rect 41152 272806 41216 272870
rect 40384 272214 40448 272278
rect 41728 270646 41792 270650
rect 41728 270590 41780 270646
rect 41780 270590 41792 270646
rect 41728 270586 41792 270590
rect 40960 269994 41024 270058
rect 42304 269254 42368 269318
rect 675328 265998 675392 266062
rect 673984 265406 674048 265470
rect 676288 261706 676352 261770
rect 675712 260966 675776 261030
rect 675520 258894 675584 258958
rect 674944 258450 675008 258514
rect 674560 257858 674624 257922
rect 674752 256378 674816 256442
rect 675904 253270 675968 253334
rect 676096 253122 676160 253186
rect 40768 252234 40832 252298
rect 41728 252012 41792 252076
rect 40576 251642 40640 251706
rect 40960 250754 41024 250818
rect 676288 250754 676352 250818
rect 41536 250310 41600 250374
rect 41920 249570 41984 249634
rect 41152 248830 41216 248894
rect 41344 248238 41408 248302
rect 40384 246758 40448 246822
rect 675520 246670 675584 246674
rect 675520 246614 675572 246670
rect 675572 246614 675584 246670
rect 675520 246610 675584 246614
rect 675712 243562 675776 243566
rect 675712 243506 675724 243562
rect 675724 243506 675776 243562
rect 675712 243502 675776 243506
rect 674560 242022 674624 242086
rect 674752 241726 674816 241790
rect 674944 240542 675008 240606
rect 676096 238618 676160 238682
rect 41728 237938 41792 237942
rect 41728 237882 41780 237938
rect 41780 237882 41792 237938
rect 41728 237878 41792 237882
rect 40768 237138 40832 237202
rect 41536 237138 41600 237202
rect 675904 236842 675968 236906
rect 409024 236694 409088 236758
rect 408640 236102 408704 236166
rect 409024 235806 409088 235870
rect 408448 235066 408512 235130
rect 41728 233350 41792 233354
rect 41728 233294 41780 233350
rect 41780 233294 41792 233350
rect 41728 233290 41792 233294
rect 40384 231070 40448 231134
rect 41344 230330 41408 230394
rect 41152 229590 41216 229654
rect 40960 228998 41024 229062
rect 41536 227370 41600 227434
rect 41920 226838 41984 226842
rect 41920 226782 41932 226838
rect 41932 226782 41984 226838
rect 41920 226778 41984 226782
rect 40576 225890 40640 225954
rect 673984 220710 674048 220774
rect 674368 219970 674432 220034
rect 673984 219230 674048 219294
rect 674176 218194 674240 218258
rect 675904 217750 675968 217814
rect 675712 216270 675776 216334
rect 675520 215678 675584 215742
rect 676288 207686 676352 207750
rect 676672 207538 676736 207602
rect 676480 207390 676544 207454
rect 41152 205910 41216 205974
rect 41344 205318 41408 205382
rect 40768 204874 40832 204938
rect 41920 203542 41984 203606
rect 675904 204430 675968 204494
rect 675712 202714 675776 202718
rect 675712 202658 675724 202714
rect 675724 202658 675776 202714
rect 675712 202654 675776 202658
rect 40960 201470 41024 201534
rect 41728 200878 41792 200942
rect 42304 200730 42368 200794
rect 42112 199990 42176 200054
rect 41536 199694 41600 199758
rect 675520 198422 675584 198426
rect 675520 198366 675572 198422
rect 675572 198366 675584 198422
rect 675520 198362 675584 198366
rect 41728 195314 41792 195318
rect 41728 195258 41780 195314
rect 41780 195258 41792 195314
rect 41728 195254 41792 195258
rect 676480 195254 676544 195318
rect 676288 193478 676352 193542
rect 676672 191554 676736 191618
rect 41536 190074 41600 190138
rect 41344 189630 41408 189694
rect 41344 189186 41408 189250
rect 41920 187914 41984 187918
rect 41920 187858 41932 187914
rect 41932 187858 41984 187914
rect 41920 187854 41984 187858
rect 40768 187114 40832 187178
rect 41344 186670 41408 186734
rect 40960 185782 41024 185846
rect 42304 184154 42368 184218
rect 41920 183622 41984 183626
rect 41920 183566 41932 183622
rect 41932 183566 41984 183622
rect 41920 183562 41984 183566
rect 42112 182882 42176 182886
rect 42112 182826 42124 182882
rect 42124 182826 42176 182882
rect 42112 182822 42176 182826
rect 674368 176162 674432 176226
rect 674368 175570 674432 175634
rect 673984 175422 674048 175486
rect 674176 174090 674240 174154
rect 674176 173942 674240 174006
rect 673984 173498 674048 173562
rect 675904 173202 675968 173266
rect 675136 171130 675200 171194
rect 674752 168614 674816 168678
rect 674944 168170 675008 168234
rect 674560 167134 674624 167198
rect 675712 161510 675776 161574
rect 676672 161362 676736 161426
rect 675904 159290 675968 159354
rect 675136 153370 675200 153434
rect 674560 152482 674624 152546
rect 674944 152186 675008 152250
rect 674752 150262 674816 150326
rect 675712 148546 675776 148550
rect 675712 148490 675764 148546
rect 675764 148490 675776 148546
rect 675712 148486 675776 148490
rect 676672 146562 676736 146626
rect 674368 130578 674432 130642
rect 674176 129394 674240 129458
rect 673984 128506 674048 128570
rect 674368 125546 674432 125610
rect 674560 123030 674624 123094
rect 673984 122142 674048 122206
rect 676480 117998 676544 118062
rect 675904 117850 675968 117914
rect 674368 108082 674432 108146
rect 673984 106602 674048 106666
rect 674560 105122 674624 105186
rect 675904 103198 675968 103262
rect 676480 101422 676544 101486
<< metal4 >>
rect 40383 813958 40449 813959
rect 40383 813894 40384 813958
rect 40448 813894 40449 813958
rect 40383 813893 40449 813894
rect 40386 774591 40446 813893
rect 40575 812774 40641 812775
rect 40575 812710 40576 812774
rect 40640 812710 40641 812774
rect 40575 812709 40641 812710
rect 40383 774590 40449 774591
rect 40383 774526 40384 774590
rect 40448 774526 40449 774590
rect 40383 774525 40449 774526
rect 40578 773999 40638 812709
rect 41535 808926 41601 808927
rect 41535 808862 41536 808926
rect 41600 808862 41601 808926
rect 41535 808861 41601 808862
rect 41151 801378 41217 801379
rect 41151 801314 41152 801378
rect 41216 801314 41217 801378
rect 41151 801313 41217 801314
rect 41154 791759 41214 801313
rect 41538 791907 41598 808861
rect 41727 800490 41793 800491
rect 41727 800426 41728 800490
rect 41792 800426 41793 800490
rect 41727 800425 41793 800426
rect 41730 792943 41790 800425
rect 41919 800342 41985 800343
rect 41919 800278 41920 800342
rect 41984 800278 41985 800342
rect 41919 800277 41985 800278
rect 42303 800342 42369 800343
rect 42303 800278 42304 800342
rect 42368 800278 42369 800342
rect 42303 800277 42369 800278
rect 41922 798123 41982 800277
rect 41919 798122 41985 798123
rect 41919 798058 41920 798122
rect 41984 798058 41985 798122
rect 41919 798057 41985 798058
rect 42306 795459 42366 800277
rect 42303 795458 42369 795459
rect 42303 795394 42304 795458
rect 42368 795394 42369 795458
rect 42303 795393 42369 795394
rect 41727 792942 41793 792943
rect 41727 792878 41728 792942
rect 41792 792878 41793 792942
rect 41727 792877 41793 792878
rect 41535 791906 41601 791907
rect 41535 791842 41536 791906
rect 41600 791842 41601 791906
rect 41535 791841 41601 791842
rect 41151 791758 41217 791759
rect 41151 791694 41152 791758
rect 41216 791694 41217 791758
rect 41151 791693 41217 791694
rect 675135 788058 675201 788059
rect 675135 787994 675136 788058
rect 675200 787994 675201 788058
rect 675135 787993 675201 787994
rect 674175 786726 674241 786727
rect 674175 786662 674176 786726
rect 674240 786662 674241 786726
rect 674175 786661 674241 786662
rect 673983 783470 674049 783471
rect 673983 783406 673984 783470
rect 674048 783406 674049 783470
rect 673983 783405 674049 783406
rect 40575 773998 40641 773999
rect 40575 773934 40576 773998
rect 40640 773934 40641 773998
rect 40575 773933 40641 773934
rect 40383 770742 40449 770743
rect 40383 770678 40384 770742
rect 40448 770678 40449 770742
rect 40383 770677 40449 770678
rect 40386 731523 40446 770677
rect 40575 769706 40641 769707
rect 40575 769642 40576 769706
rect 40640 769642 40641 769706
rect 40575 769641 40641 769642
rect 40383 731522 40449 731523
rect 40383 731458 40384 731522
rect 40448 731458 40449 731522
rect 40383 731457 40449 731458
rect 40578 731375 40638 769641
rect 40767 758902 40833 758903
rect 40767 758838 40768 758902
rect 40832 758838 40833 758902
rect 40767 758837 40833 758838
rect 40770 747211 40830 758837
rect 43071 758014 43137 758015
rect 43071 757950 43072 758014
rect 43136 757950 43137 758014
rect 43071 757949 43137 757950
rect 40959 757570 41025 757571
rect 40959 757506 40960 757570
rect 41024 757506 41025 757570
rect 40959 757505 41025 757506
rect 40767 747210 40833 747211
rect 40767 747146 40768 747210
rect 40832 747146 40833 747210
rect 40767 747145 40833 747146
rect 40962 746915 41022 757505
rect 42879 757274 42945 757275
rect 42879 757210 42880 757274
rect 42944 757210 42945 757274
rect 42879 757209 42945 757210
rect 42111 757126 42177 757127
rect 42111 757062 42112 757126
rect 42176 757062 42177 757126
rect 42111 757061 42177 757062
rect 42114 754759 42174 757061
rect 42111 754758 42177 754759
rect 42111 754694 42112 754758
rect 42176 754694 42177 754758
rect 42111 754693 42177 754694
rect 42882 751651 42942 757209
rect 42879 751650 42945 751651
rect 42879 751586 42880 751650
rect 42944 751586 42945 751650
rect 42879 751585 42945 751586
rect 43074 750467 43134 757949
rect 43071 750466 43137 750467
rect 43071 750402 43072 750466
rect 43136 750402 43137 750466
rect 43071 750401 43137 750402
rect 40959 746914 41025 746915
rect 40959 746850 40960 746914
rect 41024 746850 41025 746914
rect 40959 746849 41025 746850
rect 40575 731374 40641 731375
rect 40575 731310 40576 731374
rect 40640 731310 40641 731374
rect 40575 731309 40641 731310
rect 42687 715834 42753 715835
rect 42687 715770 42688 715834
rect 42752 715770 42753 715834
rect 42687 715769 42753 715770
rect 40383 715686 40449 715687
rect 40383 715622 40384 715686
rect 40448 715622 40449 715686
rect 40383 715621 40449 715622
rect 40386 704143 40446 715621
rect 41343 714946 41409 714947
rect 41343 714882 41344 714946
rect 41408 714882 41409 714946
rect 41343 714881 41409 714882
rect 41346 705179 41406 714881
rect 42111 714206 42177 714207
rect 42111 714142 42112 714206
rect 42176 714142 42177 714206
rect 42111 714141 42177 714142
rect 42114 707991 42174 714141
rect 42495 714058 42561 714059
rect 42495 713994 42496 714058
rect 42560 713994 42561 714058
rect 42495 713993 42561 713994
rect 42303 713910 42369 713911
rect 42303 713846 42304 713910
rect 42368 713846 42369 713910
rect 42303 713845 42369 713846
rect 42306 711099 42366 713845
rect 42303 711098 42369 711099
rect 42303 711034 42304 711098
rect 42368 711034 42369 711098
rect 42303 711033 42369 711034
rect 42498 710803 42558 713993
rect 42495 710802 42561 710803
rect 42495 710738 42496 710802
rect 42560 710738 42561 710802
rect 42495 710737 42561 710738
rect 42111 707990 42177 707991
rect 42111 707926 42112 707990
rect 42176 707926 42177 707990
rect 42111 707925 42177 707926
rect 42690 707251 42750 715769
rect 42879 714502 42945 714503
rect 42879 714438 42880 714502
rect 42944 714438 42945 714502
rect 42879 714437 42945 714438
rect 42882 708287 42942 714437
rect 42879 708286 42945 708287
rect 42879 708222 42880 708286
rect 42944 708222 42945 708286
rect 42879 708221 42945 708222
rect 42687 707250 42753 707251
rect 42687 707186 42688 707250
rect 42752 707186 42753 707250
rect 42687 707185 42753 707186
rect 673986 707103 674046 783405
rect 674178 711247 674238 786661
rect 674367 741142 674433 741143
rect 674367 741078 674368 741142
rect 674432 741078 674433 741142
rect 674367 741077 674433 741078
rect 674175 711246 674241 711247
rect 674175 711182 674176 711246
rect 674240 711182 674241 711246
rect 674175 711181 674241 711182
rect 673983 707102 674049 707103
rect 673983 707038 673984 707102
rect 674048 707038 674049 707102
rect 673983 707037 674049 707038
rect 41343 705178 41409 705179
rect 41343 705114 41344 705178
rect 41408 705114 41409 705178
rect 41343 705113 41409 705114
rect 40383 704142 40449 704143
rect 40383 704078 40384 704142
rect 40448 704078 40449 704142
rect 40383 704077 40449 704078
rect 674175 697038 674241 697039
rect 674175 696974 674176 697038
rect 674240 696974 674241 697038
rect 674175 696973 674241 696974
rect 40575 684162 40641 684163
rect 40575 684098 40576 684162
rect 40640 684098 40641 684162
rect 40575 684097 40641 684098
rect 40383 682978 40449 682979
rect 40383 682914 40384 682978
rect 40448 682914 40449 682978
rect 40383 682913 40449 682914
rect 40386 644943 40446 682913
rect 40578 645091 40638 684097
rect 41535 673654 41601 673655
rect 41535 673590 41536 673654
rect 41600 673590 41601 673654
rect 41535 673589 41601 673590
rect 41343 671138 41409 671139
rect 41343 671074 41344 671138
rect 41408 671074 41409 671138
rect 41343 671073 41409 671074
rect 41346 660335 41406 671073
rect 41343 660334 41409 660335
rect 41343 660270 41344 660334
rect 41408 660270 41409 660334
rect 41343 660269 41409 660270
rect 41538 659743 41598 673589
rect 41727 670990 41793 670991
rect 41727 670926 41728 670990
rect 41792 670926 41793 670990
rect 41727 670925 41793 670926
rect 41730 660927 41790 670925
rect 41919 670842 41985 670843
rect 41919 670778 41920 670842
rect 41984 670778 41985 670842
rect 41919 670777 41985 670778
rect 41922 666699 41982 670777
rect 42111 670694 42177 670695
rect 42111 670630 42112 670694
rect 42176 670630 42177 670694
rect 42111 670629 42177 670630
rect 41919 666698 41985 666699
rect 41919 666634 41920 666698
rect 41984 666634 41985 666698
rect 41919 666633 41985 666634
rect 42114 664775 42174 670629
rect 42111 664774 42177 664775
rect 42111 664710 42112 664774
rect 42176 664710 42177 664774
rect 42111 664709 42177 664710
rect 41727 660926 41793 660927
rect 41727 660862 41728 660926
rect 41792 660862 41793 660926
rect 41727 660861 41793 660862
rect 41535 659742 41601 659743
rect 41535 659678 41536 659742
rect 41600 659678 41601 659742
rect 41535 659677 41601 659678
rect 40575 645090 40641 645091
rect 40575 645026 40576 645090
rect 40640 645026 40641 645090
rect 40575 645025 40641 645026
rect 40383 644942 40449 644943
rect 40383 644878 40384 644942
rect 40448 644878 40449 644942
rect 40383 644877 40449 644878
rect 41727 641094 41793 641095
rect 41727 641030 41728 641094
rect 41792 641030 41793 641094
rect 41727 641029 41793 641030
rect 41535 638282 41601 638283
rect 41535 638218 41536 638282
rect 41600 638218 41601 638282
rect 41535 638217 41601 638218
rect 40383 628070 40449 628071
rect 40383 628006 40384 628070
rect 40448 628006 40449 628070
rect 40383 628005 40449 628006
rect 40386 617711 40446 628005
rect 40767 627922 40833 627923
rect 40767 627858 40768 627922
rect 40832 627858 40833 627922
rect 40767 627857 40833 627858
rect 40383 617710 40449 617711
rect 40383 617646 40384 617710
rect 40448 617646 40449 617710
rect 40383 617645 40449 617646
rect 40770 617267 40830 627857
rect 41538 625259 41598 638217
rect 41535 625258 41601 625259
rect 41535 625194 41536 625258
rect 41600 625194 41601 625258
rect 41535 625193 41601 625194
rect 40767 617266 40833 617267
rect 40767 617202 40768 617266
rect 40832 617202 40833 617266
rect 40767 617201 40833 617202
rect 41730 602171 41790 641029
rect 673983 640058 674049 640059
rect 673983 639994 673984 640058
rect 674048 639994 674049 640058
rect 673983 639993 674049 639994
rect 42303 627478 42369 627479
rect 42303 627414 42304 627478
rect 42368 627414 42369 627478
rect 42303 627413 42369 627414
rect 42306 624815 42366 627413
rect 42303 624814 42369 624815
rect 42303 624750 42304 624814
rect 42368 624750 42369 624814
rect 42303 624749 42369 624750
rect 41727 602170 41793 602171
rect 41727 602106 41728 602170
rect 41792 602106 41793 602170
rect 41727 602105 41793 602106
rect 41919 597952 41985 597953
rect 41919 597888 41920 597952
rect 41984 597888 41985 597952
rect 41919 597887 41985 597888
rect 41727 596990 41793 596991
rect 41727 596926 41728 596990
rect 41792 596926 41793 596990
rect 41727 596925 41793 596926
rect 40575 584854 40641 584855
rect 40575 584790 40576 584854
rect 40640 584790 40641 584854
rect 40575 584789 40641 584790
rect 40383 584706 40449 584707
rect 40383 584642 40384 584706
rect 40448 584642 40449 584706
rect 40383 584641 40449 584642
rect 40386 574051 40446 584641
rect 40578 574495 40638 584789
rect 41535 584558 41601 584559
rect 41535 584494 41536 584558
rect 41600 584494 41601 584558
rect 41535 584493 41601 584494
rect 41343 584262 41409 584263
rect 41343 584198 41344 584262
rect 41408 584198 41409 584262
rect 41343 584197 41409 584198
rect 40575 574494 40641 574495
rect 40575 574430 40576 574494
rect 40640 574430 40641 574494
rect 40575 574429 40641 574430
rect 40383 574050 40449 574051
rect 40383 573986 40384 574050
rect 40448 573986 40449 574050
rect 40383 573985 40449 573986
rect 41346 573459 41406 584197
rect 41538 576863 41598 584493
rect 41535 576862 41601 576863
rect 41535 576798 41536 576862
rect 41600 576798 41601 576862
rect 41535 576797 41601 576798
rect 41343 573458 41409 573459
rect 41343 573394 41344 573458
rect 41408 573394 41409 573458
rect 41343 573393 41409 573394
rect 41730 544451 41790 596925
rect 41922 547263 41982 597887
rect 42111 584706 42177 584707
rect 42111 584642 42112 584706
rect 42176 584642 42177 584706
rect 42111 584641 42177 584642
rect 42114 578195 42174 584641
rect 42303 584558 42369 584559
rect 42303 584494 42304 584558
rect 42368 584494 42369 584558
rect 42303 584493 42369 584494
rect 42306 578639 42366 584493
rect 42303 578638 42369 578639
rect 42303 578574 42304 578638
rect 42368 578574 42369 578638
rect 42303 578573 42369 578574
rect 42111 578194 42177 578195
rect 42111 578130 42112 578194
rect 42176 578130 42177 578194
rect 42111 578129 42177 578130
rect 673986 575087 674046 639993
rect 674178 620967 674238 696973
rect 674370 664627 674430 741077
rect 674943 740402 675009 740403
rect 674943 740338 674944 740402
rect 675008 740338 675009 740402
rect 674943 740337 675009 740338
rect 674559 739662 674625 739663
rect 674559 739598 674560 739662
rect 674624 739598 674625 739662
rect 674559 739597 674625 739598
rect 674367 664626 674433 664627
rect 674367 664562 674368 664626
rect 674432 664562 674433 664626
rect 674367 664561 674433 664562
rect 674562 661075 674622 739597
rect 674751 731670 674817 731671
rect 674751 731606 674752 731670
rect 674816 731606 674817 731670
rect 674751 731605 674817 731606
rect 674754 661667 674814 731605
rect 674946 663147 675006 740337
rect 675138 710507 675198 787993
rect 675711 787170 675777 787171
rect 675711 787106 675712 787170
rect 675776 787106 675777 787170
rect 675711 787105 675777 787106
rect 675327 784802 675393 784803
rect 675327 784738 675328 784802
rect 675392 784738 675393 784802
rect 675327 784737 675393 784738
rect 675135 710506 675201 710507
rect 675135 710442 675136 710506
rect 675200 710442 675201 710506
rect 675135 710441 675201 710442
rect 675330 709767 675390 784737
rect 675519 780658 675585 780659
rect 675519 780594 675520 780658
rect 675584 780594 675585 780658
rect 675519 780593 675585 780594
rect 675327 709766 675393 709767
rect 675327 709702 675328 709766
rect 675392 709702 675393 709766
rect 675327 709701 675393 709702
rect 675522 709175 675582 780593
rect 675714 771927 675774 787105
rect 676095 784210 676161 784211
rect 676095 784146 676096 784210
rect 676160 784146 676161 784210
rect 676095 784145 676161 784146
rect 675903 775478 675969 775479
rect 675903 775414 675904 775478
rect 675968 775414 675969 775478
rect 675903 775413 675969 775414
rect 675711 771926 675777 771927
rect 675711 771862 675712 771926
rect 675776 771862 675777 771926
rect 675711 771861 675777 771862
rect 675711 735518 675777 735519
rect 675711 735454 675712 735518
rect 675776 735454 675777 735518
rect 675711 735453 675777 735454
rect 675519 709174 675585 709175
rect 675519 709110 675520 709174
rect 675584 709110 675585 709174
rect 675519 709109 675585 709110
rect 675135 697926 675201 697927
rect 675135 697862 675136 697926
rect 675200 697862 675201 697926
rect 675135 697861 675201 697862
rect 674943 663146 675009 663147
rect 674943 663082 674944 663146
rect 675008 663082 675009 663146
rect 674943 663081 675009 663082
rect 674751 661666 674817 661667
rect 674751 661602 674752 661666
rect 674816 661602 674817 661666
rect 674751 661601 674817 661602
rect 674559 661074 674625 661075
rect 674559 661010 674560 661074
rect 674624 661010 674625 661074
rect 674559 661009 674625 661010
rect 674943 652638 675009 652639
rect 674943 652574 674944 652638
rect 675008 652574 675009 652638
rect 674943 652573 675009 652574
rect 674367 652194 674433 652195
rect 674367 652130 674368 652194
rect 674432 652130 674433 652194
rect 674367 652129 674433 652130
rect 674175 620966 674241 620967
rect 674175 620902 674176 620966
rect 674240 620902 674241 620966
rect 674175 620901 674241 620902
rect 674175 607794 674241 607795
rect 674175 607730 674176 607794
rect 674240 607730 674241 607794
rect 674175 607729 674241 607730
rect 673983 575086 674049 575087
rect 673983 575022 673984 575086
rect 674048 575022 674049 575086
rect 673983 575021 674049 575022
rect 41919 547262 41985 547263
rect 41919 547198 41920 547262
rect 41984 547198 41985 547262
rect 41919 547197 41985 547198
rect 41727 544450 41793 544451
rect 41727 544386 41728 544450
rect 41792 544386 41793 544450
rect 41727 544385 41793 544386
rect 41922 540307 41982 547197
rect 41919 540306 41985 540307
rect 41919 540242 41920 540306
rect 41984 540242 41985 540306
rect 41919 540241 41985 540242
rect 40575 539566 40641 539567
rect 40575 539502 40576 539566
rect 40640 539502 40641 539566
rect 40575 539501 40641 539502
rect 40578 498270 40638 539501
rect 42303 537642 42369 537643
rect 42303 537578 42304 537642
rect 42368 537578 42369 537642
rect 42303 537577 42369 537578
rect 41727 536310 41793 536311
rect 41727 536246 41728 536310
rect 41792 536246 41793 536310
rect 41727 536245 41793 536246
rect 41535 534978 41601 534979
rect 41535 534914 41536 534978
rect 41600 534914 41601 534978
rect 41535 534913 41601 534914
rect 41343 531537 41409 531538
rect 41343 531473 41344 531537
rect 41408 531473 41409 531537
rect 41343 531472 41409 531473
rect 41346 530434 41406 531472
rect 41343 530433 41409 530434
rect 41343 530369 41344 530433
rect 41408 530369 41409 530433
rect 41343 530368 41409 530369
rect 41346 525063 41406 530368
rect 41538 529651 41598 534913
rect 41730 534387 41790 536245
rect 42111 535866 42177 535867
rect 42111 535802 42112 535866
rect 42176 535802 42177 535866
rect 42111 535801 42177 535802
rect 41919 534978 41985 534979
rect 41919 534914 41920 534978
rect 41984 534914 41985 534978
rect 41919 534913 41985 534914
rect 41727 534386 41793 534387
rect 41727 534322 41728 534386
rect 41792 534322 41793 534386
rect 41727 534321 41793 534322
rect 41727 533942 41793 533943
rect 41727 533878 41728 533942
rect 41792 533878 41793 533942
rect 41727 533877 41793 533878
rect 41730 532833 41790 533877
rect 41727 532832 41793 532833
rect 41727 532768 41728 532832
rect 41792 532768 41793 532832
rect 41727 532767 41793 532768
rect 41922 532315 41982 534913
rect 41919 532314 41985 532315
rect 41919 532250 41920 532314
rect 41984 532250 41985 532314
rect 41919 532249 41985 532250
rect 42114 530687 42174 535801
rect 42306 532759 42366 537577
rect 42303 532758 42369 532759
rect 42303 532694 42304 532758
rect 42368 532694 42369 532758
rect 42303 532693 42369 532694
rect 42111 530686 42177 530687
rect 42111 530622 42112 530686
rect 42176 530622 42177 530686
rect 42111 530621 42177 530622
rect 674178 529947 674238 607729
rect 674370 572571 674430 652129
rect 674751 651454 674817 651455
rect 674751 651390 674752 651454
rect 674816 651390 674817 651454
rect 674751 651389 674817 651390
rect 674559 604834 674625 604835
rect 674559 604770 674560 604834
rect 674624 604770 674625 604834
rect 674559 604769 674625 604770
rect 674367 572570 674433 572571
rect 674367 572506 674368 572570
rect 674432 572506 674433 572570
rect 674367 572505 674433 572506
rect 674367 561470 674433 561471
rect 674367 561406 674368 561470
rect 674432 561406 674433 561470
rect 674367 561405 674433 561406
rect 674175 529946 674241 529947
rect 674175 529882 674176 529946
rect 674240 529882 674241 529946
rect 674175 529881 674241 529882
rect 41535 529650 41601 529651
rect 41535 529586 41536 529650
rect 41600 529586 41601 529650
rect 41535 529585 41601 529586
rect 41343 525062 41409 525063
rect 41343 524998 41344 525062
rect 41408 524998 41409 525062
rect 41343 524997 41409 524998
rect 40386 498210 40638 498270
rect 40386 425607 40446 498210
rect 674370 486435 674430 561405
rect 674562 529355 674622 604769
rect 674754 575827 674814 651389
rect 674751 575826 674817 575827
rect 674751 575762 674752 575826
rect 674816 575762 674817 575826
rect 674751 575761 674817 575762
rect 674946 574495 675006 652573
rect 675138 619931 675198 697861
rect 675519 694818 675585 694819
rect 675519 694754 675520 694818
rect 675584 694754 675585 694818
rect 675519 694753 675585 694754
rect 675327 649678 675393 649679
rect 675327 649614 675328 649678
rect 675392 649614 675393 649678
rect 675327 649613 675393 649614
rect 675135 619930 675201 619931
rect 675135 619866 675136 619930
rect 675200 619866 675201 619930
rect 675135 619865 675201 619866
rect 675135 606018 675201 606019
rect 675135 605954 675136 606018
rect 675200 605954 675201 606018
rect 675135 605953 675201 605954
rect 674943 574494 675009 574495
rect 674943 574430 674944 574494
rect 675008 574430 675009 574494
rect 674943 574429 675009 574430
rect 674943 562950 675009 562951
rect 674943 562886 674944 562950
rect 675008 562886 675009 562950
rect 674943 562885 675009 562886
rect 674751 558954 674817 558955
rect 674751 558890 674752 558954
rect 674816 558890 674817 558954
rect 674751 558889 674817 558890
rect 674559 529354 674625 529355
rect 674559 529290 674560 529354
rect 674624 529290 674625 529354
rect 674559 529289 674625 529290
rect 674367 486434 674433 486435
rect 674367 486370 674368 486434
rect 674432 486370 674433 486434
rect 674367 486369 674433 486370
rect 674754 482883 674814 558889
rect 674946 485695 675006 562885
rect 675138 530835 675198 605953
rect 675330 574347 675390 649613
rect 675522 619487 675582 694753
rect 675714 662555 675774 735453
rect 675906 710655 675966 775413
rect 675903 710654 675969 710655
rect 675903 710590 675904 710654
rect 675968 710590 675969 710654
rect 675903 710589 675969 710590
rect 676098 707991 676158 784145
rect 676287 779918 676353 779919
rect 676287 779854 676288 779918
rect 676352 779854 676353 779918
rect 676287 779853 676353 779854
rect 676290 745879 676350 779853
rect 676479 779178 676545 779179
rect 676479 779114 676480 779178
rect 676544 779114 676545 779178
rect 676479 779113 676545 779114
rect 676287 745878 676353 745879
rect 676287 745814 676288 745878
rect 676352 745814 676353 745878
rect 676287 745813 676353 745814
rect 676482 733003 676542 779113
rect 676671 777698 676737 777699
rect 676671 777634 676672 777698
rect 676736 777634 676737 777698
rect 676671 777633 676737 777634
rect 676479 733002 676545 733003
rect 676479 732938 676480 733002
rect 676544 732938 676545 733002
rect 676479 732937 676545 732938
rect 676287 728562 676353 728563
rect 676287 728498 676288 728562
rect 676352 728498 676353 728562
rect 676287 728497 676353 728498
rect 676095 707990 676161 707991
rect 676095 707926 676096 707990
rect 676160 707926 676161 707990
rect 676095 707925 676161 707926
rect 675903 697186 675969 697187
rect 675903 697122 675904 697186
rect 675968 697122 675969 697186
rect 675903 697121 675969 697122
rect 675711 662554 675777 662555
rect 675711 662490 675712 662554
rect 675776 662490 675777 662554
rect 675711 662489 675777 662490
rect 675711 645386 675777 645387
rect 675711 645322 675712 645386
rect 675776 645322 675777 645386
rect 675711 645321 675777 645322
rect 675519 619486 675585 619487
rect 675519 619422 675520 619486
rect 675584 619422 675585 619486
rect 675519 619421 675585 619422
rect 675519 600246 675585 600247
rect 675519 600182 675520 600246
rect 675584 600182 675585 600246
rect 675519 600181 675585 600182
rect 675327 574346 675393 574347
rect 675327 574282 675328 574346
rect 675392 574282 675393 574346
rect 675327 574281 675393 574282
rect 675327 561766 675393 561767
rect 675327 561702 675328 561766
rect 675392 561702 675393 561766
rect 675327 561701 675393 561702
rect 675135 530834 675201 530835
rect 675135 530770 675136 530834
rect 675200 530770 675201 530834
rect 675135 530769 675201 530770
rect 674943 485694 675009 485695
rect 674943 485630 674944 485694
rect 675008 485630 675009 485694
rect 674943 485629 675009 485630
rect 675330 483475 675390 561701
rect 675522 528763 675582 600181
rect 675714 573607 675774 645321
rect 675906 618007 675966 697121
rect 676290 663887 676350 728497
rect 676674 728119 676734 777633
rect 677439 745878 677505 745879
rect 677439 745814 677440 745878
rect 677504 745814 677505 745878
rect 677439 745813 677505 745814
rect 676863 738034 676929 738035
rect 676863 737970 676864 738034
rect 676928 737970 676929 738034
rect 676863 737969 676929 737970
rect 676866 732559 676926 737969
rect 677055 733002 677121 733003
rect 677055 732938 677056 733002
rect 677120 732963 677121 733002
rect 677120 732938 677310 732963
rect 677055 732937 677310 732938
rect 677058 732903 677310 732937
rect 676863 732558 676929 732559
rect 676863 732494 676864 732558
rect 676928 732494 676929 732558
rect 676863 732493 676929 732494
rect 676863 732114 676929 732115
rect 676863 732050 676864 732114
rect 676928 732050 676929 732114
rect 676863 732049 676929 732050
rect 676671 728118 676737 728119
rect 676671 728054 676672 728118
rect 676736 728054 676737 728118
rect 676671 728053 676737 728054
rect 676671 694226 676737 694227
rect 676671 694162 676672 694226
rect 676736 694162 676737 694226
rect 676671 694161 676737 694162
rect 676287 663886 676353 663887
rect 676287 663822 676288 663886
rect 676352 663822 676353 663886
rect 676287 663821 676353 663822
rect 676095 638578 676161 638579
rect 676095 638514 676096 638578
rect 676160 638514 676161 638578
rect 676095 638513 676161 638514
rect 675903 618006 675969 618007
rect 675903 617942 675904 618006
rect 675968 617942 675969 618006
rect 675903 617941 675969 617942
rect 675903 593438 675969 593439
rect 675903 593374 675904 593438
rect 675968 593374 675969 593438
rect 675903 593373 675969 593374
rect 675711 573606 675777 573607
rect 675711 573542 675712 573606
rect 675776 573542 675777 573606
rect 675711 573541 675777 573542
rect 675519 528762 675585 528763
rect 675519 528698 675520 528762
rect 675584 528698 675585 528762
rect 675519 528697 675585 528698
rect 675906 528171 675966 593373
rect 676098 572867 676158 638513
rect 676674 636655 676734 694161
rect 676866 659299 676926 732049
rect 677250 706511 677310 732903
rect 677247 706510 677313 706511
rect 677247 706446 677248 706510
rect 677312 706446 677313 706510
rect 677247 706445 677313 706446
rect 677442 705475 677502 745813
rect 677439 705474 677505 705475
rect 677439 705410 677440 705474
rect 677504 705410 677505 705474
rect 677439 705409 677505 705410
rect 677055 686530 677121 686531
rect 677055 686466 677056 686530
rect 677120 686466 677121 686530
rect 677055 686465 677121 686466
rect 676863 659298 676929 659299
rect 676863 659234 676864 659298
rect 676928 659234 676929 659298
rect 676863 659233 676929 659234
rect 676671 636654 676737 636655
rect 676671 636590 676672 636654
rect 676736 636590 676737 636654
rect 676671 636589 676737 636590
rect 677058 615787 677118 686465
rect 677055 615786 677121 615787
rect 677055 615722 677056 615786
rect 677120 615722 677121 615786
rect 677055 615721 677121 615722
rect 676287 595362 676353 595363
rect 676287 595298 676288 595362
rect 676352 595298 676353 595362
rect 676287 595297 676353 595298
rect 676095 572866 676161 572867
rect 676095 572802 676096 572866
rect 676160 572802 676161 572866
rect 676095 572801 676161 572802
rect 676290 530539 676350 595297
rect 676287 530538 676353 530539
rect 676287 530474 676288 530538
rect 676352 530474 676353 530538
rect 676287 530473 676353 530474
rect 675903 528170 675969 528171
rect 675903 528106 675904 528170
rect 675968 528106 675969 528170
rect 675903 528105 675969 528106
rect 675327 483474 675393 483475
rect 675327 483410 675328 483474
rect 675392 483410 675393 483474
rect 675327 483409 675393 483410
rect 674751 482882 674817 482883
rect 674751 482818 674752 482882
rect 674816 482818 674817 482882
rect 674751 482817 674817 482818
rect 40383 425606 40449 425607
rect 40383 425542 40384 425606
rect 40448 425542 40449 425606
rect 40383 425541 40449 425542
rect 40575 424718 40641 424719
rect 40575 424654 40576 424718
rect 40640 424654 40641 424718
rect 40575 424653 40641 424654
rect 40383 418798 40449 418799
rect 40383 418734 40384 418798
rect 40448 418734 40449 418798
rect 40383 418733 40449 418734
rect 40386 382687 40446 418733
rect 40578 400151 40638 424653
rect 41727 424422 41793 424423
rect 41727 424358 41728 424422
rect 41792 424358 41793 424422
rect 41727 424357 41793 424358
rect 40767 423682 40833 423683
rect 40767 423618 40768 423682
rect 40832 423618 40833 423682
rect 40767 423617 40833 423618
rect 40575 400150 40641 400151
rect 40575 400086 40576 400150
rect 40640 400086 40641 400150
rect 40575 400085 40641 400086
rect 40770 398819 40830 423617
rect 41343 423238 41409 423239
rect 41343 423174 41344 423238
rect 41408 423174 41409 423238
rect 41343 423173 41409 423174
rect 40959 421758 41025 421759
rect 40959 421694 40960 421758
rect 41024 421694 41025 421758
rect 40959 421693 41025 421694
rect 40962 399559 41022 421693
rect 41151 420722 41217 420723
rect 41151 420658 41152 420722
rect 41216 420658 41217 420722
rect 41151 420657 41217 420658
rect 41154 403111 41214 420657
rect 41151 403110 41217 403111
rect 41151 403046 41152 403110
rect 41216 403046 41217 403110
rect 41151 403045 41217 403046
rect 41346 401927 41406 423173
rect 41535 421166 41601 421167
rect 41535 421102 41536 421166
rect 41600 421102 41601 421166
rect 41535 421101 41601 421102
rect 41538 402667 41598 421101
rect 41730 411251 41790 424357
rect 41919 422942 41985 422943
rect 41919 422878 41920 422942
rect 41984 422878 41985 422942
rect 41919 422877 41985 422878
rect 41727 411250 41793 411251
rect 41727 411186 41728 411250
rect 41792 411186 41793 411250
rect 41727 411185 41793 411186
rect 41922 406071 41982 422877
rect 42111 419390 42177 419391
rect 42111 419326 42112 419390
rect 42176 419326 42177 419390
rect 42111 419325 42177 419326
rect 41919 406070 41985 406071
rect 41919 406006 41920 406070
rect 41984 406006 41985 406070
rect 41919 406005 41985 406006
rect 42114 403851 42174 419325
rect 42111 403850 42177 403851
rect 42111 403786 42112 403850
rect 42176 403786 42177 403850
rect 42111 403785 42177 403786
rect 41535 402666 41601 402667
rect 41535 402602 41536 402666
rect 41600 402602 41601 402666
rect 41535 402601 41601 402602
rect 41343 401926 41409 401927
rect 41343 401862 41344 401926
rect 41408 401862 41409 401926
rect 41343 401861 41409 401862
rect 40959 399558 41025 399559
rect 40959 399494 40960 399558
rect 41024 399494 41025 399558
rect 40959 399493 41025 399494
rect 40767 398818 40833 398819
rect 40767 398754 40768 398818
rect 40832 398754 40833 398818
rect 40767 398753 40833 398754
rect 675903 398226 675969 398227
rect 675903 398162 675904 398226
rect 675968 398162 675969 398226
rect 675903 398161 675969 398162
rect 673983 397634 674049 397635
rect 673983 397570 673984 397634
rect 674048 397570 674049 397634
rect 673983 397569 674049 397570
rect 40383 382686 40449 382687
rect 40383 382622 40384 382686
rect 40448 382622 40449 382686
rect 40383 382621 40449 382622
rect 41727 382390 41793 382391
rect 41727 382326 41728 382390
rect 41792 382326 41793 382390
rect 41727 382325 41793 382326
rect 39807 381206 39873 381207
rect 39807 381142 39808 381206
rect 39872 381142 39873 381206
rect 39807 381141 39873 381142
rect 39810 373323 39870 381141
rect 39999 380318 40065 380319
rect 39999 380254 40000 380318
rect 40064 380254 40065 380318
rect 39999 380253 40065 380254
rect 40002 373659 40062 380253
rect 40575 378098 40641 378099
rect 40575 378034 40576 378098
rect 40640 378034 40641 378098
rect 40575 378033 40641 378034
rect 39999 373658 40065 373659
rect 39999 373594 40000 373658
rect 40064 373594 40065 373658
rect 39999 373593 40065 373594
rect 39810 373263 40446 373323
rect 40386 368183 40446 373263
rect 40383 368182 40449 368183
rect 40383 368118 40384 368182
rect 40448 368118 40449 368182
rect 40383 368117 40449 368118
rect 40578 359895 40638 378033
rect 40767 374250 40833 374251
rect 40767 374186 40768 374250
rect 40832 374186 40833 374250
rect 40767 374185 40833 374186
rect 40575 359894 40641 359895
rect 40575 359830 40576 359894
rect 40640 359830 40641 359894
rect 40575 359829 40641 359830
rect 40770 356195 40830 374185
rect 41535 373806 41601 373807
rect 41535 373742 41536 373806
rect 41600 373742 41601 373806
rect 41535 373741 41601 373742
rect 41343 373658 41409 373659
rect 41343 373594 41344 373658
rect 41408 373594 41409 373658
rect 41343 373593 41409 373594
rect 40959 372474 41025 372475
rect 40959 372410 40960 372474
rect 41024 372410 41025 372474
rect 40959 372409 41025 372410
rect 40962 356935 41022 372409
rect 41346 358859 41406 373593
rect 41538 362855 41598 373741
rect 41535 362854 41601 362855
rect 41535 362790 41536 362854
rect 41600 362790 41601 362854
rect 41535 362789 41601 362790
rect 41343 358858 41409 358859
rect 41343 358794 41344 358858
rect 41408 358794 41409 358858
rect 41343 358793 41409 358794
rect 40959 356934 41025 356935
rect 40959 356870 40960 356934
rect 41024 356870 41025 356934
rect 40959 356869 41025 356870
rect 40767 356194 40833 356195
rect 40767 356130 40768 356194
rect 40832 356130 40833 356194
rect 40767 356129 40833 356130
rect 39807 338286 39873 338287
rect 39807 338222 39808 338286
rect 39872 338222 39873 338286
rect 39807 338221 39873 338222
rect 39810 330739 39870 338221
rect 40383 337250 40449 337251
rect 40383 337186 40384 337250
rect 40448 337186 40449 337250
rect 40383 337185 40449 337186
rect 39807 330738 39873 330739
rect 39807 330674 39808 330738
rect 39872 330674 39873 330738
rect 39807 330673 39873 330674
rect 40386 328371 40446 337185
rect 40575 336806 40641 336807
rect 40575 336742 40576 336806
rect 40640 336742 40641 336806
rect 40575 336741 40641 336742
rect 40383 328370 40449 328371
rect 40383 328306 40384 328370
rect 40448 328306 40449 328370
rect 40383 328305 40449 328306
rect 40578 319787 40638 336741
rect 40959 335770 41025 335771
rect 40959 335706 40960 335770
rect 41024 335706 41025 335770
rect 40959 335705 41025 335706
rect 40767 331182 40833 331183
rect 40767 331118 40768 331182
rect 40832 331118 40833 331182
rect 40767 331117 40833 331118
rect 40575 319786 40641 319787
rect 40575 319722 40576 319786
rect 40640 319722 40641 319786
rect 40575 319721 40641 319722
rect 40770 312387 40830 331117
rect 40962 313127 41022 335705
rect 41151 335178 41217 335179
rect 41151 335114 41152 335178
rect 41216 335114 41217 335178
rect 41151 335113 41217 335114
rect 41154 316087 41214 335113
rect 41535 330738 41601 330739
rect 41535 330674 41536 330738
rect 41600 330674 41601 330738
rect 41535 330673 41601 330674
rect 41343 328370 41409 328371
rect 41343 328306 41344 328370
rect 41408 328306 41409 328370
rect 41343 328305 41409 328306
rect 41151 316086 41217 316087
rect 41151 316022 41152 316086
rect 41216 316022 41217 316086
rect 41151 316021 41217 316022
rect 41346 315643 41406 328305
rect 41538 324967 41598 330673
rect 41535 324966 41601 324967
rect 41535 324902 41536 324966
rect 41600 324902 41601 324966
rect 41535 324901 41601 324902
rect 41343 315642 41409 315643
rect 41343 315578 41344 315642
rect 41408 315578 41409 315642
rect 41343 315577 41409 315578
rect 40959 313126 41025 313127
rect 40959 313062 40960 313126
rect 41024 313062 41025 313126
rect 40959 313061 41025 313062
rect 40767 312386 40833 312387
rect 40767 312322 40768 312386
rect 40832 312322 40833 312386
rect 40767 312321 40833 312322
rect 41535 294922 41601 294923
rect 41535 294858 41536 294922
rect 41600 294858 41601 294922
rect 41535 294857 41601 294858
rect 40383 294034 40449 294035
rect 40383 293970 40384 294034
rect 40448 293970 40449 294034
rect 40383 293969 40449 293970
rect 40386 272279 40446 293969
rect 40959 292554 41025 292555
rect 40959 292490 40960 292554
rect 41024 292490 41025 292554
rect 40959 292489 41025 292490
rect 40575 290038 40641 290039
rect 40575 289974 40576 290038
rect 40640 289974 40641 290038
rect 40575 289973 40641 289974
rect 40578 274203 40638 289973
rect 40575 274202 40641 274203
rect 40575 274138 40576 274202
rect 40640 274138 40641 274202
rect 40575 274137 40641 274138
rect 40383 272278 40449 272279
rect 40383 272214 40384 272278
rect 40448 272214 40449 272278
rect 40383 272213 40449 272214
rect 40962 270059 41022 292489
rect 41151 292110 41217 292111
rect 41151 292046 41152 292110
rect 41216 292046 41217 292110
rect 41151 292045 41217 292046
rect 41154 272871 41214 292045
rect 41343 291518 41409 291519
rect 41343 291454 41344 291518
rect 41408 291454 41409 291518
rect 41343 291453 41409 291454
rect 41346 273611 41406 291453
rect 41538 281751 41598 294857
rect 41730 286077 41790 382325
rect 41919 376470 41985 376471
rect 41919 376406 41920 376470
rect 41984 376406 41985 376470
rect 41919 376405 41985 376406
rect 41922 360635 41982 376405
rect 673986 373955 674046 397569
rect 675135 396894 675201 396895
rect 675135 396830 675136 396894
rect 675200 396830 675201 396894
rect 675135 396829 675201 396830
rect 674943 396154 675009 396155
rect 674943 396090 674944 396154
rect 675008 396090 675009 396154
rect 674943 396089 675009 396090
rect 674367 393194 674433 393195
rect 674367 393130 674368 393194
rect 674432 393130 674433 393194
rect 674367 393129 674433 393130
rect 674175 391714 674241 391715
rect 674175 391650 674176 391714
rect 674240 391650 674241 391714
rect 674175 391649 674241 391650
rect 674178 376767 674238 391649
rect 674370 377211 674430 393129
rect 674946 378839 675006 396089
rect 675138 385943 675198 396829
rect 675711 395266 675777 395267
rect 675711 395202 675712 395266
rect 675776 395202 675777 395266
rect 675711 395201 675777 395202
rect 675327 394674 675393 394675
rect 675327 394610 675328 394674
rect 675392 394610 675393 394674
rect 675327 394609 675393 394610
rect 675135 385942 675201 385943
rect 675135 385878 675136 385942
rect 675200 385878 675201 385942
rect 675135 385877 675201 385878
rect 675330 382391 675390 394609
rect 675519 392602 675585 392603
rect 675519 392538 675520 392602
rect 675584 392538 675585 392602
rect 675519 392537 675585 392538
rect 675327 382390 675393 382391
rect 675327 382326 675328 382390
rect 675392 382326 675393 382390
rect 675327 382325 675393 382326
rect 675522 381207 675582 392537
rect 675714 385647 675774 395201
rect 675711 385646 675777 385647
rect 675711 385582 675712 385646
rect 675776 385582 675777 385646
rect 675711 385581 675777 385582
rect 675906 384907 675966 398161
rect 676671 396450 676737 396451
rect 676671 396386 676672 396450
rect 676736 396386 676737 396450
rect 676671 396385 676737 396386
rect 676479 393934 676545 393935
rect 676479 393870 676480 393934
rect 676544 393870 676545 393934
rect 676479 393869 676545 393870
rect 676287 393342 676353 393343
rect 676287 393278 676288 393342
rect 676352 393278 676353 393342
rect 676287 393277 676353 393278
rect 676095 391862 676161 391863
rect 676095 391798 676096 391862
rect 676160 391798 676161 391862
rect 676095 391797 676161 391798
rect 675903 384906 675969 384907
rect 675903 384842 675904 384906
rect 675968 384842 675969 384906
rect 675903 384841 675969 384842
rect 675519 381206 675585 381207
rect 675519 381142 675520 381206
rect 675584 381142 675585 381206
rect 675519 381141 675585 381142
rect 674943 378838 675009 378839
rect 674943 378774 674944 378838
rect 675008 378774 675009 378838
rect 674943 378773 675009 378774
rect 676098 378099 676158 391797
rect 676095 378098 676161 378099
rect 676095 378034 676096 378098
rect 676160 378034 676161 378098
rect 676095 378033 676161 378034
rect 674367 377210 674433 377211
rect 674367 377146 674368 377210
rect 674432 377146 674433 377210
rect 674367 377145 674433 377146
rect 674175 376766 674241 376767
rect 674175 376702 674176 376766
rect 674240 376702 674241 376766
rect 674175 376701 674241 376702
rect 676290 375731 676350 393277
rect 676482 381799 676542 393869
rect 676674 382983 676734 396385
rect 676671 382982 676737 382983
rect 676671 382918 676672 382982
rect 676736 382918 676737 382982
rect 676671 382917 676737 382918
rect 676479 381798 676545 381799
rect 676479 381734 676480 381798
rect 676544 381734 676545 381798
rect 676479 381733 676545 381734
rect 676287 375730 676353 375731
rect 676287 375666 676288 375730
rect 676352 375666 676353 375730
rect 676287 375665 676353 375666
rect 673983 373954 674049 373955
rect 673983 373890 673984 373954
rect 674048 373890 674049 373954
rect 673983 373889 674049 373890
rect 42111 373214 42177 373215
rect 42111 373150 42112 373214
rect 42176 373150 42177 373214
rect 42111 373149 42177 373150
rect 41919 360634 41985 360635
rect 41919 360570 41920 360634
rect 41984 360570 41985 360634
rect 41919 360569 41985 360570
rect 42114 359303 42174 373149
rect 42303 372770 42369 372771
rect 42303 372706 42304 372770
rect 42368 372706 42369 372770
rect 42303 372705 42369 372706
rect 42111 359302 42177 359303
rect 42111 359238 42112 359302
rect 42176 359238 42177 359302
rect 42111 359237 42177 359238
rect 42306 355751 42366 372705
rect 42303 355750 42369 355751
rect 42303 355686 42304 355750
rect 42368 355686 42369 355750
rect 42303 355685 42369 355686
rect 673983 355454 674049 355455
rect 673983 355390 673984 355454
rect 674048 355390 674049 355454
rect 673983 355389 674049 355390
rect 41919 334882 41985 334883
rect 41919 334818 41920 334882
rect 41984 334818 41985 334882
rect 41919 334817 41985 334818
rect 41922 316827 41982 334817
rect 42111 333402 42177 333403
rect 42111 333338 42112 333402
rect 42176 333338 42177 333402
rect 42111 333337 42177 333338
rect 42114 317419 42174 333337
rect 42495 332662 42561 332663
rect 42495 332598 42496 332662
rect 42560 332598 42561 332662
rect 42495 332597 42561 332598
rect 42303 329258 42369 329259
rect 42303 329194 42304 329258
rect 42368 329194 42369 329258
rect 42303 329193 42369 329194
rect 42111 317418 42177 317419
rect 42111 317354 42112 317418
rect 42176 317354 42177 317418
rect 42111 317353 42177 317354
rect 41919 316826 41985 316827
rect 41919 316762 41920 316826
rect 41984 316762 41985 316826
rect 41919 316761 41985 316762
rect 42306 313719 42366 329193
rect 42498 320527 42558 332597
rect 42495 320526 42561 320527
rect 42495 320462 42496 320526
rect 42560 320462 42561 320526
rect 42495 320461 42561 320462
rect 42303 313718 42369 313719
rect 42303 313654 42304 313718
rect 42368 313654 42369 313718
rect 42303 313653 42369 313654
rect 673986 311055 674046 355389
rect 674175 354566 674241 354567
rect 674175 354502 674176 354566
rect 674240 354502 674241 354566
rect 674175 354501 674241 354502
rect 673983 311054 674049 311055
rect 673983 310990 673984 311054
rect 674048 310990 674049 311054
rect 673983 310989 674049 310990
rect 674178 309871 674238 354501
rect 674367 353382 674433 353383
rect 674367 353318 674368 353382
rect 674432 353318 674433 353382
rect 674367 353317 674433 353318
rect 674175 309870 674241 309871
rect 674175 309806 674176 309870
rect 674240 309806 674241 309870
rect 674175 309805 674241 309806
rect 673983 306466 674049 306467
rect 673983 306402 673984 306466
rect 674048 306402 674049 306466
rect 673983 306401 674049 306402
rect 42303 294774 42369 294775
rect 42303 294710 42304 294774
rect 42368 294710 42369 294774
rect 42303 294709 42369 294710
rect 41919 293738 41985 293739
rect 41919 293674 41920 293738
rect 41984 293674 41985 293738
rect 41919 293673 41985 293674
rect 41922 287967 41982 293673
rect 41919 287966 41985 287967
rect 41919 287902 41920 287966
rect 41984 287902 41985 287966
rect 41919 287901 41985 287902
rect 41730 286017 42174 286077
rect 41727 285154 41793 285155
rect 41727 285090 41728 285154
rect 41792 285090 41793 285154
rect 41727 285089 41793 285090
rect 41535 281750 41601 281751
rect 41535 281686 41536 281750
rect 41600 281686 41601 281750
rect 41535 281685 41601 281686
rect 41343 273610 41409 273611
rect 41343 273546 41344 273610
rect 41408 273546 41409 273610
rect 41343 273545 41409 273546
rect 41151 272870 41217 272871
rect 41151 272806 41152 272870
rect 41216 272806 41217 272870
rect 41151 272805 41217 272806
rect 41730 270651 41790 285089
rect 41919 281602 41985 281603
rect 41919 281538 41920 281602
rect 41984 281538 41985 281602
rect 41919 281537 41985 281538
rect 41922 278051 41982 281537
rect 41919 278050 41985 278051
rect 41919 277986 41920 278050
rect 41984 277986 41985 278050
rect 41919 277985 41985 277986
rect 42114 274351 42174 286017
rect 42111 274350 42177 274351
rect 42111 274286 42112 274350
rect 42176 274286 42177 274350
rect 42111 274285 42177 274286
rect 41727 270650 41793 270651
rect 41727 270586 41728 270650
rect 41792 270586 41793 270650
rect 41727 270585 41793 270586
rect 40959 270058 41025 270059
rect 40959 269994 40960 270058
rect 41024 269994 41025 270058
rect 40959 269993 41025 269994
rect 42306 269319 42366 294709
rect 673986 292851 674046 306401
rect 673983 292850 674049 292851
rect 673983 292786 673984 292850
rect 674048 292786 674049 292850
rect 673983 292785 674049 292786
rect 42495 287966 42561 287967
rect 42495 287902 42496 287966
rect 42560 287902 42561 287966
rect 42495 287901 42561 287902
rect 42498 276571 42558 287901
rect 674178 278199 674238 309805
rect 674370 308983 674430 353317
rect 675711 353012 675777 353013
rect 675711 352948 675712 353012
rect 675776 352948 675777 353012
rect 675711 352947 675777 352948
rect 674559 351014 674625 351015
rect 674559 350950 674560 351014
rect 674624 350950 674625 351014
rect 674559 350949 674625 350950
rect 674562 333551 674622 350949
rect 675519 348498 675585 348499
rect 675519 348434 675520 348498
rect 675584 348434 675585 348498
rect 675519 348433 675585 348434
rect 674559 333550 674625 333551
rect 674559 333486 674560 333550
rect 674624 333486 674625 333550
rect 674559 333485 674625 333486
rect 675522 330591 675582 348433
rect 675714 339619 675774 352947
rect 675903 351458 675969 351459
rect 675903 351394 675904 351458
rect 675968 351394 675969 351458
rect 675903 351393 675969 351394
rect 675711 339618 675777 339619
rect 675711 339554 675712 339618
rect 675776 339554 675777 339618
rect 675711 339553 675777 339554
rect 675906 337843 675966 351393
rect 676479 343022 676545 343023
rect 676479 342958 676480 343022
rect 676544 342958 676545 343022
rect 676479 342957 676545 342958
rect 675903 337842 675969 337843
rect 675903 337778 675904 337842
rect 675968 337778 675969 337842
rect 675903 337777 675969 337778
rect 675519 330590 675585 330591
rect 675519 330526 675520 330590
rect 675584 330526 675585 330590
rect 675519 330525 675585 330526
rect 676482 326891 676542 342957
rect 676671 342874 676737 342875
rect 676671 342810 676672 342874
rect 676736 342810 676737 342874
rect 676671 342809 676737 342810
rect 676674 328075 676734 342809
rect 676671 328074 676737 328075
rect 676671 328010 676672 328074
rect 676736 328010 676737 328074
rect 676671 328009 676737 328010
rect 676479 326890 676545 326891
rect 676479 326826 676480 326890
rect 676544 326826 676545 326890
rect 676479 326825 676545 326826
rect 675327 310462 675393 310463
rect 675327 310398 675328 310462
rect 675392 310398 675393 310462
rect 675327 310397 675393 310398
rect 675135 309130 675201 309131
rect 675135 309066 675136 309130
rect 675200 309066 675201 309130
rect 675135 309065 675201 309066
rect 674367 308982 674433 308983
rect 674367 308918 674368 308982
rect 674432 308918 674433 308982
rect 674367 308917 674433 308918
rect 674559 307502 674625 307503
rect 674559 307438 674560 307502
rect 674624 307438 674625 307502
rect 674559 307437 674625 307438
rect 674562 283675 674622 307437
rect 674751 306022 674817 306023
rect 674751 305958 674752 306022
rect 674816 305958 674817 306022
rect 674751 305957 674817 305958
rect 674754 288559 674814 305957
rect 674943 302618 675009 302619
rect 674943 302554 674944 302618
rect 675008 302554 675009 302618
rect 674943 302553 675009 302554
rect 674751 288558 674817 288559
rect 674751 288494 674752 288558
rect 674816 288494 674817 288558
rect 674751 288493 674817 288494
rect 674946 287375 675006 302553
rect 674943 287374 675009 287375
rect 674943 287310 674944 287374
rect 675008 287310 675009 287374
rect 674943 287309 675009 287310
rect 674559 283674 674625 283675
rect 674559 283610 674560 283674
rect 674624 283610 674625 283674
rect 674559 283609 674625 283610
rect 675138 278495 675198 309065
rect 675135 278494 675201 278495
rect 675135 278430 675136 278494
rect 675200 278430 675201 278494
rect 675135 278429 675201 278430
rect 674175 278198 674241 278199
rect 674175 278134 674176 278198
rect 674240 278134 674241 278198
rect 674175 278133 674241 278134
rect 42495 276570 42561 276571
rect 42495 276506 42496 276570
rect 42560 276506 42561 276570
rect 42495 276505 42561 276506
rect 42303 269318 42369 269319
rect 42303 269254 42304 269318
rect 42368 269254 42369 269318
rect 42303 269253 42369 269254
rect 675330 266063 675390 310397
rect 675519 308390 675585 308391
rect 675519 308326 675520 308390
rect 675584 308326 675585 308390
rect 675519 308325 675585 308326
rect 675522 278347 675582 308325
rect 675711 299214 675777 299215
rect 675711 299150 675712 299214
rect 675776 299150 675777 299214
rect 675711 299149 675777 299150
rect 675714 285303 675774 299149
rect 676671 298770 676737 298771
rect 676671 298706 676672 298770
rect 676736 298706 676737 298770
rect 676671 298705 676737 298706
rect 675711 285302 675777 285303
rect 675711 285238 675712 285302
rect 675776 285238 675777 285302
rect 675711 285237 675777 285238
rect 676674 281899 676734 298705
rect 676671 281898 676737 281899
rect 676671 281834 676672 281898
rect 676736 281834 676737 281898
rect 676671 281833 676737 281834
rect 675519 278346 675585 278347
rect 675519 278282 675520 278346
rect 675584 278282 675585 278346
rect 675519 278281 675585 278282
rect 675327 266062 675393 266063
rect 675327 265998 675328 266062
rect 675392 265998 675393 266062
rect 675327 265997 675393 265998
rect 673983 265470 674049 265471
rect 673983 265406 673984 265470
rect 674048 265406 674049 265470
rect 673983 265405 674049 265406
rect 40767 252298 40833 252299
rect 40767 252234 40768 252298
rect 40832 252234 40833 252298
rect 40767 252233 40833 252234
rect 40575 251706 40641 251707
rect 40575 251642 40576 251706
rect 40640 251642 40641 251706
rect 40575 251641 40641 251642
rect 40383 246822 40449 246823
rect 40383 246758 40384 246822
rect 40448 246758 40449 246822
rect 40383 246757 40449 246758
rect 40386 231135 40446 246757
rect 40383 231134 40449 231135
rect 40383 231070 40384 231134
rect 40448 231070 40449 231134
rect 40383 231069 40449 231070
rect 40578 225955 40638 251641
rect 40770 237203 40830 252233
rect 41727 252076 41793 252077
rect 41727 252012 41728 252076
rect 41792 252012 41793 252076
rect 41727 252011 41793 252012
rect 40959 250818 41025 250819
rect 40959 250754 40960 250818
rect 41024 250754 41025 250818
rect 40959 250753 41025 250754
rect 40767 237202 40833 237203
rect 40767 237138 40768 237202
rect 40832 237138 40833 237202
rect 40767 237137 40833 237138
rect 40962 229063 41022 250753
rect 41535 250374 41601 250375
rect 41535 250310 41536 250374
rect 41600 250310 41601 250374
rect 41535 250309 41601 250310
rect 41151 248894 41217 248895
rect 41151 248830 41152 248894
rect 41216 248830 41217 248894
rect 41151 248829 41217 248830
rect 41154 229655 41214 248829
rect 41343 248302 41409 248303
rect 41343 248238 41344 248302
rect 41408 248238 41409 248302
rect 41343 248237 41409 248238
rect 41346 230395 41406 248237
rect 41538 237459 41598 250309
rect 41730 237943 41790 252011
rect 41919 249634 41985 249635
rect 41919 249570 41920 249634
rect 41984 249570 41985 249634
rect 41919 249569 41985 249570
rect 41727 237942 41793 237943
rect 41727 237878 41728 237942
rect 41792 237878 41793 237942
rect 41727 237877 41793 237878
rect 41538 237399 41790 237459
rect 41535 237202 41601 237203
rect 41535 237138 41536 237202
rect 41600 237138 41601 237202
rect 41535 237137 41601 237138
rect 41343 230394 41409 230395
rect 41343 230330 41344 230394
rect 41408 230330 41409 230394
rect 41343 230329 41409 230330
rect 41151 229654 41217 229655
rect 41151 229590 41152 229654
rect 41216 229590 41217 229654
rect 41151 229589 41217 229590
rect 40959 229062 41025 229063
rect 40959 228998 40960 229062
rect 41024 228998 41025 229062
rect 40959 228997 41025 228998
rect 41538 227435 41598 237137
rect 41730 233355 41790 237399
rect 41727 233354 41793 233355
rect 41727 233290 41728 233354
rect 41792 233290 41793 233354
rect 41727 233289 41793 233290
rect 41535 227434 41601 227435
rect 41535 227370 41536 227434
rect 41600 227370 41601 227434
rect 41535 227369 41601 227370
rect 41922 226843 41982 249569
rect 408642 236759 409086 236793
rect 408642 236758 409089 236759
rect 408642 236733 409024 236758
rect 408642 236167 408702 236733
rect 409023 236694 409024 236733
rect 409088 236694 409089 236758
rect 409023 236693 409089 236694
rect 408639 236166 408705 236167
rect 408639 236102 408640 236166
rect 408704 236102 408705 236166
rect 408639 236101 408705 236102
rect 409023 235870 409089 235871
rect 409023 235806 409024 235870
rect 409088 235806 409089 235870
rect 409023 235805 409089 235806
rect 409026 235461 409086 235805
rect 408450 235401 409086 235461
rect 408450 235131 408510 235401
rect 408447 235130 408513 235131
rect 408447 235066 408448 235130
rect 408512 235066 408513 235130
rect 408447 235065 408513 235066
rect 41919 226842 41985 226843
rect 41919 226778 41920 226842
rect 41984 226778 41985 226842
rect 41919 226777 41985 226778
rect 40575 225954 40641 225955
rect 40575 225890 40576 225954
rect 40640 225890 40641 225954
rect 40575 225889 40641 225890
rect 673986 220775 674046 265405
rect 676287 261770 676353 261771
rect 676287 261706 676288 261770
rect 676352 261706 676353 261770
rect 676287 261705 676353 261706
rect 675711 261030 675777 261031
rect 675711 260966 675712 261030
rect 675776 260966 675777 261030
rect 675711 260965 675777 260966
rect 675519 258958 675585 258959
rect 675519 258894 675520 258958
rect 675584 258894 675585 258958
rect 675519 258893 675585 258894
rect 674943 258514 675009 258515
rect 674943 258450 674944 258514
rect 675008 258450 675009 258514
rect 674943 258449 675009 258450
rect 674559 257922 674625 257923
rect 674559 257858 674560 257922
rect 674624 257858 674625 257922
rect 674559 257857 674625 257858
rect 674562 242087 674622 257857
rect 674751 256442 674817 256443
rect 674751 256378 674752 256442
rect 674816 256378 674817 256442
rect 674751 256377 674817 256378
rect 674559 242086 674625 242087
rect 674559 242022 674560 242086
rect 674624 242022 674625 242086
rect 674559 242021 674625 242022
rect 674754 241791 674814 256377
rect 674751 241790 674817 241791
rect 674751 241726 674752 241790
rect 674816 241726 674817 241790
rect 674751 241725 674817 241726
rect 674946 240607 675006 258449
rect 675522 246675 675582 258893
rect 675519 246674 675585 246675
rect 675519 246610 675520 246674
rect 675584 246610 675585 246674
rect 675519 246609 675585 246610
rect 675714 243567 675774 260965
rect 675903 253334 675969 253335
rect 675903 253270 675904 253334
rect 675968 253270 675969 253334
rect 675903 253269 675969 253270
rect 675711 243566 675777 243567
rect 675711 243502 675712 243566
rect 675776 243502 675777 243566
rect 675711 243501 675777 243502
rect 674943 240606 675009 240607
rect 674943 240542 674944 240606
rect 675008 240542 675009 240606
rect 674943 240541 675009 240542
rect 675906 236907 675966 253269
rect 676095 253186 676161 253187
rect 676095 253122 676096 253186
rect 676160 253122 676161 253186
rect 676095 253121 676161 253122
rect 676098 238683 676158 253121
rect 676290 250819 676350 261705
rect 676287 250818 676353 250819
rect 676287 250754 676288 250818
rect 676352 250754 676353 250818
rect 676287 250753 676353 250754
rect 676095 238682 676161 238683
rect 676095 238618 676096 238682
rect 676160 238618 676161 238682
rect 676095 238617 676161 238618
rect 675903 236906 675969 236907
rect 675903 236842 675904 236906
rect 675968 236842 675969 236906
rect 675903 236841 675969 236842
rect 673983 220774 674049 220775
rect 673983 220710 673984 220774
rect 674048 220710 674049 220774
rect 673983 220709 674049 220710
rect 674367 220034 674433 220035
rect 674367 219970 674368 220034
rect 674432 219970 674433 220034
rect 674367 219969 674433 219970
rect 673983 219294 674049 219295
rect 673983 219230 673984 219294
rect 674048 219230 674049 219294
rect 673983 219229 674049 219230
rect 41151 205974 41217 205975
rect 41151 205910 41152 205974
rect 41216 205910 41217 205974
rect 41151 205909 41217 205910
rect 40767 204938 40833 204939
rect 40767 204874 40768 204938
rect 40832 204874 40833 204938
rect 40767 204873 40833 204874
rect 40770 187179 40830 204873
rect 40959 201534 41025 201535
rect 40959 201470 40960 201534
rect 41024 201470 41025 201534
rect 40959 201469 41025 201470
rect 40767 187178 40833 187179
rect 40767 187114 40768 187178
rect 40832 187114 40833 187178
rect 40767 187113 40833 187114
rect 40962 185847 41022 201469
rect 41154 189507 41214 205909
rect 41343 205382 41409 205383
rect 41343 205318 41344 205382
rect 41408 205318 41409 205382
rect 41343 205317 41409 205318
rect 41346 189695 41406 205317
rect 41919 203606 41985 203607
rect 41919 203542 41920 203606
rect 41984 203542 41985 203606
rect 41919 203541 41985 203542
rect 41727 200942 41793 200943
rect 41727 200878 41728 200942
rect 41792 200878 41793 200942
rect 41727 200877 41793 200878
rect 41535 199758 41601 199759
rect 41535 199694 41536 199758
rect 41600 199694 41601 199758
rect 41535 199693 41601 199694
rect 41538 190139 41598 199693
rect 41730 195319 41790 200877
rect 41727 195318 41793 195319
rect 41727 195254 41728 195318
rect 41792 195254 41793 195318
rect 41727 195253 41793 195254
rect 41535 190138 41601 190139
rect 41535 190074 41536 190138
rect 41600 190074 41601 190138
rect 41535 190073 41601 190074
rect 41343 189694 41409 189695
rect 41343 189630 41344 189694
rect 41408 189630 41409 189694
rect 41343 189629 41409 189630
rect 41154 189447 41598 189507
rect 41343 189250 41409 189251
rect 41343 189186 41344 189250
rect 41408 189186 41409 189250
rect 41343 189185 41409 189186
rect 41346 186735 41406 189185
rect 41538 187230 41598 189447
rect 41922 187919 41982 203541
rect 42303 200794 42369 200795
rect 42303 200730 42304 200794
rect 42368 200730 42369 200794
rect 42303 200729 42369 200730
rect 42111 200054 42177 200055
rect 42111 199990 42112 200054
rect 42176 199990 42177 200054
rect 42111 199989 42177 199990
rect 41919 187918 41985 187919
rect 41919 187854 41920 187918
rect 41984 187854 41985 187918
rect 41919 187853 41985 187854
rect 41538 187170 41982 187230
rect 41343 186734 41409 186735
rect 41343 186670 41344 186734
rect 41408 186670 41409 186734
rect 41343 186669 41409 186670
rect 40959 185846 41025 185847
rect 40959 185782 40960 185846
rect 41024 185782 41025 185846
rect 40959 185781 41025 185782
rect 41922 183627 41982 187170
rect 41919 183626 41985 183627
rect 41919 183562 41920 183626
rect 41984 183562 41985 183626
rect 41919 183561 41985 183562
rect 42114 182887 42174 199989
rect 42306 184219 42366 200729
rect 42303 184218 42369 184219
rect 42303 184154 42304 184218
rect 42368 184154 42369 184218
rect 42303 184153 42369 184154
rect 42111 182886 42177 182887
rect 42111 182822 42112 182886
rect 42176 182822 42177 182886
rect 42111 182821 42177 182822
rect 673986 175487 674046 219229
rect 674175 218258 674241 218259
rect 674175 218194 674176 218258
rect 674240 218194 674241 218258
rect 674175 218193 674241 218194
rect 673983 175486 674049 175487
rect 673983 175422 673984 175486
rect 674048 175422 674049 175486
rect 673983 175421 674049 175422
rect 674178 174155 674238 218193
rect 674370 176227 674430 219969
rect 675903 217814 675969 217815
rect 675903 217750 675904 217814
rect 675968 217750 675969 217814
rect 675903 217749 675969 217750
rect 675711 216334 675777 216335
rect 675711 216270 675712 216334
rect 675776 216270 675777 216334
rect 675711 216269 675777 216270
rect 675519 215742 675585 215743
rect 675519 215678 675520 215742
rect 675584 215678 675585 215742
rect 675519 215677 675585 215678
rect 675522 198427 675582 215677
rect 675714 202719 675774 216269
rect 675906 204495 675966 217749
rect 676287 207750 676353 207751
rect 676287 207686 676288 207750
rect 676352 207686 676353 207750
rect 676287 207685 676353 207686
rect 675903 204494 675969 204495
rect 675903 204430 675904 204494
rect 675968 204430 675969 204494
rect 675903 204429 675969 204430
rect 675711 202718 675777 202719
rect 675711 202654 675712 202718
rect 675776 202654 675777 202718
rect 675711 202653 675777 202654
rect 675519 198426 675585 198427
rect 675519 198362 675520 198426
rect 675584 198362 675585 198426
rect 675519 198361 675585 198362
rect 676290 193543 676350 207685
rect 676671 207602 676737 207603
rect 676671 207538 676672 207602
rect 676736 207538 676737 207602
rect 676671 207537 676737 207538
rect 676479 207454 676545 207455
rect 676479 207390 676480 207454
rect 676544 207390 676545 207454
rect 676479 207389 676545 207390
rect 676482 195319 676542 207389
rect 676479 195318 676545 195319
rect 676479 195254 676480 195318
rect 676544 195254 676545 195318
rect 676479 195253 676545 195254
rect 676287 193542 676353 193543
rect 676287 193478 676288 193542
rect 676352 193478 676353 193542
rect 676287 193477 676353 193478
rect 676674 191619 676734 207537
rect 676671 191618 676737 191619
rect 676671 191554 676672 191618
rect 676736 191554 676737 191618
rect 676671 191553 676737 191554
rect 674367 176226 674433 176227
rect 674367 176162 674368 176226
rect 674432 176162 674433 176226
rect 674367 176161 674433 176162
rect 674367 175634 674433 175635
rect 674367 175570 674368 175634
rect 674432 175570 674433 175634
rect 674367 175569 674433 175570
rect 674175 174154 674241 174155
rect 674175 174090 674176 174154
rect 674240 174090 674241 174154
rect 674175 174089 674241 174090
rect 674175 174006 674241 174007
rect 674175 173942 674176 174006
rect 674240 173942 674241 174006
rect 674175 173941 674241 173942
rect 673983 173562 674049 173563
rect 673983 173498 673984 173562
rect 674048 173498 674049 173562
rect 673983 173497 674049 173498
rect 673986 128571 674046 173497
rect 674178 129459 674238 173941
rect 674370 130643 674430 175569
rect 675903 173266 675969 173267
rect 675903 173202 675904 173266
rect 675968 173202 675969 173266
rect 675903 173201 675969 173202
rect 675135 171194 675201 171195
rect 675135 171130 675136 171194
rect 675200 171130 675201 171194
rect 675135 171129 675201 171130
rect 674751 168678 674817 168679
rect 674751 168614 674752 168678
rect 674816 168614 674817 168678
rect 674751 168613 674817 168614
rect 674559 167198 674625 167199
rect 674559 167134 674560 167198
rect 674624 167134 674625 167198
rect 674559 167133 674625 167134
rect 674562 152547 674622 167133
rect 674559 152546 674625 152547
rect 674559 152482 674560 152546
rect 674624 152482 674625 152546
rect 674559 152481 674625 152482
rect 674754 150327 674814 168613
rect 674943 168234 675009 168235
rect 674943 168170 674944 168234
rect 675008 168170 675009 168234
rect 674943 168169 675009 168170
rect 674946 152251 675006 168169
rect 675138 153435 675198 171129
rect 675711 161574 675777 161575
rect 675711 161510 675712 161574
rect 675776 161510 675777 161574
rect 675711 161509 675777 161510
rect 675135 153434 675201 153435
rect 675135 153370 675136 153434
rect 675200 153370 675201 153434
rect 675135 153369 675201 153370
rect 674943 152250 675009 152251
rect 674943 152186 674944 152250
rect 675008 152186 675009 152250
rect 674943 152185 675009 152186
rect 674751 150326 674817 150327
rect 674751 150262 674752 150326
rect 674816 150262 674817 150326
rect 674751 150261 674817 150262
rect 675714 148551 675774 161509
rect 675906 159355 675966 173201
rect 676671 161426 676737 161427
rect 676671 161362 676672 161426
rect 676736 161362 676737 161426
rect 676671 161361 676737 161362
rect 675903 159354 675969 159355
rect 675903 159290 675904 159354
rect 675968 159290 675969 159354
rect 675903 159289 675969 159290
rect 675711 148550 675777 148551
rect 675711 148486 675712 148550
rect 675776 148486 675777 148550
rect 675711 148485 675777 148486
rect 676674 146627 676734 161361
rect 676671 146626 676737 146627
rect 676671 146562 676672 146626
rect 676736 146562 676737 146626
rect 676671 146561 676737 146562
rect 674367 130642 674433 130643
rect 674367 130578 674368 130642
rect 674432 130578 674433 130642
rect 674367 130577 674433 130578
rect 674175 129458 674241 129459
rect 674175 129394 674176 129458
rect 674240 129394 674241 129458
rect 674175 129393 674241 129394
rect 673983 128570 674049 128571
rect 673983 128506 673984 128570
rect 674048 128506 674049 128570
rect 673983 128505 674049 128506
rect 674367 125610 674433 125611
rect 674367 125546 674368 125610
rect 674432 125546 674433 125610
rect 674367 125545 674433 125546
rect 673983 122206 674049 122207
rect 673983 122142 673984 122206
rect 674048 122142 674049 122206
rect 673983 122141 674049 122142
rect 673986 106667 674046 122141
rect 674370 108147 674430 125545
rect 674559 123094 674625 123095
rect 674559 123030 674560 123094
rect 674624 123030 674625 123094
rect 674559 123029 674625 123030
rect 674367 108146 674433 108147
rect 674367 108082 674368 108146
rect 674432 108082 674433 108146
rect 674367 108081 674433 108082
rect 673983 106666 674049 106667
rect 673983 106602 673984 106666
rect 674048 106602 674049 106666
rect 673983 106601 674049 106602
rect 674562 105187 674622 123029
rect 676479 118062 676545 118063
rect 676479 117998 676480 118062
rect 676544 117998 676545 118062
rect 676479 117997 676545 117998
rect 675903 117914 675969 117915
rect 675903 117850 675904 117914
rect 675968 117850 675969 117914
rect 675903 117849 675969 117850
rect 674559 105186 674625 105187
rect 674559 105122 674560 105186
rect 674624 105122 674625 105186
rect 674559 105121 674625 105122
rect 675906 103263 675966 117849
rect 675903 103262 675969 103263
rect 675903 103198 675904 103262
rect 675968 103198 675969 103262
rect 675903 103197 675969 103198
rect 676482 101487 676542 117997
rect 676479 101486 676545 101487
rect 676479 101422 676480 101486
rect 676544 101422 676545 101486
rect 676479 101421 676545 101422
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 283410 1018624 295578 1030788
rect 334810 1018624 346978 1030788
rect 385210 1018624 397378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 955022 710788 967190
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876180
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786620 19088 799160
rect 698512 774440 711002 786980
rect 6598 743420 19088 755960
rect 698512 729440 711002 741980
rect 6598 700220 19088 712760
rect 698512 684440 711002 696980
rect 6598 657020 19088 669560
rect 698512 639240 711002 651780
rect 6598 613820 19088 626360
rect 698512 594240 711002 606780
rect 6598 570620 19088 583160
rect 698512 549040 711002 561580
rect 6598 527420 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399820 19088 412360
rect 698512 371840 711002 384380
rect 6598 356620 19088 369160
rect 698512 326640 711002 339180
rect 6598 313420 19088 325960
rect 6598 270220 19088 282760
rect 698512 281640 711002 294180
rect 6598 227020 19088 239560
rect 698512 236640 711002 249180
rect 6598 183820 19088 196360
rect 698512 191440 711002 203980
rect 698512 146440 711002 158980
rect 6811 111610 18975 123778
rect 698512 101240 711002 113780
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use user_id_programming  user_id_value
timestamp 1625156099
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use storage  storage
timestamp 1625156099
transform 1 0 52032 0 1 53156
box 1066 70 92000 191480
use mgmt_core  soc
timestamp 1625156099
transform 1 0 190434 0 1 53602
box 0 0 450000 168026
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1625156099
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1625156099
transform 1 0 654146 0 -1 112882
box 25 11 11344 8291
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1625156099
transform -1 0 710203 0 1 164000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1625156099
transform -1 0 710203 0 1 118400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1625156099
transform 1 0 7631 0 1 243400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1625156099
transform 1 0 7631 0 1 200000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1625156099
transform 1 0 7631 0 1 286600
box -1620 -364 34000 13964
use mgmt_protect  mgmt_buffers
timestamp 1625156099
transform 1 0 192180 0 1 240036
box -2762 -2778 222734 26170
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1625156099
transform -1 0 710203 0 1 208600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1625156099
transform -1 0 710203 0 1 253800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1625156099
transform 1 0 7631 0 1 372800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1625156099
transform 1 0 7631 0 1 329800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1625156099
transform -1 0 710203 0 1 298800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1625156099
transform -1 0 710203 0 1 343800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1625156099
transform 1 0 7631 0 1 415800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1625156099
transform -1 0 710203 0 1 477200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1625156099
transform -1 0 710203 0 1 389000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1625156099
transform 1 0 7631 0 1 529600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1625156099
transform 1 0 7631 0 1 586824
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1625156099
transform 1 0 7631 0 1 630000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1625156099
transform 1 0 7631 0 1 673200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1625156099
transform -1 0 710203 0 1 655400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1625156099
transform -1 0 710203 0 1 611800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1625156099
transform -1 0 710203 0 1 566400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1625156099
transform -1 0 710203 0 1 521600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1625156099
transform 1 0 7631 0 1 716800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1625156099
transform 1 0 7631 0 1 759800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1625156099
transform 1 0 7631 0 1 803000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1625156099
transform -1 0 710203 0 1 702000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1625156099
transform -1 0 710203 0 1 880800
box -1620 -364 34000 13964
use user_analog_project_wrapper  mprj
timestamp 1625156099
transform 1 0 65308 0 1 278718
box -800 -800 584800 704000
use chip_io_alt  padframe
timestamp 1625156099
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113780 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696980 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741980 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786980 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876180 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 385210 1018624 397378 1030788 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 698624 955022 710788 967190 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030788 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030788 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030788 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 283410 1018624 295578 1030788 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158980 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231810 1018624 243978 1030788 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030788 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030788 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030788 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 956610 18975 968778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786620 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743420 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700220 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657020 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613820 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203980 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570620 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527420 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399820 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356620 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313420 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270220 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227020 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183820 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249180 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294180 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339180 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384380 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561580 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606780 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651780 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 697980 909666 711432 920546 6 vccd1
port 45 nsew signal bidirectional
rlabel metal5 s 6167 914054 19619 924934 6 vccd2
port 46 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda
port 47 nsew signal bidirectional
rlabel metal5 s 698624 819822 710788 831990 6 vdda1
port 48 nsew signal bidirectional
rlabel metal5 s 698624 505222 710788 517390 6 vdda1_2
port 49 nsew signal bidirectional
rlabel metal5 s 6811 484410 18975 496578 6 vdda2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 871210 18975 883378 6 vddio_2
port 51 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1
port 52 nsew signal bidirectional
rlabel metal5 s 698624 417022 710788 429190 6 vssa1_2
port 53 nsew signal bidirectional
rlabel metal5 s 6811 829010 18975 841178 6 vssa2
port 54 nsew signal bidirectional
rlabel metal5 s 697980 461866 711432 472746 6 vssd1
port 55 nsew signal bidirectional
rlabel metal5 s 6167 442854 19619 453734 6 vssd2
port 56 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030788 6 vssio_2
port 57 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio
port 58 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio
port 59 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa
port 60 nsew signal bidirectional
rlabel metal5 s 6167 70054 19619 80934 6 vccd
port 61 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd
port 62 nsew signal bidirectional
rlabel metal2 s 579796 53602 579852 54402 6 pwr_ctrl_out[0]
port 63 nsew signal tristate
rlabel metal2 s 597092 53602 597148 54402 6 pwr_ctrl_out[1]
port 64 nsew signal tristate
rlabel metal2 s 614388 53602 614444 54402 6 pwr_ctrl_out[2]
port 65 nsew signal tristate
rlabel metal2 s 631684 53602 631740 54402 6 pwr_ctrl_out[3]
port 66 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
