* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[45] HI[46] HI[47] HI[48] HI[49] HI[4]
+ HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58] HI[59] HI[5] HI[60]
+ HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69] HI[6] HI[70] HI[71]
+ HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7] HI[80] HI[81] HI[82]
+ HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90] HI[91] HI[92] HI[93]
+ HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_oen_core[0] la_oen_core[100] la_oen_core[101] la_oen_core[102]
+ la_oen_core[103] la_oen_core[104] la_oen_core[105] la_oen_core[106] la_oen_core[107]
+ la_oen_core[108] la_oen_core[109] la_oen_core[10] la_oen_core[110] la_oen_core[111]
+ la_oen_core[112] la_oen_core[113] la_oen_core[114] la_oen_core[115] la_oen_core[116]
+ la_oen_core[117] la_oen_core[118] la_oen_core[119] la_oen_core[11] la_oen_core[120]
+ la_oen_core[121] la_oen_core[122] la_oen_core[123] la_oen_core[124] la_oen_core[125]
+ la_oen_core[126] la_oen_core[127] la_oen_core[12] la_oen_core[13] la_oen_core[14]
+ la_oen_core[15] la_oen_core[16] la_oen_core[17] la_oen_core[18] la_oen_core[19]
+ la_oen_core[1] la_oen_core[20] la_oen_core[21] la_oen_core[22] la_oen_core[23] la_oen_core[24]
+ la_oen_core[25] la_oen_core[26] la_oen_core[27] la_oen_core[28] la_oen_core[29]
+ la_oen_core[2] la_oen_core[30] la_oen_core[31] la_oen_core[32] la_oen_core[33] la_oen_core[34]
+ la_oen_core[35] la_oen_core[36] la_oen_core[37] la_oen_core[38] la_oen_core[39]
+ la_oen_core[3] la_oen_core[40] la_oen_core[41] la_oen_core[42] la_oen_core[43] la_oen_core[44]
+ la_oen_core[45] la_oen_core[46] la_oen_core[47] la_oen_core[48] la_oen_core[49]
+ la_oen_core[4] la_oen_core[50] la_oen_core[51] la_oen_core[52] la_oen_core[53] la_oen_core[54]
+ la_oen_core[55] la_oen_core[56] la_oen_core[57] la_oen_core[58] la_oen_core[59]
+ la_oen_core[5] la_oen_core[60] la_oen_core[61] la_oen_core[62] la_oen_core[63] la_oen_core[64]
+ la_oen_core[65] la_oen_core[66] la_oen_core[67] la_oen_core[68] la_oen_core[69]
+ la_oen_core[6] la_oen_core[70] la_oen_core[71] la_oen_core[72] la_oen_core[73] la_oen_core[74]
+ la_oen_core[75] la_oen_core[76] la_oen_core[77] la_oen_core[78] la_oen_core[79]
+ la_oen_core[7] la_oen_core[80] la_oen_core[81] la_oen_core[82] la_oen_core[83] la_oen_core[84]
+ la_oen_core[85] la_oen_core[86] la_oen_core[87] la_oen_core[88] la_oen_core[89]
+ la_oen_core[8] la_oen_core[90] la_oen_core[91] la_oen_core[92] la_oen_core[93] la_oen_core[94]
+ la_oen_core[95] la_oen_core[96] la_oen_core[97] la_oen_core[98] la_oen_core[99]
+ la_oen_core[9] la_oen_mprj[0] la_oen_mprj[100] la_oen_mprj[101] la_oen_mprj[102]
+ la_oen_mprj[103] la_oen_mprj[104] la_oen_mprj[105] la_oen_mprj[106] la_oen_mprj[107]
+ la_oen_mprj[108] la_oen_mprj[109] la_oen_mprj[10] la_oen_mprj[110] la_oen_mprj[111]
+ la_oen_mprj[112] la_oen_mprj[113] la_oen_mprj[114] la_oen_mprj[115] la_oen_mprj[116]
+ la_oen_mprj[117] la_oen_mprj[118] la_oen_mprj[119] la_oen_mprj[11] la_oen_mprj[120]
+ la_oen_mprj[121] la_oen_mprj[122] la_oen_mprj[123] la_oen_mprj[124] la_oen_mprj[125]
+ la_oen_mprj[126] la_oen_mprj[127] la_oen_mprj[12] la_oen_mprj[13] la_oen_mprj[14]
+ la_oen_mprj[15] la_oen_mprj[16] la_oen_mprj[17] la_oen_mprj[18] la_oen_mprj[19]
+ la_oen_mprj[1] la_oen_mprj[20] la_oen_mprj[21] la_oen_mprj[22] la_oen_mprj[23] la_oen_mprj[24]
+ la_oen_mprj[25] la_oen_mprj[26] la_oen_mprj[27] la_oen_mprj[28] la_oen_mprj[29]
+ la_oen_mprj[2] la_oen_mprj[30] la_oen_mprj[31] la_oen_mprj[32] la_oen_mprj[33] la_oen_mprj[34]
+ la_oen_mprj[35] la_oen_mprj[36] la_oen_mprj[37] la_oen_mprj[38] la_oen_mprj[39]
+ la_oen_mprj[3] la_oen_mprj[40] la_oen_mprj[41] la_oen_mprj[42] la_oen_mprj[43] la_oen_mprj[44]
+ la_oen_mprj[45] la_oen_mprj[46] la_oen_mprj[47] la_oen_mprj[48] la_oen_mprj[49]
+ la_oen_mprj[4] la_oen_mprj[50] la_oen_mprj[51] la_oen_mprj[52] la_oen_mprj[53] la_oen_mprj[54]
+ la_oen_mprj[55] la_oen_mprj[56] la_oen_mprj[57] la_oen_mprj[58] la_oen_mprj[59]
+ la_oen_mprj[5] la_oen_mprj[60] la_oen_mprj[61] la_oen_mprj[62] la_oen_mprj[63] la_oen_mprj[64]
+ la_oen_mprj[65] la_oen_mprj[66] la_oen_mprj[67] la_oen_mprj[68] la_oen_mprj[69]
+ la_oen_mprj[6] la_oen_mprj[70] la_oen_mprj[71] la_oen_mprj[72] la_oen_mprj[73] la_oen_mprj[74]
+ la_oen_mprj[75] la_oen_mprj[76] la_oen_mprj[77] la_oen_mprj[78] la_oen_mprj[79]
+ la_oen_mprj[7] la_oen_mprj[80] la_oen_mprj[81] la_oen_mprj[82] la_oen_mprj[83] la_oen_mprj[84]
+ la_oen_mprj[85] la_oen_mprj[86] la_oen_mprj[87] la_oen_mprj[88] la_oen_mprj[89]
+ la_oen_mprj[8] la_oen_mprj[90] la_oen_mprj[91] la_oen_mprj[92] la_oen_mprj[93] la_oen_mprj[94]
+ la_oen_mprj[95] la_oen_mprj[96] la_oen_mprj[97] la_oen_mprj[98] la_oen_mprj[99]
+ la_oen_mprj[9] mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12]
+ mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16]
+ mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20]
+ mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24]
+ mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28]
+ mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3]
+ mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8]
+ mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12]
+ mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16]
+ mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20]
+ mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24]
+ mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28]
+ mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3]
+ mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8]
+ mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10]
+ mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14]
+ mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18]
+ mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22]
+ mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26]
+ mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30]
+ mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6]
+ mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10]
+ mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14]
+ mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18]
+ mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22]
+ mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26]
+ mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30]
+ mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6]
+ mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user1_vcc_powergood user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood
+ user_clock user_clock2 user_reset user_resetn vccd vssd vccd1 vssd1 vccd2 vssd2
+ vdda1 vssa1 vdda2 vssa2
XFILLER_27_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_501_ la_data_out_mprj[30] vssd vssd vccd vccd _501_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_432_ mprj_adr_o_core[25] vssd vssd vccd vccd _432_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_363_ la_oen_mprj[95] vssd vssd vccd vccd _363_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[36\] _507_/Y la_buf\[36\]/TE vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_9_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] mprj_logic_high_inst/HI[355] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[76\] _344_/Y mprj_logic_high_inst/HI[278] vssd vssd vccd
+ vccd la_oen_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_8_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[24\] _463_/Y mprj_dat_buf\[24\]/TE vssd vssd vccd vccd mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_415_ mprj_adr_o_core[8] vssd vssd vccd vccd _415_/Y sky130_fd_sc_hd__inv_2
X_346_ la_oen_mprj[78] vssd vssd vccd vccd _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] mprj_logic_high_inst/HI[422] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[109\] _377_/Y mprj_logic_high_inst/HI[311] vssd vssd vccd
+ vccd la_oen_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_28_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[39\] _638_/Y mprj_logic_high_inst/HI[241] vssd vssd vccd
+ vccd la_oen_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_18_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__402__A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vssd vccd vccd la_data_in_mprj[62]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_594_ la_data_out_mprj[123] vssd vssd vccd vccd _594_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[66\] _537_/Y la_buf\[66\]/TE vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__einvp_8
XPHY_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _593_/Y la_buf\[122\]/TE vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[70\]_B mprj_logic_high_inst/HI[400] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] mprj_logic_high_inst/HI[385] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[61\]_B mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_B mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_646_ la_oen_mprj[47] vssd vssd vccd vccd _646_/Y sky130_fd_sc_hd__inv_2
X_577_ la_data_out_mprj[106] vssd vssd vccd vccd _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[6\]_A _445_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vssd vccd vccd la_data_in_mprj[25]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[43\]_B mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[112\]_TE la_buf\[112\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_178 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[34\]_B mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__500__A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_500_ la_data_out_mprj[29] vssd vssd vccd vccd _500_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[3\] _602_/Y mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd la_oen_core[3] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[21\] _620_/Y mprj_logic_high_inst/HI[223] vssd vssd vccd
+ vccd la_oen_core[21] sky130_fd_sc_hd__einvp_8
X_431_ mprj_adr_o_core[24] vssd vssd vccd vccd _431_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_362_ la_oen_mprj[94] vssd vssd vccd vccd _362_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[29\] _500_/Y la_buf\[29\]/TE vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_13_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_A _593_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[25\]_B mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[86\]_A user_to_mprj_in_gates\[86\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_629_ la_oen_mprj[30] vssd vssd vccd vccd _629_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[124\]_A user_to_mprj_in_gates\[124\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] mprj_logic_high_inst/HI[348] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[113\]_A _584_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[77\]_A user_to_mprj_in_gates\[77\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_B mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_B mprj_logic_high_inst/HI[430] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[50\]_A _521_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[115\]_A user_to_mprj_in_gates\[115\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[104\]_A _575_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_A _512_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[69\] _337_/Y mprj_logic_high_inst/HI[271] vssd vssd vccd
+ vccd la_oen_core[69] sky130_fd_sc_hd__einvp_8
XFILLER_4_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[17\] _456_/Y mprj_dat_buf\[17\]/TE vssd vssd vccd vccd mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_414_ mprj_adr_o_core[7] vssd vssd vccd vccd _414_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_345_ la_oen_mprj[77] vssd vssd vccd vccd _345_/Y sky130_fd_sc_hd__inv_2
XANTENNA__405__A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[32\]_A _503_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[12\] _419_/Y mprj_adr_buf\[12\]/TE vssd vssd vccd vccd mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[126] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vssd vccd vccd la_data_in_mprj[92]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[99\]_A _570_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[23\]_A _494_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[14\]_A _485_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[96\] _567_/Y la_buf\[96\]/TE vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_19_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_58 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] mprj_logic_high_inst/HI[415] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[92\]_A _360_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[83\]_A _351_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _478_/Y la_buf\[7\]/TE vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_4_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[11\] _482_/Y la_buf\[11\]/TE vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__einvp_8
XFILLER_26_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[4\] _411_/Y mprj_adr_buf\[4\]/TE vssd vssd vccd vccd mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vssd vccd vccd la_data_in_mprj[55]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[74\]_A _342_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] mprj_logic_high_inst/HI[441] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[31\]_TE la_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[65\]_A _333_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__503__A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[121\] _389_/Y mprj_logic_high_inst/HI[323] vssd vssd vccd
+ vccd la_oen_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[2\] _405_/Y mprj_sel_buf\[2\]/TE vssd vssd vccd vccd mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[51\] _650_/Y mprj_logic_high_inst/HI[253] vssd vssd vccd
+ vccd la_oen_core[51] sky130_fd_sc_hd__einvp_8
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_593_ la_data_out_mprj[122] vssd vssd vccd vccd _593_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[59\] _530_/Y la_buf\[59\]/TE vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__einvp_8
XPHY_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[56\]_A _655_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__413__A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[115\] _586_/Y la_buf\[115\]/TE vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_3_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] mprj_logic_high_inst/HI[378] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_A _646_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _637_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[99\] _367_/Y mprj_logic_high_inst/HI[301] vssd vssd vccd
+ vccd la_oen_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_11_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_1_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_645_ la_oen_mprj[46] vssd vssd vccd vccd _645_/Y sky130_fd_sc_hd__inv_2
X_576_ la_data_out_mprj[105] vssd vssd vccd vccd _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__408__A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _628_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vssd vccd vccd la_data_in_mprj[18]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[25\]_A _432_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _601_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _423_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_430_ mprj_adr_o_core[23] vssd vssd vccd vccd _430_/Y sky130_fd_sc_hd__inv_2
X_361_ la_oen_mprj[93] vssd vssd vccd vccd _361_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[14\] _613_/Y mprj_logic_high_inst/HI[216] vssd vssd vccd
+ vccd la_oen_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_10_820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_628_ la_oen_mprj[29] vssd vssd vccd vccd _628_/Y sky130_fd_sc_hd__inv_2
X_559_ la_data_out_mprj[88] vssd vssd vccd vccd _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__601__A la_oen_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__511__A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_413_ mprj_adr_o_core[6] vssd vssd vccd vccd _413_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[41\] _512_/Y la_buf\[41\]/TE vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__einvp_8
X_344_ la_oen_mprj[76] vssd vssd vccd vccd _344_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__421__A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[119] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[29\]_A _468_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vssd vccd vccd la_data_in_mprj[85]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] mprj_logic_high_inst/HI[360] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[1\]_A _408_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__331__A la_oen_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_TE la_buf\[125\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__506__A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[81\] _349_/Y mprj_logic_high_inst/HI[283] vssd vssd vccd
+ vccd la_oen_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[89\] _560_/Y la_buf\[89\]/TE vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] mprj_logic_high_inst/HI[408] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[7\]_A _478_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vssd vccd vccd la_data_in_mprj[48]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] mprj_logic_high_inst/HI[434] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[1\]_B user_to_mprj_in_gates\[1\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[114\] _382_/Y mprj_logic_high_inst/HI[316] vssd vssd vccd
+ vccd la_oen_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_5_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[44\] _643_/Y mprj_logic_high_inst/HI[246] vssd vssd vccd
+ vccd la_oen_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_5_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_592_ la_data_out_mprj[121] vssd vssd vccd vccd _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[108\] _579_/Y la_buf\[108\]/TE vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[101] sky130_fd_sc_hd__inv_8
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__604__A la_oen_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[0\] _439_/Y mprj_dat_buf\[0\]/TE vssd vssd vccd vccd mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_26_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__514__A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high_inst/HI[309] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_644_ la_oen_mprj[45] vssd vssd vccd vccd _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[71\] _542_/Y la_buf\[71\]/TE vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__einvp_8
X_575_ la_data_out_mprj[104] vssd vssd vccd vccd _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__424__A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_12_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] mprj_logic_high_inst/HI[390] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__334__A la_oen_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__509__A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_360_ la_oen_mprj[92] vssd vssd vccd vccd _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[44\]_TE la_buf\[44\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__419__A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_627_ la_oen_mprj[28] vssd vssd vccd vccd _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_558_ la_data_out_mprj[87] vssd vssd vccd vccd _558_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_489_ la_data_out_mprj[18] vssd vssd vccd vccd _489_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vssd vccd vccd la_data_in_mprj[30]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[67\]_TE la_buf\[67\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_412_ mprj_adr_o_core[5] vssd vssd vccd vccd _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_343_ la_oen_mprj[75] vssd vssd vccd vccd _343_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[34\] _505_/Y la_buf\[34\]/TE vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_10_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vssd vccd vccd la_data_in_mprj[78]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] mprj_logic_high_inst/HI[353] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__612__A la_oen_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__522__A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[74\] _342_/Y mprj_logic_high_inst/HI[276] vssd vssd vccd
+ vccd la_oen_core[74] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[22\] _461_/Y mprj_dat_buf\[22\]/TE vssd vssd vccd vccd mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__432__A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__607__A la_oen_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[91\]_B mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__342__A la_oen_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__517__A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_B mprj_logic_high_inst/HI[412] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__427__A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_B mprj_logic_high_inst/HI[403] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[115\]_TE la_buf\[115\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] mprj_logic_high_inst/HI[420] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__337__A la_oen_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_B mprj_logic_high_inst/HI[394] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[107\] _375_/Y mprj_logic_high_inst/HI[309] vssd vssd vccd
+ vccd la_oen_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_5_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_660_ la_oen_mprj[61] vssd vssd vccd vccd _660_/Y sky130_fd_sc_hd__inv_2
X_591_ la_data_out_mprj[120] vssd vssd vccd vccd _591_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[37\] _636_/Y mprj_logic_high_inst/HI[239] vssd vssd vccd
+ vccd la_oen_core[37] sky130_fd_sc_hd__einvp_8
XFILLER_16_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[55\]_B mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vssd vccd vccd la_data_in_mprj[60]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[9\]_A _448_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[46\]_B mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_A _551_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__620__A la_oen_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_B mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_B mprj_logic_high_inst/HI[451] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _542_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__530__A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_643_ la_oen_mprj[44] vssd vssd vccd vccd _643_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_574_ la_data_out_mprj[103] vssd vssd vccd vccd _574_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[64\] _535_/Y la_buf\[64\]/TE vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__einvp_8
XPHY_151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[125\]_A _596_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[28\]_B mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B mprj_logic_high_inst/HI[442] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[62\]_A _533_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[28\] _435_/Y mprj_adr_buf\[28\]/TE vssd vssd vccd vccd mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[120\] _591_/Y la_buf\[120\]/TE vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_12_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__440__A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] mprj_logic_high_inst/HI[383] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[127\]_A user_to_mprj_in_gates\[127\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__615__A la_oen_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[116\]_A _587_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B mprj_logic_high_inst/HI[433] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_A _524_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__350__A la_oen_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[118\]_A user_to_mprj_in_gates\[118\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__525__A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_A _578_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[44\]_A _515_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_626_ la_oen_mprj[27] vssd vssd vccd vccd _626_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_557_ la_data_out_mprj[86] vssd vssd vccd vccd _557_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[109\]_A user_to_mprj_in_gates\[109\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_488_ la_data_out_mprj[17] vssd vssd vccd vccd _488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__435__A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vssd vccd vccd la_data_in_mprj[23]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[35\]_A _506_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[120\]_A _388_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__345__A la_oen_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_A _497_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[111\]_A _379_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_411_ mprj_adr_o_core[4] vssd vssd vccd vccd _411_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[1\] _600_/Y mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd la_oen_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_26_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_342_ la_oen_mprj[74] vssd vssd vccd vccd _342_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[11\]_TE la_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[17\]_A _488_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[27\] _498_/Y la_buf\[27\]/TE vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_13_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _370_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_609_ la_oen_mprj[10] vssd vssd vccd vccd _609_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] mprj_logic_high_inst/HI[346] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] mprj_logic_high_inst/HI[457] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_2010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[95\]_A _363_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_35 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[67\] _335_/Y mprj_logic_high_inst/HI[269] vssd vssd vccd
+ vccd la_oen_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _454_/Y mprj_dat_buf\[15\]/TE vssd vssd vccd vccd mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_A _354_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[10\] _417_/Y mprj_adr_buf\[10\]/TE vssd vssd vccd vccd mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[124] sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[10\]_A _609_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vssd vccd vccd la_data_in_mprj[90]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[77\]_A _345_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__623__A la_oen_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[68\]_A _336_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__533__A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[94\] _565_/Y la_buf\[94\]/TE vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_21_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _658_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__443__A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] mprj_logic_high_inst/HI[413] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__618__A la_oen_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__353__A la_oen_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_590_ la_data_out_mprj[119] vssd vssd vccd vccd _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[5\] _476_/Y la_buf\[5\]/TE vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[2\] _409_/Y mprj_adr_buf\[2\]/TE vssd vssd vccd vccd mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__438__A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vssd vccd vccd la_data_in_mprj[53]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_A _449_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[28\]_A _435_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__348__A la_oen_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _604_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[19\]_A _426_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_sel_buf\[0\] _403_/Y mprj_sel_buf\[0\]/TE vssd vssd vccd vccd mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_642_ la_oen_mprj[43] vssd vssd vccd vccd _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_573_ la_data_out_mprj[102] vssd vssd vccd vccd _573_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[57\] _528_/Y la_buf\[57\]/TE vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[105\]_TE la_buf\[105\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[113\] _584_/Y la_buf\[113\]/TE vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] mprj_logic_high_inst/HI[376] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__631__A la_oen_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] user_to_mprj_in_gates\[8\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[97\] _365_/Y mprj_logic_high_inst/HI[299] vssd vssd vccd
+ vccd la_oen_core[97] sky130_fd_sc_hd__einvp_8
XANTENNA__541__A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_625_ la_oen_mprj[26] vssd vssd vccd vccd _625_/Y sky130_fd_sc_hd__inv_2
X_556_ la_data_out_mprj[85] vssd vssd vccd vccd _556_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_487_ la_data_out_mprj[16] vssd vssd vccd vccd _487_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vssd vccd vccd la_data_in_mprj[16]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__451__A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__626__A la_oen_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _411_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A la_oen_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_410_ mprj_adr_o_core[3] vssd vssd vccd vccd _410_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__536__A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[12\] _611_/Y mprj_logic_high_inst/HI[214] vssd vssd vccd
+ vccd la_oen_core[12] sky130_fd_sc_hd__einvp_8
X_341_ la_oen_mprj[73] vssd vssd vccd vccd _341_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vssd vccd vccd la_data_in_mprj[8]
+ sky130_fd_sc_hd__inv_8
XFILLER_10_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_stb_buf _401_/Y mprj_stb_buf/TE vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_4_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_608_ la_oen_mprj[9] vssd vssd vccd vccd _608_/Y sky130_fd_sc_hd__inv_2
XANTENNA__446__A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_539_ la_data_out_mprj[68] vssd vssd vccd vccd _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__356__A la_oen_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_clk_buf_A _398_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[117] sky130_fd_sc_hd__inv_8
XFILLER_2_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vssd vccd vccd la_data_in_mprj[83]
+ sky130_fd_sc_hd__inv_8
XFILLER_24_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_B user_to_mprj_in_gates\[4\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[87\] _558_/Y la_buf\[87\]/TE vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_21_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_90 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] mprj_logic_high_inst/HI[406] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__634__A la_oen_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vssd vccd vccd la_data_in_mprj[46]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XPHY_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__629__A la_oen_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] mprj_logic_high_inst/HI[432] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__364__A la_oen_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[112\] _380_/Y mprj_logic_high_inst/HI[314] vssd vssd vccd
+ vccd la_oen_core[112] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[42\] _641_/Y mprj_logic_high_inst/HI[244] vssd vssd vccd
+ vccd la_oen_core[42] sky130_fd_sc_hd__einvp_8
XANTENNA__539__A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_641_ la_oen_mprj[42] vssd vssd vccd vccd _641_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_572_ la_data_out_mprj[101] vssd vssd vccd vccd _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[106\] _577_/Y la_buf\[106\]/TE vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_7_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__449__A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] mprj_logic_high_inst/HI[369] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__359__A la_oen_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_624_ la_oen_mprj[25] vssd vssd vccd vccd _624_/Y sky130_fd_sc_hd__inv_2
X_555_ la_data_out_mprj[84] vssd vssd vccd vccd _555_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_486_ la_data_out_mprj[15] vssd vssd vccd vccd _486_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_we_buf _402_/Y mprj_we_buf/TE vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_9_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_pwrgood mprj_pwrgood/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_9_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__642__A la_oen_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_340_ la_oen_mprj[72] vssd vssd vccd vccd _340_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__552__A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high_inst/HI[244] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_607_ la_oen_mprj[8] vssd vssd vccd vccd _607_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_538_ la_data_out_mprj[67] vssd vssd vccd vccd _538_/Y sky130_fd_sc_hd__inv_2
X_469_ mprj_dat_o_core[30] vssd vssd vccd vccd _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__462__A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__637__A la_oen_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__372__A la_oen_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[80\]_TE la_buf\[80\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__547__A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_we_buf_A _402_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[85\]_B mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[32\] _503_/Y la_buf\[32\]/TE vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__einvp_8
XFILLER_13_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vssd vccd vccd la_data_in_mprj[76]
+ sky130_fd_sc_hd__inv_8
XANTENNA__457__A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] mprj_logic_high_inst/HI[351] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[76\]_B mprj_logic_high_inst/HI[406] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[9\] _448_/Y mprj_dat_buf\[9\]/TE vssd vssd vccd vccd mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_25_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[61\]_A user_to_mprj_in_gates\[61\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__367__A la_oen_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[67\]_B mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[72\] _340_/Y mprj_logic_high_inst/HI[274] vssd vssd vccd
+ vccd la_oen_core[72] sky130_fd_sc_hd__einvp_8
XFILLER_8_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _459_/Y mprj_dat_buf\[20\]/TE vssd vssd vccd vccd mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[58\]_B mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[92\]_A _563_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] mprj_logic_high_inst/HI[399] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_B mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[83\]_A _554_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__650__A la_oen_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[124\]_B mprj_logic_high_inst/HI[454] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[74\]_A _545_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__560__A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[115\]_B mprj_logic_high_inst/HI[445] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vssd vccd vccd la_data_in_mprj[39]
+ sky130_fd_sc_hd__inv_8
XPHY_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[65\]_A _536_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__470__A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__645__A la_oen_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[119\]_A _590_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B mprj_logic_high_inst/HI[436] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[56\]_A _527_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__380__A la_oen_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[105\] _373_/Y mprj_logic_high_inst/HI[307] vssd vssd vccd
+ vccd la_oen_core[105] sky130_fd_sc_hd__einvp_8
X_640_ la_oen_mprj[41] vssd vssd vccd vccd _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_571_ la_data_out_mprj[100] vssd vssd vccd vccd _571_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[35\] _634_/Y mprj_logic_high_inst/HI[237] vssd vssd vccd
+ vccd la_oen_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_18_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__555__A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[47\]_A _518_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__465__A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[38\]_A _509_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[123\]_A _391_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__375__A la_oen_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[29\]_A _500_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[114\]_A _382_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_623_ la_oen_mprj[24] vssd vssd vccd vccd _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[62\] _533_/Y la_buf\[62\]/TE vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__einvp_8
X_554_ la_data_out_mprj[83] vssd vssd vccd vccd _554_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_485_ la_data_out_mprj[14] vssd vssd vccd vccd _485_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[26\] _433_/Y mprj_adr_buf\[26\]/TE vssd vssd vccd vccd mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[40\]_A _639_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_A _373_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] mprj_logic_high_inst/HI[381] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _630_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_A _366_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[22\]_A _621_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_A _357_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_606_ la_oen_mprj[7] vssd vssd vccd vccd _606_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_537_ la_data_out_mprj[66] vssd vssd vccd vccd _537_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_468_ mprj_dat_o_core[29] vssd vssd vccd vccd _468_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_399_ caravel_clk2 vssd vssd vccd vccd _399_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vssd vccd vccd la_data_in_mprj[21]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[13\]_A _612_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] mprj_logic_high_inst/HI[429] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__653__A la_oen_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__563__A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[25\] _496_/Y la_buf\[25\]/TE vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_6_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vssd vccd vccd la_data_in_mprj[69]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__473__A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] mprj_logic_high_inst/HI[344] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] mprj_logic_high_inst/HI[455] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__648__A la_oen_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[31\]_A _470_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__383__A la_oen_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[65\] _333_/Y mprj_logic_high_inst/HI[267] vssd vssd vccd
+ vccd la_oen_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_8_1020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[13\] _452_/Y mprj_dat_buf\[13\]/TE vssd vssd vccd vccd mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__558__A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[108\]_TE la_buf\[108\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[22\]_A _461_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[122] sky130_fd_sc_hd__inv_8
XFILLER_3_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__468__A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_A _452_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high_inst/HI[257] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__378__A la_oen_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _607_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[92\] _563_/Y la_buf\[92\]/TE vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[93\]_TE la_buf\[93\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] mprj_logic_high_inst/HI[411] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_570_ la_data_out_mprj[99] vssd vssd vccd vccd _570_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[28\] _627_/Y mprj_logic_high_inst/HI[230] vssd vssd vccd
+ vccd la_oen_core[28] sky130_fd_sc_hd__einvp_8
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[0\]_A _471_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__571__A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[3\] _474_/Y la_buf\[3\]/TE vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_10_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[0\] _407_/Y mprj_adr_buf\[0\]/TE vssd vssd vccd vccd mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vssd vccd vccd la_data_in_mprj[51]
+ sky130_fd_sc_hd__inv_8
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__481__A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__656__A la_oen_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[7\]_A _414_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__391__A la_oen_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_622_ la_oen_mprj[23] vssd vssd vccd vccd _622_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__566__A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_553_ la_data_out_mprj[82] vssd vssd vccd vccd _553_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_484_ la_data_out_mprj[13] vssd vssd vccd vccd _484_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[55\] _526_/Y la_buf\[55\]/TE vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__einvp_8
XFILLER_18_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[19\] _426_/Y mprj_adr_buf\[19\]/TE vssd vssd vccd vccd mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _582_/Y la_buf\[111\]/TE vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_25_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vssd vccd vccd la_data_in_mprj[99]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__476__A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] mprj_logic_high_inst/HI[374] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] user_to_mprj_in_gates\[6\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__386__A la_oen_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[95\] _363_/Y mprj_logic_high_inst/HI[297] vssd vssd vccd
+ vccd la_oen_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_5_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_81 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_605_ la_oen_mprj[6] vssd vssd vccd vccd _605_/Y sky130_fd_sc_hd__inv_2
X_536_ la_data_out_mprj[65] vssd vssd vccd vccd _536_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_467_ mprj_dat_o_core[28] vssd vssd vccd vccd _467_/Y sky130_fd_sc_hd__inv_2
X_398_ caravel_clk vssd vssd vccd vccd _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vssd vccd vccd la_data_in_mprj[14]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_B user_to_mprj_in_gates\[7\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[10\] _609_/Y mprj_logic_high_inst/HI[212] vssd vssd vccd
+ vccd la_oen_core[10] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vssd vccd vccd la_data_in_mprj[6]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[18\] _489_/Y la_buf\[18\]/TE vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_13_1498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_519_ la_data_out_mprj[48] vssd vssd vccd vccd _519_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] mprj_logic_high_inst/HI[448] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[58\] _657_/Y mprj_logic_high_inst/HI[260] vssd vssd vccd
+ vccd la_oen_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_5_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__574__A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[115] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vssd vccd vccd la_data_in_mprj[81]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__484__A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_1_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__659__A la_oen_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__394__A la_oen_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_51 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__569__A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[85\] _556_/Y la_buf\[85\]/TE vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_19_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__479__A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] mprj_logic_high_inst/HI[404] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__389__A la_oen_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high_inst/HI[247] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vssd vccd vccd la_data_in_mprj[44]
+ sky130_fd_sc_hd__inv_8
XPHY_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[1\]_A _404_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] mprj_logic_high_inst/HI[430] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[83\]_TE la_buf\[83\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high_inst/HI[270] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[110\] _378_/Y mprj_logic_high_inst/HI[312] vssd vssd vccd
+ vccd la_oen_core[110] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[40\] _639_/Y mprj_logic_high_inst/HI[242] vssd vssd vccd
+ vccd la_oen_core[40] sky130_fd_sc_hd__einvp_8
X_621_ la_oen_mprj[22] vssd vssd vccd vccd _621_/Y sky130_fd_sc_hd__inv_2
X_552_ la_data_out_mprj[81] vssd vssd vccd vccd _552_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_483_ la_data_out_mprj[12] vssd vssd vccd vccd _483_/Y sky130_fd_sc_hd__inv_2
XANTENNA__582__A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[48\] _519_/Y la_buf\[48\]/TE vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_9_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _441_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[104\] _575_/Y la_buf\[104\]/TE vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_23_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] mprj_logic_high_inst/HI[367] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__492__A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[91\]_A user_to_mprj_in_gates\[91\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[30\]_B mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _356_/Y mprj_logic_high_inst/HI[290] vssd vssd vccd
+ vccd la_oen_core[88] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[21\]_B mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[82\]_A user_to_mprj_in_gates\[82\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__577__A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_604_ la_oen_mprj[5] vssd vssd vccd vccd _604_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_535_ la_data_out_mprj[64] vssd vssd vccd vccd _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[88\]_B mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_466_ mprj_dat_o_core[27] vssd vssd vccd vccd _466_/Y sky130_fd_sc_hd__inv_2
X_397_ user_resetn vssd vssd vccd vccd user_reset sky130_fd_sc_hd__inv_2
XFILLER_9_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[31\] _438_/Y mprj_adr_buf\[31\]/TE vssd vssd vccd vccd mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[120\]_A user_to_mprj_in_gates\[120\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[73\]_A user_to_mprj_in_gates\[73\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_B mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__487__A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[79\]_B mprj_logic_high_inst/HI[409] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[111\]_A user_to_mprj_in_gates\[111\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[100\]_A _571_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[64\]_A user_to_mprj_in_gates\[64\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__397__A user_resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_518_ la_data_out_mprj[47] vssd vssd vccd vccd _518_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[95\]_A _566_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_449_ mprj_dat_o_core[10] vssd vssd vccd vccd _449_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[86\]_A _557_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[10\]_A _481_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B mprj_logic_high_inst/HI[457] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[77\]_A _548_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__590__A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[30\] _501_/Y la_buf\[30\]/TE vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[108] sky130_fd_sc_hd__inv_8
XFILLER_26_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vssd vccd vccd la_data_in_mprj[74]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[118\]_B mprj_logic_high_inst/HI[448] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[68\]_A _539_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[19\]_A user_to_mprj_in_gates\[19\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[7\] _446_/Y mprj_dat_buf\[7\]/TE vssd vssd vccd vccd mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_B mprj_logic_high_inst/HI[439] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[59\]_A _530_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[70\] _338_/Y mprj_logic_high_inst/HI[272] vssd vssd vccd
+ vccd la_oen_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_10_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[78\] _549_/Y la_buf\[78\]/TE vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__einvp_8
XANTENNA__585__A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[70\]_A _338_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] mprj_logic_high_inst/HI[397] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__495__A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[126\]_A _394_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[61\]_A _660_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[52\]_A _651_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_A _385_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vssd vccd vccd la_data_in_mprj[37]
+ sky130_fd_sc_hd__inv_8
XPHY_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[108\]_A _376_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[43\]_A _642_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _633_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[103\] _371_/Y mprj_logic_high_inst/HI[305] vssd vssd vccd
+ vccd la_oen_core[103] sky130_fd_sc_hd__einvp_8
X_620_ la_oen_mprj[21] vssd vssd vccd vccd _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_551_ la_data_out_mprj[80] vssd vssd vccd vccd _551_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[33\] _632_/Y mprj_logic_high_inst/HI[235] vssd vssd vccd
+ vccd la_oen_core[33] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[30\]_A _437_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_482_ la_data_out_mprj[11] vssd vssd vccd vccd _482_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_A _624_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[21\]_A _428_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _615_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_A _419_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[50\]_TE la_buf\[50\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[29\] _468_/Y mprj_dat_buf\[29\]/TE vssd vssd vccd vccd mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_2_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_603_ la_oen_mprj[4] vssd vssd vccd vccd _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_534_ la_data_out_mprj[63] vssd vssd vccd vccd _534_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[60\] _531_/Y la_buf\[60\]/TE vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__einvp_8
X_465_ mprj_dat_o_core[26] vssd vssd vccd vccd _465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__593__A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_396_ caravel_rstn vssd vssd vccd vccd _396_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[24\] _431_/Y mprj_adr_buf\[24\]/TE vssd vssd vccd vccd mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[73\]_TE la_buf\[73\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_TE mprj_logic_high_inst/HI[260] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__588__A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[96\]_TE la_buf\[96\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[25\]_A _464_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_517_ la_data_out_mprj[46] vssd vssd vccd vccd _517_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_448_ mprj_dat_o_core[9] vssd vssd vccd vccd _448_/Y sky130_fd_sc_hd__inv_2
X_379_ la_oen_mprj[111] vssd vssd vccd vccd _379_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] mprj_logic_high_inst/HI[427] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__498__A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[16\]_A _455_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[23\] _494_/Y la_buf\[23\]/TE vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_3_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vssd vccd vccd la_data_in_mprj[67]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] mprj_logic_high_inst/HI[342] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_11_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] mprj_logic_high_inst/HI[453] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[63\] _331_/Y mprj_logic_high_inst/HI[265] vssd vssd vccd
+ vccd la_oen_core[63] sky130_fd_sc_hd__einvp_8
XFILLER_27_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[11\] _450_/Y mprj_dat_buf\[11\]/TE vssd vssd vccd vccd mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_A _474_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[121\]_TE la_buf\[121\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[127\] _598_/Y la_buf\[127\]/TE vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[120] sky130_fd_sc_hd__inv_8
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__596__A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _561_/Y la_buf\[90\]/TE vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_21_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[1\]_A user_to_mprj_in_gates\[1\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_550_ la_data_out_mprj[79] vssd vssd vccd vccd _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[8\] _607_/Y mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd la_oen_core[8] sky130_fd_sc_hd__einvp_8
X_481_ la_data_out_mprj[10] vssd vssd vccd vccd _481_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[26\] _625_/Y mprj_logic_high_inst/HI[228] vssd vssd vccd
+ vccd la_oen_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_25_450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[1\] _472_/Y la_buf\[1\]/TE vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_10_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_602_ la_oen_mprj[3] vssd vssd vccd vccd _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_533_ la_data_out_mprj[62] vssd vssd vccd vccd _533_/Y sky130_fd_sc_hd__inv_2
X_464_ mprj_dat_o_core[25] vssd vssd vccd vccd _464_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[53\] _524_/Y la_buf\[53\]/TE vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__einvp_8
X_395_ la_oen_mprj[127] vssd vssd vccd vccd _395_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[17\] _424_/Y mprj_adr_buf\[17\]/TE vssd vssd vccd vccd mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vssd vccd vccd la_data_in_mprj[97]
+ sky130_fd_sc_hd__inv_8
XFILLER_27_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] mprj_logic_high_inst/HI[372] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_1660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] user_to_mprj_in_gates\[4\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[93\] _361_/Y mprj_logic_high_inst/HI[295] vssd vssd vccd
+ vccd la_oen_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_2_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_516_ la_data_out_mprj[45] vssd vssd vccd vccd _516_/Y sky130_fd_sc_hd__inv_2
X_447_ mprj_dat_o_core[8] vssd vssd vccd vccd _447_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_378_ la_oen_mprj[110] vssd vssd vccd vccd _378_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vssd vccd vccd la_data_in_mprj[12]
+ sky130_fd_sc_hd__inv_8
XFILLER_6_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high_inst/HI[227] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vssd vccd vccd la_data_in_mprj[4]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[63\]_TE la_buf\[63\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[16\] _487_/Y la_buf\[16\]/TE vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__599__A la_oen_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[9\] _416_/Y mprj_adr_buf\[9\]/TE vssd vssd vccd vccd mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] mprj_logic_high_inst/HI[446] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _394_/Y mprj_logic_high_inst/HI[328] vssd vssd vccd
+ vccd la_oen_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_0_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[56\] _655_/Y mprj_logic_high_inst/HI[258] vssd vssd vccd
+ vccd la_oen_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_19_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[113] sky130_fd_sc_hd__inv_8
XFILLER_26_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[60\]_B mprj_logic_high_inst/HI[390] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[51\]_B mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[83\] _554_/Y la_buf\[83\]/TE vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_21_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_dat_buf\[5\]_A _444_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[42\]_B mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] mprj_logic_high_inst/HI[402] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[33\]_B mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_480_ la_data_out_mprj[9] vssd vssd vccd vccd _480_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[19\] _618_/Y mprj_logic_high_inst/HI[221] vssd vssd vccd
+ vccd la_oen_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_25_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[121\]_A _592_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[85\]_A user_to_mprj_in_gates\[85\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[24\]_B mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__400__A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vssd vccd vccd la_data_in_mprj[42]
+ sky130_fd_sc_hd__inv_8
XPHY_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[123\]_A user_to_mprj_in_gates\[123\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[112\]_A _583_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_B mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[114\]_A user_to_mprj_in_gates\[114\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[103\]_A _574_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[67\]_A user_to_mprj_in_gates\[67\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[40\]_A _511_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_601_ la_oen_mprj[2] vssd vssd vccd vccd _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_532_ la_data_out_mprj[61] vssd vssd vccd vccd _532_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_463_ mprj_dat_o_core[24] vssd vssd vccd vccd _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_394_ la_oen_mprj[126] vssd vssd vccd vccd _394_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[46\] _517_/Y la_buf\[46\]/TE vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[31\]_A _502_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[102\] _573_/Y la_buf\[102\]/TE vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_1_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[98\]_A _569_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] mprj_logic_high_inst/HI[365] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[22\]_A _493_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[89\]_A _560_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[86\] _354_/Y mprj_logic_high_inst/HI[288] vssd vssd vccd
+ vccd la_oen_core[86] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[13\]_A _484_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_515_ la_data_out_mprj[44] vssd vssd vccd vccd _515_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_446_ mprj_dat_o_core[7] vssd vssd vccd vccd _446_/Y sky130_fd_sc_hd__inv_2
X_377_ la_oen_mprj[109] vssd vssd vccd vccd _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[91\]_A _359_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_A _350_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_429_ mprj_adr_o_core[22] vssd vssd vccd vccd _429_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[73\]_A _341_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] mprj_logic_high_inst/HI[439] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_A _332_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[119\] _387_/Y mprj_logic_high_inst/HI[321] vssd vssd vccd
+ vccd la_oen_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_0_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[49\] _648_/Y mprj_logic_high_inst/HI[251] vssd vssd vccd
+ vccd la_oen_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[55\]_A _654_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__403__A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[106] sky130_fd_sc_hd__inv_8
XFILLER_4_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vssd vccd vccd la_data_in_mprj[72]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[46\]_A _645_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[5\] _444_/Y mprj_dat_buf\[5\]/TE vssd vssd vccd vccd mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _636_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[76\] _547_/Y la_buf\[76\]/TE vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__einvp_8
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[28\]_A _627_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_A _431_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] mprj_logic_high_inst/HI[395] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[19\]_A _618_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _600_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[15\]_A _422_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vssd vccd vccd la_data_in_mprj[35]
+ sky130_fd_sc_hd__inv_8
XPHY_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__501__A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _369_/Y mprj_logic_high_inst/HI[303] vssd vssd vccd
+ vccd la_oen_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_24_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_600_ la_oen_mprj[1] vssd vssd vccd vccd _600_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[31\] _630_/Y mprj_logic_high_inst/HI[233] vssd vssd vccd
+ vccd la_oen_core[31] sky130_fd_sc_hd__einvp_8
X_531_ la_data_out_mprj[60] vssd vssd vccd vccd _531_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_462_ mprj_dat_o_core[23] vssd vssd vccd vccd _462_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_393_ la_oen_mprj[125] vssd vssd vccd vccd _393_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[39\] _510_/Y la_buf\[39\]/TE vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_12_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__411__A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[28\]_A _467_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] mprj_logic_high_inst/HI[358] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[0\]_A _407_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_A _458_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_66 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[79\] _347_/Y mprj_logic_high_inst/HI[281] vssd vssd vccd
+ vccd la_oen_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_1_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[27\] _466_/Y mprj_dat_buf\[27\]/TE vssd vssd vccd vccd mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_514_ la_data_out_mprj[43] vssd vssd vccd vccd _514_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[124\]_TE la_buf\[124\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_445_ mprj_dat_o_core[6] vssd vssd vccd vccd _445_/Y sky130_fd_sc_hd__inv_2
X_376_ la_oen_mprj[108] vssd vssd vccd vccd _376_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__406__A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[22\] _429_/Y mprj_adr_buf\[22\]/TE vssd vssd vccd vccd mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_7_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[6\]_A _477_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_428_ mprj_adr_o_core[21] vssd vssd vccd vccd _428_/Y sky130_fd_sc_hd__inv_2
X_359_ la_oen_mprj[91] vssd vssd vccd vccd _359_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] mprj_logic_high_inst/HI[425] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[0\]_B user_to_mprj_in_gates\[0\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[21\] _492_/Y la_buf\[21\]/TE vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__einvp_8
XFILLER_10_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vssd vccd vccd la_data_in_mprj[65]
+ sky130_fd_sc_hd__inv_8
XFILLER_21_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] mprj_logic_high_inst/HI[340] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] mprj_logic_high_inst/HI[451] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__504__A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_66 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[61\] _660_/Y mprj_logic_high_inst/HI[263] vssd vssd vccd
+ vccd la_oen_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_21_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[69\] _540_/Y la_buf\[69\]/TE vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__einvp_8
XPHY_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__414__A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _596_/Y la_buf\[125\]/TE vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_10_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] mprj_logic_high_inst/HI[388] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_88 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__409__A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vssd vccd vccd la_data_in_mprj[28]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_530_ la_data_out_mprj[59] vssd vssd vccd vccd _530_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[24\] _623_/Y mprj_logic_high_inst/HI[226] vssd vssd vccd
+ vccd la_oen_core[24] sky130_fd_sc_hd__einvp_8
X_461_ mprj_dat_o_core[22] vssd vssd vccd vccd _461_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[6\] _605_/Y mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd la_oen_core[6] sky130_fd_sc_hd__einvp_8
X_392_ la_oen_mprj[124] vssd vssd vccd vccd _392_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_659_ la_oen_mprj[60] vssd vssd vccd vccd _659_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__602__A la_oen_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[89\]_TE la_buf\[89\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__512__A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_513_ la_data_out_mprj[42] vssd vssd vccd vccd _513_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_444_ mprj_dat_o_core[5] vssd vssd vccd vccd _444_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[51\] _522_/Y la_buf\[51\]/TE vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__einvp_8
X_375_ la_oen_mprj[107] vssd vssd vccd vccd _375_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__422__A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[15\] _422_/Y mprj_adr_buf\[15\]/TE vssd vssd vccd vccd mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vssd vccd vccd la_data_in_mprj[95]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] mprj_logic_high_inst/HI[370] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_B mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__332__A la_oen_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] user_to_mprj_in_gates\[2\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__507__A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[81\]_B mprj_logic_high_inst/HI[411] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[91\] _359_/Y mprj_logic_high_inst/HI[293] vssd vssd vccd
+ vccd la_oen_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_26_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[99\] _570_/Y la_buf\[99\]/TE vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_24_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__417__A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_427_ mprj_adr_o_core[20] vssd vssd vccd vccd _427_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_358_ la_oen_mprj[90] vssd vssd vccd vccd _358_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[72\]_B mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vssd vccd vccd la_data_in_mprj[10]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] mprj_logic_high_inst/HI[418] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_B mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[114\]_TE la_buf\[114\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vssd vccd vccd la_data_in_mprj[2]
+ sky130_fd_sc_hd__inv_8
XPHY_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[54\]_B mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[14\] _485_/Y la_buf\[14\]/TE vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_10_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high_inst/HI[263] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[7\] _414_/Y mprj_adr_buf\[7\]/TE vssd vssd vccd vccd mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vssd vccd vccd la_data_in_mprj[58]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[8\]_A _447_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[45\]_B mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__610__A la_oen_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] mprj_logic_high_inst/HI[444] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[30\]_A user_to_mprj_in_gates\[30\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_B mprj_logic_high_inst/HI[450] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[97\]_A user_to_mprj_in_gates\[97\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[70\]_A _541_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _392_/Y mprj_logic_high_inst/HI[326] vssd vssd vccd
+ vccd la_oen_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_7_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__520__A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[54\] _653_/Y mprj_logic_high_inst/HI[256] vssd vssd vccd
+ vccd la_oen_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_21_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[21\]_A user_to_mprj_in_gates\[21\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[124\]_A _595_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B mprj_logic_high_inst/HI[441] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_B mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[61\]_A _532_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[118\] _589_/Y la_buf\[118\]/TE vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_10_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[111] sky130_fd_sc_hd__inv_8
XANTENNA__430__A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[126\]_A user_to_mprj_in_gates\[126\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__605__A la_oen_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[115\]_A _586_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[79\]_A user_to_mprj_in_gates\[79\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_B mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B mprj_logic_high_inst/HI[432] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[52\]_A _523_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__340__A la_oen_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[117\]_A user_to_mprj_in_gates\[117\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__515__A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[106\]_A _577_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_A _514_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[81\] _552_/Y la_buf\[81\]/TE vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_5_2084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__425__A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[34\]_A _505_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] mprj_logic_high_inst/HI[400] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _398_/Y mprj_clk_buf/TE vssd vssd vccd vccd user_clock sky130_fd_sc_hd__einvp_8
XFILLER_22_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__335__A la_oen_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[25\]_A _496_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[110\]_A _378_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_460_ mprj_dat_o_core[21] vssd vssd vccd vccd _460_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_391_ la_oen_mprj[123] vssd vssd vccd vccd _391_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[17\] _616_/Y mprj_logic_high_inst/HI[219] vssd vssd vccd
+ vccd la_oen_core[17] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[16\]_A _487_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _369_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_658_ la_oen_mprj[59] vssd vssd vccd vccd _658_/Y sky130_fd_sc_hd__inv_2
X_589_ la_data_out_mprj[118] vssd vssd vccd vccd _589_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[10\]_TE la_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vssd vccd vccd la_data_in_mprj[40]
+ sky130_fd_sc_hd__inv_8
XPHY_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_A _362_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_512_ la_data_out_mprj[41] vssd vssd vccd vccd _512_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_443_ mprj_dat_o_core[4] vssd vssd vccd vccd _443_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_A _353_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_374_ la_oen_mprj[106] vssd vssd vccd vccd _374_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[44\] _515_/Y la_buf\[44\]/TE vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_9_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[100\] _571_/Y la_buf\[100\]/TE vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_0_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vssd vccd vccd la_data_in_mprj[88]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] mprj_logic_high_inst/HI[363] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[76\]_A _344_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__613__A la_oen_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[67\]_A _335_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__523__A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[84\] _352_/Y mprj_logic_high_inst/HI[286] vssd vssd vccd
+ vccd la_oen_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_3_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_A _657_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_426_ mprj_adr_o_core[19] vssd vssd vccd vccd _426_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_357_ la_oen_mprj[89] vssd vssd vccd vccd _357_/Y sky130_fd_sc_hd__inv_2
XANTENNA__433__A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_TE la_buf\[79\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__A la_oen_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_A _648_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__343__A la_oen_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__428__A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_409_ mprj_adr_o_core[2] vssd vssd vccd vccd _409_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[27\]_A _434_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] mprj_logic_high_inst/HI[437] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__338__A la_oen_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _603_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[18\]_A _425_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[117\] _385_/Y mprj_logic_high_inst/HI[319] vssd vssd vccd
+ vccd la_oen_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_21_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[47\] _646_/Y mprj_logic_high_inst/HI[249] vssd vssd vccd
+ vccd la_oen_core[47] sky130_fd_sc_hd__einvp_8
XPHY_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[104] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vssd vccd vccd la_data_in_mprj[70]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__621__A la_oen_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[3\] _442_/Y mprj_dat_buf\[3\]/TE vssd vssd vccd vccd mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_22_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[51\]_TE mprj_logic_high_inst/HI[253] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__531__A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[7\]_TE mprj_dat_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[127\]_TE la_buf\[127\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[74\] _545_/Y la_buf\[74\]/TE vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_16_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__441__A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] mprj_logic_high_inst/HI[393] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__616__A la_oen_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_A _410_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__351__A la_oen_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_390_ la_oen_mprj[122] vssd vssd vccd vccd _390_/Y sky130_fd_sc_hd__inv_2
XANTENNA__526__A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_657_ la_oen_mprj[58] vssd vssd vccd vccd _657_/Y sky130_fd_sc_hd__inv_2
X_588_ la_data_out_mprj[117] vssd vssd vccd vccd _588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__436__A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vssd vccd vccd la_data_in_mprj[33]
+ sky130_fd_sc_hd__inv_8
XPHY_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__346__A la_oen_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_511_ la_data_out_mprj[40] vssd vssd vccd vccd _511_/Y sky130_fd_sc_hd__inv_2
X_442_ mprj_dat_o_core[3] vssd vssd vccd vccd _442_/Y sky130_fd_sc_hd__inv_2
X_373_ la_oen_mprj[105] vssd vssd vccd vccd _373_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[37\] _508_/Y la_buf\[37\]/TE vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_A _480_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] mprj_logic_high_inst/HI[356] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_B user_to_mprj_in_gates\[3\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[77\] _345_/Y mprj_logic_high_inst/HI[279] vssd vssd vccd
+ vccd la_oen_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_3_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[25\] _464_/Y mprj_dat_buf\[25\]/TE vssd vssd vccd vccd mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_425_ mprj_adr_o_core[18] vssd vssd vccd vccd _425_/Y sky130_fd_sc_hd__inv_2
X_356_ la_oen_mprj[88] vssd vssd vccd vccd _356_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[20\] _427_/Y mprj_adr_buf\[20\]/TE vssd vssd vccd vccd mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__624__A la_oen_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__534__A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_408_ mprj_adr_o_core[1] vssd vssd vccd vccd _408_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__444__A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_339_ la_oen_mprj[71] vssd vssd vccd vccd _339_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] mprj_logic_high_inst/HI[423] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__619__A la_oen_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__354__A la_oen_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_14_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__529__A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[69\]_TE la_buf\[69\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__439__A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vssd vccd vccd la_data_in_mprj[63]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__349__A la_oen_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[67\] _538_/Y la_buf\[67\]/TE vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__einvp_8
XPHY_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[123\] _594_/Y la_buf\[123\]/TE vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_26_1066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] mprj_logic_high_inst/HI[386] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__632__A la_oen_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__542__A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_656_ la_oen_mprj[57] vssd vssd vccd vccd _656_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_587_ la_data_out_mprj[116] vssd vssd vccd vccd _587_/Y sky130_fd_sc_hd__inv_2
XPHY_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vssd vccd vccd la_data_in_mprj[26]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__452__A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high_inst/HI[243] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__627__A la_oen_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[93\]_B mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__362__A la_oen_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[117\]_TE la_buf\[117\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_510_ la_data_out_mprj[39] vssd vssd vccd vccd _510_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[4\] _603_/Y mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd la_oen_core[4] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[22\] _621_/Y mprj_logic_high_inst/HI[224] vssd vssd vccd
+ vccd la_oen_core[22] sky130_fd_sc_hd__einvp_8
XANTENNA__537__A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_441_ mprj_dat_o_core[2] vssd vssd vccd vccd _441_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_372_ la_oen_mprj[104] vssd vssd vccd vccd _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high_inst/HI[266] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__447__A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_639_ la_oen_mprj[40] vssd vssd vccd vccd _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] mprj_logic_high_inst/HI[349] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[75\]_B mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__357__A la_oen_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_B mprj_logic_high_inst/HI[396] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[18\] _457_/Y mprj_dat_buf\[18\]/TE vssd vssd vccd vccd mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_424_ mprj_adr_o_core[17] vssd vssd vccd vccd _424_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_355_ la_oen_mprj[87] vssd vssd vccd vccd _355_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_B mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[91\]_A _562_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[13\] _420_/Y mprj_adr_buf\[13\]/TE vssd vssd vccd vccd mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[127] sky130_fd_sc_hd__inv_8
XFILLER_9_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vssd vccd vccd la_data_in_mprj[93]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_buffers\[42\]_A user_to_mprj_in_gates\[42\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_B mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[82\]_A _553_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__640__A la_oen_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] user_to_mprj_in_gates\[0\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[123\]_B mprj_logic_high_inst/HI[453] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[39\]_B mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[73\]_A _544_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__550__A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[97\] _568_/Y la_buf\[97\]/TE vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_4_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_407_ mprj_adr_o_core[0] vssd vssd vccd vccd _407_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[127\]_A _598_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B mprj_logic_high_inst/HI[444] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_338_ la_oen_mprj[70] vssd vssd vccd vccd _338_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[64\]_A _535_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__460__A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] mprj_logic_high_inst/HI[416] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__635__A la_oen_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_A _589_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_B mprj_logic_high_inst/HI[435] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_A _526_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__370__A la_oen_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__545__A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vssd vccd vccd la_data_in_mprj[0]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[109\]_A _580_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[46\]_A _517_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[8\] _479_/Y la_buf\[8\]/TE vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__einvp_8
Xla_buf\[12\] _483_/Y la_buf\[12\]/TE vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__einvp_8
XFILLER_10_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _412_/Y mprj_adr_buf\[5\]/TE vssd vssd vccd vccd mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vssd vccd vccd la_data_in_mprj[56]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__455__A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[37\]_A _508_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[122\]_A _390_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] mprj_logic_high_inst/HI[442] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__365__A la_oen_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[28\]_A _499_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[122\] _390_/Y mprj_logic_high_inst/HI[324] vssd vssd vccd
+ vccd la_oen_core[122] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[113\]_A _381_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_sel_buf\[3\] _406_/Y mprj_sel_buf\[3\]/TE vssd vssd vccd vccd mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[52\] _651_/Y mprj_logic_high_inst/HI[254] vssd vssd vccd
+ vccd la_oen_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_5_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[36\]_TE la_buf\[36\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[19\]_A _490_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[116\] _587_/Y la_buf\[116\]/TE vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[104\]_A _372_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk2_buf_A _399_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] mprj_logic_high_inst/HI[379] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _629_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_A _365_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[21\]_A _620_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_655_ la_oen_mprj[56] vssd vssd vccd vccd _655_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[88\]_A _356_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_586_ la_data_out_mprj[115] vssd vssd vccd vccd _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vssd vccd vccd la_data_in_mprj[19]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _611_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_A _347_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__643__A la_oen_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_440_ mprj_dat_o_core[1] vssd vssd vccd vccd _440_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[15\] _614_/Y mprj_logic_high_inst/HI[217] vssd vssd vccd
+ vccd la_oen_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_13_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_371_ la_oen_mprj[103] vssd vssd vccd vccd _371_/Y sky130_fd_sc_hd__inv_2
XANTENNA__553__A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_638_ la_oen_mprj[39] vssd vssd vccd vccd _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_569_ la_data_out_mprj[98] vssd vssd vccd vccd _569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__463__A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A la_oen_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_A _469_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__373__A la_oen_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__548__A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_423_ mprj_adr_o_core[16] vssd vssd vccd vccd _423_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[21\]_A _460_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[42\] _513_/Y la_buf\[42\]/TE vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__einvp_8
X_354_ la_oen_mprj[86] vssd vssd vccd vccd _354_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vssd vccd vccd la_data_in_mprj[86]
+ sky130_fd_sc_hd__inv_8
XFILLER_24_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__458__A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] mprj_logic_high_inst/HI[361] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[12\]_A _451_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__368__A la_oen_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _606_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high_inst/HI[256] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[82\] _350_/Y mprj_logic_high_inst/HI[284] vssd vssd vccd
+ vccd la_oen_core[82] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[30\] _469_/Y mprj_dat_buf\[30\]/TE vssd vssd vccd vccd mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_406_ mprj_sel_o_core[3] vssd vssd vccd vccd _406_/Y sky130_fd_sc_hd__inv_2
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_337_ la_oen_mprj[69] vssd vssd vccd vccd _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] mprj_logic_high_inst/HI[409] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__651__A la_oen_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__561__A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vssd vccd vccd la_data_in_mprj[49]
+ sky130_fd_sc_hd__inv_8
XANTENNA__471__A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] mprj_logic_high_inst/HI[435] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__646__A la_oen_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[6\]_A _413_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2 vssd2 mprj2_logic_high
XFILLER_25_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__381__A la_oen_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[115\] _383_/Y mprj_logic_high_inst/HI[317] vssd vssd vccd
+ vccd la_oen_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_28_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[45\] _644_/Y mprj_logic_high_inst/HI[247] vssd vssd vccd
+ vccd la_oen_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_5_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__556__A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[109\] _580_/Y la_buf\[109\]/TE vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_26_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[102] sky130_fd_sc_hd__inv_8
XFILLER_23_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[1\] _440_/Y mprj_dat_buf\[1\]/TE vssd vssd vccd vccd mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_22_1400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf\[26\]/TE la_buf\[27\]/TE la_buf\[28\]/TE
+ la_buf\[29\]/TE la_buf\[30\]/TE la_buf\[31\]/TE la_buf\[32\]/TE la_buf\[33\]/TE
+ la_buf\[34\]/TE la_buf\[35\]/TE mprj_adr_buf\[0\]/TE la_buf\[36\]/TE la_buf\[37\]/TE
+ la_buf\[38\]/TE la_buf\[39\]/TE la_buf\[40\]/TE la_buf\[41\]/TE la_buf\[42\]/TE
+ la_buf\[43\]/TE la_buf\[44\]/TE la_buf\[45\]/TE mprj_adr_buf\[1\]/TE la_buf\[46\]/TE
+ la_buf\[47\]/TE la_buf\[48\]/TE la_buf\[49\]/TE la_buf\[50\]/TE la_buf\[51\]/TE
+ la_buf\[52\]/TE la_buf\[53\]/TE la_buf\[54\]/TE la_buf\[55\]/TE mprj_adr_buf\[2\]/TE
+ la_buf\[56\]/TE la_buf\[57\]/TE la_buf\[58\]/TE la_buf\[59\]/TE la_buf\[60\]/TE
+ la_buf\[61\]/TE la_buf\[62\]/TE la_buf\[63\]/TE la_buf\[64\]/TE la_buf\[65\]/TE
+ mprj_adr_buf\[3\]/TE la_buf\[66\]/TE la_buf\[67\]/TE la_buf\[68\]/TE la_buf\[69\]/TE
+ la_buf\[70\]/TE la_buf\[71\]/TE la_buf\[72\]/TE la_buf\[73\]/TE la_buf\[74\]/TE
+ la_buf\[75\]/TE mprj_adr_buf\[4\]/TE la_buf\[76\]/TE la_buf\[77\]/TE la_buf\[78\]/TE
+ la_buf\[79\]/TE la_buf\[80\]/TE la_buf\[81\]/TE la_buf\[82\]/TE la_buf\[83\]/TE
+ la_buf\[84\]/TE la_buf\[85\]/TE mprj_adr_buf\[5\]/TE la_buf\[86\]/TE la_buf\[87\]/TE
+ la_buf\[88\]/TE la_buf\[89\]/TE la_buf\[90\]/TE la_buf\[91\]/TE la_buf\[92\]/TE
+ la_buf\[93\]/TE la_buf\[94\]/TE la_buf\[95\]/TE mprj_adr_buf\[6\]/TE la_buf\[96\]/TE
+ la_buf\[97\]/TE la_buf\[98\]/TE la_buf\[99\]/TE la_buf\[100\]/TE la_buf\[101\]/TE
+ la_buf\[102\]/TE la_buf\[103\]/TE la_buf\[104\]/TE la_buf\[105\]/TE mprj_adr_buf\[7\]/TE
+ la_buf\[106\]/TE la_buf\[107\]/TE la_buf\[108\]/TE la_buf\[109\]/TE la_buf\[110\]/TE
+ la_buf\[111\]/TE la_buf\[112\]/TE la_buf\[113\]/TE la_buf\[114\]/TE la_buf\[115\]/TE
+ mprj_adr_buf\[8\]/TE la_buf\[116\]/TE la_buf\[117\]/TE la_buf\[118\]/TE la_buf\[119\]/TE
+ la_buf\[120\]/TE la_buf\[121\]/TE la_buf\[122\]/TE la_buf\[123\]/TE la_buf\[124\]/TE
+ la_buf\[125\]/TE mprj_adr_buf\[9\]/TE mprj_clk_buf/TE la_buf\[126\]/TE la_buf\[127\]/TE
+ mprj_logic_high_inst/HI[202] mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204]
+ mprj_logic_high_inst/HI[205] mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207]
+ mprj_logic_high_inst/HI[208] mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE
+ mprj_logic_high_inst/HI[210] mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212]
+ mprj_logic_high_inst/HI[213] mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215]
+ mprj_logic_high_inst/HI[216] mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218]
+ mprj_logic_high_inst/HI[219] mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220]
+ mprj_logic_high_inst/HI[221] mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223]
+ mprj_logic_high_inst/HI[224] mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226]
+ mprj_logic_high_inst/HI[227] mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229]
+ mprj_adr_buf\[12\]/TE mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231]
+ mprj_logic_high_inst/HI[232] mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234]
+ mprj_logic_high_inst/HI[235] mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237]
+ mprj_logic_high_inst/HI[238] mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE
+ mprj_logic_high_inst/HI[240] mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242]
+ mprj_logic_high_inst/HI[243] mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245]
+ mprj_logic_high_inst/HI[246] mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248]
+ mprj_logic_high_inst/HI[249] mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250]
+ mprj_logic_high_inst/HI[251] mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253]
+ mprj_logic_high_inst/HI[254] mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256]
+ mprj_logic_high_inst/HI[257] mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259]
+ mprj_adr_buf\[15\]/TE mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261]
+ mprj_logic_high_inst/HI[262] mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264]
+ mprj_logic_high_inst/HI[265] mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267]
+ mprj_logic_high_inst/HI[268] mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE
+ mprj_logic_high_inst/HI[270] mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272]
+ mprj_logic_high_inst/HI[273] mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275]
+ mprj_logic_high_inst/HI[276] mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278]
+ mprj_logic_high_inst/HI[279] mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280]
+ mprj_logic_high_inst/HI[281] mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283]
+ mprj_logic_high_inst/HI[284] mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286]
+ mprj_logic_high_inst/HI[287] mprj_logic_high_inst/HI[288] mprj_logic_high_inst/HI[289]
+ mprj_adr_buf\[18\]/TE mprj_logic_high_inst/HI[290] mprj_logic_high_inst/HI[291]
+ mprj_logic_high_inst/HI[292] mprj_logic_high_inst/HI[293] mprj_logic_high_inst/HI[294]
+ mprj_logic_high_inst/HI[295] mprj_logic_high_inst/HI[296] mprj_logic_high_inst/HI[297]
+ mprj_logic_high_inst/HI[298] mprj_logic_high_inst/HI[299] mprj_adr_buf\[19\]/TE
+ mprj_clk2_buf/TE mprj_logic_high_inst/HI[300] mprj_logic_high_inst/HI[301] mprj_logic_high_inst/HI[302]
+ mprj_logic_high_inst/HI[303] mprj_logic_high_inst/HI[304] mprj_logic_high_inst/HI[305]
+ mprj_logic_high_inst/HI[306] mprj_logic_high_inst/HI[307] mprj_logic_high_inst/HI[308]
+ mprj_logic_high_inst/HI[309] mprj_adr_buf\[20\]/TE mprj_logic_high_inst/HI[310]
+ mprj_logic_high_inst/HI[311] mprj_logic_high_inst/HI[312] mprj_logic_high_inst/HI[313]
+ mprj_logic_high_inst/HI[314] mprj_logic_high_inst/HI[315] mprj_logic_high_inst/HI[316]
+ mprj_logic_high_inst/HI[317] mprj_logic_high_inst/HI[318] mprj_logic_high_inst/HI[319]
+ mprj_adr_buf\[21\]/TE mprj_logic_high_inst/HI[320] mprj_logic_high_inst/HI[321]
+ mprj_logic_high_inst/HI[322] mprj_logic_high_inst/HI[323] mprj_logic_high_inst/HI[324]
+ mprj_logic_high_inst/HI[325] mprj_logic_high_inst/HI[326] mprj_logic_high_inst/HI[327]
+ mprj_logic_high_inst/HI[328] mprj_logic_high_inst/HI[329] mprj_adr_buf\[22\]/TE
+ user_to_mprj_in_gates\[0\]/B user_to_mprj_in_gates\[1\]/B user_to_mprj_in_gates\[2\]/B
+ user_to_mprj_in_gates\[3\]/B user_to_mprj_in_gates\[4\]/B user_to_mprj_in_gates\[5\]/B
+ user_to_mprj_in_gates\[6\]/B user_to_mprj_in_gates\[7\]/B user_to_mprj_in_gates\[8\]/B
+ user_to_mprj_in_gates\[9\]/B mprj_adr_buf\[23\]/TE mprj_logic_high_inst/HI[340]
+ mprj_logic_high_inst/HI[341] mprj_logic_high_inst/HI[342] mprj_logic_high_inst/HI[343]
+ mprj_logic_high_inst/HI[344] mprj_logic_high_inst/HI[345] mprj_logic_high_inst/HI[346]
+ mprj_logic_high_inst/HI[347] mprj_logic_high_inst/HI[348] mprj_logic_high_inst/HI[349]
+ mprj_adr_buf\[24\]/TE mprj_logic_high_inst/HI[350] mprj_logic_high_inst/HI[351]
+ mprj_logic_high_inst/HI[352] mprj_logic_high_inst/HI[353] mprj_logic_high_inst/HI[354]
+ mprj_logic_high_inst/HI[355] mprj_logic_high_inst/HI[356] mprj_logic_high_inst/HI[357]
+ mprj_logic_high_inst/HI[358] mprj_logic_high_inst/HI[359] mprj_adr_buf\[25\]/TE
+ mprj_logic_high_inst/HI[360] mprj_logic_high_inst/HI[361] mprj_logic_high_inst/HI[362]
+ mprj_logic_high_inst/HI[363] mprj_logic_high_inst/HI[364] mprj_logic_high_inst/HI[365]
+ mprj_logic_high_inst/HI[366] mprj_logic_high_inst/HI[367] mprj_logic_high_inst/HI[368]
+ mprj_logic_high_inst/HI[369] mprj_adr_buf\[26\]/TE mprj_logic_high_inst/HI[370]
+ mprj_logic_high_inst/HI[371] mprj_logic_high_inst/HI[372] mprj_logic_high_inst/HI[373]
+ mprj_logic_high_inst/HI[374] mprj_logic_high_inst/HI[375] mprj_logic_high_inst/HI[376]
+ mprj_logic_high_inst/HI[377] mprj_logic_high_inst/HI[378] mprj_logic_high_inst/HI[379]
+ mprj_adr_buf\[27\]/TE mprj_logic_high_inst/HI[380] mprj_logic_high_inst/HI[381]
+ mprj_logic_high_inst/HI[382] mprj_logic_high_inst/HI[383] mprj_logic_high_inst/HI[384]
+ mprj_logic_high_inst/HI[385] mprj_logic_high_inst/HI[386] mprj_logic_high_inst/HI[387]
+ mprj_logic_high_inst/HI[388] mprj_logic_high_inst/HI[389] mprj_adr_buf\[28\]/TE
+ mprj_logic_high_inst/HI[390] mprj_logic_high_inst/HI[391] mprj_logic_high_inst/HI[392]
+ mprj_logic_high_inst/HI[393] mprj_logic_high_inst/HI[394] mprj_logic_high_inst/HI[395]
+ mprj_logic_high_inst/HI[396] mprj_logic_high_inst/HI[397] mprj_logic_high_inst/HI[398]
+ mprj_logic_high_inst/HI[399] mprj_adr_buf\[29\]/TE mprj_cyc_buf/TE mprj_logic_high_inst/HI[400]
+ mprj_logic_high_inst/HI[401] mprj_logic_high_inst/HI[402] mprj_logic_high_inst/HI[403]
+ mprj_logic_high_inst/HI[404] mprj_logic_high_inst/HI[405] mprj_logic_high_inst/HI[406]
+ mprj_logic_high_inst/HI[407] mprj_logic_high_inst/HI[408] mprj_logic_high_inst/HI[409]
+ mprj_adr_buf\[30\]/TE mprj_logic_high_inst/HI[410] mprj_logic_high_inst/HI[411]
+ mprj_logic_high_inst/HI[412] mprj_logic_high_inst/HI[413] mprj_logic_high_inst/HI[414]
+ mprj_logic_high_inst/HI[415] mprj_logic_high_inst/HI[416] mprj_logic_high_inst/HI[417]
+ mprj_logic_high_inst/HI[418] mprj_logic_high_inst/HI[419] mprj_adr_buf\[31\]/TE
+ mprj_logic_high_inst/HI[420] mprj_logic_high_inst/HI[421] mprj_logic_high_inst/HI[422]
+ mprj_logic_high_inst/HI[423] mprj_logic_high_inst/HI[424] mprj_logic_high_inst/HI[425]
+ mprj_logic_high_inst/HI[426] mprj_logic_high_inst/HI[427] mprj_logic_high_inst/HI[428]
+ mprj_logic_high_inst/HI[429] mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431]
+ mprj_logic_high_inst/HI[432] mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434]
+ mprj_logic_high_inst/HI[435] mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437]
+ mprj_logic_high_inst/HI[438] mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440]
+ mprj_logic_high_inst/HI[441] mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443]
+ mprj_logic_high_inst/HI[444] mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446]
+ mprj_logic_high_inst/HI[447] mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449]
+ mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450] mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452]
+ mprj_logic_high_inst/HI[453] mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455]
+ mprj_logic_high_inst/HI[456] mprj_logic_high_inst/HI[457] mprj_pwrgood/A mprj_dat_buf\[3\]/TE
+ mprj_dat_buf\[4\]/TE mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE mprj_dat_buf\[7\]/TE
+ mprj_stb_buf/TE mprj_dat_buf\[8\]/TE mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE
+ mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE
+ mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE mprj_dat_buf\[17\]/TE mprj_we_buf/TE
+ mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE
+ mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE
+ mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE
+ mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE mprj_dat_buf\[31\]/TE la_buf\[0\]/TE
+ la_buf\[1\]/TE la_buf\[2\]/TE la_buf\[3\]/TE la_buf\[4\]/TE la_buf\[5\]/TE mprj_sel_buf\[1\]/TE
+ la_buf\[6\]/TE la_buf\[7\]/TE la_buf\[8\]/TE la_buf\[9\]/TE la_buf\[10\]/TE la_buf\[11\]/TE
+ la_buf\[12\]/TE la_buf\[13\]/TE la_buf\[14\]/TE la_buf\[15\]/TE mprj_sel_buf\[2\]/TE
+ la_buf\[16\]/TE la_buf\[17\]/TE la_buf\[18\]/TE la_buf\[19\]/TE la_buf\[20\]/TE
+ la_buf\[21\]/TE la_buf\[22\]/TE la_buf\[23\]/TE la_buf\[24\]/TE la_buf\[25\]/TE
+ mprj_sel_buf\[3\]/TE vccd1 vssd1 mprj_logic_high
XFILLER_27_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__376__A la_oen_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_654_ la_oen_mprj[55] vssd vssd vccd vccd _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[72\] _543_/Y la_buf\[72\]/TE vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__einvp_8
X_585_ la_data_out_mprj[114] vssd vssd vccd vccd _585_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] mprj_logic_high_inst/HI[391] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_B user_to_mprj_in_gates\[6\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_370_ la_oen_mprj[102] vssd vssd vccd vccd _370_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_637_ la_oen_mprj[38] vssd vssd vccd vccd _637_/Y sky130_fd_sc_hd__inv_2
X_568_ la_data_out_mprj[97] vssd vssd vccd vccd _568_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vssd vccd vccd la_data_in_mprj[31]
+ sky130_fd_sc_hd__inv_8
X_499_ la_data_out_mprj[28] vssd vssd vccd vccd _499_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__654__A la_oen_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_422_ mprj_adr_o_core[15] vssd vssd vccd vccd _422_/Y sky130_fd_sc_hd__inv_2
XANTENNA__564__A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_353_ la_oen_mprj[85] vssd vssd vccd vccd _353_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[35\] _506_/Y la_buf\[35\]/TE vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_6_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vssd vccd vccd la_data_in_mprj[79]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__474__A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] mprj_logic_high_inst/HI[354] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__649__A la_oen_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XPHY_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__384__A la_oen_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[75\] _343_/Y mprj_logic_high_inst/HI[277] vssd vssd vccd
+ vccd la_oen_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_8_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[23\] _462_/Y mprj_dat_buf\[23\]/TE vssd vssd vccd vccd mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__559__A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_405_ mprj_sel_o_core[2] vssd vssd vccd vccd _405_/Y sky130_fd_sc_hd__inv_2
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_336_ la_oen_mprj[68] vssd vssd vccd vccd _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__469__A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__379__A la_oen_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xpowergood_check mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vdda1 vssa1 vdda2
+ vssa2 mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] mprj_logic_high_inst/HI[421] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high_inst/HI[246] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_sel_buf\[0\]_A _403_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[108\] _376_/Y mprj_logic_high_inst/HI[310] vssd vssd vccd
+ vccd la_oen_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_28_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[38\] _637_/Y mprj_logic_high_inst/HI[240] vssd vssd vccd
+ vccd la_oen_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_16_459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__572__A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[82\]_TE la_buf\[82\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_A _440_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vssd vccd vccd la_data_in_mprj[61]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__482__A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A la_oen_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__392__A la_oen_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[81\]_A user_to_mprj_in_gates\[81\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_B mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__567__A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_653_ la_oen_mprj[54] vssd vssd vccd vccd _653_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_584_ la_data_out_mprj[113] vssd vssd vccd vccd _584_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[65\] _536_/Y la_buf\[65\]/TE vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_16_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[87\]_B mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[29\] _436_/Y mprj_adr_buf\[29\]/TE vssd vssd vccd vccd mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[121\] _592_/Y la_buf\[121\]/TE vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__einvp_8
XFILLER_12_1669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[72\]_A user_to_mprj_in_gates\[72\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_B mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__477__A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] mprj_logic_high_inst/HI[384] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[78\]_B mprj_logic_high_inst/HI[408] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[110\]_A user_to_mprj_in_gates\[110\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[63\]_A user_to_mprj_in_gates\[63\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__387__A la_oen_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_B mprj_logic_high_inst/HI[399] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_636_ la_oen_mprj[37] vssd vssd vccd vccd _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_567_ la_data_out_mprj[96] vssd vssd vccd vccd _567_/Y sky130_fd_sc_hd__inv_2
X_498_ la_data_out_mprj[27] vssd vssd vccd vccd _498_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[94\]_A _565_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vssd vccd vccd la_data_in_mprj[24]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[85\]_A _556_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_421_ mprj_adr_o_core[14] vssd vssd vccd vccd _421_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[2\] _601_/Y mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd la_oen_core[2] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[20\] _619_/Y mprj_logic_high_inst/HI[222] vssd vssd vccd
+ vccd la_oen_core[20] sky130_fd_sc_hd__einvp_8
X_352_ la_oen_mprj[84] vssd vssd vccd vccd _352_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[126\]_B mprj_logic_high_inst/HI[456] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_A _547_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__580__A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _499_/Y la_buf\[28\]/TE vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__einvp_8
XFILLER_10_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_619_ la_oen_mprj[20] vssd vssd vccd vccd _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_B mprj_logic_high_inst/HI[447] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[67\]_A _538_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] mprj_logic_high_inst/HI[347] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__490__A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[108\]_B mprj_logic_high_inst/HI[438] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[58\]_A _529_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[68\] _336_/Y mprj_logic_high_inst/HI[270] vssd vssd vccd
+ vccd la_oen_core[68] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[16\] _455_/Y mprj_dat_buf\[16\]/TE vssd vssd vccd vccd mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__575__A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_404_ mprj_sel_o_core[1] vssd vssd vccd vccd _404_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[49\]_A _520_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_335_ la_oen_mprj[67] vssd vssd vccd vccd _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[11\] _418_/Y mprj_adr_buf\[11\]/TE vssd vssd vccd vccd mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[125] sky130_fd_sc_hd__inv_8
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vssd vccd vccd la_data_in_mprj[91]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__485__A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[125\]_A _393_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[60\]_A _659_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__395__A la_oen_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _650_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[116\]_A _384_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[95\] _566_/Y la_buf\[95\]/TE vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_19_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[42\]_A _641_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _375_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] mprj_logic_high_inst/HI[414] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _632_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[24\]_A _623_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high_inst/HI[314] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[6\] _477_/Y la_buf\[6\]/TE vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__einvp_8
Xla_buf\[10\] _481_/Y la_buf\[10\]/TE vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_26_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[3\] _410_/Y mprj_adr_buf\[3\]/TE vssd vssd vccd vccd mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[20\]_A _427_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vssd vccd vccd la_data_in_mprj[54]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _614_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] mprj_logic_high_inst/HI[440] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[11\]_A _418_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[120\] _388_/Y mprj_logic_high_inst/HI[322] vssd vssd vccd
+ vccd la_oen_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_1_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _404_/Y mprj_sel_buf\[1\]/TE vssd vssd vccd vccd mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[50\] _649_/Y mprj_logic_high_inst/HI[252] vssd vssd vccd
+ vccd la_oen_core[50] sky130_fd_sc_hd__einvp_8
XFILLER_5_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_652_ la_oen_mprj[53] vssd vssd vccd vccd _652_/Y sky130_fd_sc_hd__inv_2
X_583_ la_data_out_mprj[112] vssd vssd vccd vccd _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__583__A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[58\] _529_/Y la_buf\[58\]/TE vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__einvp_8
XPHY_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[114\] _585_/Y la_buf\[114\]/TE vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_3_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] mprj_logic_high_inst/HI[377] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__493__A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] user_to_mprj_in_gates\[9\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[57\]_TE mprj_logic_high_inst/HI[259] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _366_/Y mprj_logic_high_inst/HI[300] vssd vssd vccd
+ vccd la_oen_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_1_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__578__A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_635_ la_oen_mprj[36] vssd vssd vccd vccd _635_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[24\]_A _463_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_566_ la_data_out_mprj[95] vssd vssd vccd vccd _566_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_497_ la_data_out_mprj[26] vssd vssd vccd vccd _497_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vssd vccd vccd la_data_in_mprj[17]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_TE la_buf\[95\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__488__A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_A _454_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_420_ mprj_adr_o_core[13] vssd vssd vccd vccd _420_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[13\] _612_/Y mprj_logic_high_inst/HI[215] vssd vssd vccd
+ vccd la_oen_core[13] sky130_fd_sc_hd__einvp_8
X_351_ la_oen_mprj[83] vssd vssd vccd vccd _351_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vssd vccd vccd la_data_in_mprj[9]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_618_ la_oen_mprj[19] vssd vssd vccd vccd _618_/Y sky130_fd_sc_hd__inv_2
X_549_ la_data_out_mprj[78] vssd vssd vccd vccd _549_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_403_ mprj_sel_o_core[0] vssd vssd vccd vccd _403_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[2\]_A _473_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[40\] _511_/Y la_buf\[40\]/TE vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__einvp_8
X_334_ la_oen_mprj[66] vssd vssd vccd vccd _334_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__591__A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[118] sky130_fd_sc_hd__inv_8
XFILLER_2_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vssd vccd vccd la_data_in_mprj[84]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[120\]_TE la_buf\[120\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_A _416_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _348_/Y mprj_logic_high_inst/HI[282] vssd vssd vccd
+ vccd la_oen_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_11_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__586__A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[88\] _559_/Y la_buf\[88\]/TE vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_21_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[0\]_A user_to_mprj_in_gates\[0\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] mprj_logic_high_inst/HI[407] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__496__A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[29\]_TE la_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vssd vccd vccd la_data_in_mprj[47]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_2111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] mprj_logic_high_inst/HI[433] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[113\] _381_/Y mprj_logic_high_inst/HI[315] vssd vssd vccd
+ vccd la_oen_core[113] sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _399_/Y mprj_clk2_buf/TE vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[9\]_B user_to_mprj_in_gates\[9\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_651_ la_oen_mprj[52] vssd vssd vccd vccd _651_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[43\] _642_/Y mprj_logic_high_inst/HI[245] vssd vssd vccd
+ vccd la_oen_core[43] sky130_fd_sc_hd__einvp_8
XFILLER_25_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_582_ la_data_out_mprj[111] vssd vssd vccd vccd _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[107\] _578_/Y la_buf\[107\]/TE vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_27_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[100] sky130_fd_sc_hd__inv_8
XFILLER_3_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_634_ la_oen_mprj[35] vssd vssd vccd vccd _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__594__A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[70\] _541_/Y la_buf\[70\]/TE vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_2_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_565_ la_data_out_mprj[94] vssd vssd vccd vccd _565_/Y sky130_fd_sc_hd__inv_2
X_496_ la_data_out_mprj[25] vssd vssd vccd vccd _496_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_350_ la_oen_mprj[82] vssd vssd vccd vccd _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__589__A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_617_ la_oen_mprj[18] vssd vssd vccd vccd _617_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_548_ la_data_out_mprj[77] vssd vssd vccd vccd _548_/Y sky130_fd_sc_hd__inv_2
X_479_ la_data_out_mprj[8] vssd vssd vccd vccd _479_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__499__A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_402_ mprj_we_o_core vssd vssd vccd vccd _402_/Y sky130_fd_sc_hd__inv_2
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ la_oen_mprj[65] vssd vssd vccd vccd _333_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[33\] _504_/Y la_buf\[33\]/TE vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__einvp_8
XFILLER_13_1574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vssd vccd vccd la_data_in_mprj[77]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] mprj_logic_high_inst/HI[352] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_A _406_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[50\]_B mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[73\] _341_/Y mprj_logic_high_inst/HI[275] vssd vssd vccd
+ vccd la_oen_core[73] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[21\] _460_/Y mprj_dat_buf\[21\]/TE vssd vssd vccd vccd mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[4\]_A _443_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[41\]_B mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_B mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[99\]_B mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[120\]_A _591_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[84\]_A user_to_mprj_in_gates\[84\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[23\]_B mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__597__A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_TE la_buf\[110\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[122\]_A user_to_mprj_in_gates\[122\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[111\]_A _582_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[75\]_A user_to_mprj_in_gates\[75\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[113\]_A user_to_mprj_in_gates\[113\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[102\]_A _573_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _374_/Y mprj_logic_high_inst/HI[308] vssd vssd vccd
+ vccd la_oen_core[106] sky130_fd_sc_hd__einvp_8
X_650_ la_oen_mprj[51] vssd vssd vccd vccd _650_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[36\] _635_/Y mprj_logic_high_inst/HI[238] vssd vssd vccd
+ vccd la_oen_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_5_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_581_ la_data_out_mprj[110] vssd vssd vccd vccd _581_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[30\]_A _501_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[97\]_A _568_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[21\]_A _492_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_A _559_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[39\]_A user_to_mprj_in_gates\[39\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[12\]_A _483_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_51 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_633_ la_oen_mprj[34] vssd vssd vccd vccd _633_/Y sky130_fd_sc_hd__inv_2
X_564_ la_data_out_mprj[93] vssd vssd vccd vccd _564_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[79\]_A _550_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[63\] _534_/Y la_buf\[63\]/TE vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__einvp_8
X_495_ la_data_out_mprj[24] vssd vssd vccd vccd _495_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[27\] _434_/Y mprj_adr_buf\[27\]/TE vssd vssd vccd vccd mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] mprj_logic_high_inst/HI[382] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[90\]_A _358_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _349_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_616_ la_oen_mprj[17] vssd vssd vccd vccd _616_/Y sky130_fd_sc_hd__inv_2
X_547_ la_data_out_mprj[76] vssd vssd vccd vccd _547_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_478_ la_data_out_mprj[7] vssd vssd vccd vccd _478_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[72\]_A _340_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vssd vccd vccd la_data_in_mprj[22]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _331_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[0\] _599_/Y mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd la_oen_core[0] sky130_fd_sc_hd__einvp_8
X_401_ mprj_stb_o_core vssd vssd vccd vccd _401_/Y sky130_fd_sc_hd__inv_2
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ la_oen_mprj[64] vssd vssd vccd vccd _332_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _653_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_A _387_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[26\] _497_/Y la_buf\[26\]/TE vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_26_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] mprj_logic_high_inst/HI[345] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _644_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] mprj_logic_high_inst/HI[456] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _635_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _334_/Y mprj_logic_high_inst/HI[268] vssd vssd vccd
+ vccd la_oen_core[66] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[14\] _453_/Y mprj_dat_buf\[14\]/TE vssd vssd vccd vccd mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[52\]_TE la_buf\[52\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[27\]_A _626_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[123] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[23\]_A _430_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_A _599_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_A _617_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_A _421_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[93\] _564_/Y la_buf\[93\]/TE vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_5_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[98\]_TE la_buf\[98\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] mprj_logic_high_inst/HI[412] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_580_ la_data_out_mprj[109] vssd vssd vccd vccd _580_/Y sky130_fd_sc_hd__inv_2
XPHY_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_oen_buffers\[29\] _628_/Y mprj_logic_high_inst/HI[231] vssd vssd vccd
+ vccd la_oen_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_25_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[4\] _475_/Y la_buf\[4\]/TE vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_4_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__401__A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[1\] _408_/Y mprj_adr_buf\[1\]/TE vssd vssd vccd vccd mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[27\]_A _466_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vssd vccd vccd la_data_in_mprj[52]
+ sky130_fd_sc_hd__inv_8
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_A _457_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_632_ la_oen_mprj[33] vssd vssd vccd vccd _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_563_ la_data_out_mprj[92] vssd vssd vccd vccd _563_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_494_ la_data_out_mprj[23] vssd vssd vccd vccd _494_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[56\] _527_/Y la_buf\[56\]/TE vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_9_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[112\] _583_/Y la_buf\[112\]/TE vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_5_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] mprj_logic_high_inst/HI[375] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] user_to_mprj_in_gates\[7\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[96\] _364_/Y mprj_logic_high_inst/HI[298] vssd vssd vccd
+ vccd la_oen_core[96] sky130_fd_sc_hd__einvp_8
XFILLER_6_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[5\]_A _476_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_615_ la_oen_mprj[16] vssd vssd vccd vccd _615_/Y sky130_fd_sc_hd__inv_2
X_546_ la_data_out_mprj[75] vssd vssd vccd vccd _546_/Y sky130_fd_sc_hd__inv_2
X_477_ la_data_out_mprj[6] vssd vssd vccd vccd _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vssd vccd vccd la_data_in_mprj[15]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_pwrgood mprj2_pwrgood/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_28_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_400_ mprj_cyc_o_core vssd vssd vccd vccd _400_/Y sky130_fd_sc_hd__inv_2
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[11\] _610_/Y mprj_logic_high_inst/HI[213] vssd vssd vccd
+ vccd la_oen_core[11] sky130_fd_sc_hd__einvp_8
X_331_ la_oen_mprj[63] vssd vssd vccd vccd _331_/Y sky130_fd_sc_hd__inv_2
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vssd vccd vccd la_data_in_mprj[7]
+ sky130_fd_sc_hd__inv_8
XFILLER_10_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[19\] _490_/Y la_buf\[19\]/TE vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_13_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_529_ la_data_out_mprj[58] vssd vssd vccd vccd _529_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] mprj_logic_high_inst/HI[449] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[59\] _658_/Y mprj_logic_high_inst/HI[261] vssd vssd vccd
+ vccd la_oen_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_21_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[116] sky130_fd_sc_hd__inv_8
XFILLER_6_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vssd vccd vccd la_data_in_mprj[82]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_A _396_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_1200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[86\] _557_/Y la_buf\[86\]/TE vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_5_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] mprj_logic_high_inst/HI[405] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[42\]_TE la_buf\[42\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vssd vccd vccd la_data_in_mprj[45]
+ sky130_fd_sc_hd__inv_8
XPHY_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] mprj_logic_high_inst/HI[431] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_10_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__502__A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[111\] _379_/Y mprj_logic_high_inst/HI[313] vssd vssd vccd
+ vccd la_oen_core[111] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[41\] _640_/Y mprj_logic_high_inst/HI[243] vssd vssd vccd
+ vccd la_oen_core[41] sky130_fd_sc_hd__einvp_8
X_631_ la_oen_mprj[32] vssd vssd vccd vccd _631_/Y sky130_fd_sc_hd__inv_2
X_562_ la_data_out_mprj[91] vssd vssd vccd vccd _562_/Y sky130_fd_sc_hd__inv_2
X_493_ la_data_out_mprj[22] vssd vssd vccd vccd _493_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[49\] _520_/Y la_buf\[49\]/TE vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_16_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__412__A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[105\] _576_/Y la_buf\[105\]/TE vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_23_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] mprj_logic_high_inst/HI[368] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[80\]_B mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[89\] _357_/Y mprj_logic_high_inst/HI[291] vssd vssd vccd
+ vccd la_oen_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_2_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_614_ la_oen_mprj[15] vssd vssd vccd vccd _614_/Y sky130_fd_sc_hd__inv_2
X_545_ la_data_out_mprj[74] vssd vssd vccd vccd _545_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__407__A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_476_ la_data_out_mprj[5] vssd vssd vccd vccd _476_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B mprj_logic_high_inst/HI[401] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_B mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ la_oen_mprj[62] vssd vssd vccd vccd _330_/Y sky130_fd_sc_hd__inv_2
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[53\]_B mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[113\]_TE la_buf\[113\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[7\]_A _446_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_528_ la_data_out_mprj[57] vssd vssd vccd vccd _528_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_459_ mprj_dat_o_core[20] vssd vssd vccd vccd _459_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[44\]_B mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__600__A la_oen_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[96\]_A user_to_mprj_in_gates\[96\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[35\]_B mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__510__A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[31\] _502_/Y la_buf\[31\]/TE vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[123\]_A _594_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[26\]_B mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_B mprj_logic_high_inst/HI[440] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[60\]_A _531_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[109] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vssd vccd vccd la_data_in_mprj[75]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] mprj_logic_high_inst/HI[350] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[114\]_A _585_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[17\]_B mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B mprj_logic_high_inst/HI[431] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[78\]_A user_to_mprj_in_gates\[78\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_A _522_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[8\] _447_/Y mprj_dat_buf\[8\]/TE vssd vssd vccd vccd mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__330__A la_oen_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[105\]_A _576_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__505__A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[42\]_A _513_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[71\] _339_/Y mprj_logic_high_inst/HI[273] vssd vssd vccd
+ vccd la_oen_core[71] sky130_fd_sc_hd__einvp_8
XFILLER_23_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[79\] _550_/Y la_buf\[79\]/TE vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_27_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__415__A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[33\]_A _504_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] mprj_logic_high_inst/HI[398] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[24\]_A _495_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[15\]_A _486_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[100\]_A _368_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vssd vccd vccd la_data_in_mprj[38]
+ sky130_fd_sc_hd__inv_8
XPHY_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[93\]_A _361_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[104\] _372_/Y mprj_logic_high_inst/HI[306] vssd vssd vccd
+ vccd la_oen_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_28_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_630_ la_oen_mprj[31] vssd vssd vccd vccd _630_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[34\] _633_/Y mprj_logic_high_inst/HI[236] vssd vssd vccd
+ vccd la_oen_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_22_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_561_ la_data_out_mprj[90] vssd vssd vccd vccd _561_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_492_ la_data_out_mprj[21] vssd vssd vccd vccd _492_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[84\]_A _352_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[32\]_TE la_buf\[32\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_A _343_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A la_oen_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_A _334_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__513__A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_613_ la_oen_mprj[14] vssd vssd vccd vccd _613_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_544_ la_data_out_mprj[73] vssd vssd vccd vccd _544_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[61\] _532_/Y la_buf\[61\]/TE vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_18_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_475_ la_data_out_mprj[4] vssd vssd vccd vccd _475_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _656_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[25\] _432_/Y mprj_adr_buf\[25\]/TE vssd vssd vccd vccd mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__423__A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] mprj_logic_high_inst/HI[380] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _647_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__333__A la_oen_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[78\]_TE la_buf\[78\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__508__A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[39\]_A _638_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__418__A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_527_ la_data_out_mprj[56] vssd vssd vccd vccd _527_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_458_ mprj_dat_o_core[19] vssd vssd vccd vccd _458_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_389_ la_oen_mprj[121] vssd vssd vccd vccd _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vssd vccd vccd la_data_in_mprj[20]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] mprj_logic_high_inst/HI[428] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[26\]_A _433_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _602_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[17\]_A _424_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[24\] _495_/Y la_buf\[24\]/TE vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__einvp_8
XFILLER_11_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vssd vccd vccd la_data_in_mprj[68]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] mprj_logic_high_inst/HI[343] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__611__A la_oen_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] mprj_logic_high_inst/HI[454] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_TE la_buf\[103\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__521__A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[64\] _332_/Y mprj_logic_high_inst/HI[266] vssd vssd vccd
+ vccd la_oen_core[64] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[12\] _451_/Y mprj_dat_buf\[12\]/TE vssd vssd vccd vccd mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_cyc_buf_A _400_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__431__A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[121] sky130_fd_sc_hd__inv_8
XFILLER_3_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[126\]_TE la_buf\[126\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__606__A la_oen_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[2\]_A _409_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__341__A la_oen_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__516__A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[91\] _562_/Y la_buf\[91\]/TE vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_15_230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__426__A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] mprj_logic_high_inst/HI[410] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__336__A la_oen_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_560_ la_data_out_mprj[89] vssd vssd vccd vccd _560_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[27\] _626_/Y mprj_logic_high_inst/HI[229] vssd vssd vccd
+ vccd la_oen_core[27] sky130_fd_sc_hd__einvp_8
X_491_ la_data_out_mprj[20] vssd vssd vccd vccd _491_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[9\] _608_/Y mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd la_oen_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_25_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[2\] _473_/Y la_buf\[2\]/TE vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_48 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[8\]_A _479_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vssd vccd vccd la_data_in_mprj[50]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[2\]_B user_to_mprj_in_gates\[2\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_612_ la_oen_mprj[13] vssd vssd vccd vccd _612_/Y sky130_fd_sc_hd__inv_2
X_543_ la_data_out_mprj[72] vssd vssd vccd vccd _543_/Y sky130_fd_sc_hd__inv_2
X_474_ la_data_out_mprj[3] vssd vssd vccd vccd _474_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[54\] _525_/Y la_buf\[54\]/TE vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_9_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[18\] _425_/Y mprj_adr_buf\[18\]/TE vssd vssd vccd vccd mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[110\] _581_/Y la_buf\[110\]/TE vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_9_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vssd vccd vccd la_data_in_mprj[98]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] mprj_logic_high_inst/HI[373] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A la_oen_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] user_to_mprj_in_gates\[5\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__524__A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[94\] _362_/Y mprj_logic_high_inst/HI[296] vssd vssd vccd
+ vccd la_oen_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_2_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_526_ la_data_out_mprj[55] vssd vssd vccd vccd _526_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_457_ mprj_dat_o_core[18] vssd vssd vccd vccd _457_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_388_ la_oen_mprj[120] vssd vssd vccd vccd _388_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_9_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__434__A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vssd vccd vccd la_data_in_mprj[13]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__609__A la_oen_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__344__A la_oen_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[45\]_TE la_buf\[45\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__519__A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vssd vccd vccd la_data_in_mprj[5]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[17\] _488_/Y la_buf\[17\]/TE vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_26_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__429__A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_509_ la_data_out_mprj[38] vssd vssd vccd vccd _509_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] mprj_logic_high_inst/HI[447] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__339__A la_oen_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[127\] _395_/Y mprj_logic_high_inst/HI[329] vssd vssd vccd
+ vccd la_oen_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[57\] _656_/Y mprj_logic_high_inst/HI[259] vssd vssd vccd
+ vccd la_oen_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_25_1770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[114] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vssd vccd vccd la_data_in_mprj[80]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__622__A la_oen_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__532__A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[84\] _555_/Y la_buf\[84\]/TE vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_15_242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__442__A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] mprj_logic_high_inst/HI[403] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__617__A la_oen_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[92\]_B mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__352__A la_oen_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_490_ la_data_out_mprj[19] vssd vssd vccd vccd _490_/Y sky130_fd_sc_hd__inv_2
XANTENNA__527__A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[83\]_B mprj_logic_high_inst/HI[413] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_TE la_buf\[116\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vssd vccd vccd la_data_in_mprj[43]
+ sky130_fd_sc_hd__inv_8
XPHY_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[74\]_B mprj_logic_high_inst/HI[404] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[63\]_TE mprj_logic_high_inst/HI[265] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__347__A la_oen_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[65\]_B mprj_logic_high_inst/HI[395] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_611_ la_oen_mprj[12] vssd vssd vccd vccd _611_/Y sky130_fd_sc_hd__inv_2
X_542_ la_data_out_mprj[71] vssd vssd vccd vccd _542_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_473_ la_data_out_mprj[2] vssd vssd vccd vccd _473_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _518_/Y la_buf\[47\]/TE vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[56\]_B mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[90\]_A _561_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _574_/Y la_buf\[103\]/TE vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_9_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] mprj_logic_high_inst/HI[366] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[47\]_B mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[81\]_A _552_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__630__A la_oen_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[99\]_A user_to_mprj_in_gates\[99\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[38\]_B mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_B mprj_logic_high_inst/HI[452] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[72\]_A _543_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _355_/Y mprj_logic_high_inst/HI[289] vssd vssd vccd
+ vccd la_oen_core[87] sky130_fd_sc_hd__einvp_8
XANTENNA__540__A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_525_ la_data_out_mprj[54] vssd vssd vccd vccd _525_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_456_ mprj_dat_o_core[17] vssd vssd vccd vccd _456_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[126\]_A _597_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_387_ la_oen_mprj[119] vssd vssd vccd vccd _387_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[113\]_B mprj_logic_high_inst/HI[443] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_B mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[30\] _437_/Y mprj_adr_buf\[30\]/TE vssd vssd vccd vccd mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[63\]_A _534_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__450__A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[117\]_A _588_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__625__A la_oen_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B mprj_logic_high_inst/HI[434] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_A _525_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__360__A la_oen_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_A _401_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[119\]_A user_to_mprj_in_gates\[119\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[108\]_A _579_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__535__A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[45\]_A _516_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_508_ la_data_out_mprj[37] vssd vssd vccd vccd _508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__445__A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_439_ mprj_dat_o_core[0] vssd vssd vccd vccd _439_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[36\]_A _507_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_A _389_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__355__A la_oen_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[27\]_A _498_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[112\]_A _380_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[18\]_A _489_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[103\]_A _371_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[107] sky130_fd_sc_hd__inv_8
XFILLER_4_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vssd vccd vccd la_data_in_mprj[73]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[35\]_TE la_buf\[35\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _445_/Y mprj_dat_buf\[6\]/TE vssd vssd vccd vccd mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_25_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[96\]_A _364_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _619_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[77\] _548_/Y la_buf\[77\]/TE vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_28_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[87\]_A _355_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _610_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] mprj_logic_high_inst/HI[396] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[78\]_A _346_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__633__A la_oen_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[69\]_A _337_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vssd vccd vccd la_data_in_mprj[36]
+ sky130_fd_sc_hd__inv_8
XPHY_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__453__A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__628__A la_oen_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__363__A la_oen_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[102\] _370_/Y mprj_logic_high_inst/HI[304] vssd vssd vccd
+ vccd la_oen_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_4_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_610_ la_oen_mprj[11] vssd vssd vccd vccd _610_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ la_data_out_mprj[70] vssd vssd vccd vccd _541_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[32\] _631_/Y mprj_logic_high_inst/HI[234] vssd vssd vccd
+ vccd la_oen_core[32] sky130_fd_sc_hd__einvp_8
X_472_ la_data_out_mprj[1] vssd vssd vccd vccd _472_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_A _459_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_A _450_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] mprj_logic_high_inst/HI[359] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_A _436_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A la_oen_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _605_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[106\]_TE la_buf\[106\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _467_/Y mprj_dat_buf\[28\]/TE vssd vssd vccd vccd mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_524_ la_data_out_mprj[53] vssd vssd vccd vccd _524_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_455_ mprj_dat_o_core[16] vssd vssd vccd vccd _455_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_TE mprj_logic_high_inst/HI[255] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_386_ la_oen_mprj[118] vssd vssd vccd vccd _386_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_adr_buf\[23\] _430_/Y mprj_adr_buf\[23\]/TE vssd vssd vccd vccd mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__641__A la_oen_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[91\]_TE la_buf\[91\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__551__A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_507_ la_data_out_mprj[36] vssd vssd vccd vccd _507_/Y sky130_fd_sc_hd__inv_2
X_438_ mprj_adr_o_core[31] vssd vssd vccd vccd _438_/Y sky130_fd_sc_hd__inv_2
X_369_ la_oen_mprj[101] vssd vssd vccd vccd _369_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__461__A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] mprj_logic_high_inst/HI[426] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__636__A la_oen_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[5\]_A _412_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__371__A la_oen_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[22\] _493_/Y la_buf\[22\]/TE vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__einvp_8
XFILLER_13_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vssd vccd vccd la_data_in_mprj[66]
+ sky130_fd_sc_hd__inv_8
XANTENNA__456__A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] mprj_logic_high_inst/HI[341] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] mprj_logic_high_inst/HI[452] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__366__A la_oen_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[62\] _330_/Y mprj_logic_high_inst/HI[264] vssd vssd vccd
+ vccd la_oen_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_27_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[10\] _449_/Y mprj_dat_buf\[10\]/TE vssd vssd vccd vccd mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[126\] _597_/Y la_buf\[126\]/TE vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_10_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] mprj_logic_high_inst/HI[389] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_B user_to_mprj_in_gates\[5\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vssd vccd vccd la_data_in_mprj[29]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A la_oen_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_540_ la_data_out_mprj[69] vssd vssd vccd vccd _540_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[25\] _624_/Y mprj_logic_high_inst/HI[227] vssd vssd vccd
+ vccd la_oen_core[25] sky130_fd_sc_hd__einvp_8
X_471_ la_data_out_mprj[0] vssd vssd vccd vccd _471_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[7\] _606_/Y mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd la_oen_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_26_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__554__A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xla_buf\[0\] _471_/Y la_buf\[0\]/TE vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_5_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__464__A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__639__A la_oen_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__374__A la_oen_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_17_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__549__A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_523_ la_data_out_mprj[52] vssd vssd vccd vccd _523_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_454_ mprj_dat_o_core[15] vssd vssd vccd vccd _454_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[52\] _523_/Y la_buf\[52\]/TE vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__einvp_8
X_385_ la_oen_mprj[117] vssd vssd vccd vccd _385_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[16\] _423_/Y mprj_adr_buf\[16\]/TE vssd vssd vccd vccd mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vssd vccd vccd la_data_in_mprj[96]
+ sky130_fd_sc_hd__inv_8
XFILLER_27_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_rstn_buf _396_/Y mprj_rstn_buf/TE vssd vssd vccd vccd user_resetn sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] mprj_logic_high_inst/HI[371] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] user_to_mprj_in_gates\[3\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__369__A la_oen_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[92\] _360_/Y mprj_logic_high_inst/HI[294] vssd vssd vccd
+ vccd la_oen_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_24_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_506_ la_data_out_mprj[35] vssd vssd vccd vccd _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_437_ mprj_adr_o_core[30] vssd vssd vccd vccd _437_/Y sky130_fd_sc_hd__inv_2
X_368_ la_oen_mprj[100] vssd vssd vccd vccd _368_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vssd vccd vccd la_data_in_mprj[11]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] mprj_logic_high_inst/HI[419] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__652__A la_oen_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high_inst/HI[245] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_cyc_buf _400_/Y mprj_cyc_buf/TE vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
XFILLER_15_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vssd vccd vccd la_data_in_mprj[3]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__562__A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[15\] _486_/Y la_buf\[15\]/TE vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _439_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[8\] _415_/Y mprj_adr_buf\[8\]/TE vssd vssd vccd vccd mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vssd vccd vccd la_data_in_mprj[59]
+ sky130_fd_sc_hd__inv_8
XANTENNA__472__A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[81\]_TE la_buf\[81\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] mprj_logic_high_inst/HI[445] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__647__A la_oen_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[95\]_B mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__382__A la_oen_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[125\] _393_/Y mprj_logic_high_inst/HI[327] vssd vssd vccd
+ vccd la_oen_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_0_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[55\] _654_/Y mprj_logic_high_inst/HI[257] vssd vssd vccd
+ vccd la_oen_core[55] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[80\]_A user_to_mprj_in_gates\[80\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__557__A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_B mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[119\] _590_/Y la_buf\[119\]/TE vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_3_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[112] sky130_fd_sc_hd__inv_8
XFILLER_6_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[10\]_B mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__467__A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B mprj_logic_high_inst/HI[407] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__377__A la_oen_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[68\]_B mprj_logic_high_inst/HI[398] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[82\] _553_/Y la_buf\[82\]/TE vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_1_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[93\]_A _564_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[44\]_A user_to_mprj_in_gates\[44\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] mprj_logic_high_inst/HI[401] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[84\]_A _555_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__660__A la_oen_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_470_ mprj_dat_o_core[31] vssd vssd vccd vccd _470_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[18\] _617_/Y mprj_logic_high_inst/HI[220] vssd vssd vccd
+ vccd la_oen_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_25_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_B mprj_logic_high_inst/HI[455] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[75\]_A _546_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_599_ la_oen_mprj[0] vssd vssd vccd vccd _599_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vssd vccd vccd la_data_in_mprj[41]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[116\]_B mprj_logic_high_inst/HI[446] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[66\]_A _537_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__480__A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A la_oen_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[107\]_B mprj_logic_high_inst/HI[437] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[57\]_A _528_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__390__A la_oen_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_522_ la_data_out_mprj[51] vssd vssd vccd vccd _522_/Y sky130_fd_sc_hd__inv_2
X_453_ mprj_dat_o_core[14] vssd vssd vccd vccd _453_/Y sky130_fd_sc_hd__inv_2
XANTENNA__565__A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_384_ la_oen_mprj[116] vssd vssd vccd vccd _384_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[45\] _516_/Y la_buf\[45\]/TE vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[48\]_A _519_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _572_/Y la_buf\[101\]/TE vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_0_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vssd vccd vccd la_data_in_mprj[89]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[38\]_TE la_buf\[38\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] mprj_logic_high_inst/HI[364] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[39\]_A _510_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[124\]_A _392_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__385__A la_oen_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[85\] _353_/Y mprj_logic_high_inst/HI[287] vssd vssd vccd
+ vccd la_oen_core[85] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _649_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_A _383_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_505_ la_data_out_mprj[34] vssd vssd vccd vccd _505_/Y sky130_fd_sc_hd__inv_2
X_436_ mprj_adr_o_core[29] vssd vssd vccd vccd _436_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_367_ la_oen_mprj[99] vssd vssd vccd vccd _367_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _640_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _374_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _631_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[99\]_A _367_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _622_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_419_ mprj_adr_o_core[12] vssd vssd vccd vccd _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _613_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] mprj_logic_high_inst/HI[438] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[10\]_A _417_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _386_/Y mprj_logic_high_inst/HI[320] vssd vssd vccd
+ vccd la_oen_core[118] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[48\] _647_/Y mprj_logic_high_inst/HI[250] vssd vssd vccd
+ vccd la_oen_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_28_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__573__A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[105] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vssd vccd vccd la_data_in_mprj[71]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high_inst/HI[235] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_84 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[4\] _443_/Y mprj_dat_buf\[4\]/TE vssd vssd vccd vccd mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__658__A la_oen_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[109\]_TE la_buf\[109\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__393__A la_oen_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__568__A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_A _462_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[75\] _546_/Y la_buf\[75\]/TE vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high_inst/HI[258] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__478__A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] mprj_logic_high_inst/HI[394] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[14\]_A _453_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[94\]_TE la_buf\[94\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A la_oen_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _608_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_598_ la_data_out_mprj[127] vssd vssd vccd vccd _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vssd vccd vccd la_data_in_mprj[34]
+ sky130_fd_sc_hd__inv_8
XPHY_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[100\] _368_/Y mprj_logic_high_inst/HI[302] vssd vssd vccd
+ vccd la_oen_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_8_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _629_/Y mprj_logic_high_inst/HI[232] vssd vssd vccd
+ vccd la_oen_core[30] sky130_fd_sc_hd__einvp_8
X_521_ la_data_out_mprj[50] vssd vssd vccd vccd _521_/Y sky130_fd_sc_hd__inv_2
X_452_ mprj_dat_o_core[13] vssd vssd vccd vccd _452_/Y sky130_fd_sc_hd__inv_2
X_383_ la_oen_mprj[115] vssd vssd vccd vccd _383_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[1\]_A _472_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__581__A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[38\] _509_/Y la_buf\[38\]/TE vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_12_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] mprj_logic_high_inst/HI[357] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__491__A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_A _415_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[78\] _346_/Y mprj_logic_high_inst/HI[280] vssd vssd vccd
+ vccd la_oen_core[78] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[26\] _465_/Y mprj_dat_buf\[26\]/TE vssd vssd vccd vccd mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__576__A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_504_ la_data_out_mprj[33] vssd vssd vccd vccd _504_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_435_ mprj_adr_o_core[28] vssd vssd vccd vccd _435_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_366_ la_oen_mprj[98] vssd vssd vccd vccd _366_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[21\] _428_/Y mprj_adr_buf\[21\]/TE vssd vssd vccd vccd mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__486__A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__396__A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[28\]_TE la_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_418_ mprj_adr_o_core[11] vssd vssd vccd vccd _418_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_349_ la_oen_mprj[81] vssd vssd vccd vccd _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] mprj_logic_high_inst/HI[424] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[8\]_B user_to_mprj_in_gates\[8\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[20\] _491_/Y la_buf\[20\]/TE vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__einvp_8
XFILLER_3_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_87 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vssd vccd vccd la_data_in_mprj[64]
+ sky130_fd_sc_hd__inv_8
XFILLER_21_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_41 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] mprj_logic_high_inst/HI[450] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[60\] _659_/Y mprj_logic_high_inst/HI[262] vssd vssd vccd
+ vccd la_oen_core[60] sky130_fd_sc_hd__einvp_8
XFILLER_0_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__584__A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _539_/Y la_buf\[68\]/TE vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__einvp_8
XPHY_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[124\] _595_/Y la_buf\[124\]/TE vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_4_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] mprj_logic_high_inst/HI[387] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__494__A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_22_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__579__A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_597_ la_data_out_mprj[126] vssd vssd vccd vccd _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vssd vccd vccd la_data_in_mprj[27]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__489__A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__399__A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_520_ la_data_out_mprj[49] vssd vssd vccd vccd _520_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[5\] _604_/Y mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd la_oen_core[5] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[23\] _622_/Y mprj_logic_high_inst/HI[225] vssd vssd vccd
+ vccd la_oen_core[23] sky130_fd_sc_hd__einvp_8
X_451_ mprj_dat_o_core[12] vssd vssd vccd vccd _451_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_382_ la_oen_mprj[114] vssd vssd vccd vccd _382_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_649_ la_oen_mprj[50] vssd vssd vccd vccd _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_sel_buf\[2\]_A _405_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_dat_buf\[19\] _458_/Y mprj_dat_buf\[19\]/TE vssd vssd vccd vccd mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_503_ la_data_out_mprj[32] vssd vssd vccd vccd _503_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_434_ mprj_adr_o_core[27] vssd vssd vccd vccd _434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__592__A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[50\] _521_/Y la_buf\[50\]/TE vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__einvp_8
X_365_ la_oen_mprj[97] vssd vssd vccd vccd _365_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_A _442_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[14\] _421_/Y mprj_adr_buf\[14\]/TE vssd vssd vccd vccd mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[40\]_B mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vssd vccd vccd la_data_in_mprj[94]
+ sky130_fd_sc_hd__inv_8
XFILLER_3_76 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] user_to_mprj_in_gates\[1\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[92\]_A user_to_mprj_in_gates\[92\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[31\]_B mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[90\] _358_/Y mprj_logic_high_inst/HI[292] vssd vssd vccd
+ vccd la_oen_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_3_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[22\]_B mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[98\] _569_/Y la_buf\[98\]/TE vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_4_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__587__A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[89\]_B mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_417_ mprj_adr_o_core[10] vssd vssd vccd vccd _417_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_348_ la_oen_mprj[80] vssd vssd vccd vccd _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[121\]_A user_to_mprj_in_gates\[121\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[110\]_A _581_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[13\]_B mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] mprj_logic_high_inst/HI[417] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__497__A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_buffers\[112\]_A user_to_mprj_in_gates\[112\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[101\]_A _572_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[65\]_A user_to_mprj_in_gates\[65\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vssd vccd vccd la_data_in_mprj[1]
+ sky130_fd_sc_hd__inv_8
XPHY_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[103\]_A user_to_mprj_in_gates\[103\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[13\] _484_/Y la_buf\[13\]/TE vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__einvp_8
Xla_buf\[9\] _480_/Y la_buf\[9\]/TE vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_10_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[6\] _413_/Y mprj_adr_buf\[6\]/TE vssd vssd vccd vccd mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vssd vccd vccd la_data_in_mprj[57]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[96\]_A _567_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[20\]_A _491_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] mprj_logic_high_inst/HI[443] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[87\]_A _558_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[123\] _391_/Y mprj_logic_high_inst/HI[325] vssd vssd vccd
+ vccd la_oen_core[123] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[11\]_A _482_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[53\] _652_/Y mprj_logic_high_inst/HI[255] vssd vssd vccd
+ vccd la_oen_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_1_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[78\]_A _549_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[117\] _588_/Y la_buf\[117\]/TE vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[110] sky130_fd_sc_hd__inv_8
XFILLER_19_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_B mprj_logic_high_inst/HI[449] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[69\]_A _540_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[80\]_A _348_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _551_/Y la_buf\[80\]/TE vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__einvp_8
XANTENNA__595__A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_596_ la_data_out_mprj[125] vssd vssd vccd vccd _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _339_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[62\]_A _330_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[127\]_A _395_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_450_ mprj_dat_o_core[11] vssd vssd vccd vccd _450_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[16\] _615_/Y mprj_logic_high_inst/HI[218] vssd vssd vccd
+ vccd la_oen_core[16] sky130_fd_sc_hd__einvp_8
X_381_ la_oen_mprj[113] vssd vssd vccd vccd _381_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_A _652_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_A _386_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_648_ la_oen_mprj[49] vssd vssd vccd vccd _648_/Y sky130_fd_sc_hd__inv_2
X_579_ la_data_out_mprj[108] vssd vssd vccd vccd _579_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _643_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_A _377_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _634_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_A _438_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_40 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_502_ la_data_out_mprj[31] vssd vssd vccd vccd _502_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_433_ mprj_adr_o_core[26] vssd vssd vccd vccd _433_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_364_ la_oen_mprj[96] vssd vssd vccd vccd _364_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[43\] _514_/Y la_buf\[43\]/TE vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__einvp_8
XFILLER_9_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _625_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[22\]_A _429_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vssd vccd vccd la_data_in_mprj[87]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] mprj_logic_high_inst/HI[362] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _616_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_A _420_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[83\] _351_/Y mprj_logic_high_inst/HI[285] vssd vssd vccd
+ vccd la_oen_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_3_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[31\] _470_/Y mprj_dat_buf\[31\]/TE vssd vssd vccd vccd mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[59\]_TE mprj_logic_high_inst/HI[261] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_416_ mprj_adr_o_core[9] vssd vssd vccd vccd _416_/Y sky130_fd_sc_hd__inv_2
X_347_ la_oen_mprj[79] vssd vssd vccd vccd _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__598__A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_A _465_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_dat_buf\[17\]_A _456_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] mprj_logic_high_inst/HI[436] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[116\] _384_/Y mprj_logic_high_inst/HI[318] vssd vssd vccd
+ vccd la_oen_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_5_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _645_/Y mprj_logic_high_inst/HI[248] vssd vssd vccd
+ vccd la_oen_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_1_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[103] sky130_fd_sc_hd__inv_8
XFILLER_19_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[2\] _441_/Y mprj_dat_buf\[2\]/TE vssd vssd vccd vccd mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[4\]_A _475_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[73\] _544_/Y la_buf\[73\]/TE vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__einvp_8
X_595_ la_data_out_mprj[124] vssd vssd vccd vccd _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] mprj_logic_high_inst/HI[392] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_380_ la_oen_mprj[112] vssd vssd vccd vccd _380_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_647_ la_oen_mprj[48] vssd vssd vccd vccd _647_/Y sky130_fd_sc_hd__inv_2
X_578_ la_data_out_mprj[107] vssd vssd vccd vccd _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vssd vccd vccd la_data_in_mprj[32]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
.ends

