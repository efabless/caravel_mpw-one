magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1288 -1260 1385 1560
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1623348570
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 125 300 125 300 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 1788682
string GDS_START 1787762
<< end >>
