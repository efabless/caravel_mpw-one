magic
tech sky130A
magscale 1 2
timestamp 1623348513
<< locali >>
rect 185 480 192 514
rect 226 480 264 514
rect 298 480 336 514
rect 370 480 408 514
rect 442 480 480 514
rect 514 480 552 514
rect 586 480 591 514
rect 185 20 192 54
rect 226 20 264 54
rect 298 20 336 54
rect 370 20 408 54
rect 442 20 480 54
rect 514 20 552 54
rect 586 20 591 54
<< viali >>
rect 192 480 226 514
rect 264 480 298 514
rect 336 480 370 514
rect 408 480 442 514
rect 480 480 514 514
rect 552 480 586 514
rect 192 20 226 54
rect 264 20 298 54
rect 336 20 370 54
rect 408 20 442 54
rect 480 20 514 54
rect 552 20 586 54
<< obsli1 >>
rect 48 392 82 402
rect 48 320 82 358
rect 48 248 82 286
rect 48 176 82 214
rect 48 132 82 142
rect 159 98 193 436
rect 265 98 299 436
rect 371 98 405 436
rect 477 98 511 436
rect 583 98 617 436
rect 694 392 728 402
rect 694 320 728 358
rect 694 248 728 286
rect 694 176 728 214
rect 694 132 728 142
<< obsli1c >>
rect 48 358 82 392
rect 48 286 82 320
rect 48 214 82 248
rect 48 142 82 176
rect 694 358 728 392
rect 694 286 728 320
rect 694 214 728 248
rect 694 142 728 176
<< metal1 >>
rect 180 514 598 534
rect 180 480 192 514
rect 226 480 264 514
rect 298 480 336 514
rect 370 480 408 514
rect 442 480 480 514
rect 514 480 552 514
rect 586 480 598 514
rect 180 468 598 480
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 682 392 740 420
rect 682 358 694 392
rect 728 358 740 392
rect 682 320 740 358
rect 682 286 694 320
rect 728 286 740 320
rect 682 248 740 286
rect 682 214 694 248
rect 728 214 740 248
rect 682 176 740 214
rect 682 142 694 176
rect 728 142 740 176
rect 682 114 740 142
rect 180 54 598 66
rect 180 20 192 54
rect 226 20 264 54
rect 298 20 336 54
rect 370 20 408 54
rect 442 20 480 54
rect 514 20 552 54
rect 586 20 598 54
rect 180 0 598 20
<< obsm1 >>
rect 150 114 202 420
rect 256 114 308 420
rect 362 114 414 420
rect 468 114 520 420
rect 574 114 626 420
<< metal2 >>
rect 10 292 766 420
rect 10 114 766 242
<< labels >>
rlabel metal1 s 682 114 740 420 6 BULK
port 1 nsew
rlabel metal1 s 36 114 94 420 6 BULK
port 1 nsew
rlabel metal2 s 10 292 766 420 6 DRAIN
port 2 nsew
rlabel viali s 552 480 586 514 6 GATE
port 3 nsew
rlabel viali s 552 20 586 54 6 GATE
port 3 nsew
rlabel viali s 480 480 514 514 6 GATE
port 3 nsew
rlabel viali s 480 20 514 54 6 GATE
port 3 nsew
rlabel viali s 408 480 442 514 6 GATE
port 3 nsew
rlabel viali s 408 20 442 54 6 GATE
port 3 nsew
rlabel viali s 336 480 370 514 6 GATE
port 3 nsew
rlabel viali s 336 20 370 54 6 GATE
port 3 nsew
rlabel viali s 264 480 298 514 6 GATE
port 3 nsew
rlabel viali s 264 20 298 54 6 GATE
port 3 nsew
rlabel viali s 192 480 226 514 6 GATE
port 3 nsew
rlabel viali s 192 20 226 54 6 GATE
port 3 nsew
rlabel locali s 185 480 591 514 6 GATE
port 3 nsew
rlabel locali s 185 20 591 54 6 GATE
port 3 nsew
rlabel metal1 s 180 468 598 534 6 GATE
port 3 nsew
rlabel metal1 s 180 0 598 66 6 GATE
port 3 nsew
rlabel metal2 s 10 114 766 242 6 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 776 534
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9505486
string GDS_START 9494654
<< end >>
