***  
* Most models come from here:

.lib ../../../../../../../pdks/sky130A-xyce/libs.tech/xyce/sky130.lib.spice tt

.include ./sky130_fd_io__condiode.spice
.include ./sky130_fd_pr__model__parasitic__diode_ps2nw.spice 
.include ./sky130_fd_pr__model__parasitic__diode_pw2dn.spice
.include ./sky130_fd_pr__model__parasitic__diode_ps2dn.spice


*.include ./sky130_fd_pr__model__parasitic__diode_ps2nw.model.spice 
*.include ./sky130_fd_pr__model__parasitic__diode_pw2dn.model.spice
*.include ./sky130_fd_pr__model__parasitic__diode_ps2dn.model.spice


***************************************

*.include   ./sky130_ef_io__gpiov2_pad_wrapped.extracted.spice-calibre-202103-hs2ng
.include  ./sky130_ef_io__gpiov2_pad_wrapped-extracted.spice-calibre-202107-hs2ng

*** no space before the .include
*** removed subckts without any ports
*** converted calibre extracted netlist to spice with hs2ng
*** changed parasitic diodes to level=2.0
*** used sky130A-xyce PDK from MG

***************************************
Xsky130_ef_io__gpiov2_pad_wrapped 
+ VSS		; VSSD 
+ VSS		; VSSIO 
+ VSS		; VSSA 
+ VSS		; VSSIO_Q 
+ VDD3V3	; VDDIO 
+ VDD3V3	; VDDIO_Q 
+ OPEN1 	; PAD_A_ESD_1_H 
+ PAD		; PAD 
+ OPEN2		; PAD_A_ESD_0_H 
+ ZERO		; IB_MODE_SEL 
+ ONE3V3	; ENABLE_INP_H 
+ ONE3V3	; ENABLE_H 
+ VDD3V3	; VDDA 
+ ONE3V3	; ENABLE_VDDA_H 
+ VDD1V8	; VCCD 
+ ZERO		; OE_N 
+ ZERO		; VTRIP_SEL 
+ VDD1V8	; VCCHIB 
+ ZERO		; ENABLE_VSWITCH_H 
+ OUT		; OUT
+ ZERO		; HLD_OVR 
+ ONE1V8	; DM[2] 
+ ZERO		; ANALOG_SEL 
+ ONE3V3	; HLD_H_N 
+ ZERO		; ANALOG_EN 
+ ZERO		; INP_DIS 
+ ZERO		; ANALOG_POL 
+ ZERO		; DM[0] 
+ OPEN3		; PAD_A_NOESD_H 
+ ONE1V8	; DM[1] 
+ ZERO		; SLOW 
+ OPEN4		; TIE_HI_ESD 
+ IN		; IN 
+ OPEN5		; IN_H 
+ ONE1V8	; ENABLE_VDDIO 
+ OPEN6		; TIE_LO_ESD 
+ VDD3V3	; VSWITCH 
+ OPEN7		; AMUXBUS_A 
+ OPEN8		; AMUXBUS_B
+ sky130_ef_io__gpiov2_pad_wrapped


vvss		VSS		0 		dc 	0
vvdd1v8		VDD1V8		0 		pwl	0 0 3u  1.8  1m 1.8
vvdd3v3		VDD3V3		0 		pwl	0 0 2u  3.3  1m 3.3

vzero		ZERO		0		dc	0
vone1v8		ONE1V8		0		pwl	0 0 5.5u 0 5.6u 1.8  1m 1.8
vone3v3		ONE3V3		0		pwl	0 0 5.5u 0 5.6u 3.3  1m 3.3

vout		OUT		0		pwl	0 0 8u 0  8.1u 1.8 11u 1.8 11.1u 0 15u 0
rload		PAD		0		1000K


.PRINT TRAN FORMAT=RAW v(pad) v(out) i(vvdd3v3) i(vvdd1v8) v(vdd3v3) v(vdd1v8) v(ONE1V8) v(ONE3V3) i(vone1v8) i(vone3v3) i(vout) i(rload)
.TRAN 10n 15u

.END
