magic
tech sky130A
magscale 1 2
timestamp 1623348512
<< checkpaint >>
rect -1246 -1260 1888 2648
<< pwell >>
rect 15 163 627 1225
<< nmos >>
rect 171 189 201 1199
rect 257 189 293 1199
rect 349 189 385 1199
rect 441 189 471 1199
<< ndiff >>
rect 111 1187 171 1199
rect 111 1153 126 1187
rect 160 1153 171 1187
rect 111 1119 171 1153
rect 111 1085 126 1119
rect 160 1085 171 1119
rect 111 1051 171 1085
rect 111 1017 126 1051
rect 160 1017 171 1051
rect 111 983 171 1017
rect 111 949 126 983
rect 160 949 171 983
rect 111 915 171 949
rect 111 881 126 915
rect 160 881 171 915
rect 111 847 171 881
rect 111 813 126 847
rect 160 813 171 847
rect 111 779 171 813
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 1187 257 1199
rect 201 1153 212 1187
rect 246 1153 257 1187
rect 201 1119 257 1153
rect 201 1085 212 1119
rect 246 1085 257 1119
rect 201 1051 257 1085
rect 201 1017 212 1051
rect 246 1017 257 1051
rect 201 983 257 1017
rect 201 949 212 983
rect 246 949 257 983
rect 201 915 257 949
rect 201 881 212 915
rect 246 881 257 915
rect 201 847 257 881
rect 201 813 212 847
rect 246 813 257 847
rect 201 779 257 813
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 293 1187 349 1199
rect 293 1153 304 1187
rect 338 1153 349 1187
rect 293 1119 349 1153
rect 293 1085 304 1119
rect 338 1085 349 1119
rect 293 1051 349 1085
rect 293 1017 304 1051
rect 338 1017 349 1051
rect 293 983 349 1017
rect 293 949 304 983
rect 338 949 349 983
rect 293 915 349 949
rect 293 881 304 915
rect 338 881 349 915
rect 293 847 349 881
rect 293 813 304 847
rect 338 813 349 847
rect 293 779 349 813
rect 293 745 304 779
rect 338 745 349 779
rect 293 711 349 745
rect 293 677 304 711
rect 338 677 349 711
rect 293 643 349 677
rect 293 609 304 643
rect 338 609 349 643
rect 293 575 349 609
rect 293 541 304 575
rect 338 541 349 575
rect 293 507 349 541
rect 293 473 304 507
rect 338 473 349 507
rect 293 439 349 473
rect 293 405 304 439
rect 338 405 349 439
rect 293 371 349 405
rect 293 337 304 371
rect 338 337 349 371
rect 293 303 349 337
rect 293 269 304 303
rect 338 269 349 303
rect 293 235 349 269
rect 293 201 304 235
rect 338 201 349 235
rect 293 189 349 201
rect 385 1187 441 1199
rect 385 1153 396 1187
rect 430 1153 441 1187
rect 385 1119 441 1153
rect 385 1085 396 1119
rect 430 1085 441 1119
rect 385 1051 441 1085
rect 385 1017 396 1051
rect 430 1017 441 1051
rect 385 983 441 1017
rect 385 949 396 983
rect 430 949 441 983
rect 385 915 441 949
rect 385 881 396 915
rect 430 881 441 915
rect 385 847 441 881
rect 385 813 396 847
rect 430 813 441 847
rect 385 779 441 813
rect 385 745 396 779
rect 430 745 441 779
rect 385 711 441 745
rect 385 677 396 711
rect 430 677 441 711
rect 385 643 441 677
rect 385 609 396 643
rect 430 609 441 643
rect 385 575 441 609
rect 385 541 396 575
rect 430 541 441 575
rect 385 507 441 541
rect 385 473 396 507
rect 430 473 441 507
rect 385 439 441 473
rect 385 405 396 439
rect 430 405 441 439
rect 385 371 441 405
rect 385 337 396 371
rect 430 337 441 371
rect 385 303 441 337
rect 385 269 396 303
rect 430 269 441 303
rect 385 235 441 269
rect 385 201 396 235
rect 430 201 441 235
rect 385 189 441 201
rect 471 1187 531 1199
rect 471 1153 482 1187
rect 516 1153 531 1187
rect 471 1119 531 1153
rect 471 1085 482 1119
rect 516 1085 531 1119
rect 471 1051 531 1085
rect 471 1017 482 1051
rect 516 1017 531 1051
rect 471 983 531 1017
rect 471 949 482 983
rect 516 949 531 983
rect 471 915 531 949
rect 471 881 482 915
rect 516 881 531 915
rect 471 847 531 881
rect 471 813 482 847
rect 516 813 531 847
rect 471 779 531 813
rect 471 745 482 779
rect 516 745 531 779
rect 471 711 531 745
rect 471 677 482 711
rect 516 677 531 711
rect 471 643 531 677
rect 471 609 482 643
rect 516 609 531 643
rect 471 575 531 609
rect 471 541 482 575
rect 516 541 531 575
rect 471 507 531 541
rect 471 473 482 507
rect 516 473 531 507
rect 471 439 531 473
rect 471 405 482 439
rect 516 405 531 439
rect 471 371 531 405
rect 471 337 482 371
rect 516 337 531 371
rect 471 303 531 337
rect 471 269 482 303
rect 516 269 531 303
rect 471 235 531 269
rect 471 201 482 235
rect 516 201 531 235
rect 471 189 531 201
<< ndiffc >>
rect 126 1153 160 1187
rect 126 1085 160 1119
rect 126 1017 160 1051
rect 126 949 160 983
rect 126 881 160 915
rect 126 813 160 847
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 1153 246 1187
rect 212 1085 246 1119
rect 212 1017 246 1051
rect 212 949 246 983
rect 212 881 246 915
rect 212 813 246 847
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 304 1153 338 1187
rect 304 1085 338 1119
rect 304 1017 338 1051
rect 304 949 338 983
rect 304 881 338 915
rect 304 813 338 847
rect 304 745 338 779
rect 304 677 338 711
rect 304 609 338 643
rect 304 541 338 575
rect 304 473 338 507
rect 304 405 338 439
rect 304 337 338 371
rect 304 269 338 303
rect 304 201 338 235
rect 396 1153 430 1187
rect 396 1085 430 1119
rect 396 1017 430 1051
rect 396 949 430 983
rect 396 881 430 915
rect 396 813 430 847
rect 396 745 430 779
rect 396 677 430 711
rect 396 609 430 643
rect 396 541 430 575
rect 396 473 430 507
rect 396 405 430 439
rect 396 337 430 371
rect 396 269 430 303
rect 396 201 430 235
rect 482 1153 516 1187
rect 482 1085 516 1119
rect 482 1017 516 1051
rect 482 949 516 983
rect 482 881 516 915
rect 482 813 516 847
rect 482 745 516 779
rect 482 677 516 711
rect 482 609 516 643
rect 482 541 516 575
rect 482 473 516 507
rect 482 405 516 439
rect 482 337 516 371
rect 482 269 516 303
rect 482 201 516 235
<< psubdiff >>
rect 41 1187 111 1199
rect 41 1153 58 1187
rect 92 1153 111 1187
rect 41 1119 111 1153
rect 41 1085 58 1119
rect 92 1085 111 1119
rect 41 1051 111 1085
rect 41 1017 58 1051
rect 92 1017 111 1051
rect 41 983 111 1017
rect 41 949 58 983
rect 92 949 111 983
rect 41 915 111 949
rect 41 881 58 915
rect 92 881 111 915
rect 41 847 111 881
rect 41 813 58 847
rect 92 813 111 847
rect 41 779 111 813
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 531 1187 601 1199
rect 531 1153 550 1187
rect 584 1153 601 1187
rect 531 1119 601 1153
rect 531 1085 550 1119
rect 584 1085 601 1119
rect 531 1051 601 1085
rect 531 1017 550 1051
rect 584 1017 601 1051
rect 531 983 601 1017
rect 531 949 550 983
rect 584 949 601 983
rect 531 915 601 949
rect 531 881 550 915
rect 584 881 601 915
rect 531 847 601 881
rect 531 813 550 847
rect 584 813 601 847
rect 531 779 601 813
rect 531 745 550 779
rect 584 745 601 779
rect 531 711 601 745
rect 531 677 550 711
rect 584 677 601 711
rect 531 643 601 677
rect 531 609 550 643
rect 584 609 601 643
rect 531 575 601 609
rect 531 541 550 575
rect 584 541 601 575
rect 531 507 601 541
rect 531 473 550 507
rect 584 473 601 507
rect 531 439 601 473
rect 531 405 550 439
rect 584 405 601 439
rect 531 371 601 405
rect 531 337 550 371
rect 584 337 601 371
rect 531 303 601 337
rect 531 269 550 303
rect 584 269 601 303
rect 531 235 601 269
rect 531 201 550 235
rect 584 201 601 235
rect 531 189 601 201
<< psubdiffcont >>
rect 58 1153 92 1187
rect 58 1085 92 1119
rect 58 1017 92 1051
rect 58 949 92 983
rect 58 881 92 915
rect 58 813 92 847
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 550 1153 584 1187
rect 550 1085 584 1119
rect 550 1017 584 1051
rect 550 949 584 983
rect 550 881 584 915
rect 550 813 584 847
rect 550 745 584 779
rect 550 677 584 711
rect 550 609 584 643
rect 550 541 584 575
rect 550 473 584 507
rect 550 405 584 439
rect 550 337 584 371
rect 550 269 584 303
rect 550 201 584 235
<< poly >>
rect 243 1367 399 1388
rect 243 1333 264 1367
rect 298 1333 344 1367
rect 378 1333 399 1367
rect 243 1299 399 1333
rect 120 1275 201 1291
rect 120 1241 136 1275
rect 170 1241 201 1275
rect 243 1265 264 1299
rect 298 1265 344 1299
rect 378 1265 399 1299
rect 243 1249 399 1265
rect 441 1275 522 1291
rect 120 1225 201 1241
rect 171 1199 201 1225
rect 257 1199 293 1249
rect 349 1199 385 1249
rect 441 1241 472 1275
rect 506 1241 522 1275
rect 441 1225 522 1241
rect 441 1199 471 1225
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 293 189
rect 349 139 385 189
rect 441 163 471 189
rect 441 147 522 163
rect 120 97 201 113
rect 243 123 399 139
rect 243 89 264 123
rect 298 89 344 123
rect 378 89 399 123
rect 441 113 472 147
rect 506 113 522 147
rect 441 97 522 113
rect 243 55 399 89
rect 243 21 264 55
rect 298 21 344 55
rect 378 21 399 55
rect 243 0 399 21
<< polycont >>
rect 264 1333 298 1367
rect 344 1333 378 1367
rect 136 1241 170 1275
rect 264 1265 298 1299
rect 344 1265 378 1299
rect 472 1241 506 1275
rect 136 113 170 147
rect 264 89 298 123
rect 344 89 378 123
rect 472 113 506 147
rect 264 21 298 55
rect 344 21 378 55
<< locali >>
rect 248 1369 394 1388
rect 248 1335 262 1369
rect 296 1367 346 1369
rect 248 1333 264 1335
rect 298 1333 344 1367
rect 380 1335 394 1369
rect 378 1333 394 1335
rect 248 1299 394 1333
rect 248 1297 264 1299
rect 120 1275 186 1291
rect 120 1241 136 1275
rect 170 1241 186 1275
rect 248 1263 262 1297
rect 298 1265 344 1299
rect 378 1297 394 1299
rect 296 1263 346 1265
rect 380 1263 394 1297
rect 248 1249 394 1263
rect 456 1275 522 1291
rect 120 1225 186 1241
rect 456 1241 472 1275
rect 506 1241 522 1275
rect 456 1225 522 1241
rect 120 1203 160 1225
rect 482 1203 522 1225
rect 41 1187 160 1203
rect 41 1153 58 1187
rect 92 1179 126 1187
rect 94 1153 126 1179
rect 41 1145 60 1153
rect 94 1145 160 1153
rect 41 1119 160 1145
rect 41 1085 58 1119
rect 92 1107 126 1119
rect 94 1085 126 1107
rect 41 1073 60 1085
rect 94 1073 160 1085
rect 41 1051 160 1073
rect 41 1017 58 1051
rect 92 1035 126 1051
rect 94 1017 126 1035
rect 41 1001 60 1017
rect 94 1001 160 1017
rect 41 983 160 1001
rect 41 949 58 983
rect 92 963 126 983
rect 94 949 126 963
rect 41 929 60 949
rect 94 929 160 949
rect 41 915 160 929
rect 41 881 58 915
rect 92 891 126 915
rect 94 881 126 891
rect 41 857 60 881
rect 94 857 160 881
rect 41 847 160 857
rect 41 813 58 847
rect 92 819 126 847
rect 94 813 126 819
rect 41 785 60 813
rect 94 785 160 813
rect 41 779 160 785
rect 41 745 58 779
rect 92 747 126 779
rect 94 745 126 747
rect 41 713 60 745
rect 94 713 160 745
rect 41 711 160 713
rect 41 677 58 711
rect 92 677 126 711
rect 41 675 160 677
rect 41 643 60 675
rect 94 643 160 675
rect 41 609 58 643
rect 94 641 126 643
rect 92 609 126 641
rect 41 603 160 609
rect 41 575 60 603
rect 94 575 160 603
rect 41 541 58 575
rect 94 569 126 575
rect 92 541 126 569
rect 41 531 160 541
rect 41 507 60 531
rect 94 507 160 531
rect 41 473 58 507
rect 94 497 126 507
rect 92 473 126 497
rect 41 459 160 473
rect 41 439 60 459
rect 94 439 160 459
rect 41 405 58 439
rect 94 425 126 439
rect 92 405 126 425
rect 41 387 160 405
rect 41 371 60 387
rect 94 371 160 387
rect 41 337 58 371
rect 94 353 126 371
rect 92 337 126 353
rect 41 315 160 337
rect 41 303 60 315
rect 94 303 160 315
rect 41 269 58 303
rect 94 281 126 303
rect 92 269 126 281
rect 41 243 160 269
rect 41 235 60 243
rect 94 235 160 243
rect 41 201 58 235
rect 94 209 126 235
rect 92 201 126 209
rect 41 185 160 201
rect 212 1187 246 1203
rect 212 1119 246 1145
rect 212 1051 246 1073
rect 212 983 246 1001
rect 212 915 246 929
rect 212 847 246 857
rect 212 779 246 785
rect 212 711 246 713
rect 212 675 246 677
rect 212 603 246 609
rect 212 531 246 541
rect 212 459 246 473
rect 212 387 246 405
rect 212 315 246 337
rect 212 243 246 269
rect 212 185 246 201
rect 304 1187 338 1203
rect 304 1119 338 1145
rect 304 1051 338 1073
rect 304 983 338 1001
rect 304 915 338 929
rect 304 847 338 857
rect 304 779 338 785
rect 304 711 338 713
rect 304 675 338 677
rect 304 603 338 609
rect 304 531 338 541
rect 304 459 338 473
rect 304 387 338 405
rect 304 315 338 337
rect 304 243 338 269
rect 304 185 338 201
rect 396 1187 430 1203
rect 396 1119 430 1145
rect 396 1051 430 1073
rect 396 983 430 1001
rect 396 915 430 929
rect 396 847 430 857
rect 396 779 430 785
rect 396 711 430 713
rect 396 675 430 677
rect 396 603 430 609
rect 396 531 430 541
rect 396 459 430 473
rect 396 387 430 405
rect 396 315 430 337
rect 396 243 430 269
rect 396 185 430 201
rect 482 1187 601 1203
rect 516 1179 550 1187
rect 516 1153 548 1179
rect 584 1153 601 1187
rect 482 1145 548 1153
rect 582 1145 601 1153
rect 482 1119 601 1145
rect 516 1107 550 1119
rect 516 1085 548 1107
rect 584 1085 601 1119
rect 482 1073 548 1085
rect 582 1073 601 1085
rect 482 1051 601 1073
rect 516 1035 550 1051
rect 516 1017 548 1035
rect 584 1017 601 1051
rect 482 1001 548 1017
rect 582 1001 601 1017
rect 482 983 601 1001
rect 516 963 550 983
rect 516 949 548 963
rect 584 949 601 983
rect 482 929 548 949
rect 582 929 601 949
rect 482 915 601 929
rect 516 891 550 915
rect 516 881 548 891
rect 584 881 601 915
rect 482 857 548 881
rect 582 857 601 881
rect 482 847 601 857
rect 516 819 550 847
rect 516 813 548 819
rect 584 813 601 847
rect 482 785 548 813
rect 582 785 601 813
rect 482 779 601 785
rect 516 747 550 779
rect 516 745 548 747
rect 584 745 601 779
rect 482 713 548 745
rect 582 713 601 745
rect 482 711 601 713
rect 516 677 550 711
rect 584 677 601 711
rect 482 675 601 677
rect 482 643 548 675
rect 582 643 601 675
rect 516 641 548 643
rect 516 609 550 641
rect 584 609 601 643
rect 482 603 601 609
rect 482 575 548 603
rect 582 575 601 603
rect 516 569 548 575
rect 516 541 550 569
rect 584 541 601 575
rect 482 531 601 541
rect 482 507 548 531
rect 582 507 601 531
rect 516 497 548 507
rect 516 473 550 497
rect 584 473 601 507
rect 482 459 601 473
rect 482 439 548 459
rect 582 439 601 459
rect 516 425 548 439
rect 516 405 550 425
rect 584 405 601 439
rect 482 387 601 405
rect 482 371 548 387
rect 582 371 601 387
rect 516 353 548 371
rect 516 337 550 353
rect 584 337 601 371
rect 482 315 601 337
rect 482 303 548 315
rect 582 303 601 315
rect 516 281 548 303
rect 516 269 550 281
rect 584 269 601 303
rect 482 243 601 269
rect 482 235 548 243
rect 582 235 601 243
rect 516 209 548 235
rect 516 201 550 209
rect 584 201 601 235
rect 482 185 601 201
rect 120 163 160 185
rect 482 163 522 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 456 147 522 163
rect 120 97 186 113
rect 248 125 394 139
rect 248 91 262 125
rect 296 123 346 125
rect 248 89 264 91
rect 298 89 344 123
rect 380 91 394 125
rect 456 113 472 147
rect 506 113 522 147
rect 456 97 522 113
rect 378 89 394 91
rect 248 55 394 89
rect 248 53 264 55
rect 248 19 262 53
rect 298 21 344 55
rect 378 53 394 55
rect 296 19 346 21
rect 380 19 394 53
rect 248 0 394 19
<< viali >>
rect 262 1367 296 1369
rect 346 1367 380 1369
rect 262 1335 264 1367
rect 264 1335 296 1367
rect 346 1335 378 1367
rect 378 1335 380 1367
rect 262 1265 264 1297
rect 264 1265 296 1297
rect 346 1265 378 1297
rect 378 1265 380 1297
rect 262 1263 296 1265
rect 346 1263 380 1265
rect 60 1153 92 1179
rect 92 1153 94 1179
rect 60 1145 94 1153
rect 60 1085 92 1107
rect 92 1085 94 1107
rect 60 1073 94 1085
rect 60 1017 92 1035
rect 92 1017 94 1035
rect 60 1001 94 1017
rect 60 949 92 963
rect 92 949 94 963
rect 60 929 94 949
rect 60 881 92 891
rect 92 881 94 891
rect 60 857 94 881
rect 60 813 92 819
rect 92 813 94 819
rect 60 785 94 813
rect 60 745 92 747
rect 92 745 94 747
rect 60 713 94 745
rect 60 643 94 675
rect 60 641 92 643
rect 92 641 94 643
rect 60 575 94 603
rect 60 569 92 575
rect 92 569 94 575
rect 60 507 94 531
rect 60 497 92 507
rect 92 497 94 507
rect 60 439 94 459
rect 60 425 92 439
rect 92 425 94 439
rect 60 371 94 387
rect 60 353 92 371
rect 92 353 94 371
rect 60 303 94 315
rect 60 281 92 303
rect 92 281 94 303
rect 60 235 94 243
rect 60 209 92 235
rect 92 209 94 235
rect 212 1153 246 1179
rect 212 1145 246 1153
rect 212 1085 246 1107
rect 212 1073 246 1085
rect 212 1017 246 1035
rect 212 1001 246 1017
rect 212 949 246 963
rect 212 929 246 949
rect 212 881 246 891
rect 212 857 246 881
rect 212 813 246 819
rect 212 785 246 813
rect 212 745 246 747
rect 212 713 246 745
rect 212 643 246 675
rect 212 641 246 643
rect 212 575 246 603
rect 212 569 246 575
rect 212 507 246 531
rect 212 497 246 507
rect 212 439 246 459
rect 212 425 246 439
rect 212 371 246 387
rect 212 353 246 371
rect 212 303 246 315
rect 212 281 246 303
rect 212 235 246 243
rect 212 209 246 235
rect 304 1153 338 1179
rect 304 1145 338 1153
rect 304 1085 338 1107
rect 304 1073 338 1085
rect 304 1017 338 1035
rect 304 1001 338 1017
rect 304 949 338 963
rect 304 929 338 949
rect 304 881 338 891
rect 304 857 338 881
rect 304 813 338 819
rect 304 785 338 813
rect 304 745 338 747
rect 304 713 338 745
rect 304 643 338 675
rect 304 641 338 643
rect 304 575 338 603
rect 304 569 338 575
rect 304 507 338 531
rect 304 497 338 507
rect 304 439 338 459
rect 304 425 338 439
rect 304 371 338 387
rect 304 353 338 371
rect 304 303 338 315
rect 304 281 338 303
rect 304 235 338 243
rect 304 209 338 235
rect 396 1153 430 1179
rect 396 1145 430 1153
rect 396 1085 430 1107
rect 396 1073 430 1085
rect 396 1017 430 1035
rect 396 1001 430 1017
rect 396 949 430 963
rect 396 929 430 949
rect 396 881 430 891
rect 396 857 430 881
rect 396 813 430 819
rect 396 785 430 813
rect 396 745 430 747
rect 396 713 430 745
rect 396 643 430 675
rect 396 641 430 643
rect 396 575 430 603
rect 396 569 430 575
rect 396 507 430 531
rect 396 497 430 507
rect 396 439 430 459
rect 396 425 430 439
rect 396 371 430 387
rect 396 353 430 371
rect 396 303 430 315
rect 396 281 430 303
rect 396 235 430 243
rect 396 209 430 235
rect 548 1153 550 1179
rect 550 1153 582 1179
rect 548 1145 582 1153
rect 548 1085 550 1107
rect 550 1085 582 1107
rect 548 1073 582 1085
rect 548 1017 550 1035
rect 550 1017 582 1035
rect 548 1001 582 1017
rect 548 949 550 963
rect 550 949 582 963
rect 548 929 582 949
rect 548 881 550 891
rect 550 881 582 891
rect 548 857 582 881
rect 548 813 550 819
rect 550 813 582 819
rect 548 785 582 813
rect 548 745 550 747
rect 550 745 582 747
rect 548 713 582 745
rect 548 643 582 675
rect 548 641 550 643
rect 550 641 582 643
rect 548 575 582 603
rect 548 569 550 575
rect 550 569 582 575
rect 548 507 582 531
rect 548 497 550 507
rect 550 497 582 507
rect 548 439 582 459
rect 548 425 550 439
rect 550 425 582 439
rect 548 371 582 387
rect 548 353 550 371
rect 550 353 582 371
rect 548 303 582 315
rect 548 281 550 303
rect 550 281 582 303
rect 548 235 582 243
rect 548 209 550 235
rect 550 209 582 235
rect 262 123 296 125
rect 346 123 380 125
rect 262 91 264 123
rect 264 91 296 123
rect 346 91 378 123
rect 378 91 380 123
rect 262 21 264 53
rect 264 21 296 53
rect 346 21 378 53
rect 378 21 380 53
rect 262 19 296 21
rect 346 19 380 21
<< metal1 >>
rect 250 1369 392 1388
rect 250 1335 262 1369
rect 296 1335 346 1369
rect 380 1335 392 1369
rect 250 1297 392 1335
rect 250 1263 262 1297
rect 296 1263 346 1297
rect 380 1263 392 1297
rect 250 1251 392 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 203 1179 255 1191
rect 203 1145 212 1179
rect 246 1145 255 1179
rect 203 1107 255 1145
rect 203 1073 212 1107
rect 246 1073 255 1107
rect 203 1035 255 1073
rect 203 1001 212 1035
rect 246 1001 255 1035
rect 203 963 255 1001
rect 203 929 212 963
rect 246 929 255 963
rect 203 891 255 929
rect 203 857 212 891
rect 246 857 255 891
rect 203 819 255 857
rect 203 785 212 819
rect 246 785 255 819
rect 203 747 255 785
rect 203 713 212 747
rect 246 713 255 747
rect 203 675 255 713
rect 203 641 212 675
rect 246 641 255 675
rect 203 639 255 641
rect 203 575 212 587
rect 246 575 255 587
rect 203 511 212 523
rect 246 511 255 523
rect 203 447 212 459
rect 246 447 255 459
rect 203 387 255 395
rect 203 383 212 387
rect 246 383 255 387
rect 203 319 255 331
rect 203 255 255 267
rect 203 197 255 203
rect 295 1185 347 1191
rect 295 1121 347 1133
rect 295 1057 347 1069
rect 295 1001 304 1005
rect 338 1001 347 1005
rect 295 993 347 1001
rect 295 929 304 941
rect 338 929 347 941
rect 295 865 304 877
rect 338 865 347 877
rect 295 801 304 813
rect 338 801 347 813
rect 295 747 347 749
rect 295 713 304 747
rect 338 713 347 747
rect 295 675 347 713
rect 295 641 304 675
rect 338 641 347 675
rect 295 603 347 641
rect 295 569 304 603
rect 338 569 347 603
rect 295 531 347 569
rect 295 497 304 531
rect 338 497 347 531
rect 295 459 347 497
rect 295 425 304 459
rect 338 425 347 459
rect 295 387 347 425
rect 295 353 304 387
rect 338 353 347 387
rect 295 315 347 353
rect 295 281 304 315
rect 338 281 347 315
rect 295 243 347 281
rect 295 209 304 243
rect 338 209 347 243
rect 295 197 347 209
rect 387 1179 439 1191
rect 387 1145 396 1179
rect 430 1145 439 1179
rect 387 1107 439 1145
rect 387 1073 396 1107
rect 430 1073 439 1107
rect 387 1035 439 1073
rect 387 1001 396 1035
rect 430 1001 439 1035
rect 387 963 439 1001
rect 387 929 396 963
rect 430 929 439 963
rect 387 891 439 929
rect 387 857 396 891
rect 430 857 439 891
rect 387 819 439 857
rect 387 785 396 819
rect 430 785 439 819
rect 387 747 439 785
rect 387 713 396 747
rect 430 713 439 747
rect 387 675 439 713
rect 387 641 396 675
rect 430 641 439 675
rect 387 639 439 641
rect 387 575 396 587
rect 430 575 439 587
rect 387 511 396 523
rect 430 511 439 523
rect 387 447 396 459
rect 430 447 439 459
rect 387 387 439 395
rect 387 383 396 387
rect 430 383 439 387
rect 387 319 439 331
rect 387 255 439 267
rect 387 197 439 203
rect 542 1179 601 1191
rect 542 1145 548 1179
rect 582 1145 601 1179
rect 542 1107 601 1145
rect 542 1073 548 1107
rect 582 1073 601 1107
rect 542 1035 601 1073
rect 542 1001 548 1035
rect 582 1001 601 1035
rect 542 963 601 1001
rect 542 929 548 963
rect 582 929 601 963
rect 542 891 601 929
rect 542 857 548 891
rect 582 857 601 891
rect 542 819 601 857
rect 542 785 548 819
rect 582 785 601 819
rect 542 747 601 785
rect 542 713 548 747
rect 582 713 601 747
rect 542 675 601 713
rect 542 641 548 675
rect 582 641 601 675
rect 542 603 601 641
rect 542 569 548 603
rect 582 569 601 603
rect 542 531 601 569
rect 542 497 548 531
rect 582 497 601 531
rect 542 459 601 497
rect 542 425 548 459
rect 582 425 601 459
rect 542 387 601 425
rect 542 353 548 387
rect 582 353 601 387
rect 542 315 601 353
rect 542 281 548 315
rect 582 281 601 315
rect 542 243 601 281
rect 542 209 548 243
rect 582 209 601 243
rect 542 197 601 209
rect 250 125 392 137
rect 250 91 262 125
rect 296 91 346 125
rect 380 91 392 125
rect 250 53 392 91
rect 250 19 262 53
rect 296 19 346 53
rect 380 19 392 53
rect 250 0 392 19
<< via1 >>
rect 203 603 255 639
rect 203 587 212 603
rect 212 587 246 603
rect 246 587 255 603
rect 203 569 212 575
rect 212 569 246 575
rect 246 569 255 575
rect 203 531 255 569
rect 203 523 212 531
rect 212 523 246 531
rect 246 523 255 531
rect 203 497 212 511
rect 212 497 246 511
rect 246 497 255 511
rect 203 459 255 497
rect 203 425 212 447
rect 212 425 246 447
rect 246 425 255 447
rect 203 395 255 425
rect 203 353 212 383
rect 212 353 246 383
rect 246 353 255 383
rect 203 331 255 353
rect 203 315 255 319
rect 203 281 212 315
rect 212 281 246 315
rect 246 281 255 315
rect 203 267 255 281
rect 203 243 255 255
rect 203 209 212 243
rect 212 209 246 243
rect 246 209 255 243
rect 203 203 255 209
rect 295 1179 347 1185
rect 295 1145 304 1179
rect 304 1145 338 1179
rect 338 1145 347 1179
rect 295 1133 347 1145
rect 295 1107 347 1121
rect 295 1073 304 1107
rect 304 1073 338 1107
rect 338 1073 347 1107
rect 295 1069 347 1073
rect 295 1035 347 1057
rect 295 1005 304 1035
rect 304 1005 338 1035
rect 338 1005 347 1035
rect 295 963 347 993
rect 295 941 304 963
rect 304 941 338 963
rect 338 941 347 963
rect 295 891 347 929
rect 295 877 304 891
rect 304 877 338 891
rect 338 877 347 891
rect 295 857 304 865
rect 304 857 338 865
rect 338 857 347 865
rect 295 819 347 857
rect 295 813 304 819
rect 304 813 338 819
rect 338 813 347 819
rect 295 785 304 801
rect 304 785 338 801
rect 338 785 347 801
rect 295 749 347 785
rect 387 603 439 639
rect 387 587 396 603
rect 396 587 430 603
rect 430 587 439 603
rect 387 569 396 575
rect 396 569 430 575
rect 430 569 439 575
rect 387 531 439 569
rect 387 523 396 531
rect 396 523 430 531
rect 430 523 439 531
rect 387 497 396 511
rect 396 497 430 511
rect 430 497 439 511
rect 387 459 439 497
rect 387 425 396 447
rect 396 425 430 447
rect 430 425 439 447
rect 387 395 439 425
rect 387 353 396 383
rect 396 353 430 383
rect 430 353 439 383
rect 387 331 439 353
rect 387 315 439 319
rect 387 281 396 315
rect 396 281 430 315
rect 430 281 439 315
rect 387 267 439 281
rect 387 243 439 255
rect 387 209 396 243
rect 396 209 430 243
rect 430 209 439 243
rect 387 203 439 209
<< metal2 >>
rect 14 1185 628 1191
rect 14 1133 295 1185
rect 347 1133 628 1185
rect 14 1121 628 1133
rect 14 1069 295 1121
rect 347 1069 628 1121
rect 14 1057 628 1069
rect 14 1005 295 1057
rect 347 1005 628 1057
rect 14 993 628 1005
rect 14 941 295 993
rect 347 941 628 993
rect 14 929 628 941
rect 14 877 295 929
rect 347 877 628 929
rect 14 865 628 877
rect 14 813 295 865
rect 347 813 628 865
rect 14 801 628 813
rect 14 749 295 801
rect 347 749 628 801
rect 14 719 628 749
rect 14 639 628 669
rect 14 587 203 639
rect 255 587 387 639
rect 439 587 628 639
rect 14 575 628 587
rect 14 523 203 575
rect 255 523 387 575
rect 439 523 628 575
rect 14 511 628 523
rect 14 459 203 511
rect 255 459 387 511
rect 439 459 628 511
rect 14 447 628 459
rect 14 395 203 447
rect 255 395 387 447
rect 439 395 628 447
rect 14 383 628 395
rect 14 331 203 383
rect 255 331 387 383
rect 439 331 628 383
rect 14 319 628 331
rect 14 267 203 319
rect 255 267 387 319
rect 439 267 628 319
rect 14 255 628 267
rect 14 203 203 255
rect 255 203 387 255
rect 439 203 628 255
rect 14 197 628 203
<< labels >>
flabel comment s 183 749 183 749 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 453 744 453 744 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 1288 386 1339 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 255 44 386 95 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 542 683 601 713 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal2 s 14 384 35 512 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 908 35 1036 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5604528
string GDS_START 5584496
<< end >>
