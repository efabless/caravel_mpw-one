magic
tech sky130A
magscale 1 2
timestamp 1624978002
<< metal3 >>
rect 72974 992991 73774 993231
rect 72972 992989 73776 992991
rect 72972 992669 72974 992989
rect 73774 992669 73776 992989
rect 72972 992667 73776 992669
rect 72974 959024 73774 992667
rect 74374 992331 75174 993231
rect 74372 992329 75176 992331
rect 74372 992009 74374 992329
rect 75174 992009 75176 992329
rect 74372 992007 75176 992009
rect 72974 958573 72991 959024
rect 73764 958573 73774 959024
rect 72974 958558 73774 958573
rect 74374 959030 75174 992007
rect 75774 991671 76574 993231
rect 75772 991669 76576 991671
rect 75772 991349 75774 991669
rect 76574 991349 76576 991669
rect 75772 991347 76576 991349
rect 74374 958579 74394 959030
rect 75167 958579 75174 959030
rect 74374 958558 75174 958579
rect 75774 959026 76574 991347
rect 77174 991011 77974 993231
rect 124574 992991 125374 993231
rect 124572 992989 125376 992991
rect 124572 992669 124574 992989
rect 125374 992669 125376 992989
rect 124572 992667 125376 992669
rect 77172 991009 77976 991011
rect 77172 990689 77174 991009
rect 77974 990689 77976 991009
rect 77172 990687 77976 990689
rect 75774 958575 75792 959026
rect 76565 958575 76574 959026
rect 75774 958558 76574 958575
rect 77174 958558 77974 990687
rect 124574 959028 125374 992667
rect 125974 992331 126774 993231
rect 125972 992329 126776 992331
rect 125972 992009 125974 992329
rect 126774 992009 126776 992329
rect 125972 992007 126776 992009
rect 124574 958529 124589 959028
rect 125363 958529 125374 959028
rect 124574 958518 125374 958529
rect 125974 959031 126774 992007
rect 127374 991671 128174 993231
rect 127372 991669 128176 991671
rect 127372 991349 127374 991669
rect 128174 991349 128176 991669
rect 127372 991347 128176 991349
rect 125974 958532 125991 959031
rect 126765 958532 126774 959031
rect 125974 958518 126774 958532
rect 127374 959028 128174 991347
rect 128774 991011 129574 993231
rect 176174 992991 176974 993231
rect 176172 992989 176976 992991
rect 176172 992669 176174 992989
rect 176974 992669 176976 992989
rect 176172 992667 176976 992669
rect 128772 991009 129576 991011
rect 128772 990689 128774 991009
rect 129574 990689 129576 991009
rect 128772 990687 129576 990689
rect 127374 958529 127385 959028
rect 128159 958529 128174 959028
rect 127374 958518 128174 958529
rect 128774 959032 129574 990687
rect 128774 958533 128784 959032
rect 129558 958533 129574 959032
rect 176174 959022 176974 992667
rect 177574 992331 178374 993231
rect 177572 992329 178376 992331
rect 177572 992009 177574 992329
rect 178374 992009 178376 992329
rect 177572 992007 178376 992009
rect 176174 958556 176183 959022
rect 176965 958556 176974 959022
rect 176174 958544 176974 958556
rect 177574 959020 178374 992007
rect 178974 991671 179774 993231
rect 178972 991669 179776 991671
rect 178972 991349 178974 991669
rect 179774 991349 179776 991669
rect 178972 991347 179776 991349
rect 177574 958554 177584 959020
rect 178366 958554 178374 959020
rect 177574 958544 178374 958554
rect 178974 959017 179774 991347
rect 180374 991011 181174 993231
rect 227774 992991 228574 993231
rect 227772 992989 228576 992991
rect 227772 992669 227774 992989
rect 228574 992669 228576 992989
rect 227772 992667 228576 992669
rect 180372 991009 181176 991011
rect 180372 990689 180374 991009
rect 181174 990689 181176 991009
rect 180372 990687 181176 990689
rect 178974 958551 178983 959017
rect 179765 958551 179774 959017
rect 178974 958544 179774 958551
rect 180374 959021 181174 990687
rect 180374 958555 180385 959021
rect 181167 958555 181174 959021
rect 180374 958544 181174 958555
rect 227774 958978 228574 992667
rect 229174 992331 229974 993231
rect 229172 992329 229976 992331
rect 229172 992009 229174 992329
rect 229974 992009 229976 992329
rect 229172 992007 229976 992009
rect 227774 958561 227789 958978
rect 228562 958561 228574 958978
rect 227774 958545 228574 958561
rect 229174 958974 229974 992007
rect 230574 991671 231374 993231
rect 230572 991669 231376 991671
rect 230572 991349 230574 991669
rect 231374 991349 231376 991669
rect 230572 991347 231376 991349
rect 229174 958557 229185 958974
rect 229958 958557 229974 958974
rect 229174 958545 229974 958557
rect 230574 958977 231374 991347
rect 231974 991011 232774 993231
rect 279374 992991 280174 993231
rect 279372 992989 280176 992991
rect 279372 992669 279374 992989
rect 280174 992669 280176 992989
rect 279372 992667 280176 992669
rect 231972 991009 232776 991011
rect 231972 990689 231974 991009
rect 232774 990689 232776 991009
rect 231972 990687 232776 990689
rect 230574 958560 230588 958977
rect 231361 958560 231374 958977
rect 230574 958545 231374 958560
rect 231974 958976 232774 990687
rect 231974 958559 231989 958976
rect 232762 958559 232774 958976
rect 231974 958545 232774 958559
rect 279374 958993 280174 992667
rect 280774 992331 281574 993231
rect 280772 992329 281576 992331
rect 280772 992009 280774 992329
rect 281574 992009 281576 992329
rect 280772 992007 281576 992009
rect 128774 958518 129574 958533
rect 279374 958539 279382 958993
rect 280164 958539 280174 958993
rect 279374 958529 280174 958539
rect 280774 958993 281574 992007
rect 282174 991671 282974 993231
rect 282172 991669 282976 991671
rect 282172 991349 282174 991669
rect 282974 991349 282976 991669
rect 282172 991347 282976 991349
rect 280774 958539 280782 958993
rect 281564 958539 281574 958993
rect 280774 958529 281574 958539
rect 282174 958995 282974 991347
rect 283574 991011 284374 993231
rect 330974 992991 331774 993231
rect 330972 992989 331776 992991
rect 330972 992669 330974 992989
rect 331774 992669 331776 992989
rect 330972 992667 331776 992669
rect 283572 991009 284376 991011
rect 283572 990689 283574 991009
rect 284374 990689 284376 991009
rect 283572 990687 284376 990689
rect 282174 958541 282187 958995
rect 282969 958541 282974 958995
rect 282174 958529 282974 958541
rect 283574 958994 284374 990687
rect 283574 958540 283583 958994
rect 284365 958540 284374 958994
rect 283574 958529 284374 958540
rect 330974 959011 331774 992667
rect 332374 992331 333174 993231
rect 332372 992329 333176 992331
rect 332372 992009 332374 992329
rect 333174 992009 333176 992329
rect 332372 992007 333176 992009
rect 330974 958495 330988 959011
rect 331755 958495 331774 959011
rect 330974 958479 331774 958495
rect 332374 959014 333174 992007
rect 333774 991671 334574 993231
rect 333772 991669 334576 991671
rect 333772 991349 333774 991669
rect 334574 991349 334576 991669
rect 333772 991347 334576 991349
rect 332374 958498 332390 959014
rect 333157 958498 333174 959014
rect 332374 958479 333174 958498
rect 333774 959008 334574 991347
rect 335174 991011 335974 993231
rect 396974 992991 397774 993231
rect 396972 992989 397776 992991
rect 396972 992669 396974 992989
rect 397774 992669 397776 992989
rect 396972 992667 397776 992669
rect 335172 991009 335976 991011
rect 335172 990689 335174 991009
rect 335974 990689 335976 991009
rect 335172 990687 335976 990689
rect 333774 958492 333791 959008
rect 334558 958492 334574 959008
rect 333774 958479 334574 958492
rect 335174 959012 335974 990687
rect 335174 958496 335195 959012
rect 335962 958496 335974 959012
rect 396974 958982 397774 992667
rect 398374 992331 399174 993231
rect 398372 992329 399176 992331
rect 398372 992009 398374 992329
rect 399174 992009 399176 992329
rect 398372 992007 399176 992009
rect 396974 958530 396986 958982
rect 397765 958530 397774 958982
rect 396974 958517 397774 958530
rect 398374 958980 399174 992007
rect 399774 991671 400574 993231
rect 399772 991669 400576 991671
rect 399772 991349 399774 991669
rect 400574 991349 400576 991669
rect 399772 991347 400576 991349
rect 398374 958528 398383 958980
rect 399162 958528 399174 958980
rect 398374 958517 399174 958528
rect 399774 958980 400574 991347
rect 401174 991011 401974 993231
rect 474174 992991 474974 993231
rect 474172 992989 474976 992991
rect 474172 992669 474174 992989
rect 474974 992669 474976 992989
rect 474172 992667 474976 992669
rect 401172 991009 401976 991011
rect 401172 990689 401174 991009
rect 401974 990689 401976 991009
rect 401172 990687 401976 990689
rect 399774 958528 399783 958980
rect 400562 958528 400574 958980
rect 399774 958517 400574 958528
rect 401174 958982 401974 990687
rect 401174 958530 401186 958982
rect 401965 958530 401974 958982
rect 401174 958517 401974 958530
rect 474174 958993 474974 992667
rect 475574 992331 476374 993231
rect 475572 992329 476376 992331
rect 475572 992009 475574 992329
rect 476374 992009 476376 992329
rect 475572 992007 476376 992009
rect 474174 958538 474185 958993
rect 474965 958538 474974 958993
rect 474174 958529 474974 958538
rect 475574 958992 476374 992007
rect 476974 991671 477774 993231
rect 476972 991669 477776 991671
rect 476972 991349 476974 991669
rect 477774 991349 477776 991669
rect 476972 991347 477776 991349
rect 475574 958537 475583 958992
rect 476363 958537 476374 958992
rect 475574 958529 476374 958537
rect 476974 958995 477774 991347
rect 478374 991011 479174 993231
rect 525374 992991 526174 993231
rect 525372 992989 526176 992991
rect 525372 992669 525374 992989
rect 526174 992669 526176 992989
rect 525372 992667 526176 992669
rect 478372 991009 479176 991011
rect 478372 990689 478374 991009
rect 479174 990689 479176 991009
rect 478372 990687 479176 990689
rect 476974 958540 476985 958995
rect 477765 958540 477774 958995
rect 476974 958529 477774 958540
rect 478374 958994 479174 990687
rect 478374 958539 478383 958994
rect 479163 958539 479174 958994
rect 478374 958529 479174 958539
rect 525374 958959 526174 992667
rect 526774 992331 527574 993231
rect 526772 992329 527576 992331
rect 526772 992009 526774 992329
rect 527574 992009 527576 992329
rect 526772 992007 527576 992009
rect 525374 958542 525385 958959
rect 526166 958542 526174 958959
rect 525374 958532 526174 958542
rect 526774 958961 527574 992007
rect 528174 991671 528974 993231
rect 528172 991669 528976 991671
rect 528172 991349 528174 991669
rect 528974 991349 528976 991669
rect 528172 991347 528976 991349
rect 526774 958544 526784 958961
rect 527565 958544 527574 958961
rect 526774 958532 527574 958544
rect 528174 958959 528974 991347
rect 529574 991011 530374 993231
rect 529572 991009 530376 991011
rect 529572 990689 529574 991009
rect 530374 990689 530376 991009
rect 529572 990687 530376 990689
rect 528174 958542 528183 958959
rect 528964 958542 528974 958959
rect 528174 958532 528974 958542
rect 529574 958959 530374 990687
rect 529574 958542 529585 958959
rect 530366 958542 530374 958959
rect 529574 958532 530374 958542
rect 335174 958479 335974 958496
rect 537138 958512 541918 958985
rect 537138 956126 537238 958512
rect 541806 956126 541918 958512
rect 537138 955976 541918 956126
rect 547117 958490 551897 958978
rect 547117 956126 547188 958490
rect 551756 956126 551897 958490
rect 547117 955976 551897 956126
rect 533452 954559 627610 954620
rect 533452 954543 625956 954559
rect 533452 953869 533513 954543
rect 535792 953873 625956 954543
rect 627463 953873 627610 954559
rect 535792 953869 627610 953873
rect 533452 953813 627610 953869
rect 622761 953041 624394 953044
rect 533440 952980 624444 953041
rect 533440 952967 622825 952980
rect 533440 952297 533513 952967
rect 535809 952297 622825 952967
rect 533440 952296 622825 952297
rect 624330 952296 624444 952980
rect 533440 952234 624444 952296
rect 622761 952232 624394 952234
rect -31892 912054 -31568 912056
rect -32887 911254 -31890 912054
rect -31570 911987 17454 912054
rect -31570 911315 13333 911987
rect 17205 911315 17454 911987
rect -31570 911254 17454 911315
rect -31892 911252 -31568 911254
rect -32552 910654 -32228 910656
rect -32887 909854 -32550 910654
rect -32230 910585 17454 910654
rect -32230 909913 8334 910585
rect 12206 909913 17454 910585
rect -32230 909854 17454 909913
rect -32552 909852 -32228 909854
rect -30572 909152 -30248 909154
rect -32864 908352 -30570 909152
rect -30250 909069 3737 909152
rect -30250 908397 2875 909069
rect 3547 908397 3737 909069
rect 672940 908906 673254 908908
rect -30250 908352 3737 908397
rect 620554 908835 672942 908906
rect -30572 908350 -30248 908352
rect 620554 908163 625724 908835
rect 629596 908163 672942 908835
rect 620554 908106 672942 908163
rect 673252 908106 673262 908906
rect 672940 908104 673254 908106
rect -31232 907752 -30908 907754
rect -32864 906952 -31230 907752
rect -30910 907680 3737 907752
rect -30910 907008 1690 907680
rect 2362 907008 3737 907680
rect 672280 907506 672604 907508
rect -30910 906952 3737 907008
rect 620554 907447 672282 907506
rect -31232 906950 -30908 906952
rect 620554 906775 620715 907447
rect 624587 906775 672282 907447
rect 620554 906706 672282 906775
rect 672602 906706 673252 907506
rect 672280 906704 672604 906706
rect 671620 906106 671944 906108
rect 628468 906033 671622 906106
rect 628468 905361 636532 906033
rect 637204 905361 671622 906033
rect 628468 905306 671622 905361
rect 671942 905306 673252 906106
rect 671620 905304 671944 905306
rect 670960 904706 671263 904708
rect 628468 904643 670962 904706
rect 628468 903971 637932 904643
rect 638604 903971 670962 904643
rect 628468 903906 670962 903971
rect 671261 903906 673252 904706
rect 670960 903904 671263 903906
rect 781 888076 17286 888232
rect 781 883570 1793 888076
rect 17130 883570 17286 888076
rect 781 883443 17286 883570
rect 620598 883639 639620 883792
rect 620598 879190 620797 883639
rect 638082 879190 639620 883639
rect 620598 878992 639620 879190
rect 889 878028 17274 878192
rect 889 873522 1744 878028
rect 17081 873522 17274 878028
rect 889 873392 17274 873522
rect 620598 873616 639538 873741
rect 620598 869167 620810 873616
rect 638095 869167 639538 873616
rect 620598 868952 639538 869167
rect 1313 803652 5324 803750
rect 1313 799066 4359 803652
rect 5171 799066 5324 803652
rect 1313 798970 5324 799066
rect 633613 794462 639114 794593
rect 1294 793675 5299 793771
rect 1294 789089 4351 793675
rect 5163 789089 5299 793675
rect 633613 789897 633781 794462
rect 635118 789897 639114 794462
rect 633613 789813 639114 789897
rect 1294 788991 5299 789089
rect 633613 784517 639083 784614
rect -30572 783152 -30248 783154
rect -32864 782352 -30570 783152
rect -30250 783067 3784 783152
rect -30250 782395 2881 783067
rect 3553 782395 3784 783067
rect -30250 782352 3784 782395
rect -30572 782350 -30248 782352
rect -31232 781752 -30908 781754
rect -32864 780952 -31230 781752
rect -30910 781706 3784 781752
rect -30910 781034 1701 781706
rect 2373 781034 3784 781706
rect -30910 780952 3784 781034
rect -31232 780950 -30908 780952
rect 633613 779952 633749 784517
rect 635086 779952 639083 784517
rect 633613 779834 639083 779952
rect -31892 765700 -31568 765702
rect -33118 764900 -31890 765700
rect -31570 765636 17345 765700
rect -31570 764964 13329 765636
rect 17201 764964 17345 765636
rect -31570 764900 17345 764964
rect -31892 764898 -31568 764900
rect -32552 764300 -32228 764302
rect -33118 763500 -32550 764300
rect -32230 764241 17345 764300
rect -32230 763569 8334 764241
rect 12206 763569 17345 764241
rect -32230 763500 17345 763569
rect -32552 763498 -32228 763500
rect -30572 739952 -30248 739954
rect -32864 739152 -30570 739952
rect -30250 739880 3753 739952
rect -30250 739208 2886 739880
rect 3558 739208 3753 739880
rect -30250 739152 3753 739208
rect -30572 739150 -30248 739152
rect -31232 738552 -30908 738554
rect -32864 737752 -31230 738552
rect -30910 738497 3753 738552
rect -30910 737825 1690 738497
rect 2362 737825 3753 738497
rect -30910 737752 3753 737825
rect -31232 737750 -30908 737752
rect 672940 730906 673254 730908
rect 620516 730844 672942 730906
rect 620516 730172 625719 730844
rect 629591 730172 672942 730844
rect 620516 730106 672942 730172
rect 673252 730106 673262 730906
rect 672940 730104 673254 730106
rect 672280 729506 672604 729508
rect 620516 729441 672282 729506
rect 620516 728769 620720 729441
rect 624592 728769 672282 729441
rect 620516 728706 672282 728769
rect 672602 728706 673252 729506
rect 672280 728704 672604 728706
rect 671620 728106 671944 728108
rect 636151 728033 671622 728106
rect 636151 727361 636525 728033
rect 637197 727361 671622 728033
rect 636151 727306 671622 727361
rect 671942 727306 673252 728106
rect 671620 727304 671944 727306
rect 670960 726706 671284 726708
rect 636151 726647 670962 726706
rect 636151 725975 637926 726647
rect 638598 725975 670962 726647
rect 636151 725906 670962 725975
rect 671282 725906 673252 726706
rect 670960 725904 671284 725906
rect -31892 722300 -31568 722302
rect -33118 721500 -31890 722300
rect -31570 722236 17360 722300
rect -31570 721564 13337 722236
rect 17209 721564 17360 722236
rect -31570 721500 17360 721564
rect -31892 721498 -31568 721500
rect -32552 720900 -32228 720902
rect -33118 720100 -32550 720900
rect -32230 720830 17360 720900
rect -32230 720158 8330 720830
rect 12202 720158 17360 720830
rect -32230 720100 17360 720158
rect -32552 720098 -32228 720100
rect -30572 696752 -30248 696754
rect -32864 695952 -30570 696752
rect -30250 696699 3721 696752
rect -30250 696027 2892 696699
rect 3564 696027 3721 696699
rect -30250 695952 3721 696027
rect -30572 695950 -30248 695952
rect -31232 695352 -30908 695354
rect -32864 694552 -31230 695352
rect -30910 695294 3721 695352
rect -30910 694622 1695 695294
rect 2367 694622 3721 695294
rect -30910 694552 3721 694622
rect -31232 694550 -30908 694552
rect 672940 685706 673254 685708
rect 620401 685641 672942 685706
rect 620401 684969 625714 685641
rect 629586 684969 672942 685641
rect 620401 684906 672942 684969
rect 673252 684906 673262 685706
rect 672940 684904 673254 684906
rect 672280 684306 672604 684308
rect 620401 684229 672282 684306
rect 620401 683557 620720 684229
rect 624592 683557 672282 684229
rect 620401 683506 672282 683557
rect 672602 683506 673252 684306
rect 672280 683504 672604 683506
rect 671620 682906 671944 682908
rect 636325 682843 671622 682906
rect 636325 682171 636530 682843
rect 637202 682171 671622 682843
rect 636325 682106 671622 682171
rect 671942 682106 673252 682906
rect 671620 682104 671944 682106
rect 670960 681506 671284 681508
rect 636325 681433 670962 681506
rect 636325 680761 637931 681433
rect 638603 680761 670962 681433
rect 636325 680706 670962 680761
rect 671282 680706 673252 681506
rect 670960 680704 671284 680706
rect -31892 679260 -31568 679262
rect -33118 678460 -31890 679260
rect -31570 679189 17376 679260
rect -31570 678517 13348 679189
rect 17220 678517 17376 679189
rect -31570 678460 17376 678517
rect -31892 678458 -31568 678460
rect -32552 677700 -32228 677702
rect -33118 676900 -32550 677700
rect -32230 677639 17376 677700
rect -32230 676967 8334 677639
rect 12206 676967 17376 677639
rect -32230 676900 17376 676967
rect -32552 676898 -32228 676900
rect -30572 653552 -30248 653554
rect -32864 652752 -30570 653552
rect -30250 653496 3768 653552
rect -30250 652824 2886 653496
rect 3558 652824 3768 653496
rect -30250 652752 3768 652824
rect -30572 652750 -30248 652752
rect -31232 652152 -30908 652154
rect -32864 651352 -31230 652152
rect -30910 652074 3768 652152
rect -30910 651402 1684 652074
rect 2356 651402 3768 652074
rect -30910 651352 3768 651402
rect -31232 651350 -30908 651352
rect 672940 640506 673254 640508
rect 620382 640439 672942 640506
rect 620382 639767 625724 640439
rect 629596 639767 672942 640439
rect 620382 639706 672942 639767
rect 673252 639706 673262 640506
rect 672940 639704 673254 639706
rect 672280 639106 672604 639108
rect 620382 639046 672282 639106
rect 620382 638374 620725 639046
rect 624597 638374 672282 639046
rect 620382 638306 672282 638374
rect 672602 638306 673252 639106
rect 672280 638304 672604 638306
rect 671620 637706 671944 637708
rect 636306 637635 671622 637706
rect 636306 636963 636542 637635
rect 637214 636963 671622 637635
rect 636306 636906 671622 636963
rect 671942 636906 673252 637706
rect 671620 636904 671944 636906
rect 670960 636306 671284 636308
rect -31892 636300 -31568 636302
rect -33118 635500 -31890 636300
rect -31570 636226 17423 636300
rect -31570 635554 13337 636226
rect 17209 635554 17423 636226
rect -31570 635500 17423 635554
rect 636306 636237 670962 636306
rect 636306 635565 637921 636237
rect 638593 635565 670962 636237
rect 636306 635506 670962 635565
rect 671282 635506 673252 636306
rect 670960 635504 671284 635506
rect -31892 635498 -31568 635500
rect -32552 634900 -32228 634902
rect -33118 634100 -32550 634900
rect -32230 634839 17423 634900
rect -32230 634167 8342 634839
rect 12214 634167 17423 634839
rect -32230 634100 17423 634167
rect -32552 634098 -32228 634100
rect -30572 610352 -30248 610354
rect -32864 609552 -30570 610352
rect -30250 610292 3753 610352
rect -30250 609620 2903 610292
rect 3575 609620 3753 610292
rect -30250 609552 3753 609620
rect -30572 609550 -30248 609552
rect -31232 608952 -30908 608954
rect -32864 608152 -31230 608952
rect -30910 608921 3753 608952
rect -30910 608249 1690 608921
rect 2362 608249 3753 608921
rect -30910 608152 3753 608249
rect -31232 608150 -30908 608152
rect 672940 595306 673254 595308
rect 620535 595246 672942 595306
rect 620535 594574 625728 595246
rect 629600 594574 672942 595246
rect 620535 594506 672942 594574
rect 673252 594506 673262 595306
rect 672940 594504 673254 594506
rect 672280 593906 672604 593908
rect 620535 593843 672282 593906
rect 620535 593171 620715 593843
rect 624587 593171 672282 593843
rect 620535 593106 672282 593171
rect 672602 593106 673252 593906
rect 672280 593104 672604 593106
rect -31892 592700 -31568 592702
rect -33118 591900 -31890 592700
rect -31570 592638 17376 592700
rect -31570 591966 13340 592638
rect 17212 591966 17376 592638
rect 671620 592506 671944 592508
rect -31570 591900 17376 591966
rect 636171 592442 671622 592506
rect -31892 591898 -31568 591900
rect 636171 591770 636532 592442
rect 637204 591770 671622 592442
rect 636171 591706 671622 591770
rect 671942 591706 673252 592506
rect 671620 591704 671944 591706
rect -32552 591300 -32228 591302
rect -33118 590500 -32550 591300
rect -32230 591232 17376 591300
rect -32230 590560 8330 591232
rect 12202 590560 17376 591232
rect 670960 591106 671284 591108
rect -32230 590500 17376 590560
rect 636171 591039 670962 591106
rect -32552 590498 -32228 590500
rect 636171 590367 637926 591039
rect 638598 590367 670962 591039
rect 636171 590306 670962 590367
rect 671282 590306 673252 591106
rect 670960 590304 671284 590306
rect -30572 567352 -30248 567354
rect -32864 566552 -30570 567352
rect -30250 567309 3706 567352
rect -30250 566637 2897 567309
rect 3569 566637 3706 567309
rect -30250 566552 3706 566637
rect -30572 566550 -30248 566552
rect -31232 565952 -30908 565954
rect -32864 565152 -31230 565952
rect -30910 565887 3706 565952
rect -30910 565215 1684 565887
rect 2356 565215 3706 565887
rect -30910 565152 3706 565215
rect -31232 565150 -30908 565152
rect 672940 550106 673254 550108
rect 620458 550038 672942 550106
rect -31892 549500 -31568 549502
rect -33118 548700 -31890 549500
rect -31570 549436 17470 549500
rect -31570 548764 13341 549436
rect 17213 548764 17470 549436
rect 620458 549366 625728 550038
rect 629600 549366 672942 550038
rect 620458 549306 672942 549366
rect 673252 549306 673262 550106
rect 672940 549304 673254 549306
rect -31570 548700 17470 548764
rect 672280 548706 672604 548708
rect -31892 548698 -31568 548700
rect 620458 548645 672282 548706
rect -32552 548100 -32228 548102
rect -33118 547300 -32550 548100
rect -32230 548047 17470 548100
rect -32230 547375 8330 548047
rect 12202 547375 17470 548047
rect 620458 547973 620725 548645
rect 624597 547973 672282 548645
rect 620458 547906 672282 547973
rect 672602 547906 673252 548706
rect 672280 547904 672604 547906
rect -32230 547300 17470 547375
rect 671620 547306 671944 547308
rect -32552 547298 -32228 547300
rect 636364 547239 671622 547306
rect 636364 546567 636523 547239
rect 637195 546567 671622 547239
rect 636364 546506 671622 546567
rect 671942 546506 673252 547306
rect 671620 546504 671944 546506
rect 670960 545906 671284 545908
rect 636364 545845 670962 545906
rect 636364 545173 637935 545845
rect 638607 545173 670962 545845
rect 636364 545106 670962 545173
rect 671282 545106 673252 545906
rect 670960 545104 671284 545106
rect -30572 524352 -30248 524354
rect -32864 523552 -30570 524352
rect -30250 524275 3784 524352
rect -30250 523603 2903 524275
rect 3575 523603 3784 524275
rect -30250 523552 3784 523603
rect -30572 523550 -30248 523552
rect -31232 522952 -30908 522954
rect -32864 522152 -31230 522952
rect -30910 522887 3784 522952
rect -30910 522215 1673 522887
rect 2345 522215 3784 522887
rect -30910 522152 3784 522215
rect -31232 522150 -30908 522152
rect -31892 506300 -31568 506302
rect -33118 505500 -31890 506300
rect -31570 506240 17407 506300
rect -31570 505568 13337 506240
rect 17209 505568 17407 506240
rect -31570 505500 17407 505568
rect -31892 505498 -31568 505500
rect 672940 504906 673254 504908
rect -32552 504900 -32228 504902
rect -33118 504100 -32550 504900
rect -32230 504838 17407 504900
rect -32230 504166 8323 504838
rect 12195 504166 17407 504838
rect -32230 504100 17407 504166
rect 620554 504840 672942 504906
rect 620554 504168 625714 504840
rect 629586 504168 672942 504840
rect 620554 504106 672942 504168
rect 673252 504106 673262 504906
rect 672940 504104 673254 504106
rect -32552 504098 -32228 504100
rect 672280 503506 672604 503508
rect 620554 503437 672282 503506
rect 620554 502765 620729 503437
rect 624601 502765 672282 503437
rect 620554 502706 672282 502765
rect 672602 502706 673252 503506
rect 672280 502704 672604 502706
rect 671620 502106 671944 502108
rect 636248 502043 671622 502106
rect 636248 501371 636529 502043
rect 637201 501371 671622 502043
rect 636248 501306 671622 501371
rect 671942 501306 673252 502106
rect 671620 501304 671944 501306
rect 670960 500706 671284 500708
rect 636248 500647 670962 500706
rect 636248 499975 637930 500647
rect 638602 499975 670962 500647
rect 636248 499906 670962 499975
rect 671282 499906 673252 500706
rect 670960 499904 671284 499906
rect 630630 479910 639074 479993
rect 630630 475283 630713 479910
rect 632588 475283 639074 479910
rect 630630 475213 639074 475283
rect 630612 469932 639056 470014
rect 630612 465305 630706 469932
rect 632581 465305 639056 469932
rect 630612 465234 639056 465305
rect 672940 461306 673254 461308
rect 620554 461238 672942 461306
rect 620554 460566 625719 461238
rect 629591 460566 672942 461238
rect 620554 460506 672942 460566
rect 673252 460506 673262 461306
rect 672940 460504 673254 460506
rect 672280 459906 672604 459908
rect 620554 459845 672282 459906
rect 620554 459173 620715 459845
rect 624587 459173 672282 459845
rect 1282 459103 7279 459135
rect 620554 459106 672282 459173
rect 672602 459106 673252 459906
rect 672280 459104 672604 459106
rect 1282 454442 6326 459103
rect 7225 454442 7279 459103
rect 671620 458506 671944 458508
rect 636325 458440 671622 458506
rect 636325 457768 636530 458440
rect 637202 457768 671622 458440
rect 636325 457706 671622 457768
rect 671942 457706 673252 458506
rect 671620 457704 671944 457706
rect 670960 457106 671284 457108
rect 636325 457041 670962 457106
rect 636325 456369 637928 457041
rect 638600 456369 670962 457041
rect 636325 456306 670962 456369
rect 671282 456306 673252 457106
rect 670960 456304 671284 456306
rect 1282 454370 7279 454442
rect 1311 449139 7308 449171
rect 1311 444435 6315 449139
rect 7201 444435 7308 449139
rect 1311 444392 7308 444435
rect 625608 435779 639543 435992
rect 625608 431386 625855 435779
rect 638381 431386 639543 435779
rect 625608 431192 639543 431386
rect 625608 425749 639630 425941
rect 625608 421357 625811 425749
rect 638601 421357 639630 425749
rect 625608 421152 639630 421357
rect 904 416868 12379 417032
rect 904 412396 5639 416868
rect 12132 412396 12379 416868
rect 904 412243 12379 412396
rect 890 406832 12365 406992
rect 890 402360 5697 406832
rect 12190 402360 12365 406832
rect 890 402192 12365 402360
rect -30572 396352 -30248 396354
rect -32864 395552 -30570 396352
rect -30250 396279 3690 396352
rect -30250 395607 2903 396279
rect 3575 395607 3690 396279
rect -30250 395552 3690 395607
rect -30572 395550 -30248 395552
rect -31232 394952 -30908 394954
rect -32864 394152 -31230 394952
rect -30910 394896 3690 394952
rect -30910 394224 1690 394896
rect 2362 394224 3690 394896
rect -30910 394152 3690 394224
rect -31232 394150 -30908 394152
rect 633606 391672 639149 391793
rect 633606 387094 633737 391672
rect 635564 387094 639149 391672
rect 633606 387013 639149 387094
rect 633579 381734 639122 381814
rect -31892 378497 -31568 378499
rect -32747 377697 -31890 378497
rect -31570 378423 17407 378497
rect -31570 377751 13329 378423
rect 17201 377751 17407 378423
rect -31570 377697 17407 377751
rect -31892 377695 -31568 377697
rect 633579 377156 633726 381734
rect 635553 377156 639122 381734
rect -32552 377097 -32228 377099
rect -32747 376297 -32550 377097
rect -32230 377036 17407 377097
rect -32230 376364 8334 377036
rect 12206 376364 17407 377036
rect 633579 377034 639122 377156
rect -32230 376297 17407 376364
rect -32552 376295 -32228 376297
rect 672940 372906 673254 372908
rect 620535 372852 672942 372906
rect 620535 372180 625724 372852
rect 629596 372180 672942 372852
rect 620535 372106 672942 372180
rect 673252 372106 673262 372906
rect 672940 372104 673254 372106
rect 672280 371506 672604 371508
rect 620535 371449 672282 371506
rect 620535 370777 620720 371449
rect 624592 370777 672282 371449
rect 620535 370706 672282 370777
rect 672602 370706 673252 371506
rect 672280 370704 672604 370706
rect 671620 370106 671944 370108
rect 636306 370039 671622 370106
rect 636306 369367 636529 370039
rect 637201 369367 671622 370039
rect 636306 369306 671622 369367
rect 671942 369306 673252 370106
rect 671620 369304 671944 369306
rect 670960 368706 671284 368708
rect 636306 368635 670962 368706
rect 636306 367963 637929 368635
rect 638601 367963 670962 368635
rect 636306 367906 670962 367963
rect 671282 367906 673252 368706
rect 670960 367904 671284 367906
rect -30572 353352 -30248 353354
rect -32864 352552 -30570 353352
rect -30250 353296 3800 353352
rect -30250 352624 2886 353296
rect 3558 352624 3800 353296
rect -30250 352552 3800 352624
rect -30572 352550 -30248 352552
rect -31232 351952 -30908 351954
rect -32864 351152 -31230 351952
rect -30910 351879 3800 351952
rect -30910 351207 1684 351879
rect 2356 351207 3800 351879
rect -30910 351152 3800 351207
rect -31232 351150 -30908 351152
rect -31892 335297 -31568 335299
rect -32747 334497 -31890 335297
rect -31570 335232 17454 335297
rect -31570 334560 13329 335232
rect 17201 334560 17454 335232
rect -31570 334497 17454 334560
rect -31892 334495 -31568 334497
rect -32552 333897 -32228 333899
rect -32747 333097 -32550 333897
rect -32230 333829 17454 333897
rect -32230 333157 8342 333829
rect 12214 333157 17454 333829
rect -32230 333097 17454 333157
rect -32552 333095 -32228 333097
rect 672940 328106 673254 328108
rect 620554 328050 672942 328106
rect 620554 327378 625724 328050
rect 629596 327378 672942 328050
rect 620554 327306 672942 327378
rect 673252 327306 673262 328106
rect 672940 327304 673254 327306
rect 672280 326706 672604 326708
rect 620554 326666 672282 326706
rect 620554 325994 620729 326666
rect 624601 325994 672282 326666
rect 620554 325906 672282 325994
rect 672602 325906 673252 326706
rect 672280 325904 672604 325906
rect 671620 325306 671944 325308
rect 636267 325237 671622 325306
rect 636267 324565 636529 325237
rect 637201 324565 671622 325237
rect 636267 324506 671622 324565
rect 671942 324506 673252 325306
rect 671620 324504 671944 324506
rect 670960 323906 671284 323908
rect 636267 323860 670962 323906
rect 636267 323188 637924 323860
rect 638596 323188 670962 323860
rect 636267 323106 670962 323188
rect 671282 323106 673252 323906
rect 670960 323104 671284 323106
rect -30572 310352 -30248 310354
rect -32864 309552 -30570 310352
rect -30250 310312 3690 310352
rect -30250 309640 2875 310312
rect 3547 309640 3690 310312
rect -30250 309552 3690 309640
rect -30572 309550 -30248 309552
rect -31232 308952 -30908 308954
rect -32864 308152 -31230 308952
rect -30910 308884 3690 308952
rect -30910 308212 1673 308884
rect 2345 308212 3690 308884
rect -30910 308152 3690 308212
rect -31232 308150 -30908 308152
rect -31892 292097 -31568 292099
rect -32747 291297 -31890 292097
rect -31570 292032 17414 292097
rect -31570 291360 13329 292032
rect 17201 291360 17414 292032
rect -31570 291297 17414 291360
rect -31892 291295 -31568 291297
rect -32552 290697 -32228 290699
rect -32747 289897 -32550 290697
rect -32230 290622 17414 290697
rect -32230 289950 8332 290622
rect 12204 289950 17414 290622
rect -32230 289897 17414 289950
rect -32552 289895 -32228 289897
rect 672940 283306 673254 283308
rect 620592 283228 672942 283306
rect 620592 282556 625724 283228
rect 629596 282556 672942 283228
rect 620592 282506 672942 282556
rect 673252 282506 673262 283306
rect 672940 282504 673254 282506
rect 672280 281906 672604 281908
rect 620592 281849 672282 281906
rect 620592 281177 620734 281849
rect 624606 281177 672282 281849
rect 620592 281106 672282 281177
rect 672602 281106 673252 281906
rect 672280 281104 672604 281106
rect 671620 280506 671944 280508
rect 636286 280444 671622 280506
rect 636286 279772 636524 280444
rect 637196 279772 671622 280444
rect 636286 279706 671622 279772
rect 671942 279706 673252 280506
rect 671620 279704 671944 279706
rect 670960 279106 671284 279108
rect 636286 279039 670962 279106
rect 636286 278367 637915 279039
rect 638587 278367 670962 279039
rect 636286 278306 670962 278367
rect 671282 278306 673252 279106
rect 670960 278304 671284 278306
rect -30572 267352 -30248 267354
rect -32864 266552 -30570 267352
rect -30250 267292 3839 267352
rect -30250 266620 2884 267292
rect 3556 266620 3839 267292
rect -30250 266552 3839 266620
rect -30572 266550 -30248 266552
rect -31232 265952 -30908 265954
rect -32864 265152 -31230 265952
rect -30910 265891 3839 265952
rect -30910 265219 1684 265891
rect 2356 265219 3839 265891
rect -30910 265152 3839 265219
rect -31232 265150 -30908 265152
rect -31892 248897 -31568 248899
rect -32747 248097 -31890 248897
rect -31570 248824 17531 248897
rect -31570 248152 13328 248824
rect 17200 248152 17531 248824
rect -31570 248097 17531 248152
rect -31892 248095 -31568 248097
rect -32552 247497 -32228 247499
rect -32747 246697 -32550 247497
rect -32230 247417 17531 247497
rect -32230 246745 8332 247417
rect 12204 246745 17531 247417
rect -32230 246697 17531 246745
rect -32552 246695 -32228 246697
rect 672940 237906 673254 237908
rect 620482 237845 672942 237906
rect 620482 237173 625723 237845
rect 629595 237173 672942 237845
rect 620482 237106 672942 237173
rect 673252 237106 673262 237906
rect 672940 237104 673254 237106
rect 672280 236506 672604 236508
rect 620482 236448 672282 236506
rect 620482 235776 620702 236448
rect 624574 235776 672282 236448
rect 620482 235706 672282 235776
rect 672602 235706 673252 236506
rect 672280 235704 672604 235706
rect 671620 235106 671944 235108
rect 636287 235036 671622 235106
rect 636287 234364 636532 235036
rect 637204 234364 671622 235036
rect 636287 234306 671622 234364
rect 671942 234306 673252 235106
rect 671620 234304 671944 234306
rect 670960 233706 671284 233708
rect 636287 233650 670962 233706
rect 636287 232978 637933 233650
rect 638605 232978 670962 233650
rect 636287 232906 670962 232978
rect 671282 232906 673252 233706
rect 670960 232904 671284 232906
rect -30572 224352 -30248 224354
rect -32864 223552 -30570 224352
rect -30250 224294 3739 224352
rect -30250 223622 2881 224294
rect 3553 223622 3739 224294
rect -30250 223552 3739 223622
rect -30572 223550 -30248 223552
rect -31232 222952 -30908 222954
rect -32864 222152 -31230 222952
rect -30910 222893 3739 222952
rect -30910 222221 1684 222893
rect 2356 222221 3739 222893
rect -30910 222152 3739 222221
rect -31232 222150 -30908 222152
rect -31892 205697 -31568 205699
rect -32747 204897 -31890 205697
rect -31570 205628 6462 205697
rect -31570 204956 5686 205628
rect 6358 204956 6462 205628
rect -31570 204897 6462 204956
rect -31892 204895 -31568 204897
rect -32552 204297 -32228 204299
rect -32747 203497 -32550 204297
rect -32230 204225 6462 204297
rect -32230 203553 4289 204225
rect 4961 203553 6462 204225
rect -32230 203497 6462 203553
rect -32552 203495 -32228 203497
rect 629374 196101 638718 196190
rect 629374 195247 637917 196101
rect 629374 193669 629587 195247
rect 632313 193669 637917 195247
rect 629374 193295 637917 193669
rect 638627 193295 638718 196101
rect 629374 193254 638718 193295
rect 637861 193229 638663 193254
rect 672940 192506 673254 192508
rect 633429 192443 672942 192506
rect 633429 191771 635130 192443
rect 635802 191771 672942 192443
rect 633429 191706 672942 191771
rect 673252 191706 673262 192506
rect 672940 191704 673254 191706
rect 672280 191106 672604 191108
rect 633429 191042 672282 191106
rect 633429 190370 633732 191042
rect 634404 190370 672282 191042
rect 633429 190306 672282 190370
rect 672602 190306 673252 191106
rect 672280 190304 672604 190306
rect 671620 189706 671944 189708
rect 636198 189642 671622 189706
rect 636198 188970 636525 189642
rect 637197 188970 671622 189642
rect 636198 188906 671622 188970
rect 671942 188906 673252 189706
rect 671620 188904 671944 188906
rect 670960 188306 671284 188308
rect 636198 188248 670962 188306
rect 636198 187576 637919 188248
rect 638591 187576 670962 188248
rect 636198 187506 670962 187576
rect 671282 187506 673252 188306
rect 670960 187504 671284 187506
rect -30572 181352 -30248 181354
rect -32864 180552 -30570 181352
rect -30250 181286 3814 181352
rect -30250 180614 2887 181286
rect 3561 180614 3814 181286
rect -30250 180552 3814 180614
rect -30572 180550 -30248 180552
rect -31232 179952 -30908 179954
rect -32864 179152 -31230 179952
rect -30910 179924 3814 179952
rect -30910 179188 1653 179924
rect 2388 179188 3814 179924
rect -30910 179152 3814 179188
rect -31232 179150 -30908 179152
rect -31892 162497 -31568 162499
rect -32747 161697 -31890 162497
rect -31570 162450 6497 162497
rect -31570 161736 5662 162450
rect 6387 161736 6497 162450
rect -31570 161697 6497 161736
rect -31892 161695 -31568 161697
rect -32552 161097 -32228 161099
rect -32747 160297 -32550 161097
rect -32230 161066 5094 161097
rect -32230 160352 4258 161066
rect 4983 160352 5094 161066
rect -32230 160297 5094 160352
rect -32552 160295 -32228 160297
rect 672940 147106 673254 147108
rect 633446 147047 672942 147106
rect 633446 146375 635130 147047
rect 635802 146375 672942 147047
rect 633446 146306 672942 146375
rect 673252 146306 673262 147106
rect 672940 146304 673254 146306
rect 672280 145706 672604 145708
rect 633446 145639 672282 145706
rect 633446 144967 633731 145639
rect 634403 144967 672282 145639
rect 633446 144906 672282 144967
rect 672602 144906 673252 145706
rect 672280 144904 672604 144906
rect 671620 144306 671944 144308
rect 636325 144235 671622 144306
rect 636325 143563 636523 144235
rect 637195 143563 671622 144235
rect 636325 143506 671622 143563
rect 671942 143506 673252 144306
rect 671620 143504 671944 143506
rect 670960 142906 671284 142908
rect 636325 142842 670962 142906
rect 636325 142170 637930 142842
rect 638602 142170 670962 142842
rect 636325 142106 670962 142170
rect 671282 142106 673252 142906
rect 670960 142104 671284 142106
rect 672940 101706 673254 101708
rect 633407 101637 672942 101706
rect 633407 100965 635134 101637
rect 635806 100965 672942 101637
rect 633407 100906 672942 100965
rect 673252 100906 673272 101706
rect 672940 100904 673254 100906
rect 672280 100306 672604 100308
rect 633407 100241 672282 100306
rect 633407 99569 633728 100241
rect 634400 99569 672282 100241
rect 633407 99506 672282 99569
rect 672602 99506 673252 100306
rect 672280 99504 672604 99506
rect 671620 98906 671944 98908
rect 636364 98843 671622 98906
rect 636364 98171 636533 98843
rect 637205 98171 671622 98843
rect 636364 98106 671622 98171
rect 671942 98106 673252 98906
rect 671620 98104 671944 98106
rect 670960 97506 671284 97508
rect 636364 97439 670962 97506
rect 636364 96767 637931 97439
rect 638603 96767 670962 97439
rect 636364 96706 670962 96767
rect 671282 96706 673252 97506
rect 670960 96704 671284 96706
rect 1333 86219 13326 86350
rect 1333 81681 10344 86219
rect 13143 81681 13326 86219
rect 1333 81570 13326 81681
rect 1333 76201 13326 76371
rect 1333 71741 10357 76201
rect 13169 71741 13326 76201
rect 1333 71591 13326 71741
rect 770 44026 9140 44232
rect 770 39587 1813 44026
rect 8962 39587 9140 44026
rect 770 39443 9140 39587
rect 583 34000 9140 34192
rect 583 29539 1559 34000
rect 8951 29539 9140 34000
rect 583 29392 9140 29539
rect 202699 14752 207488 15025
rect 202699 9725 202830 14752
rect 207269 9725 207488 14752
rect 104417 8932 104782 8947
rect 104417 8494 104438 8932
rect 104417 8473 104782 8494
rect 104421 8407 104782 8473
rect 104421 7931 108616 8407
rect 107896 3755 108610 7931
rect 107896 1861 107928 3755
rect 108561 1861 108610 3755
rect 107896 1818 108610 1861
rect 202699 620 207488 9725
rect 212739 14720 217539 15025
rect 212739 9693 212909 14720
rect 217348 9693 217539 14720
rect 212739 599 217539 9693
rect 530581 6582 535361 6705
rect 530581 2784 530645 6582
rect 535200 2784 535361 6582
rect 530581 1218 535361 2784
rect 540560 6573 545340 6714
rect 540560 2775 540643 6573
rect 545198 2775 545340 6573
rect 540560 1227 545340 2775
<< via3 >>
rect 72974 992669 73774 992989
rect 74374 992009 75174 992329
rect 72991 958573 73764 959024
rect 75774 991349 76574 991669
rect 74394 958579 75167 959030
rect 124574 992669 125374 992989
rect 77174 990689 77974 991009
rect 75792 958575 76565 959026
rect 125974 992009 126774 992329
rect 124589 958529 125363 959028
rect 127374 991349 128174 991669
rect 125991 958532 126765 959031
rect 176174 992669 176974 992989
rect 128774 990689 129574 991009
rect 127385 958529 128159 959028
rect 128784 958533 129558 959032
rect 177574 992009 178374 992329
rect 176183 958556 176965 959022
rect 178974 991349 179774 991669
rect 177584 958554 178366 959020
rect 227774 992669 228574 992989
rect 180374 990689 181174 991009
rect 178983 958551 179765 959017
rect 180385 958555 181167 959021
rect 229174 992009 229974 992329
rect 227789 958561 228562 958978
rect 230574 991349 231374 991669
rect 229185 958557 229958 958974
rect 279374 992669 280174 992989
rect 231974 990689 232774 991009
rect 230588 958560 231361 958977
rect 231989 958559 232762 958976
rect 280774 992009 281574 992329
rect 279382 958539 280164 958993
rect 282174 991349 282974 991669
rect 280782 958539 281564 958993
rect 330974 992669 331774 992989
rect 283574 990689 284374 991009
rect 282187 958541 282969 958995
rect 283583 958540 284365 958994
rect 332374 992009 333174 992329
rect 330988 958495 331755 959011
rect 333774 991349 334574 991669
rect 332390 958498 333157 959014
rect 396974 992669 397774 992989
rect 335174 990689 335974 991009
rect 333791 958492 334558 959008
rect 335195 958496 335962 959012
rect 398374 992009 399174 992329
rect 396986 958530 397765 958982
rect 399774 991349 400574 991669
rect 398383 958528 399162 958980
rect 474174 992669 474974 992989
rect 401174 990689 401974 991009
rect 399783 958528 400562 958980
rect 401186 958530 401965 958982
rect 475574 992009 476374 992329
rect 474185 958538 474965 958993
rect 476974 991349 477774 991669
rect 475583 958537 476363 958992
rect 525374 992669 526174 992989
rect 478374 990689 479174 991009
rect 476985 958540 477765 958995
rect 478383 958539 479163 958994
rect 526774 992009 527574 992329
rect 525385 958542 526166 958959
rect 528174 991349 528974 991669
rect 526784 958544 527565 958961
rect 529574 990689 530374 991009
rect 528183 958542 528964 958959
rect 529585 958542 530366 958959
rect 537238 956126 541806 958512
rect 547188 956126 551756 958490
rect 533513 953869 535792 954543
rect 625956 953873 627463 954559
rect 533513 952297 535809 952967
rect 622825 952296 624330 952980
rect -31890 911254 -31570 912054
rect 13333 911315 17205 911987
rect -32550 909854 -32230 910654
rect 8334 909913 12206 910585
rect -30570 908352 -30250 909152
rect 2875 908397 3547 909069
rect 625724 908163 629596 908835
rect 672942 908106 673252 908906
rect -31230 906952 -30910 907752
rect 1690 907008 2362 907680
rect 620715 906775 624587 907447
rect 672282 906706 672602 907506
rect 636532 905361 637204 906033
rect 671622 905306 671942 906106
rect 637932 903971 638604 904643
rect 670962 903906 671261 904706
rect 1793 883570 17130 888076
rect 620797 879190 638082 883639
rect 1744 873522 17081 878028
rect 620810 869167 638095 873616
rect 4359 799066 5171 803652
rect 4351 789089 5163 793675
rect 633781 789897 635118 794462
rect -30570 782352 -30250 783152
rect 2881 782395 3553 783067
rect -31230 780952 -30910 781752
rect 1701 781034 2373 781706
rect 633749 779952 635086 784517
rect -31890 764900 -31570 765700
rect 13329 764964 17201 765636
rect -32550 763500 -32230 764300
rect 8334 763569 12206 764241
rect -30570 739152 -30250 739952
rect 2886 739208 3558 739880
rect -31230 737752 -30910 738552
rect 1690 737825 2362 738497
rect 625719 730172 629591 730844
rect 672942 730106 673252 730906
rect 620720 728769 624592 729441
rect 672282 728706 672602 729506
rect 636525 727361 637197 728033
rect 671622 727306 671942 728106
rect 637926 725975 638598 726647
rect 670962 725906 671282 726706
rect -31890 721500 -31570 722300
rect 13337 721564 17209 722236
rect -32550 720100 -32230 720900
rect 8330 720158 12202 720830
rect -30570 695952 -30250 696752
rect 2892 696027 3564 696699
rect -31230 694552 -30910 695352
rect 1695 694622 2367 695294
rect 625714 684969 629586 685641
rect 672942 684906 673252 685706
rect 620720 683557 624592 684229
rect 672282 683506 672602 684306
rect 636530 682171 637202 682843
rect 671622 682106 671942 682906
rect 637931 680761 638603 681433
rect 670962 680706 671282 681506
rect -31890 678460 -31570 679260
rect 13348 678517 17220 679189
rect -32550 676900 -32230 677700
rect 8334 676967 12206 677639
rect -30570 652752 -30250 653552
rect 2886 652824 3558 653496
rect -31230 651352 -30910 652152
rect 1684 651402 2356 652074
rect 625724 639767 629596 640439
rect 672942 639706 673252 640506
rect 620725 638374 624597 639046
rect 672282 638306 672602 639106
rect 636542 636963 637214 637635
rect 671622 636906 671942 637706
rect -31890 635500 -31570 636300
rect 13337 635554 17209 636226
rect 637921 635565 638593 636237
rect 670962 635506 671282 636306
rect -32550 634100 -32230 634900
rect 8342 634167 12214 634839
rect -30570 609552 -30250 610352
rect 2903 609620 3575 610292
rect -31230 608152 -30910 608952
rect 1690 608249 2362 608921
rect 625728 594574 629600 595246
rect 672942 594506 673252 595306
rect 620715 593171 624587 593843
rect 672282 593106 672602 593906
rect -31890 591900 -31570 592700
rect 13340 591966 17212 592638
rect 636532 591770 637204 592442
rect 671622 591706 671942 592506
rect -32550 590500 -32230 591300
rect 8330 590560 12202 591232
rect 637926 590367 638598 591039
rect 670962 590306 671282 591106
rect -30570 566552 -30250 567352
rect 2897 566637 3569 567309
rect -31230 565152 -30910 565952
rect 1684 565215 2356 565887
rect -31890 548700 -31570 549500
rect 13341 548764 17213 549436
rect 625728 549366 629600 550038
rect 672942 549306 673252 550106
rect -32550 547300 -32230 548100
rect 8330 547375 12202 548047
rect 620725 547973 624597 548645
rect 672282 547906 672602 548706
rect 636523 546567 637195 547239
rect 671622 546506 671942 547306
rect 637935 545173 638607 545845
rect 670962 545106 671282 545906
rect -30570 523552 -30250 524352
rect 2903 523603 3575 524275
rect -31230 522152 -30910 522952
rect 1673 522215 2345 522887
rect -31890 505500 -31570 506300
rect 13337 505568 17209 506240
rect -32550 504100 -32230 504900
rect 8323 504166 12195 504838
rect 625714 504168 629586 504840
rect 672942 504106 673252 504906
rect 620729 502765 624601 503437
rect 672282 502706 672602 503506
rect 636529 501371 637201 502043
rect 671622 501306 671942 502106
rect 637930 499975 638602 500647
rect 670962 499906 671282 500706
rect 630713 475283 632588 479910
rect 630706 465305 632581 469932
rect 625719 460566 629591 461238
rect 672942 460506 673252 461306
rect 620715 459173 624587 459845
rect 672282 459106 672602 459906
rect 6326 454442 7225 459103
rect 636530 457768 637202 458440
rect 671622 457706 671942 458506
rect 637928 456369 638600 457041
rect 670962 456306 671282 457106
rect 6315 444435 7201 449139
rect 625855 431386 638381 435779
rect 625811 421357 638601 425749
rect 5639 412396 12132 416868
rect 5697 402360 12190 406832
rect -30570 395552 -30250 396352
rect 2903 395607 3575 396279
rect -31230 394152 -30910 394952
rect 1690 394224 2362 394896
rect 633737 387094 635564 391672
rect -31890 377697 -31570 378497
rect 13329 377751 17201 378423
rect 633726 377156 635553 381734
rect -32550 376297 -32230 377097
rect 8334 376364 12206 377036
rect 625724 372180 629596 372852
rect 672942 372106 673252 372906
rect 620720 370777 624592 371449
rect 672282 370706 672602 371506
rect 636529 369367 637201 370039
rect 671622 369306 671942 370106
rect 637929 367963 638601 368635
rect 670962 367906 671282 368706
rect -30570 352552 -30250 353352
rect 2886 352624 3558 353296
rect -31230 351152 -30910 351952
rect 1684 351207 2356 351879
rect -31890 334497 -31570 335297
rect 13329 334560 17201 335232
rect -32550 333097 -32230 333897
rect 8342 333157 12214 333829
rect 625724 327378 629596 328050
rect 672942 327306 673252 328106
rect 620729 325994 624601 326666
rect 672282 325906 672602 326706
rect 636529 324565 637201 325237
rect 671622 324506 671942 325306
rect 637924 323188 638596 323860
rect 670962 323106 671282 323906
rect -30570 309552 -30250 310352
rect 2875 309640 3547 310312
rect -31230 308152 -30910 308952
rect 1673 308212 2345 308884
rect -31890 291297 -31570 292097
rect 13329 291360 17201 292032
rect -32550 289897 -32230 290697
rect 8332 289950 12204 290622
rect 625724 282556 629596 283228
rect 672942 282506 673252 283306
rect 620734 281177 624606 281849
rect 672282 281106 672602 281906
rect 636524 279772 637196 280444
rect 671622 279706 671942 280506
rect 637915 278367 638587 279039
rect 670962 278306 671282 279106
rect -30570 266552 -30250 267352
rect 2884 266620 3556 267292
rect -31230 265152 -30910 265952
rect 1684 265219 2356 265891
rect -31890 248097 -31570 248897
rect 13328 248152 17200 248824
rect -32550 246697 -32230 247497
rect 8332 246745 12204 247417
rect 625723 237173 629595 237845
rect 672942 237106 673252 237906
rect 620702 235776 624574 236448
rect 672282 235706 672602 236506
rect 636532 234364 637204 235036
rect 671622 234306 671942 235106
rect 637933 232978 638605 233650
rect 670962 232906 671282 233706
rect -30570 223552 -30250 224352
rect 2881 223622 3553 224294
rect -31230 222152 -30910 222952
rect 1684 222221 2356 222893
rect -31890 204897 -31570 205697
rect 5686 204956 6358 205628
rect -32550 203497 -32230 204297
rect 4289 203553 4961 204225
rect 629587 193669 632313 195247
rect 637917 193295 638627 196101
rect 635130 191771 635802 192443
rect 672942 191706 673252 192506
rect 633732 190370 634404 191042
rect 672282 190306 672602 191106
rect 636525 188970 637197 189642
rect 671622 188906 671942 189706
rect 637919 187576 638591 188248
rect 670962 187506 671282 188306
rect -30570 180552 -30250 181352
rect 2887 180614 3561 181286
rect -31230 179152 -30910 179952
rect 1653 179188 2388 179924
rect -31890 161697 -31570 162497
rect 5662 161736 6387 162450
rect -32550 160297 -32230 161097
rect 4258 160352 4983 161066
rect 635130 146375 635802 147047
rect 672942 146306 673252 147106
rect 633731 144967 634403 145639
rect 672282 144906 672602 145706
rect 636523 143563 637195 144235
rect 671622 143506 671942 144306
rect 637930 142170 638602 142842
rect 670962 142106 671282 142906
rect 635134 100965 635806 101637
rect 672942 100906 673252 101706
rect 633728 99569 634400 100241
rect 672282 99506 672602 100306
rect 636533 98171 637205 98843
rect 671622 98106 671942 98906
rect 637931 96767 638603 97439
rect 670962 96706 671282 97506
rect 10344 81681 13143 86219
rect 10357 71741 13169 76201
rect 1813 39587 8962 44026
rect 1559 29539 8951 34000
rect 202830 9725 207269 14752
rect 104438 8494 104782 8932
rect 107928 1861 108561 3755
rect 212909 9693 217348 14720
rect 530645 2784 535200 6582
rect 540643 2775 545198 6573
<< metal4 >>
rect 72972 992989 73776 992991
rect 124572 992989 125376 992991
rect 176172 992989 176976 992991
rect 227772 992989 228576 992991
rect 279372 992989 280176 992991
rect 330972 992989 331776 992991
rect 396972 992989 397776 992991
rect 474172 992989 474976 992991
rect 525372 992989 526176 992991
rect 71723 992669 72974 992989
rect 73774 992669 78092 992989
rect 123275 992669 124574 992989
rect 125374 992669 129653 992989
rect 174659 992669 176174 992989
rect 176974 992669 181283 992989
rect 226182 992669 227774 992989
rect 228574 992669 232884 992989
rect 277805 992669 279374 992989
rect 280174 992669 284465 992989
rect 328183 992669 330974 992989
rect 331774 992669 336125 992989
rect 395605 992669 396974 992989
rect 397774 992669 402054 992989
rect 472492 992669 474174 992989
rect 474974 992669 479264 992989
rect 523827 992669 525374 992989
rect 526174 992669 530491 992989
rect 72972 992667 73776 992669
rect 124572 992667 125376 992669
rect 176172 992667 176976 992669
rect 227772 992667 228576 992669
rect 279372 992667 280176 992669
rect 330972 992667 331776 992669
rect 396972 992667 397776 992669
rect 474172 992667 474976 992669
rect 525372 992667 526176 992669
rect 74372 992329 75176 992331
rect 125972 992329 126776 992331
rect 177572 992329 178376 992331
rect 229172 992329 229976 992331
rect 280772 992329 281576 992331
rect 332372 992329 333176 992331
rect 398372 992329 399176 992331
rect 475572 992329 476376 992331
rect 526772 992329 527576 992331
rect 71242 992009 74374 992329
rect 75174 992009 78111 992329
rect 122745 992009 125974 992329
rect 126774 992009 129663 992329
rect 174050 992009 177574 992329
rect 178374 992009 181293 992329
rect 225545 992009 229174 992329
rect 229974 992009 232864 992329
rect 277145 992009 280774 992329
rect 281574 992009 284485 992329
rect 327436 992009 332374 992329
rect 333174 992009 336115 992329
rect 394919 992009 398374 992329
rect 399174 992009 402074 992329
rect 471912 992009 475574 992329
rect 476374 992009 479244 992329
rect 523159 992009 526774 992329
rect 527574 992009 530461 992329
rect 74372 992007 75176 992009
rect 125972 992007 126776 992009
rect 177572 992007 178376 992009
rect 229172 992007 229976 992009
rect 280772 992007 281576 992009
rect 332372 992007 333176 992009
rect 398372 992007 399176 992009
rect 475572 992007 476376 992009
rect 526772 992007 527576 992009
rect 75772 991669 76576 991671
rect 127372 991669 128176 991671
rect 178972 991669 179776 991671
rect 230572 991669 231376 991671
rect 282172 991669 282976 991671
rect 333772 991669 334576 991671
rect 399772 991669 400576 991671
rect 476972 991669 477776 991671
rect 528172 991669 528976 991671
rect 70602 991349 75774 991669
rect 76574 991349 78121 991669
rect 122085 991349 127374 991669
rect 128174 991349 129663 991669
rect 173440 991349 178974 991669
rect 179774 991349 181323 991669
rect 224854 991349 230574 991669
rect 231374 991349 232854 991669
rect 276376 991349 282174 991669
rect 282974 991349 284475 991669
rect 326757 991349 333774 991669
rect 334574 991349 336105 991669
rect 394162 991349 399774 991669
rect 400574 991349 402074 991669
rect 471285 991349 476974 991669
rect 477774 991349 479244 991669
rect 522578 991349 528174 991669
rect 528974 991349 530500 991669
rect 75772 991347 76576 991349
rect 127372 991347 128176 991349
rect 178972 991347 179776 991349
rect 230572 991347 231376 991349
rect 282172 991347 282976 991349
rect 333772 991347 334576 991349
rect 399772 991347 400576 991349
rect 476972 991347 477776 991349
rect 528172 991347 528976 991349
rect 77172 991009 77976 991011
rect 128772 991009 129576 991011
rect 180372 991009 181176 991011
rect 231972 991009 232776 991011
rect 283572 991009 284376 991011
rect 335172 991009 335976 991011
rect 401172 991009 401976 991011
rect 478372 991009 479176 991011
rect 529572 991009 530376 991011
rect 70025 990689 77174 991009
rect 77974 990689 78131 991009
rect 121387 990689 128774 991009
rect 129574 990689 129712 991009
rect 172820 990689 180374 991009
rect 181174 990689 181332 991009
rect 224225 990689 231974 991009
rect 232774 990689 232874 991009
rect 275825 990689 283574 991009
rect 284374 990689 284534 991009
rect 326225 990689 335174 991009
rect 335974 990689 336095 991009
rect 393625 990689 401174 991009
rect 401974 990689 402064 991009
rect 470594 990689 478374 991009
rect 479174 990689 479254 991009
rect 521988 990689 529574 991009
rect 530374 990689 530461 991009
rect 77172 990687 77976 990689
rect 128772 990687 129576 990689
rect 180372 990687 181176 990689
rect 231972 990687 232776 990689
rect 283572 990687 284376 990689
rect 335172 990687 335976 990689
rect 401172 990687 401976 990689
rect 478372 990687 479176 990689
rect 529572 990687 530376 990689
rect 72974 959024 73774 959038
rect 72974 958573 72991 959024
rect 73764 958573 73774 959024
rect 9771 955176 10560 955289
rect 9771 947452 10560 954376
rect 72974 955115 73774 958573
rect 72974 954443 73036 955115
rect 73708 954443 73774 955115
rect 14566 953659 15343 953844
rect 14566 946390 15343 952859
rect 72974 952631 73774 954443
rect 74374 959030 75174 959038
rect 74374 958579 74394 959030
rect 75167 958579 75174 959030
rect 74374 953598 75174 958579
rect 74374 952926 74441 953598
rect 75113 952926 75174 953598
rect 74374 952631 75174 952926
rect 75774 959026 76574 959038
rect 75774 958575 75792 959026
rect 76565 958575 76574 959026
rect 75774 958188 76574 958575
rect 75774 957516 75849 958188
rect 76521 957516 76574 958188
rect 75774 952631 76574 957516
rect 77174 956684 77974 959038
rect 77174 956012 77228 956684
rect 77900 956012 77974 956684
rect 77174 952631 77974 956012
rect 124574 959028 125374 959039
rect 124574 958529 124589 959028
rect 125363 958529 125374 959028
rect 124574 955113 125374 958529
rect 124574 954441 124635 955113
rect 125307 954441 125374 955113
rect 124574 952631 125374 954441
rect 125974 959031 126774 959039
rect 125974 958532 125991 959031
rect 126765 958532 126774 959031
rect 125974 953592 126774 958532
rect 125974 952920 126040 953592
rect 126712 952920 126774 953592
rect 125974 952631 126774 952920
rect 127374 959028 128174 959039
rect 127374 958529 127385 959028
rect 128159 958529 128174 959028
rect 127374 958192 128174 958529
rect 127374 957520 127441 958192
rect 128113 957520 128174 958192
rect 127374 952631 128174 957520
rect 128774 959032 129574 959039
rect 128774 958533 128784 959032
rect 129558 958533 129574 959032
rect 128774 956698 129574 958533
rect 128774 956026 128823 956698
rect 129495 956026 129574 956698
rect 128774 952631 129574 956026
rect 176174 959022 176974 959034
rect 176174 958556 176183 959022
rect 176965 958556 176974 959022
rect 176174 955114 176974 958556
rect 176174 954442 176246 955114
rect 176918 954442 176974 955114
rect 176174 952631 176974 954442
rect 177574 959020 178374 959034
rect 177574 958554 177584 959020
rect 178366 958554 178374 959020
rect 177574 953588 178374 958554
rect 177574 952916 177636 953588
rect 178308 952916 178374 953588
rect 177574 952631 178374 952916
rect 178974 959017 179774 959034
rect 178974 958551 178983 959017
rect 179765 958551 179774 959017
rect 178974 958198 179774 958551
rect 178974 957526 179045 958198
rect 179717 957526 179774 958198
rect 178974 952631 179774 957526
rect 180374 959021 181174 959034
rect 180374 958555 180385 959021
rect 181167 958555 181174 959021
rect 330974 959011 331774 959027
rect 180374 956687 181174 958555
rect 180374 956015 180427 956687
rect 181099 956015 181174 956687
rect 180374 952631 181174 956015
rect 227774 958978 228574 958995
rect 227774 958561 227789 958978
rect 228562 958561 228574 958978
rect 227774 955118 228574 958561
rect 227774 954446 227824 955118
rect 228496 954446 228574 955118
rect 227774 952631 228574 954446
rect 229174 958974 229974 958995
rect 229174 958557 229185 958974
rect 229958 958557 229974 958974
rect 229174 953587 229974 958557
rect 229174 952915 229234 953587
rect 229906 952915 229974 953587
rect 229174 952631 229974 952915
rect 230574 958977 231374 958995
rect 230574 958560 230588 958977
rect 231361 958560 231374 958977
rect 230574 958196 231374 958560
rect 230574 957524 230640 958196
rect 231312 957524 231374 958196
rect 230574 952631 231374 957524
rect 231974 958976 232774 958995
rect 231974 958559 231989 958976
rect 232762 958559 232774 958976
rect 231974 956688 232774 958559
rect 231974 956016 232030 956688
rect 232702 956016 232774 956688
rect 231974 952631 232774 956016
rect 279374 958993 280174 959001
rect 279374 958539 279382 958993
rect 280164 958539 280174 958993
rect 279374 955108 280174 958539
rect 279374 954436 279439 955108
rect 280111 954436 280174 955108
rect 279374 952631 280174 954436
rect 280774 958993 281574 959001
rect 280774 958539 280782 958993
rect 281564 958539 281574 958993
rect 280774 953608 281574 958539
rect 280774 952936 280845 953608
rect 281517 952936 281574 953608
rect 280774 952631 281574 952936
rect 282174 958995 282974 959001
rect 282174 958541 282187 958995
rect 282969 958541 282974 958995
rect 282174 958183 282974 958541
rect 282174 957511 282251 958183
rect 282923 957511 282974 958183
rect 282174 952631 282974 957511
rect 283574 958994 284374 959001
rect 283574 958540 283583 958994
rect 284365 958540 284374 958994
rect 283574 956679 284374 958540
rect 283574 956007 283650 956679
rect 284322 956007 284374 956679
rect 283574 952631 284374 956007
rect 330974 958495 330988 959011
rect 331755 958495 331774 959011
rect 330974 955109 331774 958495
rect 330974 954437 331038 955109
rect 331710 954437 331774 955109
rect 330974 952631 331774 954437
rect 332374 959014 333174 959027
rect 332374 958498 332390 959014
rect 333157 958498 333174 959014
rect 332374 953594 333174 958498
rect 332374 952922 332434 953594
rect 333106 952922 333174 953594
rect 332374 952631 333174 952922
rect 333774 959008 334574 959027
rect 333774 958492 333791 959008
rect 334558 958492 334574 959008
rect 333774 958208 334574 958492
rect 333774 957536 333842 958208
rect 334514 957536 334574 958208
rect 333774 952631 334574 957536
rect 335174 959012 335974 959027
rect 335174 958496 335195 959012
rect 335962 958496 335974 959012
rect 474174 958993 474974 959003
rect 335174 956697 335974 958496
rect 335174 956025 335231 956697
rect 335903 956025 335974 956697
rect 335174 952631 335974 956025
rect 396974 958982 397774 958993
rect 396974 958530 396986 958982
rect 397765 958530 397774 958982
rect 396974 955110 397774 958530
rect 396974 954438 397037 955110
rect 397709 954438 397774 955110
rect 396974 952631 397774 954438
rect 398374 958980 399174 958993
rect 398374 958528 398383 958980
rect 399162 958528 399174 958980
rect 398374 953600 399174 958528
rect 398374 952928 398454 953600
rect 399126 952928 399174 953600
rect 398374 952631 399174 952928
rect 399774 958980 400574 958993
rect 399774 958528 399783 958980
rect 400562 958528 400574 958980
rect 399774 958180 400574 958528
rect 399774 957508 399823 958180
rect 400495 957508 400574 958180
rect 399774 952631 400574 957508
rect 401174 958982 401974 958993
rect 401174 958530 401186 958982
rect 401965 958530 401974 958982
rect 401174 956698 401974 958530
rect 401174 956026 401248 956698
rect 401920 956026 401974 956698
rect 401174 952631 401974 956026
rect 474174 958538 474185 958993
rect 474965 958538 474974 958993
rect 474174 955118 474974 958538
rect 474174 954446 474244 955118
rect 474916 954446 474974 955118
rect 474174 952631 474974 954446
rect 475574 958992 476374 959003
rect 475574 958537 475583 958992
rect 476363 958537 476374 958992
rect 475574 953592 476374 958537
rect 475574 952920 475644 953592
rect 476316 952920 476374 953592
rect 475574 952631 476374 952920
rect 476974 958995 477774 959003
rect 476974 958540 476985 958995
rect 477765 958540 477774 958995
rect 476974 958188 477774 958540
rect 476974 957516 477030 958188
rect 477702 957516 477774 958188
rect 476974 952631 477774 957516
rect 478374 958994 479174 959003
rect 478374 958539 478383 958994
rect 479163 958539 479174 958994
rect 478374 956690 479174 958539
rect 478374 956018 478446 956690
rect 479118 956018 479174 956690
rect 478374 952631 479174 956018
rect 525374 958959 526174 958973
rect 525374 958542 525385 958959
rect 526166 958542 526174 958959
rect 525374 955114 526174 958542
rect 525374 954442 525432 955114
rect 526104 954442 526174 955114
rect 525374 952631 526174 954442
rect 526774 958961 527574 958973
rect 526774 958544 526784 958961
rect 527565 958544 527574 958961
rect 526774 953596 527574 958544
rect 526774 952924 526844 953596
rect 527516 952924 527574 953596
rect 526774 952631 527574 952924
rect 528174 958959 528974 958973
rect 528174 958542 528183 958959
rect 528964 958542 528974 958959
rect 528174 958196 528974 958542
rect 528174 957524 528241 958196
rect 528913 957524 528974 958196
rect 528174 952631 528974 957524
rect 529574 958959 530374 958973
rect 529574 958542 529585 958959
rect 530366 958542 530374 958959
rect 529574 956682 530374 958542
rect 529574 956010 529646 956682
rect 530318 956010 530374 956682
rect 529574 952631 530374 956010
rect 537142 958512 541910 958586
rect 537142 956126 537238 958512
rect 541806 956126 541910 958512
rect 537142 955220 541910 956126
rect 533449 954543 535856 954607
rect 533449 953869 533513 954543
rect 535792 953869 535856 954543
rect 533449 953805 535856 953869
rect 533449 952967 535873 953031
rect 533449 952297 533513 952967
rect 535809 952297 535873 952967
rect 537142 952456 537238 955220
rect 541828 952456 541910 955220
rect 537142 952337 541910 952456
rect 547106 958490 551874 958572
rect 547106 956126 547188 958490
rect 551756 956126 551874 958490
rect 547106 955205 551874 956126
rect 547106 952441 547180 955205
rect 551770 952441 551874 955205
rect 625896 954559 627525 954835
rect 625896 953873 625956 954559
rect 627463 953873 627525 954559
rect 622767 953044 624396 953061
rect 547106 952323 551874 952441
rect 622761 952980 624396 953044
rect 533449 952233 535873 952297
rect 622761 952296 622825 952980
rect 624330 952296 624396 952980
rect 622761 952232 624396 952296
rect 622767 944801 624396 952232
rect 622767 943225 622828 944801
rect 624321 943225 624396 944801
rect 625896 945737 627525 953873
rect 625896 943324 625971 945737
rect 627460 943324 627525 945737
rect 625896 943242 627525 943324
rect 622767 943148 624396 943225
rect -32550 910656 -32230 912124
rect -31890 912056 -31570 912124
rect -31892 912054 -31568 912056
rect -31892 911254 -31890 912054
rect -31570 911254 -31568 912054
rect -31892 911252 -31568 911254
rect 13269 911987 17269 912051
rect 13269 911315 13333 911987
rect 17205 911315 17269 911987
rect -32552 910654 -32228 910656
rect -32552 909854 -32550 910654
rect -32230 909854 -32228 910654
rect -32552 909852 -32228 909854
rect -32550 905848 -32230 909852
rect -31890 905124 -31570 911252
rect 13269 911251 17269 911315
rect 8270 910585 12270 910649
rect 8270 909913 8334 910585
rect 12206 909913 12270 910585
rect 8270 909849 12270 909913
rect -31230 907754 -30910 909263
rect -30570 909154 -30250 909273
rect -30572 909152 -30248 909154
rect -30572 908352 -30570 909152
rect -30250 908352 -30248 909152
rect -30572 908350 -30248 908352
rect 2811 909069 3611 909133
rect 2811 908397 2875 909069
rect 3547 908397 3611 909069
rect -31232 907752 -30908 907754
rect -31232 906952 -31230 907752
rect -30910 906952 -30908 907752
rect -31232 906950 -30908 906952
rect -31230 904562 -30910 906950
rect -30570 903892 -30250 908350
rect 2811 908333 3611 908397
rect 625660 908835 629660 908899
rect 625660 908163 625724 908835
rect 629596 908163 629660 908835
rect 625660 908099 629660 908163
rect 1626 907680 2426 907744
rect 1626 907008 1690 907680
rect 2362 907008 2426 907680
rect 1626 906944 2426 907008
rect 620651 907447 624651 907511
rect 620651 906775 620715 907447
rect 624587 906775 624651 907447
rect 620651 906711 624651 906775
rect 636468 906033 637268 906097
rect 636468 905361 636532 906033
rect 637204 905361 637268 906033
rect 636468 905297 637268 905361
rect 670962 904708 671282 909088
rect 671622 906108 671942 909039
rect 672282 907508 672602 908999
rect 672942 908908 673262 909019
rect 672940 908906 673262 908908
rect 672940 908106 672942 908906
rect 673252 908106 673262 908906
rect 672940 908104 673262 908106
rect 672280 907506 672604 907508
rect 672280 906706 672282 907506
rect 672602 906706 672604 907506
rect 672280 906704 672604 906706
rect 671620 906106 671944 906108
rect 671620 905306 671622 906106
rect 671942 905306 671944 906106
rect 671620 905304 671944 905306
rect 637868 904643 638668 904707
rect 637868 903971 637932 904643
rect 638604 903971 638668 904643
rect 637868 903907 638668 903971
rect 670960 904706 671282 904708
rect 670960 903906 670962 904706
rect 671261 903906 671282 904706
rect 670960 903904 671282 903906
rect 670962 900216 671282 903904
rect 671622 900907 671942 905304
rect 672282 901598 672602 906704
rect 672942 902258 673262 908104
rect 1648 888076 17286 888256
rect 1648 883570 1793 888076
rect 17130 883570 17286 888076
rect 1648 883473 17286 883570
rect 620660 883639 638402 883817
rect 620660 879190 620797 883639
rect 638082 879190 638402 883639
rect 620660 879028 638402 879190
rect 1612 878028 17250 878185
rect 1612 873522 1744 878028
rect 17081 878016 17250 878028
rect 17165 873619 17250 878016
rect 17081 873522 17250 873619
rect 1612 873402 17250 873522
rect 620598 873616 638332 873741
rect 620598 869167 620810 873616
rect 638095 869167 638332 873616
rect 620598 868952 638332 869167
rect 4270 803652 5272 803759
rect 4270 799066 4359 803652
rect 5171 799066 5272 803652
rect 4270 798985 5272 799066
rect 633661 794462 635232 794563
rect 4269 793675 5271 793760
rect 4269 789089 4351 793675
rect 5163 789089 5271 793675
rect 633661 789897 633781 794462
rect 635118 789897 635232 794462
rect 633661 789817 635232 789897
rect 4269 788986 5271 789089
rect 633673 784517 635244 784599
rect -31230 781754 -30910 783212
rect -30570 783154 -30250 783192
rect -30572 783152 -30248 783154
rect -30572 782352 -30570 783152
rect -30250 782352 -30248 783152
rect -30572 782350 -30248 782352
rect 2817 783067 3617 783131
rect 2817 782395 2881 783067
rect 3553 782395 3617 783067
rect -31232 781752 -30908 781754
rect -31232 780952 -31230 781752
rect -30910 780952 -30908 781752
rect -31232 780950 -30908 780952
rect -31230 778738 -30910 780950
rect -30570 778078 -30250 782350
rect 2817 782331 3617 782395
rect 1637 781706 2437 781770
rect 1637 781034 1701 781706
rect 2373 781034 2437 781706
rect 1637 780970 2437 781034
rect 633673 779952 633749 784517
rect 635086 779952 635244 784517
rect 633673 779853 635244 779952
rect -32550 764302 -32230 767013
rect -31890 765702 -31570 767609
rect -31892 765700 -31568 765702
rect -31892 764900 -31890 765700
rect -31570 764900 -31568 765700
rect 13265 765636 17265 765700
rect 13265 764964 13329 765636
rect 17201 764964 17265 765636
rect 13265 764900 17265 764964
rect -31892 764898 -31568 764900
rect -32552 764300 -32228 764302
rect -32552 763500 -32550 764300
rect -32230 763500 -32228 764300
rect -32552 763498 -32228 763500
rect -32550 763464 -32230 763498
rect -31890 763406 -31570 764898
rect 8270 764241 12270 764305
rect 8270 763569 8334 764241
rect 12206 763569 12270 764241
rect 8270 763505 12270 763569
rect -31230 738554 -30910 740010
rect -30570 739954 -30250 740068
rect -30572 739952 -30248 739954
rect -30572 739152 -30570 739952
rect -30250 739152 -30248 739952
rect -30572 739150 -30248 739152
rect 2822 739880 3622 739944
rect 2822 739208 2886 739880
rect 3558 739208 3622 739880
rect -31232 738552 -30908 738554
rect -31232 737752 -31230 738552
rect -30910 737752 -30908 738552
rect -31232 737750 -30908 737752
rect -31230 735508 -30910 737750
rect -30570 734878 -30250 739150
rect 2822 739144 3622 739208
rect 1626 738497 2426 738561
rect 1626 737825 1690 738497
rect 2362 737825 2426 738497
rect 1626 737761 2426 737825
rect 625655 730844 629655 730908
rect 625655 730172 625719 730844
rect 629591 730172 629655 730844
rect 625655 730108 629655 730172
rect 620656 729441 624656 729505
rect 620656 728769 620720 729441
rect 624592 728769 624656 729441
rect 620656 728705 624656 728769
rect 636461 728033 637261 728097
rect 636461 727361 636525 728033
rect 637197 727361 637261 728033
rect 636461 727297 637261 727361
rect 637862 726647 638662 726711
rect 670962 726708 671282 731017
rect 671622 728108 671942 731007
rect 672282 729508 672602 730978
rect 672942 730908 673262 730978
rect 672940 730906 673262 730908
rect 672940 730106 672942 730906
rect 673252 730106 673262 730906
rect 672940 730104 673262 730106
rect 672280 729506 672604 729508
rect 672280 728706 672282 729506
rect 672602 728706 672604 729506
rect 672280 728704 672604 728706
rect 671620 728106 671944 728108
rect 671620 727306 671622 728106
rect 671942 727306 671944 728106
rect 671620 727304 671944 727306
rect 637862 725975 637926 726647
rect 638598 725975 638662 726647
rect 637862 725911 638662 725975
rect 670960 726706 671284 726708
rect 670960 725906 670962 726706
rect 671282 725906 671284 726706
rect 670960 725904 671284 725906
rect -32550 720902 -32230 723726
rect -31890 722302 -31570 724427
rect -31892 722300 -31568 722302
rect -31892 721500 -31890 722300
rect -31570 721500 -31568 722300
rect 13273 722236 17273 722300
rect 13273 721564 13337 722236
rect 17209 721564 17273 722236
rect 670962 721878 671282 725904
rect 671622 722538 671942 727304
rect 672282 723198 672602 728704
rect 672942 723804 673262 730104
rect 13273 721500 17273 721564
rect -31892 721498 -31568 721500
rect -32552 720900 -32228 720902
rect -32552 720100 -32550 720900
rect -32230 720100 -32228 720900
rect -32552 720098 -32228 720100
rect -32550 719964 -32230 720098
rect -31890 719974 -31570 721498
rect 8266 720830 12266 720894
rect 8266 720158 8330 720830
rect 12202 720158 12266 720830
rect 8266 720094 12266 720158
rect -31230 695354 -30910 696847
rect -30570 696754 -30250 696905
rect -30572 696752 -30248 696754
rect -30572 695952 -30570 696752
rect -30250 695952 -30248 696752
rect 2828 696699 3628 696763
rect 2828 696027 2892 696699
rect 3564 696027 3628 696699
rect 2828 695963 3628 696027
rect -30572 695950 -30248 695952
rect -31232 695352 -30908 695354
rect -31232 694552 -31230 695352
rect -30910 694552 -30908 695352
rect -31232 694550 -30908 694552
rect -31230 692335 -30910 694550
rect -30570 691678 -30250 695950
rect 1631 695294 2431 695358
rect 1631 694622 1695 695294
rect 2367 694622 2431 695294
rect 1631 694558 2431 694622
rect 625650 685641 629650 685705
rect 625650 684969 625714 685641
rect 629586 684969 629650 685641
rect 625650 684905 629650 684969
rect 620656 684229 624656 684293
rect 620656 683557 620720 684229
rect 624592 683557 624656 684229
rect 620656 683493 624656 683557
rect 636466 682843 637266 682907
rect 636466 682171 636530 682843
rect 637202 682171 637266 682843
rect 636466 682107 637266 682171
rect 670962 681508 671282 685796
rect 671622 682908 671942 685825
rect 672282 684308 672602 685845
rect 672942 685708 673262 685865
rect 672940 685706 673262 685708
rect 672940 684906 672942 685706
rect 673252 684906 673262 685706
rect 672940 684904 673262 684906
rect 672280 684306 672604 684308
rect 672280 683506 672282 684306
rect 672602 683506 672604 684306
rect 672280 683504 672604 683506
rect 671620 682906 671944 682908
rect 671620 682106 671622 682906
rect 671942 682106 671944 682906
rect 671620 682104 671944 682106
rect 670960 681506 671284 681508
rect 637867 681433 638667 681497
rect -32550 677702 -32230 680526
rect -31890 679262 -31570 681186
rect 637867 680761 637931 681433
rect 638603 680761 638667 681433
rect 637867 680697 638667 680761
rect 670960 680706 670962 681506
rect 671282 680706 671284 681506
rect 670960 680704 671284 680706
rect -31892 679260 -31568 679262
rect -31892 678460 -31890 679260
rect -31570 678460 -31568 679260
rect -31892 678458 -31568 678460
rect 13284 679189 17284 679253
rect 13284 678517 13348 679189
rect 17220 678517 17284 679189
rect -32552 677700 -32228 677702
rect -32552 676900 -32550 677700
rect -32230 676900 -32228 677700
rect -32552 676898 -32228 676900
rect -32550 676840 -32230 676898
rect -31890 676821 -31570 678458
rect 13284 678453 17284 678517
rect 8270 677639 12270 677703
rect 8270 676967 8334 677639
rect 12206 676967 12270 677639
rect 8270 676903 12270 676967
rect 670962 676878 671282 680704
rect 671622 677476 671942 682104
rect 672282 678009 672602 683504
rect 672942 678760 673262 684904
rect -31230 652154 -30910 653644
rect -30570 653554 -30250 653635
rect -30572 653552 -30248 653554
rect -30572 652752 -30570 653552
rect -30250 652752 -30248 653552
rect 2822 653496 3622 653560
rect 2822 652824 2886 653496
rect 3558 652824 3622 653496
rect 2822 652760 3622 652824
rect -30572 652750 -30248 652752
rect -31232 652152 -30908 652154
rect -31232 651352 -31230 652152
rect -30910 651352 -30908 652152
rect -31232 651350 -30908 651352
rect -31230 649138 -30910 651350
rect -30570 648478 -30250 652750
rect 1620 652074 2420 652138
rect 1620 651402 1684 652074
rect 2356 651402 2420 652074
rect 1620 651338 2420 651402
rect 625660 640439 629660 640503
rect 625660 639767 625724 640439
rect 629596 639767 629660 640439
rect 625660 639703 629660 639767
rect 620661 639046 624661 639110
rect 620661 638374 620725 639046
rect 624597 638374 624661 639046
rect 620661 638310 624661 638374
rect -32550 634902 -32230 637326
rect -31890 636302 -31570 637986
rect 636478 637635 637278 637699
rect 636478 636963 636542 637635
rect 637214 636963 637278 637635
rect 636478 636899 637278 636963
rect 670962 636308 671282 640604
rect 671622 637708 671942 640624
rect 672282 639108 672602 640584
rect 672942 640508 673262 640584
rect 672940 640506 673262 640508
rect 672940 639706 672942 640506
rect 673252 639706 673262 640506
rect 672940 639704 673262 639706
rect 672280 639106 672604 639108
rect 672280 638306 672282 639106
rect 672602 638306 672604 639106
rect 672280 638304 672604 638306
rect 671620 637706 671944 637708
rect 671620 636906 671622 637706
rect 671942 636906 671944 637706
rect 671620 636904 671944 636906
rect 670960 636306 671284 636308
rect -31892 636300 -31568 636302
rect -31892 635500 -31890 636300
rect -31570 635500 -31568 636300
rect -31892 635498 -31568 635500
rect 13273 636226 17273 636290
rect 13273 635554 13337 636226
rect 17209 635554 17273 636226
rect -32552 634900 -32228 634902
rect -32552 634100 -32550 634900
rect -32230 634100 -32228 634900
rect -32552 634098 -32228 634100
rect -32550 634009 -32230 634098
rect -31890 633970 -31570 635498
rect 13273 635490 17273 635554
rect 637857 636237 638657 636301
rect 637857 635565 637921 636237
rect 638593 635565 638657 636237
rect 637857 635501 638657 635565
rect 670960 635506 670962 636306
rect 671282 635506 671284 636306
rect 670960 635504 671284 635506
rect 8278 634839 12278 634903
rect 8278 634167 8342 634839
rect 12214 634167 12278 634839
rect 8278 634103 12278 634167
rect 670962 631613 671282 635504
rect 671622 632176 671942 636904
rect 672282 632946 672602 638304
rect 672942 633647 673262 639704
rect -31230 608954 -30910 610452
rect -30570 610354 -30250 610511
rect -30572 610352 -30248 610354
rect -30572 609552 -30570 610352
rect -30250 609552 -30248 610352
rect 2839 610292 3639 610356
rect 2839 609620 2903 610292
rect 3575 609620 3639 610292
rect 2839 609556 3639 609620
rect -30572 609550 -30248 609552
rect -31232 608952 -30908 608954
rect -31232 608152 -31230 608952
rect -30910 608152 -30908 608952
rect -31232 608150 -30908 608152
rect -31230 605938 -30910 608150
rect -30570 605278 -30250 609550
rect 1626 608921 2426 608985
rect 1626 608249 1690 608921
rect 2362 608249 2426 608921
rect 1626 608185 2426 608249
rect 625664 595246 629664 595310
rect -32550 591302 -32230 594126
rect -31890 592702 -31570 594859
rect 625664 594574 625728 595246
rect 629600 594574 629664 595246
rect 625664 594510 629664 594574
rect 620651 593843 624651 593907
rect 620651 593171 620715 593843
rect 624587 593171 624651 593843
rect 620651 593107 624651 593171
rect -31892 592700 -31568 592702
rect -31892 591900 -31890 592700
rect -31570 591900 -31568 592700
rect 13276 592638 17276 592702
rect 13276 591966 13340 592638
rect 17212 591966 17276 592638
rect 13276 591902 17276 591966
rect 636468 592442 637268 592506
rect -31892 591898 -31568 591900
rect -32552 591300 -32228 591302
rect -32552 590500 -32550 591300
rect -32230 590500 -32228 591300
rect -32552 590498 -32228 590500
rect -32550 590377 -32230 590498
rect -31890 590387 -31570 591898
rect 636468 591770 636532 592442
rect 637204 591770 637268 592442
rect 636468 591706 637268 591770
rect 8266 591232 12266 591296
rect 8266 590560 8330 591232
rect 12202 590560 12266 591232
rect 670962 591108 671282 595392
rect 671622 592508 671942 595461
rect 672282 593908 672602 595461
rect 672942 595308 673262 595412
rect 672940 595306 673262 595308
rect 672940 594506 672942 595306
rect 673252 594506 673262 595306
rect 672940 594504 673262 594506
rect 672280 593906 672604 593908
rect 672280 593106 672282 593906
rect 672602 593106 672604 593906
rect 672280 593104 672604 593106
rect 671620 592506 671944 592508
rect 671620 591706 671622 592506
rect 671942 591706 671944 592506
rect 671620 591704 671944 591706
rect 670960 591106 671284 591108
rect 8266 590496 12266 590560
rect 637862 591039 638662 591103
rect 637862 590367 637926 591039
rect 638598 590367 638662 591039
rect 637862 590303 638662 590367
rect 670960 590306 670962 591106
rect 671282 590306 671284 591106
rect 670960 590304 671284 590306
rect 670962 586678 671282 590304
rect 671622 587191 671942 591704
rect 672282 587922 672602 593104
rect 672942 588505 673262 594504
rect -31230 565954 -30910 567455
rect -30570 567354 -30250 567455
rect -30572 567352 -30248 567354
rect -30572 566552 -30570 567352
rect -30250 566552 -30248 567352
rect 2833 567309 3633 567373
rect 2833 566637 2897 567309
rect 3569 566637 3633 567309
rect 2833 566573 3633 566637
rect -30572 566550 -30248 566552
rect -31232 565952 -30908 565954
rect -31232 565152 -31230 565952
rect -30910 565152 -30908 565952
rect -31232 565150 -30908 565152
rect -31230 562738 -30910 565150
rect -30570 562074 -30250 566550
rect 1620 565887 2420 565951
rect 1620 565215 1684 565887
rect 2356 565215 2420 565887
rect 1620 565151 2420 565215
rect -32550 548102 -32230 550926
rect -31890 549502 -31570 551586
rect 625664 550038 629664 550102
rect -31892 549500 -31568 549502
rect -31892 548700 -31890 549500
rect -31570 548700 -31568 549500
rect 13277 549436 17277 549500
rect 13277 548764 13341 549436
rect 17213 548764 17277 549436
rect 625664 549366 625728 550038
rect 629600 549366 629664 550038
rect 625664 549302 629664 549366
rect 13277 548700 17277 548764
rect -31892 548698 -31568 548700
rect -32552 548100 -32228 548102
rect -32552 547300 -32550 548100
rect -32230 547300 -32228 548100
rect -32552 547298 -32228 547300
rect -32550 547185 -32230 547298
rect -31890 547234 -31570 548698
rect 620661 548645 624661 548709
rect 8266 548047 12266 548111
rect 8266 547375 8330 548047
rect 12202 547375 12266 548047
rect 620661 547973 620725 548645
rect 624597 547973 624661 548645
rect 620661 547909 624661 547973
rect 8266 547311 12266 547375
rect 636459 547239 637259 547303
rect 636459 546567 636523 547239
rect 637195 546567 637259 547239
rect 636459 546503 637259 546567
rect 637871 545845 638671 545909
rect 670962 545908 671282 550161
rect 671622 547308 671942 550181
rect 672282 548708 672602 550200
rect 672942 550108 673262 550220
rect 672940 550106 673262 550108
rect 672940 549306 672942 550106
rect 673252 549306 673262 550106
rect 672940 549304 673262 549306
rect 672280 548706 672604 548708
rect 672280 547906 672282 548706
rect 672602 547906 672604 548706
rect 672280 547904 672604 547906
rect 671620 547306 671944 547308
rect 671620 546506 671622 547306
rect 671942 546506 671944 547306
rect 671620 546504 671944 546506
rect 637871 545173 637935 545845
rect 638607 545173 638671 545845
rect 637871 545109 638671 545173
rect 670960 545906 671284 545908
rect 670960 545106 670962 545906
rect 671282 545106 671284 545906
rect 670960 545104 671284 545106
rect 670962 541367 671282 545104
rect 671622 542138 671942 546504
rect 672282 542711 672602 547904
rect 672942 543353 673262 549304
rect -31230 522954 -30910 524450
rect -30570 524354 -30250 524460
rect -30572 524352 -30248 524354
rect -30572 523552 -30570 524352
rect -30250 523552 -30248 524352
rect -30572 523550 -30248 523552
rect 2839 524275 3639 524339
rect 2839 523603 2903 524275
rect 3575 523603 3639 524275
rect -31232 522952 -30908 522954
rect -31232 522152 -31230 522952
rect -30910 522152 -30908 522952
rect -31232 522150 -30908 522152
rect -31230 519538 -30910 522150
rect -30570 518878 -30250 523550
rect 2839 523539 3639 523603
rect 1609 522887 2409 522951
rect 1609 522215 1673 522887
rect 2345 522215 2409 522887
rect 1609 522151 2409 522215
rect -32550 504902 -32230 507755
rect -31890 506302 -31570 508436
rect -31892 506300 -31568 506302
rect -31892 505500 -31890 506300
rect -31570 505500 -31568 506300
rect 13273 506240 17273 506304
rect 13273 505568 13337 506240
rect 17209 505568 17273 506240
rect 13273 505504 17273 505568
rect -31892 505498 -31568 505500
rect -32552 504900 -32228 504902
rect -32552 504100 -32550 504900
rect -32230 504100 -32228 504900
rect -32552 504098 -32228 504100
rect -32550 503986 -32230 504098
rect -31890 503957 -31570 505498
rect 8259 504838 12259 504902
rect 8259 504166 8323 504838
rect 12195 504166 12259 504838
rect 8259 504102 12259 504166
rect 625650 504840 629650 504904
rect 625650 504168 625714 504840
rect 629586 504168 629650 504840
rect 625650 504104 629650 504168
rect 620665 503437 624665 503501
rect 620665 502765 620729 503437
rect 624601 502765 624665 503437
rect 620665 502701 624665 502765
rect 636465 502043 637265 502107
rect 636465 501371 636529 502043
rect 637201 501371 637265 502043
rect 636465 501307 637265 501371
rect 637866 500647 638666 500711
rect 670962 500708 671282 505048
rect 671622 502108 671942 504999
rect 672282 503508 672602 504979
rect 672942 504908 673262 504949
rect 672940 504906 673262 504908
rect 672940 504106 672942 504906
rect 673252 504106 673262 504906
rect 672940 504104 673262 504106
rect 672280 503506 672604 503508
rect 672280 502706 672282 503506
rect 672602 502706 672604 503506
rect 672280 502704 672604 502706
rect 671620 502106 671944 502108
rect 671620 501306 671622 502106
rect 671942 501306 671944 502106
rect 671620 501304 671944 501306
rect 637866 499975 637930 500647
rect 638602 499975 638666 500647
rect 637866 499911 638666 499975
rect 670960 500706 671284 500708
rect 670960 499906 670962 500706
rect 671282 499906 671284 500706
rect 670960 499904 671284 499906
rect 670962 496478 671282 499904
rect 671622 497084 671942 501304
rect 672282 497798 672602 502704
rect 672942 498418 673262 504104
rect 630652 479910 632660 479992
rect 630652 475283 630713 479910
rect 632588 475283 632660 479910
rect 630652 475222 632660 475283
rect 630648 469932 632656 470000
rect 630648 465305 630706 469932
rect 632581 465305 632656 469932
rect 630648 465230 632656 465305
rect 625655 461238 629655 461302
rect 625655 460566 625719 461238
rect 629591 460566 629655 461238
rect 625655 460502 629655 460566
rect 620651 459845 624651 459909
rect 6245 459103 7322 459189
rect 620651 459173 620715 459845
rect 624587 459173 624651 459845
rect 620651 459109 624651 459173
rect 6245 454442 6326 459103
rect 7225 454442 7322 459103
rect 636466 458440 637266 458504
rect 636466 457768 636530 458440
rect 637202 457768 637266 458440
rect 636466 457704 637266 457768
rect 670962 457108 671282 461427
rect 671622 458508 671942 461387
rect 672282 459908 672602 461466
rect 672942 461308 673262 461456
rect 672940 461306 673262 461308
rect 672940 460506 672942 461306
rect 673252 460506 673262 461306
rect 672940 460504 673262 460506
rect 672280 459906 672604 459908
rect 672280 459106 672282 459906
rect 672602 459106 672604 459906
rect 672280 459104 672604 459106
rect 671620 458506 671944 458508
rect 671620 457706 671622 458506
rect 671942 457706 671944 458506
rect 671620 457704 671944 457706
rect 670960 457106 671284 457108
rect 637864 457041 638664 457105
rect 637864 456369 637928 457041
rect 638600 456369 638664 457041
rect 637864 456305 638664 456369
rect 670960 456306 670962 457106
rect 671282 456306 671284 457106
rect 670960 456304 671284 456306
rect 6245 454364 7322 454442
rect 670962 452478 671282 456304
rect 671622 453087 671942 457704
rect 672282 453739 672602 459104
rect 672942 454458 673262 460504
rect 6220 449139 7297 449200
rect 6220 444435 6315 449139
rect 7201 444435 7297 449139
rect 6220 444375 7297 444435
rect 625608 435866 638675 435998
rect 625608 431326 625815 435866
rect 629491 435779 638675 435866
rect 638381 431386 638675 435779
rect 629491 431326 638675 431386
rect 625608 431192 638675 431326
rect 625608 425749 638807 425935
rect 625608 421357 625811 425749
rect 638601 421357 638807 425749
rect 625608 421152 638807 421357
rect 5551 416912 12278 417071
rect 5551 416868 8417 416912
rect 5551 412396 5639 416868
rect 12175 412440 12278 416912
rect 12132 412396 12278 412440
rect 5551 412250 12278 412396
rect 5551 406832 12278 407006
rect 5551 402360 5697 406832
rect 12190 402360 12278 406832
rect 5551 402185 12278 402360
rect -31230 394954 -30910 396456
rect -30570 396354 -30250 396437
rect -30572 396352 -30248 396354
rect -30572 395552 -30570 396352
rect -30250 395552 -30248 396352
rect -30572 395550 -30248 395552
rect 2839 396279 3639 396343
rect 2839 395607 2903 396279
rect 3575 395607 3639 396279
rect -31232 394952 -30908 394954
rect -31232 394152 -31230 394952
rect -30910 394152 -30908 394952
rect -31232 394150 -30908 394152
rect -31230 391915 -30910 394150
rect -30570 391278 -30250 395550
rect 2839 395543 3639 395607
rect 1626 394896 2426 394960
rect 1626 394224 1690 394896
rect 2362 394224 2426 394896
rect 1626 394160 2426 394224
rect 633661 391672 635651 391772
rect 633661 387094 633737 391672
rect 635564 387094 635651 391672
rect 633661 386987 635651 387094
rect 633639 381734 635651 381821
rect -32550 377099 -32230 380174
rect -31890 378499 -31570 380786
rect -31892 378497 -31568 378499
rect -31892 377697 -31890 378497
rect -31570 377697 -31568 378497
rect -31892 377695 -31568 377697
rect 13265 378423 17265 378487
rect 13265 377751 13329 378423
rect 17201 377751 17265 378423
rect -32552 377097 -32228 377099
rect -32552 376297 -32550 377097
rect -32230 376297 -32228 377097
rect -32552 376295 -32228 376297
rect -32550 376137 -32230 376295
rect -31890 376098 -31570 377695
rect 13265 377687 17265 377751
rect 633639 377156 633726 381734
rect 635553 377156 635651 381734
rect 8270 377036 12270 377100
rect 633639 377052 635651 377156
rect 8270 376364 8334 377036
rect 12206 376364 12270 377036
rect 8270 376300 12270 376364
rect 625660 372852 629660 372916
rect 625660 372180 625724 372852
rect 629596 372180 629660 372852
rect 625660 372116 629660 372180
rect 620656 371449 624656 371513
rect 620656 370777 620720 371449
rect 624592 370777 624656 371449
rect 620656 370713 624656 370777
rect 636465 370039 637265 370103
rect 636465 369367 636529 370039
rect 637201 369367 637265 370039
rect 636465 369303 637265 369367
rect 670962 368708 671282 373048
rect 671622 370108 671942 373068
rect 672282 371508 672602 373008
rect 672942 372908 673262 373018
rect 672940 372906 673262 372908
rect 672940 372106 672942 372906
rect 673252 372106 673262 372906
rect 672940 372104 673262 372106
rect 672280 371506 672604 371508
rect 672280 370706 672282 371506
rect 672602 370706 672604 371506
rect 672280 370704 672604 370706
rect 671620 370106 671944 370108
rect 671620 369306 671622 370106
rect 671942 369306 671944 370106
rect 671620 369304 671944 369306
rect 670960 368706 671284 368708
rect 637865 368635 638665 368699
rect 637865 367963 637929 368635
rect 638601 367963 638665 368635
rect 637865 367899 638665 367963
rect 670960 367906 670962 368706
rect 671282 367906 671284 368706
rect 670960 367904 671284 367906
rect 670962 364156 671282 367904
rect 671622 364896 671942 369304
rect 672282 365598 672602 370704
rect 672942 366258 673262 372104
rect -31230 351954 -30910 353417
rect -30570 353354 -30250 353475
rect -30572 353352 -30248 353354
rect -30572 352552 -30570 353352
rect -30250 352552 -30248 353352
rect 2822 353296 3622 353360
rect 2822 352624 2886 353296
rect 3558 352624 3622 353296
rect 2822 352560 3622 352624
rect -30572 352550 -30248 352552
rect -31232 351952 -30908 351954
rect -31232 351152 -31230 351952
rect -30910 351152 -30908 351952
rect -31232 351150 -30908 351152
rect -31230 348722 -30910 351150
rect -30570 348044 -30250 352550
rect 1620 351879 2420 351943
rect 1620 351207 1684 351879
rect 2356 351207 2420 351879
rect 1620 351143 2420 351207
rect -32550 333899 -32230 337019
rect -31890 335299 -31570 337696
rect -31892 335297 -31568 335299
rect -31892 334497 -31890 335297
rect -31570 334497 -31568 335297
rect -31892 334495 -31568 334497
rect 13265 335232 17265 335296
rect 13265 334560 13329 335232
rect 17201 334560 17265 335232
rect 13265 334496 17265 334560
rect -32552 333897 -32228 333899
rect -32552 333097 -32550 333897
rect -32230 333097 -32228 333897
rect -32552 333095 -32228 333097
rect -32550 332943 -32230 333095
rect -31890 332865 -31570 334495
rect 8278 333829 12278 333893
rect 8278 333157 8342 333829
rect 12214 333157 12278 333829
rect 8278 333093 12278 333157
rect 625660 328050 629660 328114
rect 625660 327378 625724 328050
rect 629596 327378 629660 328050
rect 625660 327314 629660 327378
rect 620665 326666 624665 326730
rect 620665 325994 620729 326666
rect 624601 325994 624665 326666
rect 620665 325930 624665 325994
rect 636465 325237 637265 325301
rect 636465 324565 636529 325237
rect 637201 324565 637265 325237
rect 636465 324501 637265 324565
rect 637860 323860 638660 323924
rect 670962 323908 671282 328202
rect 671622 325308 671942 328202
rect 672282 326708 672602 328271
rect 672942 328108 673262 328192
rect 672940 328106 673262 328108
rect 672940 327306 672942 328106
rect 673252 327306 673262 328106
rect 672940 327304 673262 327306
rect 672280 326706 672604 326708
rect 672280 325906 672282 326706
rect 672602 325906 672604 326706
rect 672280 325904 672604 325906
rect 671620 325306 671944 325308
rect 671620 324506 671622 325306
rect 671942 324506 671944 325306
rect 671620 324504 671944 324506
rect 637860 323188 637924 323860
rect 638596 323188 638660 323860
rect 637860 323124 638660 323188
rect 670960 323906 671284 323908
rect 670960 323106 670962 323906
rect 671282 323106 671284 323906
rect 670960 323104 671284 323106
rect 670962 319063 671282 323104
rect 671622 319738 671942 324504
rect 672282 320398 672602 325904
rect 672942 320929 673262 327304
rect -31230 308954 -30910 310437
rect -30570 310354 -30250 310514
rect -30572 310352 -30248 310354
rect -30572 309552 -30570 310352
rect -30250 309552 -30248 310352
rect 2811 310312 3611 310376
rect 2811 309640 2875 310312
rect 3547 309640 3611 310312
rect 2811 309576 3611 309640
rect -30572 309550 -30248 309552
rect -31232 308952 -30908 308954
rect -31232 308152 -31230 308952
rect -30910 308152 -30908 308952
rect -31232 308150 -30908 308152
rect -31230 305528 -30910 308150
rect -30570 304850 -30250 309550
rect 1609 308884 2409 308948
rect 1609 308212 1673 308884
rect 2345 308212 2409 308884
rect 1609 308148 2409 308212
rect -32550 290699 -32230 293728
rect -31890 292099 -31570 294386
rect -31892 292097 -31568 292099
rect -31892 291297 -31890 292097
rect -31570 291297 -31568 292097
rect -31892 291295 -31568 291297
rect 13265 292032 17265 292096
rect 13265 291360 13329 292032
rect 17201 291360 17265 292032
rect 13265 291296 17265 291360
rect -32552 290697 -32228 290699
rect -32552 289897 -32550 290697
rect -32230 289897 -32228 290697
rect -32552 289895 -32228 289897
rect -32550 289807 -32230 289895
rect -31890 289768 -31570 291295
rect 8268 290622 12268 290686
rect 8268 289950 8332 290622
rect 12204 289950 12268 290622
rect 8268 289886 12268 289950
rect 625660 283228 629660 283292
rect 625660 282556 625724 283228
rect 629596 282556 629660 283228
rect 625660 282492 629660 282556
rect 620670 281849 624670 281913
rect 620670 281177 620734 281849
rect 624606 281177 624670 281849
rect 620670 281113 624670 281177
rect 636460 280444 637260 280508
rect 636460 279772 636524 280444
rect 637196 279772 637260 280444
rect 636460 279708 637260 279772
rect 670962 279108 671282 283385
rect 671622 280508 671942 283395
rect 672282 281908 672602 283425
rect 672942 283308 673262 283435
rect 672940 283306 673262 283308
rect 672940 282506 672942 283306
rect 673252 282506 673262 283306
rect 672940 282504 673262 282506
rect 672280 281906 672604 281908
rect 672280 281106 672282 281906
rect 672602 281106 672604 281906
rect 672280 281104 672604 281106
rect 671620 280506 671944 280508
rect 671620 279706 671622 280506
rect 671942 279706 671944 280506
rect 671620 279704 671944 279706
rect 670960 279106 671284 279108
rect 637851 279039 638651 279103
rect 637851 278367 637915 279039
rect 638587 278367 638651 279039
rect 637851 278303 638651 278367
rect 670960 278306 670962 279106
rect 671282 278306 671284 279106
rect 670960 278304 671284 278306
rect 670962 274078 671282 278304
rect 671622 274738 671942 279704
rect 672282 275283 672602 281104
rect 672942 276058 673262 282504
rect -31230 265954 -30910 267456
rect -30570 267354 -30250 267514
rect -30572 267352 -30248 267354
rect -30572 266552 -30570 267352
rect -30250 266552 -30248 267352
rect 2820 267292 3620 267356
rect 2820 266620 2884 267292
rect 3556 266620 3620 267292
rect 2820 266556 3620 266620
rect -30572 266550 -30248 266552
rect -31232 265952 -30908 265954
rect -31232 265152 -31230 265952
rect -30910 265152 -30908 265952
rect -31232 265150 -30908 265152
rect -31230 262334 -30910 265150
rect -30570 261637 -30250 266550
rect 1620 265891 2420 265955
rect 1620 265219 1684 265891
rect 2356 265219 2420 265891
rect 1620 265155 2420 265219
rect -32550 247499 -32230 250747
rect -31890 248899 -31570 251290
rect -31892 248897 -31568 248899
rect -31892 248097 -31890 248897
rect -31570 248097 -31568 248897
rect -31892 248095 -31568 248097
rect 13264 248824 17264 248888
rect 13264 248152 13328 248824
rect 17200 248152 17264 248824
rect -32552 247497 -32228 247499
rect -32552 246697 -32550 247497
rect -32230 246697 -32228 247497
rect -32552 246695 -32228 246697
rect -32550 246652 -32230 246695
rect -31890 246594 -31570 248095
rect 13264 248088 17264 248152
rect 8268 247417 12268 247481
rect 8268 246745 8332 247417
rect 12204 246745 12268 247417
rect 8268 246681 12268 246745
rect 620641 242438 624668 242587
rect 8286 240968 12286 241061
rect 6237 238811 7262 238942
rect 6237 233558 6344 238811
rect 7160 233558 7262 238811
rect 6237 231502 7262 233558
rect 6237 227791 6355 231502
rect 7149 227791 7262 231502
rect 6237 227659 7262 227791
rect 8286 234855 8378 240968
rect 12145 234855 12286 240968
rect 8286 231501 12286 234855
rect 8286 227903 8423 231501
rect 12144 227903 12286 231501
rect 8286 227701 12286 227903
rect 13282 240911 17282 241061
rect 13282 237313 13396 240911
rect 17117 237313 17282 240911
rect 13282 231468 17282 237313
rect 13282 227870 13419 231468
rect 17140 227870 17282 231468
rect 620641 239279 620804 242438
rect 624519 239279 624668 242438
rect 620641 236448 624668 239279
rect 620641 235776 620702 236448
rect 624574 235776 624668 236448
rect 620641 233434 624668 235776
rect 620641 230071 620817 233434
rect 624505 230071 624668 233434
rect 620641 229841 624668 230071
rect 625658 242425 629685 242587
rect 625658 237845 625807 242425
rect 629455 237845 629685 242425
rect 625658 237173 625723 237845
rect 629595 237173 629685 237845
rect 625658 236391 625807 237173
rect 629455 236391 629685 237173
rect 625658 233407 629685 236391
rect 625658 230044 625848 233407
rect 629536 230044 629685 233407
rect 625658 229841 629685 230044
rect 630635 242425 632682 242547
rect 630635 235468 630784 242425
rect 632547 235468 632682 242425
rect 630635 233461 632682 235468
rect 636468 235036 637268 235100
rect 636468 234364 636532 235036
rect 637204 234364 637268 235036
rect 636468 234300 637268 234364
rect 630635 230058 630865 233461
rect 632506 230058 632682 233461
rect 637869 233650 638669 233714
rect 670962 233708 671282 238006
rect 671622 235108 671942 238006
rect 672282 236508 672602 237986
rect 672942 237908 673262 238045
rect 672940 237906 673262 237908
rect 672940 237106 672942 237906
rect 673252 237106 673262 237906
rect 672940 237104 673262 237106
rect 672280 236506 672604 236508
rect 672280 235706 672282 236506
rect 672602 235706 672604 236506
rect 672280 235704 672604 235706
rect 671620 235106 671944 235108
rect 671620 234306 671622 235106
rect 671942 234306 671944 235106
rect 671620 234304 671944 234306
rect 637869 232978 637933 233650
rect 638605 232978 638669 233650
rect 637869 232914 638669 232978
rect 670960 233706 671284 233708
rect 670960 232906 670962 233706
rect 671282 232906 671284 233706
rect 670960 232904 671284 232906
rect 630635 229868 632682 230058
rect 13282 227701 17282 227870
rect -31230 222954 -30910 224591
rect -30570 224354 -30250 224572
rect -30572 224352 -30248 224354
rect -30572 223552 -30570 224352
rect -30250 223552 -30248 224352
rect 2817 224294 3617 224358
rect 2817 223622 2881 224294
rect 3553 223622 3617 224294
rect 2817 223558 3617 223622
rect -30572 223550 -30248 223552
rect -31232 222952 -30908 222954
rect -31232 222152 -31230 222952
rect -30910 222152 -30908 222952
rect -31232 222150 -30908 222152
rect -31230 219063 -30910 222150
rect -30570 218478 -30250 223550
rect 1620 222893 2420 222957
rect 1620 222221 1684 222893
rect 2356 222221 2420 222893
rect 1620 222157 2420 222221
rect 8953 216654 9757 227701
rect 4228 215850 9757 216654
rect 4228 213801 5032 215850
rect 4228 211917 4272 213801
rect 4958 211917 5032 213801
rect 4228 211808 5032 211917
rect 5629 215113 6433 215119
rect 14228 215113 15032 227701
rect 159182 225528 159543 225563
rect 159182 224103 159217 225528
rect 159507 224103 159543 225528
rect 159182 224066 159543 224103
rect 189282 225528 189643 225563
rect 189282 224103 189317 225528
rect 189607 224103 189643 225528
rect 189282 224066 189643 224103
rect 219382 225528 219743 225563
rect 219382 224103 219417 225528
rect 219707 224103 219743 225528
rect 219382 224066 219743 224103
rect 249482 225528 249843 225563
rect 249482 224103 249517 225528
rect 249807 224103 249843 225528
rect 249482 224066 249843 224103
rect 279582 225528 279943 225563
rect 279582 224103 279617 225528
rect 279907 224103 279943 225528
rect 279582 224066 279943 224103
rect 309682 225528 310043 225563
rect 309682 224103 309717 225528
rect 310007 224103 310043 225528
rect 309682 224066 310043 224103
rect 339782 225528 340143 225563
rect 339782 224103 339817 225528
rect 340107 224103 340143 225528
rect 339782 224066 340143 224103
rect 369882 225528 370243 225563
rect 369882 224103 369917 225528
rect 370207 224103 370243 225528
rect 369882 224066 370243 224103
rect 174229 223017 174620 223066
rect 174229 221605 174274 223017
rect 174572 221605 174620 223017
rect 174229 221563 174620 221605
rect 204329 223017 204720 223066
rect 204329 221605 204374 223017
rect 204672 221605 204720 223017
rect 204329 221563 204720 221605
rect 234429 223017 234820 223066
rect 234429 221605 234474 223017
rect 234772 221605 234820 223017
rect 234429 221563 234820 221605
rect 264529 223017 264920 223066
rect 264529 221605 264574 223017
rect 264872 221605 264920 223017
rect 264529 221563 264920 221605
rect 294629 223017 295020 223066
rect 294629 221605 294674 223017
rect 294972 221605 295020 223017
rect 294629 221563 295020 221605
rect 324729 223017 325120 223066
rect 324729 221605 324774 223017
rect 325072 221605 325120 223017
rect 324729 221563 325120 221605
rect 354829 223017 355220 223066
rect 354829 221605 354874 223017
rect 355172 221605 355220 223017
rect 354829 221563 355220 221605
rect 159984 220516 160416 220561
rect 159984 219105 160027 220516
rect 160382 219105 160416 220516
rect 159984 219067 160416 219105
rect 190084 220516 190516 220561
rect 190084 219105 190127 220516
rect 190482 219105 190516 220516
rect 190084 219067 190516 219105
rect 220184 220516 220616 220561
rect 220184 219105 220227 220516
rect 220582 219105 220616 220516
rect 220184 219067 220616 219105
rect 250224 220516 250576 220561
rect 250224 219105 250267 220516
rect 250542 219105 250576 220516
rect 250224 219067 250576 219105
rect 280384 220516 280816 220561
rect 280384 219105 280427 220516
rect 280782 219105 280816 220516
rect 280384 219067 280816 219105
rect 310484 220516 310916 220561
rect 310484 219105 310527 220516
rect 310882 219105 310916 220516
rect 310484 219067 310916 219105
rect 340584 220516 341016 220561
rect 340584 219105 340627 220516
rect 340982 219105 341016 220516
rect 340584 219067 341016 219105
rect 370684 220516 371116 220561
rect 370684 219105 370727 220516
rect 371082 219105 371116 220516
rect 370684 219067 371116 219105
rect 175882 218030 176215 218067
rect 175882 216618 175919 218030
rect 176178 216618 176215 218030
rect 175882 216577 176215 216618
rect 205982 218030 206315 218067
rect 205982 216618 206019 218030
rect 206278 216618 206315 218030
rect 205982 216577 206315 216618
rect 236082 218030 236415 218067
rect 236082 216618 236119 218030
rect 236378 216618 236415 218030
rect 236082 216577 236415 216618
rect 266182 218030 266515 218067
rect 266182 216613 266219 218030
rect 266478 216613 266515 218030
rect 266182 216572 266515 216613
rect 296282 218030 296615 218067
rect 296282 216618 296319 218030
rect 296578 216618 296615 218030
rect 296282 216577 296615 216618
rect 326382 218030 326715 218067
rect 326382 216618 326419 218030
rect 326678 216618 326715 218030
rect 326382 216577 326715 216618
rect 356482 218030 356815 218067
rect 356482 216618 356519 218030
rect 356778 216618 356815 218030
rect 356482 216577 356815 216618
rect 5629 214309 15032 215113
rect 158364 215526 158733 215566
rect 5629 213781 6433 214309
rect 158364 214096 158407 215526
rect 158695 214096 158733 215526
rect 158364 214066 158733 214096
rect 188464 215526 188833 215566
rect 188464 214096 188507 215526
rect 188795 214096 188833 215526
rect 188464 214066 188833 214096
rect 218564 215526 218933 215566
rect 218564 214096 218607 215526
rect 218895 214096 218933 215526
rect 218564 214066 218933 214096
rect 248754 215526 249113 215566
rect 248754 214096 248797 215526
rect 249075 214096 249113 215526
rect 248754 214066 249113 214096
rect 278764 215526 279083 215566
rect 278764 214096 278807 215526
rect 279045 214096 279083 215526
rect 278764 214066 279083 214096
rect 308864 215526 309233 215566
rect 308864 214096 308907 215526
rect 309195 214096 309233 215526
rect 308864 214066 309233 214096
rect 338964 215526 339333 215566
rect 338964 214096 339007 215526
rect 339295 214096 339333 215526
rect 338964 214066 339333 214096
rect 369064 215526 369433 215566
rect 369064 214096 369107 215526
rect 369395 214096 369433 215526
rect 623095 214972 623904 229841
rect 627551 216651 628360 229841
rect 670962 229078 671282 232904
rect 671622 229738 671942 234304
rect 672282 230378 672602 235704
rect 672942 230990 673262 237104
rect 627551 215842 633959 216651
rect 623095 214163 631298 214972
rect 369064 214066 369433 214096
rect 5629 211897 5673 213781
rect 6359 211897 6433 213781
rect 5629 211828 6433 211897
rect 109921 213365 116936 213753
rect -32550 204299 -32230 207825
rect -31890 205699 -31570 208425
rect 109921 207012 110403 213365
rect 116528 207012 116936 213365
rect -31892 205697 -31568 205699
rect -31892 204897 -31890 205697
rect -31570 204897 -31568 205697
rect -31892 204895 -31568 204897
rect 5622 205628 6422 205692
rect 5622 204956 5686 205628
rect 6358 204956 6422 205628
rect -32552 204297 -32228 204299
rect -32552 203497 -32550 204297
rect -32230 203497 -32228 204297
rect -32552 203495 -32228 203497
rect -32550 203284 -32230 203495
rect -31890 203226 -31570 204895
rect 5622 204892 6422 204956
rect 4225 204225 5025 204289
rect 4225 203553 4289 204225
rect 4961 203553 5025 204225
rect 4225 203489 5025 203553
rect 109921 200162 116936 207012
rect 109921 199698 110021 200162
rect 116816 199698 116936 200162
rect 109921 197631 116936 199698
rect 109936 190162 116936 197631
rect 129936 213365 136936 213574
rect 129936 207012 130322 213365
rect 136447 207012 136936 213365
rect 173422 213029 173760 213061
rect 173422 211601 173451 213029
rect 173725 211601 173760 213029
rect 173422 211564 173760 211601
rect 203522 213029 203860 213061
rect 203522 211601 203551 213029
rect 203825 211601 203860 213029
rect 203522 211564 203860 211601
rect 233672 213029 234010 213061
rect 233672 211601 233701 213029
rect 233975 211601 234010 213029
rect 293822 213029 294160 213061
rect 233672 211564 234010 211601
rect 263662 212949 264000 212981
rect 263662 211601 263691 212949
rect 263965 211601 264000 212949
rect 263662 211564 264000 211601
rect 293822 211601 293851 213029
rect 294125 211601 294160 213029
rect 293822 211564 294160 211601
rect 323922 213029 324260 213061
rect 323922 211601 323951 213029
rect 324225 211601 324260 213029
rect 323922 211564 324260 211601
rect 354022 213029 354360 213061
rect 354022 211601 354051 213029
rect 354325 211601 354360 213029
rect 354022 211564 354360 211601
rect 160062 210533 160393 210565
rect 160062 209096 160095 210533
rect 160347 209096 160393 210533
rect 160062 209060 160393 209096
rect 190162 210533 190493 210565
rect 190162 209096 190195 210533
rect 190447 209096 190493 210533
rect 190162 209060 190493 209096
rect 220262 210533 220593 210565
rect 220262 209096 220295 210533
rect 220547 209096 220593 210533
rect 220262 209060 220593 209096
rect 250242 210533 250573 210565
rect 250242 209096 250275 210533
rect 250527 209096 250573 210533
rect 250242 209060 250573 209096
rect 280462 210533 280793 210565
rect 280462 209096 280495 210533
rect 280747 209096 280793 210533
rect 280462 209060 280793 209096
rect 310562 210533 310893 210565
rect 310562 209096 310595 210533
rect 310847 209096 310893 210533
rect 310562 209060 310893 209096
rect 340662 210533 340993 210565
rect 340662 209096 340695 210533
rect 340947 209096 340993 210533
rect 340662 209060 340993 209096
rect 370762 210533 371093 210565
rect 370762 209096 370795 210533
rect 371047 209096 371093 210533
rect 370762 209060 371093 209096
rect 109936 189698 110021 190162
rect 116816 189698 116936 190162
rect -31230 179954 -30910 181591
rect -30570 181354 -30250 181610
rect -30572 181352 -30248 181354
rect -30572 180552 -30570 181352
rect -30250 180552 -30248 181352
rect -30572 180550 -30248 180552
rect 2823 181286 3625 181350
rect 2823 180614 2887 181286
rect 3561 180614 3625 181286
rect 2823 180550 3625 180614
rect -31232 179952 -30908 179954
rect -31232 179152 -31230 179952
rect -30910 179152 -30908 179952
rect -31232 179150 -30908 179152
rect -31230 175889 -30910 179150
rect -30570 175211 -30250 180550
rect 109936 180162 116936 189698
rect 1621 179924 2423 179951
rect 1621 179188 1653 179924
rect 2388 179188 2423 179924
rect 1621 179151 2423 179188
rect 109936 179698 110021 180162
rect 116816 179698 116936 180162
rect 109936 170162 116936 179698
rect 109936 169698 110021 170162
rect 116816 169698 116936 170162
rect -32550 161099 -32230 164379
rect -31890 162499 -31570 164825
rect -31892 162497 -31568 162499
rect -31892 161697 -31890 162497
rect -31570 161697 -31568 162497
rect 5633 162450 6433 162497
rect 5633 161736 5662 162450
rect 6387 161736 6433 162450
rect 5633 161697 6433 161736
rect -31892 161695 -31568 161697
rect -32552 161097 -32228 161099
rect -32552 160297 -32550 161097
rect -32230 160297 -32228 161097
rect -32552 160295 -32228 160297
rect -32550 160168 -32230 160295
rect -31890 160110 -31570 161695
rect 4217 161066 5017 161113
rect 4217 160352 4258 161066
rect 4983 160352 5017 161066
rect 4217 160313 5017 160352
rect 109936 160162 116936 169698
rect 109936 159698 110021 160162
rect 116816 159698 116936 160162
rect 109936 150162 116936 159698
rect 109936 149698 110021 150162
rect 116816 149698 116936 150162
rect 109936 140162 116936 149698
rect 109936 139698 110021 140162
rect 116816 139698 116936 140162
rect 109936 130162 116936 139698
rect 109936 129698 110021 130162
rect 116816 129698 116936 130162
rect 109936 120162 116936 129698
rect 109936 119698 110021 120162
rect 116816 119698 116936 120162
rect 109936 110162 116936 119698
rect 109936 109698 110021 110162
rect 116816 109698 116936 110162
rect 109936 100162 116936 109698
rect 109936 99698 110021 100162
rect 116816 99698 116936 100162
rect 109936 90162 116936 99698
rect 109936 89698 110021 90162
rect 116816 89698 116936 90162
rect 10265 86219 13265 86428
rect 10265 81681 10344 86219
rect 13143 81681 13265 86219
rect 10265 76201 13265 81681
rect 10265 71741 10357 76201
rect 13169 71741 13265 76201
rect 1687 44026 9128 44216
rect 1687 39587 1813 44026
rect 8962 39587 9128 44026
rect 1687 39426 9128 39587
rect 1399 34000 9121 34185
rect 1399 29539 1559 34000
rect 8951 29539 9121 34000
rect 1399 29395 9121 29539
rect 10265 8084 13265 71741
rect 109936 80162 116936 89698
rect 109936 79698 110021 80162
rect 116816 79698 116936 80162
rect 109936 70162 116936 79698
rect 109936 69698 110021 70162
rect 116816 69698 116936 70162
rect 109936 60162 116936 69698
rect 109936 59698 110021 60162
rect 116816 59698 116936 60162
rect 109936 50162 116936 59698
rect 109936 49698 110021 50162
rect 116816 49698 116936 50162
rect 109936 40162 116936 49698
rect 109936 39698 110021 40162
rect 116816 39698 116936 40162
rect 109936 30162 116936 39698
rect 109936 29698 110021 30162
rect 116816 29698 116936 30162
rect 109936 20162 116936 29698
rect 119936 195145 126936 195210
rect 119936 194628 119991 195145
rect 126852 194628 126936 195145
rect 119936 188265 126936 194628
rect 119936 183580 120133 188265
rect 126688 183580 126936 188265
rect 119936 175168 126936 183580
rect 119936 174631 120020 175168
rect 126822 174631 126936 175168
rect 119936 165168 126936 174631
rect 119936 164631 120020 165168
rect 126822 164631 126936 165168
rect 119936 155168 126936 164631
rect 119936 154631 120020 155168
rect 126822 154631 126936 155168
rect 119936 145168 126936 154631
rect 119936 144631 120020 145168
rect 126822 144631 126936 145168
rect 119936 135168 126936 144631
rect 119936 134631 120020 135168
rect 126822 134631 126936 135168
rect 119936 125168 126936 134631
rect 119936 124631 120020 125168
rect 126822 124631 126936 125168
rect 119936 115168 126936 124631
rect 119936 114631 120020 115168
rect 126822 114631 126936 115168
rect 119936 105168 126936 114631
rect 119936 104631 120020 105168
rect 126822 104631 126936 105168
rect 119936 95168 126936 104631
rect 119936 94631 120020 95168
rect 126822 94631 126936 95168
rect 119936 85168 126936 94631
rect 119936 84631 120020 85168
rect 126822 84631 126936 85168
rect 119936 75168 126936 84631
rect 119936 74631 120020 75168
rect 126822 74631 126936 75168
rect 119936 65168 126936 74631
rect 119936 64631 120020 65168
rect 126822 64631 126936 65168
rect 119936 55168 126936 64631
rect 119936 54631 120020 55168
rect 126822 54631 126936 55168
rect 119936 45168 126936 54631
rect 119936 44631 120020 45168
rect 126822 44631 126936 45168
rect 119936 35168 126936 44631
rect 119936 34631 120020 35168
rect 126822 34631 126936 35168
rect 119936 26772 126936 34631
rect 119936 22141 120212 26772
rect 126733 22141 126936 26772
rect 119936 21906 126936 22141
rect 129936 176657 136936 207012
rect 175073 208037 175402 208065
rect 175073 206605 175100 208037
rect 175364 206605 175402 208037
rect 175073 206567 175402 206605
rect 205173 208037 205502 208065
rect 205173 206605 205200 208037
rect 205464 206605 205502 208037
rect 205173 206567 205502 206605
rect 235333 208037 235662 208065
rect 235333 206605 235360 208037
rect 235624 206605 235662 208037
rect 235333 206567 235662 206605
rect 265323 208037 265652 208065
rect 265323 206605 265350 208037
rect 265614 206605 265652 208037
rect 265323 206567 265652 206605
rect 295473 208037 295802 208065
rect 295473 206605 295500 208037
rect 295764 206605 295802 208037
rect 295473 206567 295802 206605
rect 325573 208037 325902 208065
rect 325573 206605 325600 208037
rect 325864 206605 325902 208037
rect 325573 206567 325902 206605
rect 355673 208037 356002 208065
rect 355673 206605 355700 208037
rect 355964 206605 356002 208037
rect 355673 206567 356002 206605
rect 157538 205533 157910 205564
rect 157538 204093 157566 205533
rect 157877 204093 157910 205533
rect 157538 204068 157910 204093
rect 187638 205533 188010 205564
rect 187638 204093 187666 205533
rect 187977 204093 188010 205533
rect 187638 204068 188010 204093
rect 217738 205533 218110 205564
rect 217738 204093 217766 205533
rect 218077 204093 218110 205533
rect 217738 204068 218110 204093
rect 247788 205533 248160 205564
rect 247788 204093 247816 205533
rect 248127 204093 248160 205533
rect 247788 204068 248160 204093
rect 278018 205533 278340 205564
rect 278018 204093 278046 205533
rect 278307 204093 278340 205533
rect 278018 204068 278340 204093
rect 308038 205533 308410 205564
rect 308038 204093 308066 205533
rect 308377 204093 308410 205533
rect 308038 204068 308410 204093
rect 338138 205533 338510 205564
rect 338138 204093 338166 205533
rect 338477 204093 338510 205533
rect 338138 204068 338510 204093
rect 368238 205533 368610 205564
rect 368238 204093 368266 205533
rect 368577 204093 368610 205533
rect 368238 204068 368610 204093
rect 630489 204214 631298 214163
rect 172596 203026 172965 203066
rect 172596 201601 172628 203026
rect 172929 201601 172965 203026
rect 172596 201566 172965 201601
rect 202696 203026 203065 203066
rect 202696 201601 202728 203026
rect 203029 201601 203065 203026
rect 202696 201566 203065 201601
rect 232796 203026 233165 203066
rect 232796 201601 232828 203026
rect 233129 201601 233165 203026
rect 232796 201566 233165 201601
rect 262896 203026 263265 203066
rect 262896 201601 262928 203026
rect 263229 201601 263265 203026
rect 262896 201566 263265 201601
rect 292886 203026 293255 203066
rect 292886 201601 292918 203026
rect 293219 201601 293255 203026
rect 292886 201566 293255 201601
rect 323096 203026 323465 203066
rect 323096 201601 323128 203026
rect 323429 201601 323465 203026
rect 323096 201566 323465 201601
rect 353196 203026 353565 203066
rect 353196 201601 353228 203026
rect 353529 201601 353565 203026
rect 353196 201566 353565 201601
rect 387736 202845 394099 203087
rect 387736 201297 387985 202845
rect 393910 201297 394099 202845
rect 630489 202234 630549 204214
rect 631216 202234 631298 204214
rect 630489 202148 631298 202234
rect 633150 204351 633959 215842
rect 633150 202289 633219 204351
rect 633869 202289 633959 204351
rect 633150 202216 633959 202289
rect 129936 176107 130009 176657
rect 136855 176107 136936 176657
rect 129936 150657 136936 176107
rect 129936 150107 130009 150657
rect 136855 150107 136936 150657
rect 129936 124657 136936 150107
rect 129936 124107 130009 124657
rect 136855 124107 136936 124657
rect 129936 98657 136936 124107
rect 129936 98107 130009 98657
rect 136855 98107 136936 98657
rect 129936 72657 136936 98107
rect 129936 72107 130009 72657
rect 136855 72107 136936 72657
rect 129936 46657 136936 72107
rect 129936 46107 130009 46657
rect 136855 46107 136936 46657
rect 129936 29832 136936 46107
rect 129936 29243 129997 29832
rect 136890 29243 136936 29832
rect 109936 19698 110021 20162
rect 116816 19698 116936 20162
rect 103995 16262 104641 16287
rect 103995 15523 104025 16262
rect 104608 15523 104641 16262
rect 103995 15490 104641 15523
rect 103999 8961 104179 15490
rect 109936 14272 116936 19698
rect 105009 13315 105775 13367
rect 105009 12252 105051 13315
rect 105711 12252 105775 13315
rect 105009 12187 105775 12252
rect 105299 10514 105479 12187
rect 109936 9641 110144 14272
rect 116665 9641 116936 14272
rect 109936 9338 116936 9641
rect 129936 14174 136936 29243
rect 138936 188234 145936 188621
rect 138936 183549 139135 188234
rect 145690 183549 145936 188234
rect 138936 163654 145936 183549
rect 387736 188204 394099 201297
rect 637861 196101 638663 196153
rect 608559 195168 613559 195344
rect 608559 190557 608763 195168
rect 613356 190557 613559 195168
rect 629447 195247 632454 195413
rect 629447 193669 629587 195247
rect 632313 193669 632454 195247
rect 629447 193511 632454 193669
rect 637861 193295 637917 196101
rect 638627 193295 638663 196101
rect 637861 193229 638663 193295
rect 635066 192443 635866 192507
rect 635066 191771 635130 192443
rect 635802 191771 635866 192443
rect 635066 191707 635866 191771
rect 387736 183649 388000 188204
rect 393895 183649 394099 188204
rect 387736 183011 394099 183649
rect 602559 188229 607559 188383
rect 602559 183618 602772 188229
rect 607365 183618 607559 188229
rect 138936 163065 138995 163654
rect 145878 163065 145936 163654
rect 138936 137654 145936 163065
rect 138936 137065 138995 137654
rect 145878 137065 145936 137654
rect 138936 111654 145936 137065
rect 138936 111065 138995 111654
rect 145878 111065 145936 111654
rect 138936 85654 145936 111065
rect 138936 85065 138995 85654
rect 145878 85065 145936 85654
rect 138936 59654 145936 85065
rect 138936 59065 138995 59654
rect 145878 59065 145936 59654
rect 138936 33654 145936 59065
rect 138936 33065 138995 33654
rect 145878 33065 145936 33654
rect 138936 26804 145936 33065
rect 138936 22173 139167 26804
rect 145688 22173 145936 26804
rect 138936 21906 145936 22173
rect 602559 163571 607559 183618
rect 602559 163148 602628 163571
rect 607445 163148 607559 163571
rect 602559 137571 607559 163148
rect 602559 137148 602628 137571
rect 607445 137148 607559 137571
rect 602559 111571 607559 137148
rect 602559 111148 602628 111571
rect 607445 111148 607559 111571
rect 602559 85571 607559 111148
rect 602559 85148 602628 85571
rect 607445 85148 607559 85571
rect 602559 59571 607559 85148
rect 602559 59148 602628 59571
rect 607445 59148 607559 59571
rect 602559 46757 607559 59148
rect 602559 46284 602636 46757
rect 607470 46284 607559 46757
rect 602559 45120 607559 46284
rect 602559 44647 602600 45120
rect 607434 44647 607559 45120
rect 602559 33615 607559 44647
rect 602559 33085 602623 33615
rect 607495 33085 607559 33615
rect 602559 18529 607559 33085
rect 129936 9543 130166 14174
rect 136687 9543 136936 14174
rect 129936 9207 136936 9543
rect 202686 14832 207477 15041
rect 202686 10234 202782 14832
rect 207285 10234 207477 14832
rect 202686 9725 202830 10234
rect 207269 9725 207477 10234
rect 202686 9501 207477 9725
rect 212765 14800 217556 14993
rect 212765 10202 212877 14800
rect 217380 10202 217556 14800
rect 602559 14168 602693 18529
rect 607423 14168 607559 18529
rect 608559 176601 613559 190557
rect 633668 191042 634468 191106
rect 633668 190370 633732 191042
rect 634404 190370 634468 191042
rect 633668 190306 634468 190370
rect 636461 189642 637261 189706
rect 636461 188970 636525 189642
rect 637197 188970 637261 189642
rect 636461 188906 637261 188970
rect 637855 188248 638655 188312
rect 670962 188308 671282 192626
rect 671622 189708 671942 192616
rect 672282 191108 672602 192577
rect 672942 192508 673262 192587
rect 672940 192506 673262 192508
rect 672940 191706 672942 192506
rect 673252 191706 673262 192506
rect 672940 191704 673262 191706
rect 672280 191106 672604 191108
rect 672280 190306 672282 191106
rect 672602 190306 672604 191106
rect 672280 190304 672604 190306
rect 671620 189706 671944 189708
rect 671620 188906 671622 189706
rect 671942 188906 671944 189706
rect 671620 188904 671944 188906
rect 637855 187576 637919 188248
rect 638591 187576 638655 188248
rect 637855 187512 638655 187576
rect 670960 188306 671284 188308
rect 670960 187506 670962 188306
rect 671282 187506 671284 188306
rect 670960 187504 671284 187506
rect 670962 183853 671282 187504
rect 671622 184514 671942 188904
rect 672282 185048 672602 190304
rect 672942 185551 673262 191704
rect 608559 176153 608613 176601
rect 613500 176153 613559 176601
rect 608559 150601 613559 176153
rect 608559 150153 608613 150601
rect 613500 150153 613559 150601
rect 608559 124601 613559 150153
rect 635066 147047 635866 147111
rect 635066 146375 635130 147047
rect 635802 146375 635866 147047
rect 635066 146311 635866 146375
rect 633667 145639 634467 145703
rect 633667 144967 633731 145639
rect 634403 144967 634467 145639
rect 633667 144903 634467 144967
rect 636459 144235 637259 144299
rect 636459 143563 636523 144235
rect 637195 143563 637259 144235
rect 636459 143499 637259 143563
rect 670962 142908 671282 147196
rect 671622 144308 671942 147255
rect 672282 145708 672602 147265
rect 672942 147108 673262 147255
rect 672940 147106 673262 147108
rect 672940 146306 672942 147106
rect 673252 146306 673262 147106
rect 672940 146304 673262 146306
rect 672280 145706 672604 145708
rect 672280 144906 672282 145706
rect 672602 144906 672604 145706
rect 672280 144904 672604 144906
rect 671620 144306 671944 144308
rect 671620 143506 671622 144306
rect 671942 143506 671944 144306
rect 671620 143504 671944 143506
rect 670960 142906 671284 142908
rect 637866 142842 638666 142906
rect 637866 142170 637930 142842
rect 638602 142170 638666 142842
rect 637866 142106 638666 142170
rect 670960 142106 670962 142906
rect 671282 142106 671284 142906
rect 670960 142104 671284 142106
rect 670962 138863 671282 142104
rect 671622 139538 671942 143504
rect 672282 140151 672602 144904
rect 672942 140815 673262 146304
rect 608559 124153 608613 124601
rect 613500 124153 613559 124601
rect 608559 98601 613559 124153
rect 635070 101637 635870 101701
rect 635070 100965 635134 101637
rect 635806 100965 635870 101637
rect 635070 100901 635870 100965
rect 633664 100241 634464 100305
rect 633664 99569 633728 100241
rect 634400 99569 634464 100241
rect 633664 99505 634464 99569
rect 608559 98153 608613 98601
rect 613500 98153 613559 98601
rect 608559 72601 613559 98153
rect 636469 98843 637269 98907
rect 636469 98171 636533 98843
rect 637205 98171 637269 98843
rect 636469 98107 637269 98171
rect 670962 97508 671282 101864
rect 671622 98908 671942 101845
rect 672282 100308 672602 101815
rect 672942 101708 673262 101775
rect 672940 101706 673262 101708
rect 672940 100906 672942 101706
rect 673252 100906 673262 101706
rect 672940 100904 673262 100906
rect 672280 100306 672604 100308
rect 672280 99506 672282 100306
rect 672602 99506 672604 100306
rect 672280 99504 672604 99506
rect 671620 98906 671944 98908
rect 671620 98106 671622 98906
rect 671942 98106 671944 98906
rect 671620 98104 671944 98106
rect 670960 97506 671284 97508
rect 637867 97439 638667 97503
rect 637867 96767 637931 97439
rect 638603 96767 638667 97439
rect 637867 96703 638667 96767
rect 670960 96706 670962 97506
rect 671282 96706 671284 97506
rect 670960 96704 671284 96706
rect 670962 93621 671282 96704
rect 671622 94338 671942 98104
rect 672282 94998 672602 99504
rect 672942 95602 673262 100904
rect 608559 72153 608613 72601
rect 613500 72153 613559 72601
rect 608559 65265 613559 72153
rect 614123 75734 615417 75779
rect 614123 74690 614156 75734
rect 615367 74690 615417 75734
rect 614123 66919 615417 74690
rect 614123 66521 616130 66919
rect 614173 66519 616130 66521
rect 608559 64636 608612 65265
rect 613504 64636 613559 65265
rect 608559 47558 613559 64636
rect 614106 65891 615647 66209
rect 622876 66145 626729 66212
rect 614106 63098 615400 65891
rect 622870 65883 626729 66145
rect 622870 65118 624708 65883
rect 622870 64798 622897 65118
rect 624672 64798 624708 65118
rect 622870 64757 624708 64798
rect 614106 61750 614165 63098
rect 615335 61750 615400 63098
rect 614106 61685 615400 61750
rect 608559 47085 608618 47558
rect 613452 47085 613559 47558
rect 608559 45911 613559 47085
rect 608559 45438 608633 45911
rect 613467 45438 613559 45911
rect 608559 44256 613559 45438
rect 608559 43861 608607 44256
rect 613498 43861 613559 44256
rect 608559 20655 613559 43861
rect 608559 16294 608661 20655
rect 613391 16294 613559 20655
rect 608559 16161 613559 16294
rect 602559 14061 607559 14168
rect 222286 11866 631506 11878
rect 222231 11854 631506 11866
rect 212765 9693 212909 10202
rect 217348 9693 217556 10202
rect 212765 9453 217556 9693
rect 222053 11787 631506 11854
rect 104417 8932 104879 8947
rect 104417 8494 104438 8932
rect 104782 8494 104879 8932
rect 104417 8473 104879 8494
rect 106179 8084 106359 8902
rect 222053 8084 628597 11787
rect 10265 7973 628597 8084
rect 631428 7973 631506 11787
rect 10265 7878 631506 7973
rect 10265 4775 225362 7878
rect 229032 6588 635531 6686
rect 229032 6582 632642 6588
rect 10265 3815 106953 4775
rect 229032 3803 530645 6582
rect 107864 3755 530645 3803
rect 107864 1861 107928 3755
rect 108561 2784 530645 3755
rect 535200 6573 632642 6582
rect 535200 2784 540643 6573
rect 108561 2775 540643 2784
rect 545198 2815 632642 6573
rect 635402 2815 635531 6588
rect 545198 2775 635531 2815
rect 108561 2686 635531 2775
rect 108561 1861 231437 2686
rect 107864 1803 231437 1861
<< via4 >>
rect 9771 954376 10560 955176
rect 73036 954443 73708 955115
rect 9771 945799 10560 947452
rect 14566 952859 15343 953659
rect 74441 952926 75113 953598
rect 75849 957516 76521 958188
rect 77228 956012 77900 956684
rect 124635 954441 125307 955113
rect 126040 952920 126712 953592
rect 127441 957520 128113 958192
rect 128823 956026 129495 956698
rect 176246 954442 176918 955114
rect 177636 952916 178308 953588
rect 179045 957526 179717 958198
rect 180427 956015 181099 956687
rect 227824 954446 228496 955118
rect 229234 952915 229906 953587
rect 230640 957524 231312 958196
rect 232030 956016 232702 956688
rect 279439 954436 280111 955108
rect 280845 952936 281517 953608
rect 282251 957511 282923 958183
rect 283650 956007 284322 956679
rect 331038 954437 331710 955109
rect 332434 952922 333106 953594
rect 333842 957536 334514 958208
rect 335231 956025 335903 956697
rect 397037 954438 397709 955110
rect 398454 952928 399126 953600
rect 399823 957508 400495 958180
rect 401248 956026 401920 956698
rect 474244 954446 474916 955118
rect 475644 952920 476316 953592
rect 477030 957516 477702 958188
rect 478446 956018 479118 956690
rect 525432 954442 526104 955114
rect 526844 952924 527516 953596
rect 528241 957524 528913 958196
rect 529646 956010 530318 956682
rect 533513 953869 535792 954543
rect 533513 952297 535809 952967
rect 537238 952456 541828 955220
rect 547180 952441 551770 955205
rect 14566 944562 15343 946390
rect 622828 943225 624321 944801
rect 625971 943324 627460 945737
rect 2875 908397 3547 909069
rect 625724 908163 629596 908835
rect 1690 907008 2362 907680
rect 620715 906775 624587 907447
rect 636532 905361 637204 906033
rect 637932 903971 638604 904643
rect 13382 883618 17116 888015
rect 620860 879253 624447 883577
rect 13431 873619 17081 878016
rect 17081 873619 17165 878016
rect 620810 869167 624397 873491
rect 4359 799066 5171 803652
rect 4351 789089 5163 793675
rect 633781 789897 635118 794462
rect 2881 782395 3553 783067
rect 1701 781034 2373 781706
rect 633749 779952 635086 784517
rect 13329 764964 17201 765636
rect 8334 763569 12206 764241
rect 2886 739208 3558 739880
rect 1690 737825 2362 738497
rect 625719 730172 629591 730844
rect 620720 728769 624592 729441
rect 636525 727361 637197 728033
rect 637926 725975 638598 726647
rect 13337 721564 17209 722236
rect 8330 720158 12202 720830
rect 2892 696027 3564 696699
rect 1695 694622 2367 695294
rect 625714 684969 629586 685641
rect 620720 683557 624592 684229
rect 636530 682171 637202 682843
rect 637931 680761 638603 681433
rect 13348 678517 17220 679189
rect 8334 676967 12206 677639
rect 2886 652824 3558 653496
rect 1684 651402 2356 652074
rect 625724 639767 629596 640439
rect 620725 638374 624597 639046
rect 636542 636963 637214 637635
rect 13337 635554 17209 636226
rect 637921 635565 638593 636237
rect 8342 634167 12214 634839
rect 2903 609620 3575 610292
rect 1690 608249 2362 608921
rect 625728 594574 629600 595246
rect 620715 593171 624587 593843
rect 13340 591966 17212 592638
rect 636532 591770 637204 592442
rect 8330 590560 12202 591232
rect 637926 590367 638598 591039
rect 2897 566637 3569 567309
rect 1684 565215 2356 565887
rect 13341 548764 17213 549436
rect 625728 549366 629600 550038
rect 8330 547375 12202 548047
rect 620725 547973 624597 548645
rect 636523 546567 637195 547239
rect 637935 545173 638607 545845
rect 2903 523603 3575 524275
rect 1673 522215 2345 522887
rect 13337 505568 17209 506240
rect 8323 504166 12195 504838
rect 625714 504168 629586 504840
rect 620729 502765 624601 503437
rect 636529 501371 637201 502043
rect 637930 499975 638602 500647
rect 630713 475283 632588 479910
rect 630706 465305 632581 469932
rect 625719 460566 629591 461238
rect 620715 459173 624587 459845
rect 6326 454442 7225 459103
rect 636530 457768 637202 458440
rect 637928 456369 638600 457041
rect 6315 444435 7201 449139
rect 625815 435779 629491 435866
rect 625815 431386 625855 435779
rect 625855 431386 629491 435779
rect 625815 431326 629491 431386
rect 625811 421357 629472 425749
rect 8417 416868 12175 416912
rect 8417 412440 12132 416868
rect 12132 412440 12175 416868
rect 8374 402360 12132 406832
rect 2903 395607 3575 396279
rect 1690 394224 2362 394896
rect 633737 387094 635564 391672
rect 13329 377751 17201 378423
rect 633726 377156 635553 381734
rect 8334 376364 12206 377036
rect 625724 372180 629596 372852
rect 620720 370777 624592 371449
rect 636529 369367 637201 370039
rect 637929 367963 638601 368635
rect 2886 352624 3558 353296
rect 1684 351207 2356 351879
rect 13329 334560 17201 335232
rect 8342 333157 12214 333829
rect 625724 327378 629596 328050
rect 620729 325994 624601 326666
rect 636529 324565 637201 325237
rect 637924 323188 638596 323860
rect 2875 309640 3547 310312
rect 1673 308212 2345 308884
rect 13329 291360 17201 292032
rect 8332 289950 12204 290622
rect 625724 282556 629596 283228
rect 620734 281177 624606 281849
rect 636524 279772 637196 280444
rect 637915 278367 638587 279039
rect 2884 266620 3556 267292
rect 1684 265219 2356 265891
rect 13328 248152 17200 248824
rect 8332 246745 12204 247417
rect 6344 233558 7160 238811
rect 6355 227791 7149 231502
rect 8378 234855 12145 240968
rect 8423 227903 12144 231501
rect 13396 237313 17117 240911
rect 13419 227870 17140 231468
rect 620804 239279 624519 242438
rect 620817 230071 624505 233434
rect 625807 237845 629455 242425
rect 625807 237173 629455 237845
rect 625807 236391 629455 237173
rect 625848 230044 629536 233407
rect 630784 235468 632547 242425
rect 636532 234364 637204 235036
rect 630865 230058 632506 233461
rect 637933 232978 638605 233650
rect 2881 223622 3553 224294
rect 1684 222221 2356 222893
rect 4272 211917 4958 213801
rect 159217 224103 159507 225528
rect 189317 224103 189607 225528
rect 219417 224103 219707 225528
rect 249517 224103 249807 225528
rect 279617 224103 279907 225528
rect 309717 224103 310007 225528
rect 339817 224103 340107 225528
rect 369917 224103 370207 225528
rect 174274 221605 174572 223017
rect 204374 221605 204672 223017
rect 234474 221605 234772 223017
rect 264574 221605 264872 223017
rect 294674 221605 294972 223017
rect 324774 221605 325072 223017
rect 354874 221605 355172 223017
rect 160027 219105 160382 220516
rect 190127 219105 190482 220516
rect 220227 219105 220582 220516
rect 250267 219105 250542 220516
rect 280427 219105 280782 220516
rect 310527 219105 310882 220516
rect 340627 219105 340982 220516
rect 370727 219105 371082 220516
rect 175919 216618 176178 218030
rect 206019 216618 206278 218030
rect 236119 216618 236378 218030
rect 266219 216613 266478 218030
rect 296319 216618 296578 218030
rect 326419 216618 326678 218030
rect 356519 216618 356778 218030
rect 158407 214096 158695 215526
rect 188507 214096 188795 215526
rect 218607 214096 218895 215526
rect 248797 214096 249075 215526
rect 278807 214096 279045 215526
rect 308907 214096 309195 215526
rect 339007 214096 339295 215526
rect 369107 214096 369395 215526
rect 5673 211897 6359 213781
rect 110403 207012 116528 213365
rect 5686 204956 6358 205628
rect 4289 203553 4961 204225
rect 110021 199698 116816 200162
rect 130322 207012 136447 213365
rect 173451 211601 173725 213029
rect 203551 211601 203825 213029
rect 233701 211601 233975 213029
rect 263691 211601 263965 212949
rect 293851 211601 294125 213029
rect 323951 211601 324225 213029
rect 354051 211601 354325 213029
rect 160095 209096 160347 210533
rect 190195 209096 190447 210533
rect 220295 209096 220547 210533
rect 250275 209096 250527 210533
rect 280495 209096 280747 210533
rect 310595 209096 310847 210533
rect 340695 209096 340947 210533
rect 370795 209096 371047 210533
rect 110021 189698 116816 190162
rect 2887 180614 3561 181286
rect 1653 179188 2388 179924
rect 110021 179698 116816 180162
rect 110021 169698 116816 170162
rect 5662 161736 6387 162450
rect 4258 160352 4983 161066
rect 110021 159698 116816 160162
rect 110021 149698 116816 150162
rect 110021 139698 116816 140162
rect 110021 129698 116816 130162
rect 110021 119698 116816 120162
rect 110021 109698 116816 110162
rect 110021 99698 116816 100162
rect 110021 89698 116816 90162
rect 4302 39598 8940 43927
rect 4280 30314 8918 33967
rect 4280 29638 8917 30314
rect 110021 79698 116816 80162
rect 110021 69698 116816 70162
rect 110021 59698 116816 60162
rect 110021 49698 116816 50162
rect 110021 39698 116816 40162
rect 110021 29698 116816 30162
rect 119991 194628 126852 195145
rect 120133 183580 126688 188265
rect 120020 174631 126822 175168
rect 120020 164631 126822 165168
rect 120020 154631 126822 155168
rect 120020 144631 126822 145168
rect 120020 134631 126822 135168
rect 120020 124631 126822 125168
rect 120020 114631 126822 115168
rect 120020 104631 126822 105168
rect 120020 94631 126822 95168
rect 120020 84631 126822 85168
rect 120020 74631 126822 75168
rect 120020 64631 126822 65168
rect 120020 54631 126822 55168
rect 120020 44631 126822 45168
rect 120020 34631 126822 35168
rect 120212 22141 126733 26772
rect 175100 206605 175364 208037
rect 205200 206605 205464 208037
rect 235360 206605 235624 208037
rect 265350 206605 265614 208037
rect 295500 206605 295764 208037
rect 325600 206605 325864 208037
rect 355700 206605 355964 208037
rect 157566 204093 157877 205533
rect 187666 204093 187977 205533
rect 217766 204093 218077 205533
rect 247816 204093 248127 205533
rect 278046 204093 278307 205533
rect 308066 204093 308377 205533
rect 338166 204093 338477 205533
rect 368266 204093 368577 205533
rect 172628 201601 172929 203026
rect 202728 201601 203029 203026
rect 232828 201601 233129 203026
rect 262928 201601 263229 203026
rect 292918 201601 293219 203026
rect 323128 201601 323429 203026
rect 353228 201601 353529 203026
rect 387985 201297 393910 202845
rect 630549 202234 631216 204214
rect 633219 202289 633869 204351
rect 130009 176107 136855 176657
rect 130009 150107 136855 150657
rect 130009 124107 136855 124657
rect 130009 98107 136855 98657
rect 130009 72107 136855 72657
rect 130009 46107 136855 46657
rect 129997 29243 136890 29832
rect 110021 19698 116816 20162
rect 104025 15523 104608 16262
rect 105051 12252 105711 13315
rect 110144 9641 116665 14272
rect 139135 183549 145690 188234
rect 608763 190557 613356 195168
rect 629587 193669 632313 195247
rect 637917 193295 638627 196101
rect 635130 191771 635802 192443
rect 388000 183649 393895 188204
rect 602772 183618 607365 188229
rect 138995 163065 145878 163654
rect 138995 137065 145878 137654
rect 138995 111065 145878 111654
rect 138995 85065 145878 85654
rect 138995 59065 145878 59654
rect 138995 33065 145878 33654
rect 139167 22173 145688 26804
rect 602628 163148 607445 163571
rect 602628 137148 607445 137571
rect 602628 111148 607445 111571
rect 602628 85148 607445 85571
rect 602628 59148 607445 59571
rect 602636 46284 607470 46757
rect 602600 44647 607434 45120
rect 602623 33085 607495 33615
rect 130166 9543 136687 14174
rect 202782 14752 207285 14832
rect 202782 10234 202830 14752
rect 202830 10234 207269 14752
rect 207269 10234 207285 14752
rect 212877 14720 217380 14800
rect 212877 10202 212909 14720
rect 212909 10202 217348 14720
rect 217348 10202 217380 14720
rect 602693 14168 607423 18529
rect 633732 190370 634404 191042
rect 636525 188970 637197 189642
rect 637919 187576 638591 188248
rect 608613 176153 613500 176601
rect 608613 150153 613500 150601
rect 635130 146375 635802 147047
rect 633731 144967 634403 145639
rect 636523 143563 637195 144235
rect 637930 142170 638602 142842
rect 608613 124153 613500 124601
rect 635134 100965 635806 101637
rect 633728 99569 634400 100241
rect 608613 98153 613500 98601
rect 636533 98171 637205 98843
rect 637931 96767 638603 97439
rect 608613 72153 613500 72601
rect 614156 74690 615367 75734
rect 608612 64636 613504 65265
rect 622897 64798 624672 65118
rect 614165 61750 615335 63098
rect 608618 47085 613452 47558
rect 608633 45438 613467 45911
rect 608607 43861 613498 44256
rect 608661 16294 613391 20655
rect 628597 7973 631428 11787
rect 632642 2815 635402 6588
<< metal5 >>
rect 1623 958255 2423 958257
rect 1623 958208 638667 958255
rect 1623 958198 333842 958208
rect 1623 958192 179045 958198
rect 1623 958188 127441 958192
rect 1623 957516 75849 958188
rect 76521 957520 127441 958188
rect 128113 957526 179045 958192
rect 179717 958196 333842 958198
rect 179717 957526 230640 958196
rect 128113 957524 230640 957526
rect 231312 958183 333842 958196
rect 231312 957524 282251 958183
rect 128113 957520 282251 957524
rect 76521 957516 282251 957520
rect 1623 957511 282251 957516
rect 282923 957536 333842 958183
rect 334514 958196 638667 958208
rect 334514 958188 528241 958196
rect 334514 958180 477030 958188
rect 334514 957536 399823 958180
rect 282923 957511 399823 957536
rect 1623 957508 399823 957511
rect 400495 957516 477030 958180
rect 477702 957524 528241 958188
rect 528913 957524 638667 958196
rect 477702 957516 638667 957524
rect 400495 957508 638667 957516
rect 1623 957455 638667 957508
rect 1623 907680 2423 957455
rect 1623 907008 1690 907680
rect 2362 907008 2423 907680
rect 1623 781706 2423 907008
rect 1623 781034 1701 781706
rect 2373 781034 2423 781706
rect 1623 738497 2423 781034
rect 1623 737825 1690 738497
rect 2362 737825 2423 738497
rect 1623 695294 2423 737825
rect 1623 694622 1695 695294
rect 2367 694622 2423 695294
rect 1623 652074 2423 694622
rect 1623 651402 1684 652074
rect 2356 651402 2423 652074
rect 1623 608921 2423 651402
rect 1623 608249 1690 608921
rect 2362 608249 2423 608921
rect 1623 565887 2423 608249
rect 1623 565215 1684 565887
rect 2356 565215 2423 565887
rect 1623 522887 2423 565215
rect 1623 522215 1673 522887
rect 2345 522215 2423 522887
rect 1623 394896 2423 522215
rect 1623 394224 1690 394896
rect 2362 394224 2423 394896
rect 1623 351879 2423 394224
rect 1623 351207 1684 351879
rect 2356 351207 2423 351879
rect 1623 308884 2423 351207
rect 1623 308212 1673 308884
rect 2345 308212 2423 308884
rect 1623 265891 2423 308212
rect 1623 265219 1684 265891
rect 2356 265219 2423 265891
rect 1623 222893 2423 265219
rect 1623 222221 1684 222893
rect 2356 222221 2423 222893
rect 1623 179924 2423 222221
rect 1623 179188 1653 179924
rect 2388 179188 2423 179924
rect 1623 107739 2423 179188
rect 2823 956758 3623 956762
rect 2823 956698 637267 956758
rect 2823 956684 128823 956698
rect 2823 956012 77228 956684
rect 77900 956026 128823 956684
rect 129495 956697 401248 956698
rect 129495 956688 335231 956697
rect 129495 956687 232030 956688
rect 129495 956026 180427 956687
rect 77900 956015 180427 956026
rect 181099 956016 232030 956687
rect 232702 956679 335231 956688
rect 232702 956016 283650 956679
rect 181099 956015 283650 956016
rect 77900 956012 283650 956015
rect 2823 956007 283650 956012
rect 284322 956025 335231 956679
rect 335903 956026 401248 956697
rect 401920 956690 637267 956698
rect 401920 956026 478446 956690
rect 335903 956025 478446 956026
rect 284322 956018 478446 956025
rect 479118 956682 637267 956690
rect 479118 956018 529646 956682
rect 284322 956010 529646 956018
rect 530318 956010 637267 956682
rect 284322 956007 637267 956010
rect 2823 955958 637267 956007
rect 2823 909069 3623 955958
rect 633657 955325 635657 955329
rect 537099 955220 635657 955325
rect 9747 955176 10584 955200
rect 9445 954376 9771 955176
rect 10560 955118 285188 955176
rect 10560 955115 227824 955118
rect 10560 954443 73036 955115
rect 73708 955114 227824 955115
rect 73708 955113 176246 955114
rect 73708 954443 124635 955113
rect 10560 954441 124635 954443
rect 125307 954442 176246 955113
rect 176918 954446 227824 955114
rect 228496 955108 285188 955118
rect 228496 954446 279439 955108
rect 176918 954442 279439 954446
rect 125307 954441 279439 954442
rect 10560 954436 279439 954441
rect 280111 954436 285188 955108
rect 10560 954376 285188 954436
rect 329924 955118 531466 955176
rect 329924 955110 474244 955118
rect 329924 955109 397037 955110
rect 329924 954437 331038 955109
rect 331710 954438 397037 955109
rect 397709 954446 474244 955110
rect 474916 955114 531466 955118
rect 474916 954446 525432 955114
rect 397709 954442 525432 954446
rect 526104 954606 531466 955114
rect 526104 954543 535861 954606
rect 526104 954442 533513 954543
rect 397709 954438 533513 954442
rect 331710 954437 533513 954438
rect 329924 954376 533513 954437
rect 9747 954352 10584 954376
rect 530666 953869 533513 954376
rect 535792 953869 535861 954543
rect 530666 953806 535861 953869
rect 14542 953659 15367 953683
rect 14423 952859 14566 953659
rect 15343 953608 285188 953659
rect 15343 953598 280845 953608
rect 15343 952926 74441 953598
rect 75113 953592 280845 953598
rect 75113 952926 126040 953592
rect 15343 952920 126040 952926
rect 126712 953588 280845 953592
rect 126712 952920 177636 953588
rect 15343 952916 177636 952920
rect 178308 953587 280845 953588
rect 178308 952916 229234 953587
rect 15343 952915 229234 952916
rect 229906 952936 280845 953587
rect 281517 952936 285188 953608
rect 229906 952915 285188 952936
rect 15343 952859 285188 952915
rect 329924 953600 530027 953659
rect 329924 953594 398454 953600
rect 329924 952922 332434 953594
rect 333106 952928 398454 953594
rect 399126 953596 530027 953600
rect 399126 953592 526844 953596
rect 399126 952928 475644 953592
rect 333106 952922 475644 952928
rect 329924 952920 475644 952922
rect 476316 952924 526844 953592
rect 527516 953032 530027 953596
rect 527516 952967 535876 953032
rect 527516 952924 533513 952967
rect 476316 952920 533513 952924
rect 329924 952859 533513 952920
rect 14542 952835 15367 952859
rect 529227 952297 533513 952859
rect 535809 952297 535876 952967
rect 537099 952456 537238 955220
rect 541828 955205 635657 955220
rect 541828 952456 547180 955205
rect 537099 952441 547180 952456
rect 551770 952441 635657 955205
rect 537099 952325 635657 952441
rect 529227 952232 535876 952297
rect 2823 908397 2875 909069
rect 3547 908397 3623 909069
rect 2823 783067 3623 908397
rect 2823 782395 2881 783067
rect 3553 782395 3623 783067
rect 2823 739880 3623 782395
rect 2823 739208 2886 739880
rect 3558 739208 3623 739880
rect 2823 696699 3623 739208
rect 2823 696027 2892 696699
rect 3564 696027 3623 696699
rect 2823 653496 3623 696027
rect 2823 652824 2886 653496
rect 3558 652824 3623 653496
rect 2823 610292 3623 652824
rect 2823 609620 2903 610292
rect 3575 609620 3623 610292
rect 2823 567309 3623 609620
rect 2823 566637 2897 567309
rect 3569 566637 3623 567309
rect 2823 524275 3623 566637
rect 2823 523603 2903 524275
rect 3575 523603 3623 524275
rect 2823 396279 3623 523603
rect 2823 395607 2903 396279
rect 3575 395607 3623 396279
rect 2823 353296 3623 395607
rect 2823 352624 2886 353296
rect 3558 352624 3623 353296
rect 2823 310312 3623 352624
rect 2823 309640 2875 310312
rect 3547 309640 3623 310312
rect 2823 267292 3623 309640
rect 2823 266620 2884 267292
rect 3556 266620 3623 267292
rect 2823 224294 3623 266620
rect 2823 223622 2881 224294
rect 3553 223622 3623 224294
rect 2823 181286 3623 223622
rect 4273 950850 18820 951450
rect 4273 803652 5273 950850
rect 4273 799066 4359 803652
rect 5171 799066 5273 803652
rect 4273 793675 5273 799066
rect 4273 789089 4351 793675
rect 5163 789089 5273 793675
rect 4273 233106 5273 789089
rect 6273 949910 19792 950510
rect 6273 459103 7273 949910
rect 633657 949570 635657 952325
rect 616645 948970 635657 949570
rect 615787 948030 632657 948630
rect 6273 454442 6326 459103
rect 7225 454442 7273 459103
rect 6273 449139 7273 454442
rect 6273 444435 6315 449139
rect 7201 444435 7273 449139
rect 6273 238811 7273 444435
rect 6273 233558 6344 238811
rect 7160 234046 7273 238811
rect 8273 947452 22611 947690
rect 8273 945799 9771 947452
rect 10560 947090 22611 947452
rect 10560 945799 12273 947090
rect 8273 910585 12273 945799
rect 8273 910513 8334 910585
rect 12206 910513 12273 910585
rect 8273 764241 12273 910513
rect 8273 763569 8334 764241
rect 12206 763569 12273 764241
rect 8273 720830 12273 763569
rect 8273 720158 8330 720830
rect 12202 720158 12273 720830
rect 8273 677639 12273 720158
rect 8273 676967 8334 677639
rect 12206 676967 12273 677639
rect 8273 634839 12273 676967
rect 8273 634167 8342 634839
rect 12214 634167 12273 634839
rect 8273 591232 12273 634167
rect 8273 590560 8330 591232
rect 12202 590560 12273 591232
rect 8273 548047 12273 590560
rect 8273 547375 8330 548047
rect 12202 547375 12273 548047
rect 8273 504838 12273 547375
rect 8273 504166 8323 504838
rect 12195 504166 12273 504838
rect 8273 416912 12273 504166
rect 8273 412440 8417 416912
rect 12175 412440 12273 416912
rect 8273 406832 12273 412440
rect 8273 402360 8374 406832
rect 12132 402360 12273 406832
rect 8273 377036 12273 402360
rect 8273 376364 8334 377036
rect 12206 376364 12273 377036
rect 8273 333829 12273 376364
rect 8273 333157 8342 333829
rect 12214 333157 12273 333829
rect 8273 290622 12273 333157
rect 8273 289950 8332 290622
rect 12204 289950 12273 290622
rect 8273 247417 12273 289950
rect 8273 246745 8332 247417
rect 12204 246745 12273 247417
rect 8273 240968 12273 246745
rect 8273 234855 8378 240968
rect 12145 236866 12273 240968
rect 13273 946390 23511 946750
rect 13273 944562 14566 946390
rect 15343 946150 23511 946390
rect 15343 944562 17273 946150
rect 625657 945810 629657 945814
rect 612964 945737 629657 945810
rect 612964 945210 625971 945737
rect 13273 911987 17273 944562
rect 612016 944847 624648 944870
rect 612016 944801 624657 944847
rect 612016 944270 622828 944801
rect 13273 911915 13333 911987
rect 17205 911915 17273 911987
rect 13273 888015 17273 911915
rect 13273 883618 13382 888015
rect 17116 883618 17273 888015
rect 13273 878016 17273 883618
rect 13273 873619 13431 878016
rect 17165 873619 17273 878016
rect 13273 765636 17273 873619
rect 13273 764964 13329 765636
rect 17201 764964 17273 765636
rect 13273 722236 17273 764964
rect 13273 721564 13337 722236
rect 17209 721564 17273 722236
rect 13273 679189 17273 721564
rect 13273 678517 13348 679189
rect 17220 678517 17273 679189
rect 13273 636226 17273 678517
rect 13273 635554 13337 636226
rect 17209 635554 17273 636226
rect 13273 592638 17273 635554
rect 13273 591966 13340 592638
rect 17212 591966 17273 592638
rect 13273 549436 17273 591966
rect 13273 548764 13341 549436
rect 17213 548764 17273 549436
rect 13273 506240 17273 548764
rect 13273 505568 13337 506240
rect 17209 505568 17273 506240
rect 13273 378423 17273 505568
rect 13273 377751 13329 378423
rect 17201 377751 17273 378423
rect 13273 335232 17273 377751
rect 13273 334560 13329 335232
rect 17201 334560 17273 335232
rect 13273 292032 17273 334560
rect 13273 291360 13329 292032
rect 17201 291360 17273 292032
rect 13273 248824 17273 291360
rect 13273 248152 13328 248824
rect 17200 248152 17273 248824
rect 13273 240911 17273 248152
rect 13273 237313 13396 240911
rect 17117 237806 17273 240911
rect 620657 943225 622828 944270
rect 624321 943225 624657 944801
rect 620657 907447 624657 943225
rect 620657 906775 620715 907447
rect 624587 906775 624657 907447
rect 620657 883577 624657 906775
rect 620657 879253 620860 883577
rect 624447 879253 624657 883577
rect 620657 873491 624657 879253
rect 620657 869167 620810 873491
rect 624397 869167 624657 873491
rect 620657 729441 624657 869167
rect 620657 728769 620720 729441
rect 624592 728769 624657 729441
rect 620657 684229 624657 728769
rect 620657 683557 620720 684229
rect 624592 683557 624657 684229
rect 620657 639046 624657 683557
rect 620657 638374 620725 639046
rect 624597 638374 624657 639046
rect 620657 593843 624657 638374
rect 620657 593171 620715 593843
rect 624587 593171 624657 593843
rect 620657 548645 624657 593171
rect 620657 547973 620725 548645
rect 624597 547973 624657 548645
rect 620657 503437 624657 547973
rect 620657 502765 620729 503437
rect 624601 502765 624657 503437
rect 620657 459845 624657 502765
rect 620657 459173 620715 459845
rect 624587 459173 624657 459845
rect 620657 371449 624657 459173
rect 620657 370777 620720 371449
rect 624592 370777 624657 371449
rect 620657 326666 624657 370777
rect 620657 325994 620729 326666
rect 624601 325994 624657 326666
rect 620657 281849 624657 325994
rect 620657 281177 620734 281849
rect 624606 281177 624657 281849
rect 620657 242438 624657 281177
rect 620657 239686 620804 242438
rect 611967 239279 620804 239686
rect 624519 239279 624657 242438
rect 611967 239093 624657 239279
rect 625657 943324 625971 945210
rect 627460 943324 629657 945737
rect 625657 908835 629657 943324
rect 625657 908163 625724 908835
rect 629596 908163 629657 908835
rect 625657 730844 629657 908163
rect 625657 730172 625719 730844
rect 629591 730172 629657 730844
rect 625657 685641 629657 730172
rect 625657 684969 625714 685641
rect 629586 684969 629657 685641
rect 625657 640439 629657 684969
rect 625657 639767 625724 640439
rect 629596 639767 629657 640439
rect 625657 595246 629657 639767
rect 625657 594574 625728 595246
rect 629600 594574 629657 595246
rect 625657 550038 629657 594574
rect 625657 549366 625728 550038
rect 629600 549366 629657 550038
rect 625657 504840 629657 549366
rect 625657 504168 625714 504840
rect 629586 504168 629657 504840
rect 625657 461238 629657 504168
rect 625657 460566 625719 461238
rect 629591 460566 629657 461238
rect 625657 435866 629657 460566
rect 625657 431326 625815 435866
rect 629491 431326 629657 435866
rect 625657 425749 629657 431326
rect 625657 421357 625811 425749
rect 629472 421357 629657 425749
rect 625657 372852 629657 421357
rect 625657 372180 625724 372852
rect 629596 372180 629657 372852
rect 625657 328050 629657 372180
rect 625657 327378 625724 328050
rect 629596 327378 629657 328050
rect 625657 283228 629657 327378
rect 625657 282556 625724 283228
rect 629596 282556 629657 283228
rect 625657 242425 629657 282556
rect 611967 239086 624610 239093
rect 625657 238746 625807 242425
rect 612951 238146 625807 238746
rect 17117 237313 23509 237806
rect 13273 237206 23509 237313
rect 12145 236266 22611 236866
rect 625657 236391 625807 238146
rect 629455 238746 629657 242425
rect 630657 479910 632657 948030
rect 630657 475283 630713 479910
rect 632588 475283 632657 479910
rect 630657 469932 632657 475283
rect 630657 465305 630706 469932
rect 632581 465305 632657 469932
rect 630657 242425 632657 465305
rect 629455 238146 629686 238746
rect 629455 236391 629657 238146
rect 625657 236278 629657 236391
rect 12145 234855 12273 236266
rect 630657 235926 630784 242425
rect 615700 235468 630784 235926
rect 632547 235468 632657 242425
rect 615700 235326 632657 235468
rect 630657 235323 632657 235326
rect 633657 794462 635657 948970
rect 633657 789897 633781 794462
rect 635118 789897 635657 794462
rect 633657 784517 635657 789897
rect 633657 779952 633749 784517
rect 635086 779952 635657 784517
rect 633657 391672 635657 779952
rect 633657 387094 633737 391672
rect 635564 387094 635657 391672
rect 633657 381734 635657 387094
rect 633657 377156 633726 381734
rect 635553 377156 635657 381734
rect 630657 235315 632621 235323
rect 633657 234986 635657 377156
rect 8273 234697 12273 234855
rect 616560 234386 635657 234986
rect 7160 233558 19774 234046
rect 6273 233446 19774 233558
rect 6273 233435 7273 233446
rect 620657 233434 624657 233624
rect 4273 232506 18789 233106
rect 4273 217854 5273 232506
rect 6273 231502 7273 231631
rect 6273 227791 6355 231502
rect 7149 227791 7273 231502
rect 6273 220854 7273 227791
rect 8273 231501 12273 231631
rect 8273 227903 8423 231501
rect 12144 227903 12273 231501
rect 8273 224854 12273 227903
rect 13273 231468 17273 231631
rect 13273 227870 13419 231468
rect 17140 229854 17273 231468
rect 620657 230071 620817 233434
rect 624505 230071 624657 233434
rect 17140 227870 144995 229854
rect 13273 226854 144995 227870
rect 620657 227074 624657 230071
rect 143495 225564 144995 226854
rect 143495 225528 372157 225564
rect 8273 223064 141281 224854
rect 143495 224103 159217 225528
rect 159507 224103 189317 225528
rect 189607 224103 219417 225528
rect 219707 224103 249517 225528
rect 249807 224103 279617 225528
rect 279907 224103 309717 225528
rect 310007 224103 339817 225528
rect 340107 224103 369917 225528
rect 370207 224103 372157 225528
rect 143495 224064 372157 224103
rect 383256 223074 624657 227074
rect 625657 233407 629657 233624
rect 625657 230044 625848 233407
rect 629536 230044 629657 233407
rect 8273 223017 372157 223064
rect 8273 221854 174274 223017
rect 139781 221605 174274 221854
rect 174572 221605 204374 223017
rect 204672 221605 234474 223017
rect 234772 221605 264574 223017
rect 264872 221605 294674 223017
rect 294972 221605 324774 223017
rect 325072 221605 354874 223017
rect 355172 221605 372157 223017
rect 139781 221564 372157 221605
rect 6273 220564 137328 220854
rect 6273 220516 372157 220564
rect 6273 219105 160027 220516
rect 160382 219105 190127 220516
rect 190482 219105 220227 220516
rect 220582 219105 250267 220516
rect 250542 219105 280427 220516
rect 280782 219105 310527 220516
rect 310882 219105 340627 220516
rect 340982 219105 370727 220516
rect 371082 219105 372157 220516
rect 6273 219064 372157 219105
rect 6273 218854 137328 219064
rect 138364 218030 357099 218064
rect 138364 217854 175919 218030
rect 4273 216618 175919 217854
rect 176178 216618 206019 218030
rect 206278 216618 236119 218030
rect 236378 216618 266219 218030
rect 4273 216613 266219 216618
rect 266478 216618 296319 218030
rect 296578 216618 326419 218030
rect 326678 216618 356519 218030
rect 356778 216618 357099 218030
rect 266478 216613 357099 216618
rect 4273 216564 357099 216613
rect 4273 215854 140993 216564
rect 383256 215564 387256 223074
rect 625657 221074 629657 230044
rect 158192 215526 387256 215564
rect 158192 214096 158407 215526
rect 158695 214096 188507 215526
rect 188795 214096 218607 215526
rect 218895 214096 248797 215526
rect 249075 214096 278807 215526
rect 279045 214096 308907 215526
rect 309195 214096 339007 215526
rect 339295 214096 369107 215526
rect 369395 214096 387256 215526
rect 158192 214064 387256 214096
rect 389353 217074 629657 221074
rect 630657 233461 632657 233624
rect 630657 230058 630865 233461
rect 632506 230058 632657 233461
rect 2823 180614 2887 181286
rect 3561 180614 3623 181286
rect 2823 103255 3623 180614
rect 4223 213801 5023 213859
rect 4223 211917 4272 213801
rect 4958 211917 5023 213801
rect 4223 204225 5023 211917
rect 4223 203553 4289 204225
rect 4961 203553 5023 204225
rect 4223 161066 5023 203553
rect 5623 213781 6423 213859
rect 5623 211897 5673 213781
rect 6359 211897 6423 213781
rect 5623 205628 6423 211897
rect 5623 204956 5686 205628
rect 6358 204956 6423 205628
rect 5623 162450 6423 204956
rect 5623 161736 5662 162450
rect 6387 161736 6423 162450
rect 5623 161637 6423 161736
rect 7506 213365 145906 213604
rect 7506 207012 110403 213365
rect 116528 207012 130322 213365
rect 136447 207012 145906 213365
rect 389353 213064 393353 217074
rect 630657 213074 632657 230058
rect 173291 213029 393353 213064
rect 173291 211601 173451 213029
rect 173725 211601 203551 213029
rect 203825 211601 233701 213029
rect 233975 212949 293851 213029
rect 233975 211601 263691 212949
rect 263965 211601 293851 212949
rect 294125 211601 323951 213029
rect 324225 211601 354051 213029
rect 354325 211601 393353 213029
rect 173291 211564 393353 211601
rect 395119 210564 632657 213074
rect 159813 210533 632657 210564
rect 159813 209096 160095 210533
rect 160347 209096 190195 210533
rect 190447 209096 220295 210533
rect 220547 209096 250275 210533
rect 250527 209096 280495 210533
rect 280747 209096 310595 210533
rect 310847 209096 340695 210533
rect 340947 209096 370795 210533
rect 371047 210074 632657 210533
rect 371047 209096 398119 210074
rect 159813 209064 398119 209096
rect 633657 209074 635657 234386
rect 401055 208064 635657 209074
rect 7506 206604 145906 207012
rect 7506 200066 12506 206604
rect 138906 205564 145906 206604
rect 174811 208037 635657 208064
rect 174811 206605 175100 208037
rect 175364 206605 205200 208037
rect 205464 206605 235360 208037
rect 235624 206605 265350 208037
rect 265614 206605 295500 208037
rect 295764 206605 325600 208037
rect 325864 206605 355700 208037
rect 355964 206605 635657 208037
rect 174811 206564 635657 206605
rect 401055 206074 635657 206564
rect 636467 906033 637267 955958
rect 636467 905361 636532 906033
rect 637204 905361 637267 906033
rect 636467 728033 637267 905361
rect 636467 727361 636525 728033
rect 637197 727361 637267 728033
rect 636467 682843 637267 727361
rect 636467 682171 636530 682843
rect 637202 682171 637267 682843
rect 636467 637635 637267 682171
rect 636467 636963 636542 637635
rect 637214 636963 637267 637635
rect 636467 592442 637267 636963
rect 636467 591770 636532 592442
rect 637204 591770 637267 592442
rect 636467 547239 637267 591770
rect 636467 546567 636523 547239
rect 637195 546567 637267 547239
rect 636467 502043 637267 546567
rect 636467 501371 636529 502043
rect 637201 501371 637267 502043
rect 636467 458440 637267 501371
rect 636467 457768 636530 458440
rect 637202 457768 637267 458440
rect 636467 370039 637267 457768
rect 636467 369367 636529 370039
rect 637201 369367 637267 370039
rect 636467 325237 637267 369367
rect 636467 324565 636529 325237
rect 637201 324565 637267 325237
rect 636467 280444 637267 324565
rect 636467 279772 636524 280444
rect 637196 279772 637267 280444
rect 636467 235036 637267 279772
rect 636467 234364 636532 235036
rect 637204 234364 637267 235036
rect 138906 205533 368771 205564
rect 138906 204093 157566 205533
rect 157877 204093 187666 205533
rect 187977 204093 217766 205533
rect 218077 204093 247816 205533
rect 248127 204093 278046 205533
rect 278307 204093 308066 205533
rect 308377 204093 338166 205533
rect 338477 204093 368266 205533
rect 368577 204093 368771 205533
rect 633146 204351 633946 204430
rect 138906 204064 368771 204093
rect 630491 204214 631291 204293
rect 109924 200162 116943 200253
rect 109924 200066 110021 200162
rect 7506 199746 14895 200066
rect 104047 199746 110021 200066
rect 7506 190066 12506 199746
rect 109924 199698 110021 199746
rect 116816 200066 116943 200162
rect 116816 199746 116961 200066
rect 116816 199698 116943 199746
rect 109924 199612 116943 199698
rect 119975 195272 126969 195687
rect 138906 195370 145906 204064
rect 172379 203026 394268 203064
rect 172379 201601 172628 203026
rect 172929 201601 202728 203026
rect 203029 201601 232828 203026
rect 233129 201601 262928 203026
rect 263229 201601 292918 203026
rect 293219 201601 323128 203026
rect 323429 201601 353228 203026
rect 353529 202845 394268 203026
rect 353529 201601 387985 202845
rect 172379 201564 387985 201601
rect 387723 201297 387985 201564
rect 393910 201297 394268 202845
rect 387723 201064 394268 201297
rect 630491 202234 630549 204214
rect 631216 202234 631291 204214
rect 387741 201053 394235 201064
rect 630491 198246 631291 202234
rect 633146 202289 633219 204351
rect 633869 202289 633946 204351
rect 633146 200815 633946 202289
rect 633146 200015 635867 200815
rect 630491 197446 634467 198246
rect 119933 195145 126973 195272
rect 119933 195066 119991 195145
rect 104047 194746 119991 195066
rect 119933 194628 119991 194746
rect 126852 195066 126973 195145
rect 138906 195247 632476 195370
rect 138906 195168 629587 195247
rect 126852 194746 126975 195066
rect 126852 194628 126973 194746
rect 119933 194559 126973 194628
rect 109924 190162 116943 190253
rect 109924 190066 110021 190162
rect 7506 189746 14884 190066
rect 104047 189746 110021 190066
rect 7506 180066 12506 189746
rect 109924 189698 110021 189746
rect 116816 189698 116943 190162
rect 109924 189612 116943 189698
rect 119975 188370 126969 194559
rect 138906 190557 608763 195168
rect 613356 193669 629587 195168
rect 632313 193669 632476 195247
rect 613356 193545 632476 193669
rect 613356 190557 613608 193545
rect 138906 190370 613608 190557
rect 633667 191042 634467 197446
rect 633667 190370 633732 191042
rect 634404 190370 634467 191042
rect 138906 190347 145906 190370
rect 119975 188265 607566 188370
rect 119975 185066 120133 188265
rect 104047 184746 120133 185066
rect 119975 183580 120133 184746
rect 126688 188234 607566 188265
rect 126688 183580 139135 188234
rect 119975 183549 139135 183580
rect 145690 188229 607566 188234
rect 145690 188204 602772 188229
rect 145690 183649 388000 188204
rect 393895 183649 602772 188204
rect 145690 183618 602772 183649
rect 607365 183618 607566 188229
rect 145690 183549 607566 183618
rect 119975 183370 607566 183549
rect 109924 180162 116943 180253
rect 109924 180066 110021 180162
rect 7506 179746 14884 180066
rect 104047 179746 110021 180066
rect 7506 170066 12506 179746
rect 109924 179698 110021 179746
rect 116816 179698 116943 180162
rect 109924 179612 116943 179698
rect 129802 176657 136933 176729
rect 129802 176107 130009 176657
rect 136855 176512 136933 176657
rect 608556 176601 613582 176652
rect 608556 176512 608613 176601
rect 136855 176192 153297 176512
rect 600378 176192 608613 176512
rect 136855 176107 136933 176192
rect 129802 176012 136933 176107
rect 608556 176153 608613 176192
rect 613500 176512 613582 176601
rect 613500 176192 613584 176512
rect 613500 176153 613582 176192
rect 608556 176088 613582 176153
rect 119938 175168 126930 175245
rect 119938 175066 120020 175168
rect 104047 174746 120020 175066
rect 119938 174631 120020 174746
rect 126822 175066 126930 175168
rect 126822 174746 126933 175066
rect 126822 174631 126930 174746
rect 119938 174555 126930 174631
rect 109924 170162 116943 170253
rect 109924 170066 110021 170162
rect 7506 169746 14884 170066
rect 104005 169746 110021 170066
rect 4223 160352 4258 161066
rect 4983 160352 5023 161066
rect 4223 160094 5023 160352
rect 7506 160066 12506 169746
rect 109924 169698 110021 169746
rect 116816 169698 116943 170162
rect 109924 169612 116943 169698
rect 119938 165168 126930 165245
rect 119938 165066 120020 165168
rect 104047 164746 120020 165066
rect 119938 164631 120020 164746
rect 126822 165066 126930 165168
rect 126822 164746 126968 165066
rect 126822 164631 126930 164746
rect 119938 164555 126930 164631
rect 138925 163654 145941 163717
rect 138925 163065 138995 163654
rect 145878 163512 145941 163654
rect 602550 163571 607549 163646
rect 602550 163512 602628 163571
rect 145878 163192 153297 163512
rect 600421 163192 602628 163512
rect 145878 163065 145941 163192
rect 602550 163148 602628 163192
rect 607445 163512 607549 163571
rect 607445 163192 607587 163512
rect 607445 163148 607549 163192
rect 602550 163065 607549 163148
rect 138925 163012 145941 163065
rect 109924 160162 116943 160253
rect 109924 160066 110021 160162
rect 7506 159746 14884 160066
rect 104047 159746 110021 160066
rect 7506 150066 12506 159746
rect 109924 159698 110021 159746
rect 116816 159698 116943 160162
rect 109924 159612 116943 159698
rect 119938 155168 126930 155245
rect 119938 155066 120020 155168
rect 104006 154746 120020 155066
rect 119938 154631 120020 154746
rect 126822 155066 126930 155168
rect 126822 154746 126947 155066
rect 126822 154631 126930 154746
rect 119938 154555 126930 154631
rect 129802 150657 136933 150729
rect 109924 150162 116943 150253
rect 109924 150066 110021 150162
rect 7506 149746 14884 150066
rect 104047 149746 110021 150066
rect 7506 140066 12506 149746
rect 109924 149698 110021 149746
rect 116816 150066 116943 150162
rect 129802 150107 130009 150657
rect 136855 150512 136933 150657
rect 608556 150601 613582 150652
rect 608556 150512 608613 150601
rect 136855 150192 153297 150512
rect 600420 150192 608613 150512
rect 136855 150107 136933 150192
rect 116816 149746 116951 150066
rect 129802 150012 136933 150107
rect 608556 150153 608613 150192
rect 613500 150512 613582 150601
rect 613500 150192 613584 150512
rect 613500 150153 613582 150192
rect 608556 150088 613582 150153
rect 116816 149698 116943 149746
rect 109924 149612 116943 149698
rect 633667 145639 634467 190370
rect 119938 145168 126930 145245
rect 119938 145066 120020 145168
rect 104017 144746 120020 145066
rect 119938 144631 120020 144746
rect 126822 145066 126930 145168
rect 126822 144746 126958 145066
rect 633667 144967 633731 145639
rect 634403 144967 634467 145639
rect 126822 144631 126930 144746
rect 119938 144555 126930 144631
rect 109924 140162 116943 140253
rect 109924 140066 110021 140162
rect 7506 139746 14884 140066
rect 104047 139746 110021 140066
rect 7506 130066 12506 139746
rect 109924 139698 110021 139746
rect 116816 139698 116943 140162
rect 109924 139612 116943 139698
rect 138925 137654 145941 137717
rect 138925 137065 138995 137654
rect 145878 137512 145941 137654
rect 602550 137571 607549 137646
rect 602550 137512 602628 137571
rect 145878 137192 153327 137512
rect 600392 137192 602628 137512
rect 145878 137065 145941 137192
rect 602550 137148 602628 137192
rect 607445 137512 607549 137571
rect 607445 137192 607573 137512
rect 607445 137148 607549 137192
rect 602550 137065 607549 137148
rect 138925 137012 145941 137065
rect 119938 135168 126930 135245
rect 119938 135066 120020 135168
rect 104047 134746 120020 135066
rect 119938 134631 120020 134746
rect 126822 135066 126930 135168
rect 126822 134746 126937 135066
rect 126822 134631 126930 134746
rect 119938 134555 126930 134631
rect 109924 130162 116943 130253
rect 109924 130066 110021 130162
rect 7506 129746 14884 130066
rect 104047 129746 110021 130066
rect 7506 120066 12506 129746
rect 109924 129698 110021 129746
rect 116816 130066 116943 130162
rect 116816 129746 116951 130066
rect 116816 129698 116943 129746
rect 109924 129612 116943 129698
rect 119938 125168 126930 125245
rect 119938 125066 120020 125168
rect 104047 124746 120020 125066
rect 119938 124631 120020 124746
rect 126822 125066 126930 125168
rect 126822 124746 126979 125066
rect 126822 124631 126930 124746
rect 119938 124555 126930 124631
rect 129802 124657 136933 124729
rect 129802 124107 130009 124657
rect 136855 124512 136933 124657
rect 608556 124601 613582 124652
rect 608556 124512 608613 124601
rect 136855 124192 153297 124512
rect 600421 124192 608613 124512
rect 136855 124107 136933 124192
rect 129802 124012 136933 124107
rect 608556 124153 608613 124192
rect 613500 124512 613582 124601
rect 613500 124192 613612 124512
rect 613500 124153 613582 124192
rect 608556 124088 613582 124153
rect 109924 120162 116943 120253
rect 109924 120066 110021 120162
rect 7506 119746 14884 120066
rect 104047 119746 110021 120066
rect 7506 110066 12506 119746
rect 109924 119698 110021 119746
rect 116816 119698 116943 120162
rect 109924 119612 116943 119698
rect 119938 115168 126930 115245
rect 119938 115066 120020 115168
rect 104047 114746 120020 115066
rect 119938 114631 120020 114746
rect 126822 115066 126930 115168
rect 126822 114746 126958 115066
rect 126822 114631 126930 114746
rect 119938 114555 126930 114631
rect 138925 111654 145941 111717
rect 138925 111512 138995 111654
rect 138912 111192 138995 111512
rect 138925 111065 138995 111192
rect 145878 111512 145941 111654
rect 602550 111571 607549 111646
rect 602550 111512 602628 111571
rect 145878 111192 153297 111512
rect 600421 111192 602628 111512
rect 145878 111065 145941 111192
rect 602550 111148 602628 111192
rect 607445 111148 607549 111571
rect 602550 111065 607549 111148
rect 138925 111012 145941 111065
rect 109924 110162 116943 110253
rect 109924 110066 110021 110162
rect 7506 109746 14884 110066
rect 104047 109746 110021 110066
rect 7506 103255 12506 109746
rect 109924 109698 110021 109746
rect 116816 110066 116943 110162
rect 116816 109746 116972 110066
rect 116816 109698 116943 109746
rect 109924 109612 116943 109698
rect 119938 105168 126930 105245
rect 119938 105066 120020 105168
rect 104047 104746 120020 105066
rect 119938 104631 120020 104746
rect 126822 105066 126930 105168
rect 126822 104746 126947 105066
rect 126822 104631 126930 104746
rect 119938 104555 126930 104631
rect 2823 102455 12506 103255
rect 4106 100066 12506 102455
rect 109924 100162 116943 100253
rect 109924 100066 110021 100162
rect 4106 99746 14884 100066
rect 104047 99746 110021 100066
rect 4106 93783 12506 99746
rect 109924 99698 110021 99746
rect 116816 99698 116943 100162
rect 109924 99612 116943 99698
rect 633667 100241 634467 144967
rect 633667 99569 633728 100241
rect 634400 99569 634467 100241
rect 633667 99320 634467 99569
rect 635067 192443 635867 200015
rect 635067 191771 635130 192443
rect 635802 191771 635867 192443
rect 635067 147047 635867 191771
rect 635067 146375 635130 147047
rect 635802 146375 635867 147047
rect 635067 101637 635867 146375
rect 635067 100965 635134 101637
rect 635806 100965 635867 101637
rect 635067 99320 635867 100965
rect 636467 189642 637267 234364
rect 636467 188970 636525 189642
rect 637197 188970 637267 189642
rect 636467 144235 637267 188970
rect 636467 143563 636523 144235
rect 637195 143563 637267 144235
rect 636467 98843 637267 143563
rect 129802 98657 136933 98729
rect 129802 98107 130009 98657
rect 136855 98512 136933 98657
rect 608556 98601 613582 98652
rect 608556 98512 608613 98601
rect 136855 98192 153344 98512
rect 600421 98192 608613 98512
rect 136855 98107 136933 98192
rect 129802 98012 136933 98107
rect 608556 98153 608613 98192
rect 613500 98512 613582 98601
rect 613500 98192 613584 98512
rect 613500 98153 613582 98192
rect 608556 98088 613582 98153
rect 636467 98171 636533 98843
rect 637205 98171 637267 98843
rect 636467 96386 637267 98171
rect 637867 904643 638667 957455
rect 637867 903971 637932 904643
rect 638604 903971 638667 904643
rect 637867 726647 638667 903971
rect 637867 725975 637926 726647
rect 638598 725975 638667 726647
rect 637867 681433 638667 725975
rect 637867 680761 637931 681433
rect 638603 680761 638667 681433
rect 637867 636237 638667 680761
rect 637867 635565 637921 636237
rect 638593 635565 638667 636237
rect 637867 591039 638667 635565
rect 637867 590367 637926 591039
rect 638598 590367 638667 591039
rect 637867 545845 638667 590367
rect 637867 545173 637935 545845
rect 638607 545173 638667 545845
rect 637867 500647 638667 545173
rect 637867 499975 637930 500647
rect 638602 499975 638667 500647
rect 637867 457041 638667 499975
rect 637867 456369 637928 457041
rect 638600 456369 638667 457041
rect 637867 368635 638667 456369
rect 637867 367963 637929 368635
rect 638601 367963 638667 368635
rect 637867 323860 638667 367963
rect 637867 323188 637924 323860
rect 638596 323188 638667 323860
rect 637867 279039 638667 323188
rect 637867 278367 637915 279039
rect 638587 278367 638667 279039
rect 637867 233650 638667 278367
rect 637867 232978 637933 233650
rect 638605 232978 638667 233650
rect 637867 196101 638667 232978
rect 637867 193295 637917 196101
rect 638627 193295 638667 196101
rect 637867 188248 638667 193295
rect 637867 187576 637919 188248
rect 638591 187576 638667 188248
rect 637867 142842 638667 187576
rect 637867 142170 637930 142842
rect 638602 142170 638667 142842
rect 637867 97439 638667 142170
rect 637867 96767 637931 97439
rect 638603 96767 638667 97439
rect 637867 96386 638667 96767
rect 119938 95168 126930 95245
rect 119938 95066 120020 95168
rect 103996 94746 120020 95066
rect 119938 94631 120020 94746
rect 126822 95066 126930 95168
rect 126822 94746 126958 95066
rect 126822 94631 126930 94746
rect 119938 94555 126930 94631
rect 4106 90066 9106 93783
rect 109924 90162 116943 90253
rect 109924 90066 110021 90162
rect 4106 89746 14884 90066
rect 104047 89746 110021 90066
rect 4106 80066 9106 89746
rect 109924 89698 110021 89746
rect 116816 90066 116943 90162
rect 116816 89746 116983 90066
rect 116816 89698 116943 89746
rect 109924 89612 116943 89698
rect 138925 85654 145941 85717
rect 138925 85512 138995 85654
rect 119938 85168 126930 85245
rect 138878 85192 138995 85512
rect 119938 85066 120020 85168
rect 104047 84746 120020 85066
rect 119938 84631 120020 84746
rect 126822 85066 126930 85168
rect 126822 84746 126958 85066
rect 138925 85065 138995 85192
rect 145878 85512 145941 85654
rect 602550 85571 607549 85646
rect 602550 85512 602628 85571
rect 145878 85192 153327 85512
rect 600421 85192 602628 85512
rect 145878 85065 145941 85192
rect 602550 85148 602628 85192
rect 607445 85512 607549 85571
rect 607445 85192 607593 85512
rect 607445 85148 607549 85192
rect 602550 85065 607549 85148
rect 138925 85012 145941 85065
rect 126822 84631 126930 84746
rect 119938 84555 126930 84631
rect 109924 80162 116943 80253
rect 109924 80066 110021 80162
rect 4106 79746 14854 80066
rect 104047 79746 110021 80066
rect 4106 70066 9106 79746
rect 109924 79698 110021 79746
rect 116816 79698 116943 80162
rect 109924 79612 116943 79698
rect 628513 75779 631513 75781
rect 614103 75734 635513 75779
rect 119938 75168 126930 75245
rect 119938 75066 120020 75168
rect 104047 74746 120020 75066
rect 119938 74631 120020 74746
rect 126822 75066 126930 75168
rect 126822 74746 126958 75066
rect 126822 74631 126930 74746
rect 614103 74690 614156 75734
rect 615367 74690 635513 75734
rect 614103 74653 635513 74690
rect 628513 74650 631513 74653
rect 119938 74555 126930 74631
rect 129802 72657 136933 72729
rect 129802 72107 130009 72657
rect 136855 72512 136933 72657
rect 608556 72601 613582 72652
rect 608556 72512 608613 72601
rect 136855 72192 153297 72512
rect 600395 72192 608613 72512
rect 136855 72107 136933 72192
rect 129802 72012 136933 72107
rect 608556 72153 608613 72192
rect 613500 72512 613582 72601
rect 613500 72192 613584 72512
rect 613500 72153 613582 72192
rect 608556 72088 613582 72153
rect 109924 70162 116943 70253
rect 109924 70066 110021 70162
rect 4106 69746 14854 70066
rect 104047 69746 110021 70066
rect 4106 60066 9106 69746
rect 109924 69698 110021 69746
rect 116816 69698 116943 70162
rect 109924 69612 116943 69698
rect 608537 65265 613556 65312
rect 119938 65168 126930 65245
rect 119938 65066 120020 65168
rect 104027 64746 120020 65066
rect 119938 64631 120020 64746
rect 126822 65066 126930 65168
rect 126822 64746 126947 65066
rect 126822 64631 126930 64746
rect 119938 64555 126930 64631
rect 608537 64636 608612 65265
rect 613504 65160 613556 65265
rect 613504 65118 624709 65160
rect 613504 64798 622897 65118
rect 624672 64798 624709 65118
rect 613504 64760 624709 64798
rect 613504 64636 613556 64760
rect 608537 64599 613556 64636
rect 614106 63098 631513 63171
rect 614106 61750 614165 63098
rect 615335 61750 631513 63098
rect 614106 61685 631513 61750
rect 109924 60162 116943 60253
rect 109924 60066 110021 60162
rect 4106 59746 14854 60066
rect 104047 59746 110021 60066
rect 4106 50066 9106 59746
rect 109924 59698 110021 59746
rect 116816 60066 116943 60162
rect 116816 59746 116983 60066
rect 116816 59698 116943 59746
rect 109924 59612 116943 59698
rect 138925 59654 145941 59717
rect 138925 59065 138995 59654
rect 145878 59512 145941 59654
rect 602550 59571 607549 59646
rect 602550 59512 602628 59571
rect 145878 59192 153302 59512
rect 600406 59192 602628 59512
rect 145878 59065 145941 59192
rect 602550 59148 602628 59192
rect 607445 59148 607549 59571
rect 602550 59065 607549 59148
rect 138925 59012 145941 59065
rect 119938 55168 126930 55245
rect 119938 55066 120020 55168
rect 104047 54746 120020 55066
rect 119938 54631 120020 54746
rect 126822 55066 126930 55168
rect 126822 54746 126979 55066
rect 126822 54631 126930 54746
rect 119938 54555 126930 54631
rect 109924 50162 116943 50253
rect 109924 50066 110021 50162
rect 4106 49746 14854 50066
rect 103996 49746 110021 50066
rect 4106 43927 9106 49746
rect 109924 49698 110021 49746
rect 116816 49698 116943 50162
rect 109924 49612 116943 49698
rect 608557 47558 613537 47628
rect 608557 47498 608618 47558
rect 601533 47418 608618 47498
rect 601528 47178 608618 47418
rect 129802 46657 136933 46729
rect 129802 46107 130009 46657
rect 136855 46512 136933 46657
rect 601528 46512 601848 47178
rect 608557 47085 608618 47178
rect 613452 47498 613537 47558
rect 613452 47178 619487 47498
rect 613452 47085 613537 47178
rect 608557 47039 613537 47085
rect 136855 46192 153355 46512
rect 600421 46192 601848 46512
rect 602565 46757 607545 46812
rect 602565 46284 602636 46757
rect 607470 46682 607545 46757
rect 607470 46362 619530 46682
rect 607470 46284 607545 46362
rect 602565 46223 607545 46284
rect 136855 46107 136933 46192
rect 129802 46012 136933 46107
rect 608567 45911 613547 45972
rect 608567 45438 608633 45911
rect 613467 45866 613547 45911
rect 613467 45546 619512 45866
rect 613467 45438 613547 45546
rect 608567 45383 613547 45438
rect 119938 45168 126930 45245
rect 119938 45066 120020 45168
rect 103967 44746 120020 45066
rect 119938 44631 120020 44746
rect 126822 45066 126930 45168
rect 602560 45120 607540 45171
rect 126822 44746 126933 45066
rect 126822 44631 126930 44746
rect 119938 44555 126930 44631
rect 602560 44647 602600 45120
rect 607434 45050 607540 45120
rect 607434 44730 619487 45050
rect 607434 44647 607540 44730
rect 602560 44582 607540 44647
rect 608552 44256 613571 44314
rect 608552 44234 608607 44256
rect 4106 39598 4302 43927
rect 8940 40066 9106 43927
rect 608551 43914 608607 44234
rect 608552 43861 608607 43914
rect 613498 44234 613571 44256
rect 613498 43914 619487 44234
rect 613498 43861 613571 43914
rect 608552 43813 613571 43861
rect 109924 40162 116943 40253
rect 109924 40066 110021 40162
rect 8940 39746 14854 40066
rect 103764 39746 110021 40066
rect 8940 39598 9106 39746
rect 109924 39698 110021 39746
rect 116816 40066 116943 40162
rect 116816 39746 116988 40066
rect 116816 39698 116943 39746
rect 109924 39612 116943 39698
rect 4106 33967 9106 39598
rect 119938 35168 126930 35245
rect 119938 35066 120020 35168
rect 103906 34746 120020 35066
rect 119938 34631 120020 34746
rect 126822 35066 126930 35168
rect 126822 34746 126933 35066
rect 126822 34631 126930 34746
rect 119938 34555 126930 34631
rect 4106 29638 4280 33967
rect 8918 30314 9106 33967
rect 138925 33654 145941 33717
rect 138925 33065 138995 33654
rect 145878 33512 145941 33654
rect 602565 33615 607553 33681
rect 602565 33512 602623 33615
rect 145878 33192 153446 33512
rect 600415 33192 602623 33512
rect 145878 33065 145941 33192
rect 138925 33012 145941 33065
rect 602565 33085 602623 33192
rect 607495 33512 607553 33615
rect 607495 33192 607560 33512
rect 607495 33085 607553 33192
rect 602565 33039 607553 33085
rect 8917 30066 9106 30314
rect 109924 30162 116943 30253
rect 109924 30066 110021 30162
rect 8917 29746 14854 30066
rect 104047 29746 110021 30066
rect 8917 29638 9106 29746
rect 4106 20066 9106 29638
rect 109924 29698 110021 29746
rect 116816 29698 116943 30162
rect 109924 29612 116943 29698
rect 129908 29832 136938 29895
rect 129908 29243 129997 29832
rect 136890 29708 136938 29832
rect 136890 29388 149780 29708
rect 136890 29243 136938 29388
rect 129908 29189 136938 29243
rect 119814 26804 145999 26947
rect 119814 26772 139167 26804
rect 119814 25066 120212 26772
rect 103886 24746 120212 25066
rect 119814 22141 120212 24746
rect 126733 22173 139167 26772
rect 145688 22173 145999 26804
rect 126733 22141 145999 22173
rect 119814 21947 145999 22141
rect 109924 20162 116943 20253
rect 109924 20066 110021 20162
rect 4106 19746 14854 20066
rect 104021 19746 110021 20066
rect 4106 14415 9106 19746
rect 109924 19698 110021 19746
rect 116816 19698 116943 20162
rect 109924 19612 116943 19698
rect 140999 16289 145999 21947
rect 149460 20512 149780 29388
rect 608551 20655 613551 20812
rect 608551 20512 608661 20655
rect 149460 20192 153471 20512
rect 600421 20192 608661 20512
rect 104033 16287 145999 16289
rect 103984 16262 145999 16287
rect 103984 15523 104025 16262
rect 104608 15523 145999 16262
rect 103984 15490 145999 15523
rect 104033 15489 145999 15490
rect 140999 15015 145999 15489
rect 602560 18529 607560 18653
rect 602560 15015 602693 18529
rect 140999 14832 602693 15015
rect 131993 14415 136993 14418
rect 4106 14272 136993 14415
rect 4106 13315 110144 14272
rect 4106 12252 105051 13315
rect 105711 12252 110144 13315
rect 4106 9641 110144 12252
rect 116665 14174 136993 14272
rect 116665 9641 130166 14174
rect 4106 9543 130166 9641
rect 136687 9543 136993 14174
rect 140999 10234 202782 14832
rect 207285 14800 602693 14832
rect 207285 10234 212877 14800
rect 140999 10202 212877 10234
rect 217380 14168 602693 14800
rect 607423 14168 607560 18529
rect 217380 10202 607560 14168
rect 140999 10015 607560 10202
rect 608551 16294 608661 20192
rect 613391 16294 613551 20655
rect 4106 9415 136993 9543
rect 131993 8415 136993 9415
rect 608551 8415 613551 16294
rect 131993 3415 613551 8415
rect 628513 11787 631513 61685
rect 628513 7973 628597 11787
rect 631428 7973 631513 11787
rect 628513 7887 631513 7973
rect 632513 6588 635513 74653
rect 632513 2815 632642 6588
rect 635402 2815 635513 6588
rect 632513 2669 635513 2815
<< labels >>
flabel metal5 145438 217320 145438 217320 0 FreeSans 8000 0 0 0 VSSA2
flabel metal5 144640 219774 144640 219774 0 FreeSans 8000 0 0 0 VDDA2
flabel metal5 144395 222474 144395 222474 0 FreeSans 8000 0 0 0 VSSD2
flabel metal5 146359 224867 146359 224867 0 FreeSans 8000 0 0 0 VCCD2
flabel metal5 147893 204740 147893 204740 0 FreeSans 8000 0 0 0 VCCD
flabel metal5 379355 202224 379355 202224 0 FreeSans 8000 0 0 0 VSSD
flabel metal5 379539 207256 379539 207256 0 FreeSans 8000 0 0 0 VSSA1
flabel metal5 379232 209895 379232 209895 0 FreeSans 8000 0 0 0 VDDA1
flabel metal5 378925 212288 378925 212288 0 FreeSans 8000 0 0 0 VSSD1
flabel metal5 378557 214804 378557 214804 0 FreeSans 8000 0 0 0 VCCD1
<< end >>
