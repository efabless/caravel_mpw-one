magic
tech sky130A
magscale 1 2
timestamp 1624271966
<< viali >>
rect 1961 1377 1995 1411
<< metal1 >>
rect 0 2746 2392 2768
rect 0 2694 742 2746
rect 794 2694 806 2746
rect 858 2694 1542 2746
rect 1594 2694 1606 2746
rect 1658 2694 2392 2746
rect 0 2672 2392 2694
rect 0 2202 2392 2224
rect 0 2150 342 2202
rect 394 2150 406 2202
rect 458 2150 1142 2202
rect 1194 2150 1206 2202
rect 1258 2150 1942 2202
rect 1994 2150 2006 2202
rect 2058 2150 2392 2202
rect 0 2128 2392 2150
rect 0 1658 2392 1680
rect 0 1606 742 1658
rect 794 1606 806 1658
rect 858 1606 1542 1658
rect 1594 1606 1606 1658
rect 1658 1606 2392 1658
rect 0 1584 2392 1606
rect 1394 1368 1400 1420
rect 1452 1408 1458 1420
rect 1949 1411 2007 1417
rect 1949 1408 1961 1411
rect 1452 1380 1961 1408
rect 1452 1368 1458 1380
rect 1949 1377 1961 1380
rect 1995 1377 2007 1411
rect 1949 1371 2007 1377
rect 0 1114 2392 1136
rect 0 1062 342 1114
rect 394 1062 406 1114
rect 458 1062 1142 1114
rect 1194 1062 1206 1114
rect 1258 1062 1942 1114
rect 1994 1062 2006 1114
rect 2058 1062 2392 1114
rect 0 1040 2392 1062
rect 0 570 2392 592
rect 0 518 742 570
rect 794 518 806 570
rect 858 518 1542 570
rect 1594 518 1606 570
rect 1658 518 2392 570
rect 0 496 2392 518
rect 0 26 2392 48
rect 0 -26 342 26
rect 394 -26 406 26
rect 458 -26 1142 26
rect 1194 -26 1206 26
rect 1258 -26 1942 26
rect 1994 -26 2006 26
rect 2058 -26 2392 26
rect 0 -48 2392 -26
<< via1 >>
rect 742 2694 794 2746
rect 806 2694 858 2746
rect 1542 2694 1594 2746
rect 1606 2694 1658 2746
rect 342 2150 394 2202
rect 406 2150 458 2202
rect 1142 2150 1194 2202
rect 1206 2150 1258 2202
rect 1942 2150 1994 2202
rect 2006 2150 2058 2202
rect 742 1606 794 1658
rect 806 1606 858 1658
rect 1542 1606 1594 1658
rect 1606 1606 1658 1658
rect 1400 1368 1452 1420
rect 342 1062 394 1114
rect 406 1062 458 1114
rect 1142 1062 1194 1114
rect 1206 1062 1258 1114
rect 1942 1062 1994 1114
rect 2006 1062 2058 1114
rect 742 518 794 570
rect 806 518 858 570
rect 1542 518 1594 570
rect 1606 518 1658 570
rect 342 -26 394 26
rect 406 -26 458 26
rect 1142 -26 1194 26
rect 1206 -26 1258 26
rect 1942 -26 1994 26
rect 2006 -26 2058 26
<< metal2 >>
rect 732 2748 868 2768
rect 788 2746 812 2748
rect 794 2694 806 2746
rect 788 2692 812 2694
rect 732 2672 868 2692
rect 1532 2748 1668 2768
rect 1588 2746 1612 2748
rect 1594 2694 1606 2746
rect 1588 2692 1612 2694
rect 1532 2672 1668 2692
rect 332 2204 468 2224
rect 388 2202 412 2204
rect 394 2150 406 2202
rect 388 2148 412 2150
rect 332 2128 468 2148
rect 1132 2204 1268 2224
rect 1188 2202 1212 2204
rect 1194 2150 1206 2202
rect 1188 2148 1212 2150
rect 1132 2128 1268 2148
rect 1932 2204 2068 2224
rect 1988 2202 2012 2204
rect 1994 2150 2006 2202
rect 1988 2148 2012 2150
rect 1932 2128 2068 2148
rect 732 1660 868 1680
rect 788 1658 812 1660
rect 794 1606 806 1658
rect 788 1604 812 1606
rect 732 1584 868 1604
rect 1532 1660 1668 1680
rect 1588 1658 1612 1660
rect 1594 1606 1606 1658
rect 1588 1604 1612 1606
rect 1532 1584 1668 1604
rect 1398 1456 1454 1465
rect 1398 1391 1400 1400
rect 1452 1391 1454 1400
rect 1400 1362 1452 1368
rect 332 1116 468 1136
rect 388 1114 412 1116
rect 394 1062 406 1114
rect 388 1060 412 1062
rect 332 1040 468 1060
rect 1132 1116 1268 1136
rect 1188 1114 1212 1116
rect 1194 1062 1206 1114
rect 1188 1060 1212 1062
rect 1132 1040 1268 1060
rect 1932 1116 2068 1136
rect 1988 1114 2012 1116
rect 1994 1062 2006 1114
rect 1988 1060 2012 1062
rect 1932 1040 2068 1060
rect 732 572 868 592
rect 788 570 812 572
rect 794 518 806 570
rect 788 516 812 518
rect 732 496 868 516
rect 1532 572 1668 592
rect 1588 570 1612 572
rect 1594 518 1606 570
rect 1588 516 1612 518
rect 1532 496 1668 516
rect 332 28 468 48
rect 388 26 412 28
rect 394 -26 406 26
rect 388 -28 412 -26
rect 332 -48 468 -28
rect 1132 28 1268 48
rect 1188 26 1212 28
rect 1194 -26 1206 26
rect 1188 -28 1212 -26
rect 1132 -48 1268 -28
rect 1932 28 2068 48
rect 1988 26 2012 28
rect 1994 -26 2006 26
rect 1988 -28 2012 -26
rect 1932 -48 2068 -28
<< via2 >>
rect 732 2746 788 2748
rect 812 2746 868 2748
rect 732 2694 742 2746
rect 742 2694 788 2746
rect 812 2694 858 2746
rect 858 2694 868 2746
rect 732 2692 788 2694
rect 812 2692 868 2694
rect 1532 2746 1588 2748
rect 1612 2746 1668 2748
rect 1532 2694 1542 2746
rect 1542 2694 1588 2746
rect 1612 2694 1658 2746
rect 1658 2694 1668 2746
rect 1532 2692 1588 2694
rect 1612 2692 1668 2694
rect 332 2202 388 2204
rect 412 2202 468 2204
rect 332 2150 342 2202
rect 342 2150 388 2202
rect 412 2150 458 2202
rect 458 2150 468 2202
rect 332 2148 388 2150
rect 412 2148 468 2150
rect 1132 2202 1188 2204
rect 1212 2202 1268 2204
rect 1132 2150 1142 2202
rect 1142 2150 1188 2202
rect 1212 2150 1258 2202
rect 1258 2150 1268 2202
rect 1132 2148 1188 2150
rect 1212 2148 1268 2150
rect 1932 2202 1988 2204
rect 2012 2202 2068 2204
rect 1932 2150 1942 2202
rect 1942 2150 1988 2202
rect 2012 2150 2058 2202
rect 2058 2150 2068 2202
rect 1932 2148 1988 2150
rect 2012 2148 2068 2150
rect 732 1658 788 1660
rect 812 1658 868 1660
rect 732 1606 742 1658
rect 742 1606 788 1658
rect 812 1606 858 1658
rect 858 1606 868 1658
rect 732 1604 788 1606
rect 812 1604 868 1606
rect 1532 1658 1588 1660
rect 1612 1658 1668 1660
rect 1532 1606 1542 1658
rect 1542 1606 1588 1658
rect 1612 1606 1658 1658
rect 1658 1606 1668 1658
rect 1532 1604 1588 1606
rect 1612 1604 1668 1606
rect 1398 1420 1454 1456
rect 1398 1400 1400 1420
rect 1400 1400 1452 1420
rect 1452 1400 1454 1420
rect 332 1114 388 1116
rect 412 1114 468 1116
rect 332 1062 342 1114
rect 342 1062 388 1114
rect 412 1062 458 1114
rect 458 1062 468 1114
rect 332 1060 388 1062
rect 412 1060 468 1062
rect 1132 1114 1188 1116
rect 1212 1114 1268 1116
rect 1132 1062 1142 1114
rect 1142 1062 1188 1114
rect 1212 1062 1258 1114
rect 1258 1062 1268 1114
rect 1132 1060 1188 1062
rect 1212 1060 1268 1062
rect 1932 1114 1988 1116
rect 2012 1114 2068 1116
rect 1932 1062 1942 1114
rect 1942 1062 1988 1114
rect 2012 1062 2058 1114
rect 2058 1062 2068 1114
rect 1932 1060 1988 1062
rect 2012 1060 2068 1062
rect 732 570 788 572
rect 812 570 868 572
rect 732 518 742 570
rect 742 518 788 570
rect 812 518 858 570
rect 858 518 868 570
rect 732 516 788 518
rect 812 516 868 518
rect 1532 570 1588 572
rect 1612 570 1668 572
rect 1532 518 1542 570
rect 1542 518 1588 570
rect 1612 518 1658 570
rect 1658 518 1668 570
rect 1532 516 1588 518
rect 1612 516 1668 518
rect 332 26 388 28
rect 412 26 468 28
rect 332 -26 342 26
rect 342 -26 388 26
rect 412 -26 458 26
rect 458 -26 468 26
rect 332 -28 388 -26
rect 412 -28 468 -26
rect 1132 26 1188 28
rect 1212 26 1268 28
rect 1132 -26 1142 26
rect 1142 -26 1188 26
rect 1212 -26 1258 26
rect 1258 -26 1268 26
rect 1132 -28 1188 -26
rect 1212 -28 1268 -26
rect 1932 26 1988 28
rect 2012 26 2068 28
rect 1932 -26 1942 26
rect 1942 -26 1988 26
rect 2012 -26 2058 26
rect 2058 -26 2068 26
rect 1932 -28 1988 -26
rect 2012 -28 2068 -26
<< metal3 >>
rect 720 2752 880 2753
rect 720 2688 728 2752
rect 792 2688 808 2752
rect 872 2688 880 2752
rect 720 2687 880 2688
rect 1520 2752 1680 2753
rect 1520 2688 1528 2752
rect 1592 2688 1608 2752
rect 1672 2688 1680 2752
rect 1520 2687 1680 2688
rect 320 2208 480 2209
rect 320 2144 328 2208
rect 392 2144 408 2208
rect 472 2144 480 2208
rect 320 2143 480 2144
rect 1120 2208 1280 2209
rect 1120 2144 1128 2208
rect 1192 2144 1208 2208
rect 1272 2144 1280 2208
rect 1120 2143 1280 2144
rect 1920 2208 2080 2209
rect 1920 2144 1928 2208
rect 1992 2144 2008 2208
rect 2072 2144 2080 2208
rect 1920 2143 2080 2144
rect 720 1664 880 1665
rect 720 1600 728 1664
rect 792 1600 808 1664
rect 872 1600 880 1664
rect 720 1599 880 1600
rect 1520 1664 1680 1665
rect 1520 1600 1528 1664
rect 1592 1600 1608 1664
rect 1672 1600 1680 1664
rect 1520 1599 1680 1600
rect 1393 1458 1459 1461
rect 1600 1458 2400 1488
rect 1393 1456 2400 1458
rect 1393 1400 1398 1456
rect 1454 1400 2400 1456
rect 1393 1398 2400 1400
rect 1393 1395 1459 1398
rect 1600 1368 2400 1398
rect 320 1120 480 1121
rect 320 1056 328 1120
rect 392 1056 408 1120
rect 472 1056 480 1120
rect 320 1055 480 1056
rect 1120 1120 1280 1121
rect 1120 1056 1128 1120
rect 1192 1056 1208 1120
rect 1272 1056 1280 1120
rect 1120 1055 1280 1056
rect 1920 1120 2080 1121
rect 1920 1056 1928 1120
rect 1992 1056 2008 1120
rect 2072 1056 2080 1120
rect 1920 1055 2080 1056
rect 720 576 880 577
rect 720 512 728 576
rect 792 512 808 576
rect 872 512 880 576
rect 720 511 880 512
rect 1520 576 1680 577
rect 1520 512 1528 576
rect 1592 512 1608 576
rect 1672 512 1680 576
rect 1520 511 1680 512
rect 320 32 480 33
rect 320 -32 328 32
rect 392 -32 408 32
rect 472 -32 480 32
rect 320 -33 480 -32
rect 1120 32 1280 33
rect 1120 -32 1128 32
rect 1192 -32 1208 32
rect 1272 -32 1280 32
rect 1120 -33 1280 -32
rect 1920 32 2080 33
rect 1920 -32 1928 32
rect 1992 -32 2008 32
rect 2072 -32 2080 32
rect 1920 -33 2080 -32
<< via3 >>
rect 728 2748 792 2752
rect 728 2692 732 2748
rect 732 2692 788 2748
rect 788 2692 792 2748
rect 728 2688 792 2692
rect 808 2748 872 2752
rect 808 2692 812 2748
rect 812 2692 868 2748
rect 868 2692 872 2748
rect 808 2688 872 2692
rect 1528 2748 1592 2752
rect 1528 2692 1532 2748
rect 1532 2692 1588 2748
rect 1588 2692 1592 2748
rect 1528 2688 1592 2692
rect 1608 2748 1672 2752
rect 1608 2692 1612 2748
rect 1612 2692 1668 2748
rect 1668 2692 1672 2748
rect 1608 2688 1672 2692
rect 328 2204 392 2208
rect 328 2148 332 2204
rect 332 2148 388 2204
rect 388 2148 392 2204
rect 328 2144 392 2148
rect 408 2204 472 2208
rect 408 2148 412 2204
rect 412 2148 468 2204
rect 468 2148 472 2204
rect 408 2144 472 2148
rect 1128 2204 1192 2208
rect 1128 2148 1132 2204
rect 1132 2148 1188 2204
rect 1188 2148 1192 2204
rect 1128 2144 1192 2148
rect 1208 2204 1272 2208
rect 1208 2148 1212 2204
rect 1212 2148 1268 2204
rect 1268 2148 1272 2204
rect 1208 2144 1272 2148
rect 1928 2204 1992 2208
rect 1928 2148 1932 2204
rect 1932 2148 1988 2204
rect 1988 2148 1992 2204
rect 1928 2144 1992 2148
rect 2008 2204 2072 2208
rect 2008 2148 2012 2204
rect 2012 2148 2068 2204
rect 2068 2148 2072 2204
rect 2008 2144 2072 2148
rect 728 1660 792 1664
rect 728 1604 732 1660
rect 732 1604 788 1660
rect 788 1604 792 1660
rect 728 1600 792 1604
rect 808 1660 872 1664
rect 808 1604 812 1660
rect 812 1604 868 1660
rect 868 1604 872 1660
rect 808 1600 872 1604
rect 1528 1660 1592 1664
rect 1528 1604 1532 1660
rect 1532 1604 1588 1660
rect 1588 1604 1592 1660
rect 1528 1600 1592 1604
rect 1608 1660 1672 1664
rect 1608 1604 1612 1660
rect 1612 1604 1668 1660
rect 1668 1604 1672 1660
rect 1608 1600 1672 1604
rect 328 1116 392 1120
rect 328 1060 332 1116
rect 332 1060 388 1116
rect 388 1060 392 1116
rect 328 1056 392 1060
rect 408 1116 472 1120
rect 408 1060 412 1116
rect 412 1060 468 1116
rect 468 1060 472 1116
rect 408 1056 472 1060
rect 1128 1116 1192 1120
rect 1128 1060 1132 1116
rect 1132 1060 1188 1116
rect 1188 1060 1192 1116
rect 1128 1056 1192 1060
rect 1208 1116 1272 1120
rect 1208 1060 1212 1116
rect 1212 1060 1268 1116
rect 1268 1060 1272 1116
rect 1208 1056 1272 1060
rect 1928 1116 1992 1120
rect 1928 1060 1932 1116
rect 1932 1060 1988 1116
rect 1988 1060 1992 1116
rect 1928 1056 1992 1060
rect 2008 1116 2072 1120
rect 2008 1060 2012 1116
rect 2012 1060 2068 1116
rect 2068 1060 2072 1116
rect 2008 1056 2072 1060
rect 728 572 792 576
rect 728 516 732 572
rect 732 516 788 572
rect 788 516 792 572
rect 728 512 792 516
rect 808 572 872 576
rect 808 516 812 572
rect 812 516 868 572
rect 868 516 872 572
rect 808 512 872 516
rect 1528 572 1592 576
rect 1528 516 1532 572
rect 1532 516 1588 572
rect 1588 516 1592 572
rect 1528 512 1592 516
rect 1608 572 1672 576
rect 1608 516 1612 572
rect 1612 516 1668 572
rect 1668 516 1672 572
rect 1608 512 1672 516
rect 328 28 392 32
rect 328 -28 332 28
rect 332 -28 388 28
rect 388 -28 392 28
rect 328 -32 392 -28
rect 408 28 472 32
rect 408 -28 412 28
rect 412 -28 468 28
rect 468 -28 472 28
rect 408 -32 472 -28
rect 1128 28 1192 32
rect 1128 -28 1132 28
rect 1132 -28 1188 28
rect 1188 -28 1192 28
rect 1128 -32 1192 -28
rect 1208 28 1272 32
rect 1208 -28 1212 28
rect 1212 -28 1268 28
rect 1268 -28 1272 28
rect 1208 -32 1272 -28
rect 1928 28 1992 32
rect 1928 -28 1932 28
rect 1932 -28 1988 28
rect 1988 -28 1992 28
rect 1928 -32 1992 -28
rect 2008 28 2072 32
rect 2008 -28 2012 28
rect 2012 -28 2068 28
rect 2068 -28 2072 28
rect 2008 -32 2072 -28
<< metal4 >>
rect 320 2208 480 2768
rect 320 2144 328 2208
rect 392 2144 408 2208
rect 472 2144 480 2208
rect 320 1120 480 2144
rect 320 1056 328 1120
rect 392 1056 408 1120
rect 472 1056 480 1120
rect 320 32 480 1056
rect 320 -32 328 32
rect 392 -32 408 32
rect 472 -32 480 32
rect 320 -48 480 -32
rect 720 2752 880 2768
rect 720 2688 728 2752
rect 792 2688 808 2752
rect 872 2688 880 2752
rect 720 1664 880 2688
rect 720 1600 728 1664
rect 792 1600 808 1664
rect 872 1600 880 1664
rect 720 576 880 1600
rect 720 512 728 576
rect 792 512 808 576
rect 872 512 880 576
rect 720 -48 880 512
rect 1120 2208 1280 2768
rect 1120 2144 1128 2208
rect 1192 2144 1208 2208
rect 1272 2144 1280 2208
rect 1120 1120 1280 2144
rect 1120 1056 1128 1120
rect 1192 1056 1208 1120
rect 1272 1056 1280 1120
rect 1120 32 1280 1056
rect 1120 -32 1128 32
rect 1192 -32 1208 32
rect 1272 -32 1280 32
rect 1120 -48 1280 -32
rect 1520 2752 1680 2768
rect 1520 2688 1528 2752
rect 1592 2688 1608 2752
rect 1672 2688 1680 2752
rect 1520 1664 1680 2688
rect 1520 1600 1528 1664
rect 1592 1600 1608 1664
rect 1672 1600 1680 1664
rect 1520 576 1680 1600
rect 1520 512 1528 576
rect 1592 512 1608 576
rect 1672 512 1680 576
rect 1520 -48 1680 512
rect 1920 2208 2080 2768
rect 1920 2144 1928 2208
rect 1992 2144 2008 2208
rect 2072 2144 2080 2208
rect 1920 1120 2080 2144
rect 1920 1056 1928 1120
rect 1992 1056 2008 1120
rect 2072 1056 2080 1120
rect 1920 32 2080 1056
rect 1920 -32 1928 32
rect 1992 -32 2008 32
rect 2072 -32 2080 32
rect 1920 -48 2080 -32
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 0 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624015447
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 828 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 276 0 -1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 920 0 -1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 276 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624015447
transform -1 0 2392 0 -1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624015447
transform -1 0 2392 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_11
timestamp 1624015447
transform 1 0 1656 0 -1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_12
timestamp 1624015447
transform 1 0 1656 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 1748 0 -1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp 1624015447
transform 1 0 1380 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1624015447
transform 1 0 1748 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624015447
transform 1 0 0 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_13
timestamp 1624015447
transform 1 0 828 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1624015447
transform 1 0 276 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_10
timestamp 1624015447
transform 1 0 920 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform -1 0 2024 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624015447
transform -1 0 2392 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624015447
transform 1 0 1656 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_22
timestamp 1624015447
transform 1 0 2024 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624015447
transform 1 0 0 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624015447
transform 1 0 276 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624015447
transform -1 0 2392 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_14
timestamp 1624015447
transform 1 0 1656 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp 1624015447
transform 1 0 1380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1624015447
transform 1 0 1748 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624015447
transform 1 0 0 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_15
timestamp 1624015447
transform 1 0 828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1624015447
transform 1 0 276 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_10
timestamp 1624015447
transform 1 0 920 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624015447
transform -1 0 2392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16
timestamp 1624015447
transform 1 0 1656 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_19
timestamp 1624015447
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
<< labels >>
rlabel metal3 s 1600 1368 2400 1488 6 gpio_logic1
port 0 nsew signal tristate
rlabel metal4 s 1920 -48 2080 2768 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 1120 -48 1280 2768 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 320 -48 480 2768 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 1520 -48 1680 2768 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 720 -48 880 2768 6 vssd1
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2400 2800
<< end >>
