magic
tech sky130A
magscale 1 2
timestamp 1605576936
<< error_s >>
rect 61041 1037419 62959 1037501
rect 60828 1036284 60910 1037318
rect 61120 1036454 61202 1037148
rect 61342 1037137 62648 1037219
rect 61510 1036943 62452 1036993
rect 61365 1036900 61405 1036940
rect 62485 1036900 62525 1036940
rect 61395 1036860 61489 1036900
rect 62401 1036860 62495 1036900
rect 61395 1036700 61489 1036740
rect 62401 1036700 62495 1036740
rect 61365 1036660 61405 1036700
rect 62485 1036660 62525 1036700
rect 61510 1036599 62452 1036649
rect 61342 1036385 62648 1036467
rect 62688 1036454 62770 1037148
rect 62980 1036284 63062 1037318
rect 63881 1036417 63931 1037417
rect 64031 1036417 64159 1037417
rect 64187 1036417 64237 1037417
rect 64303 1036417 64353 1037417
rect 64513 1036417 64569 1037417
rect 64729 1036417 64785 1037417
rect 64885 1036417 65013 1037417
rect 65041 1036417 65091 1037417
rect 65207 1036417 65257 1037417
rect 65417 1036417 65473 1037417
rect 65573 1036417 65701 1037417
rect 65729 1036417 65785 1037417
rect 65885 1036417 66013 1037417
rect 66041 1036417 66097 1037417
rect 66197 1036417 66247 1037417
rect 66313 1036417 66363 1037017
rect 66463 1036417 66513 1037017
rect 66579 1036417 66629 1037417
rect 66729 1036417 66785 1037417
rect 66885 1036417 66935 1037417
rect 67825 1036413 67883 1036447
rect 68665 1036425 68715 1037425
rect 68815 1036425 68943 1037425
rect 68971 1036425 69099 1037425
rect 69127 1036425 69255 1037425
rect 69283 1036425 69411 1037425
rect 69439 1036425 69489 1037425
rect 69555 1036425 69605 1037425
rect 69705 1036425 69761 1037425
rect 69861 1036425 69911 1037425
rect 69977 1036425 70027 1037425
rect 70127 1036425 70255 1037425
rect 70283 1036425 70339 1037425
rect 70439 1036425 70567 1037425
rect 70595 1036425 70645 1037425
rect 70711 1036425 70761 1037425
rect 70861 1036425 70989 1037425
rect 71017 1036425 71073 1037425
rect 71173 1036425 71301 1037425
rect 71329 1036797 71379 1037425
rect 109041 1037419 110959 1037501
rect 161041 1037419 162959 1037501
rect 71329 1036725 71382 1036797
rect 71329 1036425 71379 1036725
rect 71442 1036425 71454 1036725
rect 75030 1036262 76030 1036312
rect 108828 1036284 108910 1037318
rect 109120 1036454 109202 1037148
rect 109342 1037137 110648 1037219
rect 109510 1036943 110452 1036993
rect 109365 1036900 109405 1036940
rect 109395 1036860 109489 1036900
rect 109395 1036700 109489 1036740
rect 109365 1036660 109405 1036700
rect 109510 1036599 110452 1036649
rect 109342 1036385 110648 1036467
rect 110688 1036454 110770 1037148
rect 110980 1036284 111062 1037318
rect 123030 1036262 124030 1036312
rect 160828 1036284 160910 1037318
rect 161120 1036454 161202 1037148
rect 161342 1037137 162648 1037219
rect 161510 1036943 162452 1036993
rect 161365 1036900 161405 1036940
rect 162485 1036900 162525 1036940
rect 161395 1036860 161489 1036900
rect 162401 1036860 162495 1036900
rect 161395 1036700 161489 1036740
rect 162401 1036700 162495 1036740
rect 161365 1036660 161405 1036700
rect 162485 1036660 162525 1036700
rect 161510 1036599 162452 1036649
rect 161342 1036385 162648 1036467
rect 162688 1036454 162770 1037148
rect 162980 1036284 163062 1037318
rect 163881 1036417 163931 1037417
rect 164031 1036417 164159 1037417
rect 164187 1036417 164237 1037417
rect 164303 1036417 164353 1037417
rect 164513 1036417 164569 1037417
rect 164729 1036417 164785 1037417
rect 164885 1036417 165013 1037417
rect 165041 1036417 165091 1037417
rect 165207 1036417 165257 1037417
rect 165417 1036417 165473 1037417
rect 165573 1036417 165701 1037417
rect 165729 1036417 165785 1037417
rect 165885 1036417 166013 1037417
rect 166041 1036417 166097 1037417
rect 166197 1036417 166247 1037417
rect 166313 1036417 166363 1037017
rect 166463 1036417 166513 1037017
rect 166579 1036417 166629 1037417
rect 166729 1036417 166785 1037417
rect 166885 1036417 166935 1037417
rect 167825 1036413 167883 1036447
rect 168665 1036425 168715 1037425
rect 168815 1036425 168943 1037425
rect 168971 1036425 169099 1037425
rect 169127 1036425 169255 1037425
rect 169283 1036425 169411 1037425
rect 169439 1036425 169489 1037425
rect 169555 1036425 169605 1037425
rect 169705 1036425 169761 1037425
rect 169861 1036425 169911 1037425
rect 169977 1036425 170027 1037425
rect 170127 1036425 170255 1037425
rect 170283 1036425 170339 1037425
rect 170439 1036425 170567 1037425
rect 170595 1036425 170645 1037425
rect 170711 1036425 170761 1037425
rect 170861 1036425 170989 1037425
rect 171017 1036425 171073 1037425
rect 171173 1036425 171301 1037425
rect 171329 1036797 171379 1037425
rect 213041 1037419 214959 1037501
rect 261041 1037419 262080 1037501
rect 313041 1037419 314959 1037501
rect 365041 1037419 366959 1037501
rect 171329 1036725 171382 1036797
rect 171329 1036425 171379 1036725
rect 171442 1036425 171454 1036725
rect 175030 1036262 176030 1036312
rect 212828 1036284 212910 1037318
rect 213120 1036454 213202 1037148
rect 213342 1037137 214648 1037219
rect 213510 1036943 214452 1036993
rect 213365 1036900 213405 1036940
rect 213395 1036860 213489 1036900
rect 213395 1036700 213489 1036740
rect 213365 1036660 213405 1036700
rect 213510 1036599 214452 1036649
rect 213342 1036385 214648 1036467
rect 214688 1036454 214770 1037148
rect 214980 1036284 215062 1037318
rect 227030 1036262 228030 1036312
rect 260828 1036284 260910 1037318
rect 261120 1036454 261202 1037148
rect 261342 1037137 262080 1037219
rect 261510 1036943 262080 1036993
rect 261365 1036900 261405 1036940
rect 261395 1036860 261489 1036900
rect 261395 1036700 261489 1036740
rect 261365 1036660 261405 1036700
rect 261510 1036599 262080 1036649
rect 261342 1036385 262080 1036467
rect 275030 1036262 276030 1036312
rect 312828 1036284 312910 1037318
rect 313120 1036454 313202 1037148
rect 313342 1037137 314648 1037219
rect 313510 1036943 314452 1036993
rect 313365 1036900 313405 1036940
rect 313395 1036860 313489 1036900
rect 313395 1036700 313489 1036740
rect 313365 1036660 313405 1036700
rect 313510 1036599 314452 1036649
rect 313342 1036385 314648 1036467
rect 314688 1036454 314770 1037148
rect 314980 1036284 315062 1037318
rect 327030 1036262 328030 1036312
rect 364828 1036284 364910 1037318
rect 365120 1036454 365202 1037148
rect 365342 1037137 366648 1037219
rect 365510 1036943 366452 1036993
rect 365365 1036900 365405 1036940
rect 366485 1036900 366525 1036940
rect 365395 1036860 365489 1036900
rect 366401 1036860 366495 1036900
rect 365395 1036700 365489 1036740
rect 366401 1036700 366495 1036740
rect 365365 1036660 365405 1036700
rect 366485 1036660 366525 1036700
rect 365510 1036599 366452 1036649
rect 365342 1036385 366648 1036467
rect 366688 1036454 366770 1037148
rect 366980 1036284 367062 1037318
rect 367881 1036417 367931 1037417
rect 368031 1036417 368159 1037417
rect 368187 1036417 368237 1037417
rect 368303 1036417 368353 1037417
rect 368513 1036417 368569 1037417
rect 368729 1036417 368785 1037417
rect 368885 1036417 369013 1037417
rect 369041 1036417 369091 1037417
rect 369207 1036417 369257 1037417
rect 369417 1036417 369473 1037417
rect 369573 1036417 369701 1037417
rect 369729 1036417 369785 1037417
rect 369885 1036417 370013 1037417
rect 370041 1036417 370097 1037417
rect 370197 1036417 370247 1037417
rect 370313 1036417 370363 1037017
rect 370463 1036417 370513 1037017
rect 370579 1036417 370629 1037417
rect 370729 1036417 370785 1037417
rect 370885 1036417 370935 1037417
rect 371825 1036413 371883 1036447
rect 372665 1036425 372715 1037425
rect 372815 1036425 372943 1037425
rect 372971 1036425 373099 1037425
rect 373127 1036425 373255 1037425
rect 373283 1036425 373411 1037425
rect 373439 1036425 373489 1037425
rect 373555 1036425 373605 1037425
rect 373705 1036425 373761 1037425
rect 373861 1036425 373911 1037425
rect 373977 1036425 374027 1037425
rect 374127 1036425 374255 1037425
rect 374283 1036425 374339 1037425
rect 374439 1036425 374567 1037425
rect 374595 1036425 374645 1037425
rect 374711 1036425 374761 1037425
rect 374861 1036425 374989 1037425
rect 375017 1036425 375073 1037425
rect 375173 1036425 375301 1037425
rect 375329 1036797 375379 1037425
rect 413041 1037419 414959 1037501
rect 465041 1037419 466959 1037501
rect 375329 1036725 375382 1036797
rect 375329 1036425 375379 1036725
rect 375442 1036425 375454 1036725
rect 379030 1036262 380030 1036312
rect 412828 1036284 412910 1037318
rect 413120 1036454 413202 1037148
rect 413342 1037137 414648 1037219
rect 413510 1036943 414452 1036993
rect 413365 1036900 413405 1036940
rect 413395 1036860 413489 1036900
rect 413395 1036700 413489 1036740
rect 413365 1036660 413405 1036700
rect 413510 1036599 414452 1036649
rect 413342 1036385 414648 1036467
rect 414688 1036454 414770 1037148
rect 414980 1036284 415062 1037318
rect 427030 1036262 428030 1036312
rect 464828 1036284 464910 1037318
rect 465120 1036454 465202 1037148
rect 465342 1037137 466648 1037219
rect 465510 1036943 466452 1036993
rect 465365 1036900 465405 1036940
rect 466485 1036900 466525 1036940
rect 465395 1036860 465489 1036900
rect 466401 1036860 466495 1036900
rect 465395 1036700 465489 1036740
rect 466401 1036700 466495 1036740
rect 465365 1036660 465405 1036700
rect 466485 1036660 466525 1036700
rect 465510 1036599 466452 1036649
rect 465342 1036385 466648 1036467
rect 466688 1036454 466770 1037148
rect 466980 1036284 467062 1037318
rect 467881 1036417 467931 1037417
rect 468031 1036417 468159 1037417
rect 468187 1036417 468237 1037417
rect 468303 1036417 468353 1037417
rect 468513 1036417 468569 1037417
rect 468729 1036417 468785 1037417
rect 468885 1036417 469013 1037417
rect 469041 1036417 469091 1037417
rect 469207 1036417 469257 1037417
rect 469417 1036417 469473 1037417
rect 469573 1036417 469701 1037417
rect 469729 1036417 469785 1037417
rect 469885 1036417 470013 1037417
rect 470041 1036417 470097 1037417
rect 470197 1036417 470247 1037417
rect 470313 1036417 470363 1037017
rect 470463 1036417 470513 1037017
rect 470579 1036417 470629 1037417
rect 470729 1036417 470785 1037417
rect 470885 1036417 470935 1037417
rect 471825 1036413 471883 1036447
rect 472665 1036425 472715 1037425
rect 472815 1036425 472943 1037425
rect 472971 1036425 473099 1037425
rect 473127 1036425 473255 1037425
rect 473283 1036425 473411 1037425
rect 473439 1036425 473489 1037425
rect 473555 1036425 473605 1037425
rect 473705 1036425 473761 1037425
rect 473861 1036425 473911 1037425
rect 473977 1036425 474027 1037425
rect 474127 1036425 474255 1037425
rect 474283 1036425 474339 1037425
rect 474439 1036425 474567 1037425
rect 474595 1036425 474645 1037425
rect 474711 1036425 474761 1037425
rect 474861 1036425 474989 1037425
rect 475017 1036425 475073 1037425
rect 475173 1036425 475301 1037425
rect 475329 1036797 475379 1037425
rect 517041 1037419 518959 1037501
rect 569041 1037419 570959 1037501
rect 475329 1036725 475382 1036797
rect 475329 1036425 475379 1036725
rect 475442 1036425 475454 1036725
rect 479030 1036262 480030 1036312
rect 516828 1036284 516910 1037318
rect 517120 1036454 517202 1037148
rect 517342 1037137 518648 1037219
rect 517510 1036943 518452 1036993
rect 517365 1036900 517405 1036940
rect 517395 1036860 517489 1036900
rect 517395 1036700 517489 1036740
rect 517365 1036660 517405 1036700
rect 517510 1036599 518452 1036649
rect 517342 1036385 518648 1036467
rect 518688 1036454 518770 1037148
rect 518980 1036284 519062 1037318
rect 531030 1036262 532030 1036312
rect 568828 1036284 568910 1037318
rect 569120 1036454 569202 1037148
rect 569342 1037137 570648 1037219
rect 569510 1036943 570452 1036993
rect 569365 1036900 569405 1036940
rect 570485 1036900 570525 1036940
rect 569395 1036860 569489 1036900
rect 570401 1036860 570495 1036900
rect 569395 1036700 569489 1036740
rect 570401 1036700 570495 1036740
rect 569365 1036660 569405 1036700
rect 570485 1036660 570525 1036700
rect 569510 1036599 570452 1036649
rect 569342 1036385 570648 1036467
rect 570688 1036454 570770 1037148
rect 570980 1036284 571062 1037318
rect 571881 1036417 571931 1037417
rect 572031 1036417 572159 1037417
rect 572187 1036417 572237 1037417
rect 572303 1036417 572353 1037417
rect 572513 1036417 572569 1037417
rect 572729 1036417 572785 1037417
rect 572885 1036417 573013 1037417
rect 573041 1036417 573091 1037417
rect 573207 1036417 573257 1037417
rect 573417 1036417 573473 1037417
rect 573573 1036417 573701 1037417
rect 573729 1036417 573785 1037417
rect 573885 1036417 574013 1037417
rect 574041 1036417 574097 1037417
rect 574197 1036417 574247 1037417
rect 574313 1036417 574363 1037017
rect 574463 1036417 574513 1037017
rect 574579 1036417 574629 1037417
rect 574729 1036417 574785 1037417
rect 574885 1036417 574935 1037417
rect 575825 1036413 575883 1036447
rect 576665 1036425 576715 1037425
rect 576815 1036425 576943 1037425
rect 576971 1036425 577099 1037425
rect 577127 1036425 577255 1037425
rect 577283 1036425 577411 1037425
rect 577439 1036425 577489 1037425
rect 577555 1036425 577605 1037425
rect 577705 1036425 577761 1037425
rect 577861 1036425 577911 1037425
rect 577977 1036425 578027 1037425
rect 578127 1036425 578255 1037425
rect 578283 1036425 578339 1037425
rect 578439 1036425 578567 1037425
rect 578595 1036425 578645 1037425
rect 578711 1036425 578761 1037425
rect 578861 1036425 578989 1037425
rect 579017 1036425 579073 1037425
rect 579173 1036425 579301 1037425
rect 579329 1036797 579379 1037425
rect 579329 1036725 579382 1036797
rect 579329 1036425 579379 1036725
rect 579442 1036425 579454 1036725
rect 583030 1036262 584030 1036312
rect 63088 1036210 63091 1036211
rect 63088 1036209 63089 1036210
rect 63090 1036209 63091 1036210
rect 63088 1036208 63091 1036209
rect 61041 1036100 62959 1036182
rect 75030 1036106 76030 1036234
rect 111088 1036210 111091 1036211
rect 111088 1036209 111089 1036210
rect 111090 1036209 111091 1036210
rect 111088 1036208 111091 1036209
rect 109041 1036100 110959 1036182
rect 123473 1036106 124030 1036234
rect 163088 1036210 163091 1036211
rect 163088 1036209 163089 1036210
rect 163090 1036209 163091 1036210
rect 163088 1036208 163091 1036209
rect 161041 1036100 162959 1036182
rect 175030 1036106 176030 1036234
rect 215088 1036210 215091 1036211
rect 215088 1036209 215089 1036210
rect 215090 1036209 215091 1036210
rect 215088 1036208 215091 1036209
rect 213041 1036100 214959 1036182
rect 227473 1036106 228030 1036234
rect 261041 1036100 262080 1036182
rect 275473 1036106 276030 1036234
rect 315088 1036210 315091 1036211
rect 315088 1036209 315089 1036210
rect 315090 1036209 315091 1036210
rect 315088 1036208 315091 1036209
rect 313041 1036100 314959 1036182
rect 327473 1036106 328030 1036234
rect 367088 1036210 367091 1036211
rect 367088 1036209 367089 1036210
rect 367090 1036209 367091 1036210
rect 367088 1036208 367091 1036209
rect 365041 1036100 366959 1036182
rect 379030 1036106 380030 1036234
rect 415088 1036210 415091 1036211
rect 415088 1036209 415089 1036210
rect 415090 1036209 415091 1036210
rect 415088 1036208 415091 1036209
rect 413041 1036100 414959 1036182
rect 427473 1036106 428030 1036234
rect 467088 1036210 467091 1036211
rect 467088 1036209 467089 1036210
rect 467090 1036209 467091 1036210
rect 467088 1036208 467091 1036209
rect 465041 1036100 466959 1036182
rect 479030 1036106 480030 1036234
rect 519088 1036210 519091 1036211
rect 519088 1036209 519089 1036210
rect 519090 1036209 519091 1036210
rect 519088 1036208 519091 1036209
rect 517041 1036100 518959 1036182
rect 531473 1036106 532030 1036234
rect 571088 1036210 571091 1036211
rect 571088 1036209 571089 1036210
rect 571090 1036209 571091 1036210
rect 571088 1036208 571091 1036209
rect 569041 1036100 570959 1036182
rect 583030 1036106 584030 1036234
rect 63088 1036073 63091 1036074
rect 63088 1036072 63089 1036073
rect 63090 1036072 63091 1036073
rect 63088 1036071 63091 1036072
rect 111088 1036073 111091 1036074
rect 111088 1036072 111089 1036073
rect 111090 1036072 111091 1036073
rect 111088 1036071 111091 1036072
rect 163088 1036073 163091 1036074
rect 163088 1036072 163089 1036073
rect 163090 1036072 163091 1036073
rect 163088 1036071 163091 1036072
rect 215088 1036073 215091 1036074
rect 215088 1036072 215089 1036073
rect 215090 1036072 215091 1036073
rect 215088 1036071 215091 1036072
rect 315088 1036073 315091 1036074
rect 315088 1036072 315089 1036073
rect 315090 1036072 315091 1036073
rect 315088 1036071 315091 1036072
rect 367088 1036073 367091 1036074
rect 367088 1036072 367089 1036073
rect 367090 1036072 367091 1036073
rect 367088 1036071 367091 1036072
rect 415088 1036073 415091 1036074
rect 415088 1036072 415089 1036073
rect 415090 1036072 415091 1036073
rect 415088 1036071 415091 1036072
rect 467088 1036073 467091 1036074
rect 467088 1036072 467089 1036073
rect 467090 1036072 467091 1036073
rect 467088 1036071 467091 1036072
rect 519088 1036073 519091 1036074
rect 519088 1036072 519089 1036073
rect 519090 1036072 519091 1036073
rect 519088 1036071 519091 1036072
rect 571088 1036073 571091 1036074
rect 571088 1036072 571089 1036073
rect 571090 1036072 571091 1036073
rect 571088 1036071 571091 1036072
rect 60828 1034964 60910 1035998
rect 61120 1035134 61202 1035828
rect 61342 1035815 62648 1035897
rect 61510 1035633 62452 1035683
rect 61365 1035582 61405 1035622
rect 62485 1035582 62525 1035622
rect 61395 1035560 61489 1035582
rect 61395 1035542 61405 1035560
rect 61427 1035542 61489 1035560
rect 62401 1035560 62495 1035582
rect 62401 1035542 62463 1035560
rect 62485 1035542 62495 1035560
rect 61395 1035404 61405 1035422
rect 61427 1035404 61489 1035422
rect 61395 1035382 61489 1035404
rect 62401 1035404 62463 1035422
rect 62485 1035404 62495 1035422
rect 62401 1035382 62495 1035404
rect 61374 1035351 61405 1035382
rect 62485 1035351 62516 1035382
rect 61365 1035342 61374 1035351
rect 62516 1035342 62525 1035351
rect 61510 1035289 62452 1035339
rect 61342 1035063 62648 1035145
rect 62688 1035134 62770 1035828
rect 62980 1034964 63062 1035998
rect 68924 1035972 69924 1036022
rect 70320 1035972 70920 1036022
rect 68924 1035816 69924 1035944
rect 72664 1035912 73664 1035962
rect 75030 1035956 76030 1036006
rect 70320 1035816 70920 1035872
rect 68924 1035660 69924 1035788
rect 70320 1035660 70920 1035716
rect 72664 1035696 73664 1035824
rect 68924 1035510 69924 1035560
rect 70320 1035504 70920 1035560
rect 72664 1035486 73664 1035536
rect 70320 1035354 70920 1035404
rect 108828 1034964 108910 1035998
rect 109120 1035134 109202 1035828
rect 109342 1035815 110648 1035897
rect 109510 1035633 110452 1035683
rect 109365 1035582 109405 1035622
rect 109395 1035542 109489 1035582
rect 109395 1035382 109489 1035422
rect 109365 1035342 109405 1035382
rect 109510 1035289 110452 1035339
rect 109342 1035063 110648 1035145
rect 110688 1035134 110770 1035828
rect 110980 1034964 111062 1035998
rect 123030 1035956 124030 1036006
rect 160828 1034964 160910 1035998
rect 161120 1035134 161202 1035828
rect 161342 1035815 162648 1035897
rect 161510 1035633 162452 1035683
rect 161365 1035582 161405 1035622
rect 162485 1035582 162525 1035622
rect 161395 1035560 161489 1035582
rect 161395 1035542 161405 1035560
rect 161427 1035542 161489 1035560
rect 162401 1035560 162495 1035582
rect 162401 1035542 162463 1035560
rect 162485 1035542 162495 1035560
rect 161395 1035404 161405 1035422
rect 161427 1035404 161489 1035422
rect 161395 1035382 161489 1035404
rect 162401 1035404 162463 1035422
rect 162485 1035404 162495 1035422
rect 162401 1035382 162495 1035404
rect 161374 1035351 161405 1035382
rect 162485 1035351 162516 1035382
rect 161365 1035342 161374 1035351
rect 162516 1035342 162525 1035351
rect 161510 1035289 162452 1035339
rect 161342 1035063 162648 1035145
rect 162688 1035134 162770 1035828
rect 162980 1034964 163062 1035998
rect 168924 1035972 169924 1036022
rect 170320 1035972 170920 1036022
rect 168924 1035816 169924 1035944
rect 172664 1035912 173664 1035962
rect 175030 1035956 176030 1036006
rect 170320 1035816 170920 1035872
rect 168924 1035660 169924 1035788
rect 170320 1035660 170920 1035716
rect 172664 1035696 173664 1035824
rect 168924 1035510 169924 1035560
rect 170320 1035504 170920 1035560
rect 172664 1035486 173664 1035536
rect 170320 1035354 170920 1035404
rect 212828 1034964 212910 1035998
rect 213120 1035134 213202 1035828
rect 213342 1035815 214648 1035897
rect 213510 1035633 214452 1035683
rect 213365 1035582 213405 1035622
rect 213395 1035542 213489 1035582
rect 213395 1035382 213489 1035422
rect 213365 1035342 213405 1035382
rect 213510 1035289 214452 1035339
rect 213342 1035063 214648 1035145
rect 214688 1035134 214770 1035828
rect 214980 1034964 215062 1035998
rect 227030 1035956 228030 1036006
rect 260828 1034964 260910 1035998
rect 275030 1035956 276030 1036006
rect 261120 1035134 261202 1035828
rect 261342 1035815 262080 1035897
rect 261510 1035633 262080 1035683
rect 261365 1035582 261405 1035622
rect 261395 1035542 261489 1035582
rect 261395 1035382 261489 1035422
rect 261365 1035342 261405 1035382
rect 261510 1035289 262080 1035339
rect 261342 1035063 262080 1035145
rect 312828 1034964 312910 1035998
rect 313120 1035134 313202 1035828
rect 313342 1035815 314648 1035897
rect 313510 1035633 314452 1035683
rect 313365 1035582 313405 1035622
rect 313395 1035542 313489 1035582
rect 313395 1035382 313489 1035422
rect 313365 1035342 313405 1035382
rect 313510 1035289 314452 1035339
rect 313342 1035063 314648 1035145
rect 314688 1035134 314770 1035828
rect 314980 1034964 315062 1035998
rect 327030 1035956 328030 1036006
rect 364828 1034964 364910 1035998
rect 365120 1035134 365202 1035828
rect 365342 1035815 366648 1035897
rect 365510 1035633 366452 1035683
rect 365365 1035582 365405 1035622
rect 366485 1035582 366525 1035622
rect 365395 1035560 365489 1035582
rect 365395 1035542 365405 1035560
rect 365427 1035542 365489 1035560
rect 366401 1035560 366495 1035582
rect 366401 1035542 366463 1035560
rect 366485 1035542 366495 1035560
rect 365395 1035404 365405 1035422
rect 365427 1035404 365489 1035422
rect 365395 1035382 365489 1035404
rect 366401 1035404 366463 1035422
rect 366485 1035404 366495 1035422
rect 366401 1035382 366495 1035404
rect 365374 1035351 365405 1035382
rect 366485 1035351 366516 1035382
rect 365365 1035342 365374 1035351
rect 366516 1035342 366525 1035351
rect 365510 1035289 366452 1035339
rect 365342 1035063 366648 1035145
rect 366688 1035134 366770 1035828
rect 366980 1034964 367062 1035998
rect 372924 1035972 373924 1036022
rect 374320 1035972 374920 1036022
rect 372924 1035816 373924 1035944
rect 376664 1035912 377664 1035962
rect 379030 1035956 380030 1036006
rect 374320 1035816 374920 1035872
rect 372924 1035660 373924 1035788
rect 374320 1035660 374920 1035716
rect 376664 1035696 377664 1035824
rect 372924 1035510 373924 1035560
rect 374320 1035504 374920 1035560
rect 376664 1035486 377664 1035536
rect 374320 1035354 374920 1035404
rect 412828 1034964 412910 1035998
rect 413120 1035134 413202 1035828
rect 413342 1035815 414648 1035897
rect 413510 1035633 414452 1035683
rect 413365 1035582 413405 1035622
rect 413395 1035542 413489 1035582
rect 413395 1035382 413489 1035422
rect 413365 1035342 413405 1035382
rect 413510 1035289 414452 1035339
rect 413342 1035063 414648 1035145
rect 414688 1035134 414770 1035828
rect 414980 1034964 415062 1035998
rect 427030 1035956 428030 1036006
rect 464828 1034964 464910 1035998
rect 465120 1035134 465202 1035828
rect 465342 1035815 466648 1035897
rect 465510 1035633 466452 1035683
rect 465365 1035582 465405 1035622
rect 466485 1035582 466525 1035622
rect 465395 1035560 465489 1035582
rect 465395 1035542 465405 1035560
rect 465427 1035542 465489 1035560
rect 466401 1035560 466495 1035582
rect 466401 1035542 466463 1035560
rect 466485 1035542 466495 1035560
rect 465395 1035404 465405 1035422
rect 465427 1035404 465489 1035422
rect 465395 1035382 465489 1035404
rect 466401 1035404 466463 1035422
rect 466485 1035404 466495 1035422
rect 466401 1035382 466495 1035404
rect 465374 1035351 465405 1035382
rect 466485 1035351 466516 1035382
rect 465365 1035342 465374 1035351
rect 466516 1035342 466525 1035351
rect 465510 1035289 466452 1035339
rect 465342 1035063 466648 1035145
rect 466688 1035134 466770 1035828
rect 466980 1034964 467062 1035998
rect 472924 1035972 473924 1036022
rect 474320 1035972 474920 1036022
rect 472924 1035816 473924 1035944
rect 476664 1035912 477664 1035962
rect 479030 1035956 480030 1036006
rect 474320 1035816 474920 1035872
rect 472924 1035660 473924 1035788
rect 474320 1035660 474920 1035716
rect 476664 1035696 477664 1035824
rect 472924 1035510 473924 1035560
rect 474320 1035504 474920 1035560
rect 476664 1035486 477664 1035536
rect 474320 1035354 474920 1035404
rect 516828 1034964 516910 1035998
rect 517120 1035134 517202 1035828
rect 517342 1035815 518648 1035897
rect 517510 1035633 518452 1035683
rect 517365 1035582 517405 1035622
rect 517395 1035542 517489 1035582
rect 517395 1035382 517489 1035422
rect 517365 1035342 517405 1035382
rect 517510 1035289 518452 1035339
rect 517342 1035063 518648 1035145
rect 518688 1035134 518770 1035828
rect 518980 1034964 519062 1035998
rect 531030 1035956 532030 1036006
rect 568828 1034964 568910 1035998
rect 569120 1035134 569202 1035828
rect 569342 1035815 570648 1035897
rect 569510 1035633 570452 1035683
rect 569365 1035582 569405 1035622
rect 570485 1035582 570525 1035622
rect 569395 1035560 569489 1035582
rect 569395 1035542 569405 1035560
rect 569427 1035542 569489 1035560
rect 570401 1035560 570495 1035582
rect 570401 1035542 570463 1035560
rect 570485 1035542 570495 1035560
rect 569395 1035404 569405 1035422
rect 569427 1035404 569489 1035422
rect 569395 1035382 569489 1035404
rect 570401 1035404 570463 1035422
rect 570485 1035404 570495 1035422
rect 570401 1035382 570495 1035404
rect 569374 1035351 569405 1035382
rect 570485 1035351 570516 1035382
rect 569365 1035342 569374 1035351
rect 570516 1035342 570525 1035351
rect 569510 1035289 570452 1035339
rect 569342 1035063 570648 1035145
rect 570688 1035134 570770 1035828
rect 570980 1034964 571062 1035998
rect 576924 1035972 577924 1036022
rect 578320 1035972 578920 1036022
rect 576924 1035816 577924 1035944
rect 580664 1035912 581664 1035962
rect 583030 1035956 584030 1036006
rect 578320 1035816 578920 1035872
rect 576924 1035660 577924 1035788
rect 578320 1035660 578920 1035716
rect 580664 1035696 581664 1035824
rect 576924 1035510 577924 1035560
rect 578320 1035504 578920 1035560
rect 580664 1035486 581664 1035536
rect 578320 1035354 578920 1035404
rect 61041 1034781 62959 1034863
rect 61754 1034726 61924 1034781
rect 62988 1034726 63157 1034794
rect 109041 1034781 110959 1034863
rect 161041 1034781 162959 1034863
rect 61822 1034686 61924 1034726
rect 63056 1034686 63157 1034726
rect 61822 1034645 61856 1034686
rect 63056 1034645 63090 1034686
rect 62131 1034425 62731 1034475
rect 62131 1034175 62731 1034225
rect 63851 1033750 63901 1034750
rect 64061 1033750 64189 1034750
rect 64277 1033750 64405 1034750
rect 64493 1033750 64621 1034750
rect 64709 1033750 64837 1034750
rect 64925 1033750 64981 1034750
rect 65141 1033750 65197 1034750
rect 65357 1033750 65485 1034750
rect 65573 1033750 65701 1034750
rect 65789 1033750 65917 1034750
rect 66005 1033750 66133 1034750
rect 66221 1033750 66277 1034750
rect 66437 1033750 66565 1034750
rect 66653 1033750 66781 1034750
rect 66869 1033750 66997 1034750
rect 67085 1033750 67135 1034750
rect 67201 1033750 67251 1034750
rect 67411 1033750 67461 1034750
rect 67527 1033750 67577 1034750
rect 67737 1033750 67787 1034750
rect 67853 1033750 67903 1034750
rect 68063 1033750 68113 1034750
rect 68176 1034565 68188 1034765
rect 68179 1033750 68229 1034350
rect 68429 1033750 68485 1034350
rect 68585 1033750 68713 1034350
rect 68741 1033750 68797 1034350
rect 68897 1033750 69025 1034350
rect 69053 1033750 69103 1034350
rect 69169 1033750 69219 1034750
rect 69319 1033750 69375 1034750
rect 69475 1033750 69525 1034750
rect 69603 1033750 69653 1034750
rect 69753 1033750 69881 1034750
rect 69909 1033750 70037 1034750
rect 70065 1033750 70121 1034750
rect 70221 1033750 70349 1034750
rect 70377 1033750 70505 1034750
rect 70533 1033750 70661 1034750
rect 70689 1033750 70739 1034750
rect 70805 1033750 70855 1034750
rect 70955 1033750 71083 1034750
rect 71111 1033750 71239 1034750
rect 71267 1033750 71395 1034750
rect 71423 1033750 71479 1034750
rect 71579 1033750 71707 1034750
rect 71735 1033750 71863 1034750
rect 71891 1033750 71947 1034750
rect 72047 1033750 72097 1034750
rect 73318 1034550 73371 1034750
rect 73321 1033750 73371 1034550
rect 73531 1033750 73659 1034750
rect 73747 1033750 73803 1034750
rect 73963 1033750 74091 1034750
rect 74179 1033750 74229 1034750
rect 74295 1033750 74345 1034750
rect 74505 1033750 74555 1034750
rect 109754 1034726 109924 1034781
rect 109822 1034686 109924 1034726
rect 109822 1034645 109856 1034686
rect 111056 1034645 111090 1034752
rect 110131 1034425 110731 1034475
rect 110131 1034175 110731 1034225
rect 122213 1033750 122229 1034750
rect 122295 1033750 122345 1034750
rect 122505 1033750 122555 1034750
rect 161754 1034726 161924 1034781
rect 162988 1034726 163157 1034794
rect 213041 1034781 214959 1034863
rect 261041 1034781 262080 1034863
rect 313041 1034781 314959 1034863
rect 365041 1034781 366959 1034863
rect 161822 1034686 161924 1034726
rect 163056 1034686 163157 1034726
rect 161822 1034645 161856 1034686
rect 163056 1034645 163090 1034686
rect 162131 1034425 162731 1034475
rect 162131 1034175 162731 1034225
rect 163851 1033750 163901 1034750
rect 164061 1033750 164189 1034750
rect 164277 1033750 164405 1034750
rect 164493 1033750 164621 1034750
rect 164709 1033750 164837 1034750
rect 164925 1033750 164981 1034750
rect 165141 1033750 165197 1034750
rect 165357 1033750 165485 1034750
rect 165573 1033750 165701 1034750
rect 165789 1033750 165917 1034750
rect 166005 1033750 166133 1034750
rect 166221 1033750 166277 1034750
rect 166437 1033750 166565 1034750
rect 166653 1033750 166781 1034750
rect 166869 1033750 166997 1034750
rect 167085 1033750 167135 1034750
rect 167201 1033750 167251 1034750
rect 167411 1033750 167461 1034750
rect 167527 1033750 167577 1034750
rect 167737 1033750 167787 1034750
rect 167853 1033750 167903 1034750
rect 168063 1033750 168113 1034750
rect 168176 1034565 168188 1034765
rect 168179 1033750 168229 1034350
rect 168429 1033750 168485 1034350
rect 168585 1033750 168713 1034350
rect 168741 1033750 168797 1034350
rect 168897 1033750 169025 1034350
rect 169053 1033750 169103 1034350
rect 169169 1033750 169219 1034750
rect 169319 1033750 169375 1034750
rect 169475 1033750 169525 1034750
rect 169603 1033750 169653 1034750
rect 169753 1033750 169881 1034750
rect 169909 1033750 170037 1034750
rect 170065 1033750 170121 1034750
rect 170221 1033750 170349 1034750
rect 170377 1033750 170505 1034750
rect 170533 1033750 170661 1034750
rect 170689 1033750 170739 1034750
rect 170805 1033750 170855 1034750
rect 170955 1033750 171083 1034750
rect 171111 1033750 171239 1034750
rect 171267 1033750 171395 1034750
rect 171423 1033750 171479 1034750
rect 171579 1033750 171707 1034750
rect 171735 1033750 171863 1034750
rect 171891 1033750 171947 1034750
rect 172047 1033750 172097 1034750
rect 173318 1034550 173371 1034750
rect 173321 1033750 173371 1034550
rect 173531 1033750 173659 1034750
rect 173747 1033750 173803 1034750
rect 173963 1033750 174091 1034750
rect 174179 1033750 174229 1034750
rect 174295 1033750 174345 1034750
rect 174505 1033750 174555 1034750
rect 213754 1034726 213924 1034781
rect 213822 1034686 213924 1034726
rect 213822 1034645 213856 1034686
rect 215056 1034645 215090 1034752
rect 214131 1034425 214731 1034475
rect 214131 1034175 214731 1034225
rect 226213 1033750 226229 1034750
rect 226295 1033750 226345 1034750
rect 226505 1033750 226555 1034750
rect 261754 1034726 261924 1034781
rect 261822 1034686 261924 1034726
rect 261822 1034645 261856 1034686
rect 274213 1033750 274229 1034750
rect 274295 1033750 274345 1034750
rect 274505 1033750 274555 1034750
rect 313754 1034726 313924 1034781
rect 313822 1034686 313924 1034726
rect 313822 1034645 313856 1034686
rect 315056 1034645 315090 1034752
rect 314131 1034425 314731 1034475
rect 314131 1034175 314731 1034225
rect 326213 1033750 326229 1034750
rect 326295 1033750 326345 1034750
rect 326505 1033750 326555 1034750
rect 365754 1034726 365924 1034781
rect 366988 1034726 367157 1034794
rect 413041 1034781 414959 1034863
rect 465041 1034781 466959 1034863
rect 365822 1034686 365924 1034726
rect 367056 1034686 367157 1034726
rect 365822 1034645 365856 1034686
rect 367056 1034645 367090 1034686
rect 366131 1034425 366731 1034475
rect 366131 1034175 366731 1034225
rect 367851 1033750 367901 1034750
rect 368061 1033750 368189 1034750
rect 368277 1033750 368405 1034750
rect 368493 1033750 368621 1034750
rect 368709 1033750 368837 1034750
rect 368925 1033750 368981 1034750
rect 369141 1033750 369197 1034750
rect 369357 1033750 369485 1034750
rect 369573 1033750 369701 1034750
rect 369789 1033750 369917 1034750
rect 370005 1033750 370133 1034750
rect 370221 1033750 370277 1034750
rect 370437 1033750 370565 1034750
rect 370653 1033750 370781 1034750
rect 370869 1033750 370997 1034750
rect 371085 1033750 371135 1034750
rect 371201 1033750 371251 1034750
rect 371411 1033750 371461 1034750
rect 371527 1033750 371577 1034750
rect 371737 1033750 371787 1034750
rect 371853 1033750 371903 1034750
rect 372063 1033750 372113 1034750
rect 372176 1034565 372188 1034765
rect 372179 1033750 372229 1034350
rect 372429 1033750 372485 1034350
rect 372585 1033750 372713 1034350
rect 372741 1033750 372797 1034350
rect 372897 1033750 373025 1034350
rect 373053 1033750 373103 1034350
rect 373169 1033750 373219 1034750
rect 373319 1033750 373375 1034750
rect 373475 1033750 373525 1034750
rect 373603 1033750 373653 1034750
rect 373753 1033750 373881 1034750
rect 373909 1033750 374037 1034750
rect 374065 1033750 374121 1034750
rect 374221 1033750 374349 1034750
rect 374377 1033750 374505 1034750
rect 374533 1033750 374661 1034750
rect 374689 1033750 374739 1034750
rect 374805 1033750 374855 1034750
rect 374955 1033750 375083 1034750
rect 375111 1033750 375239 1034750
rect 375267 1033750 375395 1034750
rect 375423 1033750 375479 1034750
rect 375579 1033750 375707 1034750
rect 375735 1033750 375863 1034750
rect 375891 1033750 375947 1034750
rect 376047 1033750 376097 1034750
rect 377318 1034550 377371 1034750
rect 377321 1033750 377371 1034550
rect 377531 1033750 377659 1034750
rect 377747 1033750 377803 1034750
rect 377963 1033750 378091 1034750
rect 378179 1033750 378229 1034750
rect 378295 1033750 378345 1034750
rect 378505 1033750 378555 1034750
rect 413754 1034726 413924 1034781
rect 413822 1034686 413924 1034726
rect 413822 1034645 413856 1034686
rect 415056 1034645 415090 1034752
rect 414131 1034425 414731 1034475
rect 414131 1034175 414731 1034225
rect 426213 1033750 426229 1034750
rect 426295 1033750 426345 1034750
rect 426505 1033750 426555 1034750
rect 465754 1034726 465924 1034781
rect 466988 1034726 467157 1034794
rect 517041 1034781 518959 1034863
rect 569041 1034781 570959 1034863
rect 465822 1034686 465924 1034726
rect 467056 1034686 467157 1034726
rect 465822 1034645 465856 1034686
rect 467056 1034645 467090 1034686
rect 466131 1034425 466731 1034475
rect 466131 1034175 466731 1034225
rect 467851 1033750 467901 1034750
rect 468061 1033750 468189 1034750
rect 468277 1033750 468405 1034750
rect 468493 1033750 468621 1034750
rect 468709 1033750 468837 1034750
rect 468925 1033750 468981 1034750
rect 469141 1033750 469197 1034750
rect 469357 1033750 469485 1034750
rect 469573 1033750 469701 1034750
rect 469789 1033750 469917 1034750
rect 470005 1033750 470133 1034750
rect 470221 1033750 470277 1034750
rect 470437 1033750 470565 1034750
rect 470653 1033750 470781 1034750
rect 470869 1033750 470997 1034750
rect 471085 1033750 471135 1034750
rect 471201 1033750 471251 1034750
rect 471411 1033750 471461 1034750
rect 471527 1033750 471577 1034750
rect 471737 1033750 471787 1034750
rect 471853 1033750 471903 1034750
rect 472063 1033750 472113 1034750
rect 472176 1034565 472188 1034765
rect 472179 1033750 472229 1034350
rect 472429 1033750 472485 1034350
rect 472585 1033750 472713 1034350
rect 472741 1033750 472797 1034350
rect 472897 1033750 473025 1034350
rect 473053 1033750 473103 1034350
rect 473169 1033750 473219 1034750
rect 473319 1033750 473375 1034750
rect 473475 1033750 473525 1034750
rect 473603 1033750 473653 1034750
rect 473753 1033750 473881 1034750
rect 473909 1033750 474037 1034750
rect 474065 1033750 474121 1034750
rect 474221 1033750 474349 1034750
rect 474377 1033750 474505 1034750
rect 474533 1033750 474661 1034750
rect 474689 1033750 474739 1034750
rect 474805 1033750 474855 1034750
rect 474955 1033750 475083 1034750
rect 475111 1033750 475239 1034750
rect 475267 1033750 475395 1034750
rect 475423 1033750 475479 1034750
rect 475579 1033750 475707 1034750
rect 475735 1033750 475863 1034750
rect 475891 1033750 475947 1034750
rect 476047 1033750 476097 1034750
rect 477318 1034550 477371 1034750
rect 477321 1033750 477371 1034550
rect 477531 1033750 477659 1034750
rect 477747 1033750 477803 1034750
rect 477963 1033750 478091 1034750
rect 478179 1033750 478229 1034750
rect 478295 1033750 478345 1034750
rect 478505 1033750 478555 1034750
rect 517754 1034726 517924 1034781
rect 517822 1034686 517924 1034726
rect 517822 1034645 517856 1034686
rect 519056 1034645 519090 1034752
rect 518131 1034425 518731 1034475
rect 518131 1034175 518731 1034225
rect 530213 1033750 530229 1034750
rect 530295 1033750 530345 1034750
rect 530505 1033750 530555 1034750
rect 569754 1034726 569924 1034781
rect 570988 1034726 571157 1034794
rect 569822 1034686 569924 1034726
rect 571056 1034686 571157 1034726
rect 569822 1034645 569856 1034686
rect 571056 1034645 571090 1034686
rect 570131 1034425 570731 1034475
rect 570131 1034175 570731 1034225
rect 571851 1033750 571901 1034750
rect 572061 1033750 572189 1034750
rect 572277 1033750 572405 1034750
rect 572493 1033750 572621 1034750
rect 572709 1033750 572837 1034750
rect 572925 1033750 572981 1034750
rect 573141 1033750 573197 1034750
rect 573357 1033750 573485 1034750
rect 573573 1033750 573701 1034750
rect 573789 1033750 573917 1034750
rect 574005 1033750 574133 1034750
rect 574221 1033750 574277 1034750
rect 574437 1033750 574565 1034750
rect 574653 1033750 574781 1034750
rect 574869 1033750 574997 1034750
rect 575085 1033750 575135 1034750
rect 575201 1033750 575251 1034750
rect 575411 1033750 575461 1034750
rect 575527 1033750 575577 1034750
rect 575737 1033750 575787 1034750
rect 575853 1033750 575903 1034750
rect 576063 1033750 576113 1034750
rect 576176 1034565 576188 1034765
rect 576179 1033750 576229 1034350
rect 576429 1033750 576485 1034350
rect 576585 1033750 576713 1034350
rect 576741 1033750 576797 1034350
rect 576897 1033750 577025 1034350
rect 577053 1033750 577103 1034350
rect 577169 1033750 577219 1034750
rect 577319 1033750 577375 1034750
rect 577475 1033750 577525 1034750
rect 577603 1033750 577653 1034750
rect 577753 1033750 577881 1034750
rect 577909 1033750 578037 1034750
rect 578065 1033750 578121 1034750
rect 578221 1033750 578349 1034750
rect 578377 1033750 578505 1034750
rect 578533 1033750 578661 1034750
rect 578689 1033750 578739 1034750
rect 578805 1033750 578855 1034750
rect 578955 1033750 579083 1034750
rect 579111 1033750 579239 1034750
rect 579267 1033750 579395 1034750
rect 579423 1033750 579479 1034750
rect 579579 1033750 579707 1034750
rect 579735 1033750 579863 1034750
rect 579891 1033750 579947 1034750
rect 580047 1033750 580097 1034750
rect 581318 1034550 581371 1034750
rect 581321 1033750 581371 1034550
rect 581531 1033750 581659 1034750
rect 581747 1033750 581803 1034750
rect 581963 1033750 582091 1034750
rect 582179 1033750 582229 1034750
rect 582295 1033750 582345 1034750
rect 582505 1033750 582555 1034750
rect 72042 1033663 72078 1033674
rect 72194 1033663 74518 1033674
rect 72042 1033641 74518 1033663
rect 172042 1033663 172078 1033674
rect 172194 1033663 174518 1033674
rect 172042 1033641 174518 1033663
rect 376042 1033663 376078 1033674
rect 376194 1033663 378518 1033674
rect 376042 1033641 378518 1033663
rect 476042 1033663 476078 1033674
rect 476194 1033663 478518 1033674
rect 476042 1033641 478518 1033663
rect 580042 1033663 580078 1033674
rect 580194 1033663 582518 1033674
rect 580042 1033641 582518 1033663
rect 72042 1033640 72078 1033641
rect 72194 1033640 74518 1033641
rect 122213 1033640 122518 1033641
rect 172042 1033640 172078 1033641
rect 172194 1033640 174518 1033641
rect 226213 1033640 226518 1033641
rect 274213 1033640 274518 1033641
rect 326213 1033640 326518 1033641
rect 376042 1033640 376078 1033641
rect 376194 1033640 378518 1033641
rect 426213 1033640 426518 1033641
rect 476042 1033640 476078 1033641
rect 476194 1033640 478518 1033641
rect 530213 1033640 530518 1033641
rect 580042 1033640 580078 1033641
rect 580194 1033640 582518 1033641
rect 67104 1032409 74218 1032431
rect 62430 1032062 63430 1032112
rect 63540 1032062 64540 1032112
rect 64661 1032062 65661 1032112
rect 65782 1032062 66782 1032112
rect 67339 1032062 68339 1032112
rect 68460 1032062 69460 1032112
rect 69581 1032062 70581 1032112
rect 70691 1032062 71691 1032112
rect 71812 1032062 72812 1032112
rect 72933 1032062 73933 1032112
rect 62430 1031892 63430 1031942
rect 63540 1031892 64540 1031942
rect 64661 1031892 65661 1031942
rect 65782 1031892 66782 1031942
rect 67339 1031892 68339 1031942
rect 68460 1031892 69460 1031942
rect 69581 1031892 70581 1031942
rect 70691 1031892 71691 1031942
rect 71812 1031892 72812 1031942
rect 72933 1031892 73933 1031942
rect 62035 1031629 62170 1031633
rect 67044 1031629 67078 1031633
rect 74147 1031629 74286 1031663
rect 62035 1031605 74286 1031629
rect 76050 1031619 76064 1032463
rect 122213 1032409 122218 1032431
rect 110430 1032062 111253 1032112
rect 110430 1031892 111253 1031942
rect 124050 1031619 124064 1032463
rect 167104 1032409 174218 1032431
rect 162430 1032062 163430 1032112
rect 163540 1032062 164540 1032112
rect 164661 1032062 165661 1032112
rect 165782 1032062 166782 1032112
rect 167339 1032062 168339 1032112
rect 168460 1032062 169460 1032112
rect 169581 1032062 170581 1032112
rect 170691 1032062 171691 1032112
rect 171812 1032062 172812 1032112
rect 172933 1032062 173933 1032112
rect 162430 1031892 163430 1031942
rect 163540 1031892 164540 1031942
rect 164661 1031892 165661 1031942
rect 165782 1031892 166782 1031942
rect 167339 1031892 168339 1031942
rect 168460 1031892 169460 1031942
rect 169581 1031892 170581 1031942
rect 170691 1031892 171691 1031942
rect 171812 1031892 172812 1031942
rect 172933 1031892 173933 1031942
rect 76040 1031605 76064 1031619
rect 124040 1031605 124064 1031619
rect 62035 1031595 76064 1031605
rect 62034 1031579 76064 1031595
rect 110034 1031579 111253 1031595
rect 122213 1031579 122228 1031595
rect 122258 1031579 124064 1031605
rect 162035 1031629 162170 1031633
rect 167044 1031629 167078 1031633
rect 174147 1031629 174286 1031663
rect 162035 1031605 174286 1031629
rect 176050 1031619 176064 1032463
rect 226213 1032409 226218 1032431
rect 214430 1032062 215253 1032112
rect 214430 1031892 215253 1031942
rect 228050 1031619 228064 1032463
rect 274213 1032409 274218 1032431
rect 276050 1031619 276064 1032463
rect 326213 1032409 326218 1032431
rect 314430 1032062 315253 1032112
rect 314430 1031892 315253 1031942
rect 328050 1031619 328064 1032463
rect 371104 1032409 378218 1032431
rect 366430 1032062 367430 1032112
rect 367540 1032062 368540 1032112
rect 368661 1032062 369661 1032112
rect 369782 1032062 370782 1032112
rect 371339 1032062 372339 1032112
rect 372460 1032062 373460 1032112
rect 373581 1032062 374581 1032112
rect 374691 1032062 375691 1032112
rect 375812 1032062 376812 1032112
rect 376933 1032062 377933 1032112
rect 366430 1031892 367430 1031942
rect 367540 1031892 368540 1031942
rect 368661 1031892 369661 1031942
rect 369782 1031892 370782 1031942
rect 371339 1031892 372339 1031942
rect 372460 1031892 373460 1031942
rect 373581 1031892 374581 1031942
rect 374691 1031892 375691 1031942
rect 375812 1031892 376812 1031942
rect 376933 1031892 377933 1031942
rect 176040 1031605 176064 1031619
rect 228040 1031605 228064 1031619
rect 276040 1031605 276064 1031619
rect 328040 1031605 328064 1031619
rect 162035 1031595 176064 1031605
rect 162034 1031579 176064 1031595
rect 214034 1031579 215253 1031595
rect 226213 1031579 226228 1031595
rect 226258 1031579 228064 1031605
rect 262034 1031579 262080 1031595
rect 274213 1031579 274228 1031595
rect 274258 1031579 276064 1031605
rect 314034 1031579 315253 1031595
rect 326213 1031579 326228 1031595
rect 326258 1031579 328064 1031605
rect 366035 1031629 366170 1031633
rect 371044 1031629 371078 1031633
rect 378147 1031629 378286 1031663
rect 366035 1031605 378286 1031629
rect 380050 1031619 380064 1032463
rect 426213 1032409 426218 1032431
rect 414430 1032062 415253 1032112
rect 414430 1031892 415253 1031942
rect 428050 1031619 428064 1032463
rect 471104 1032409 478218 1032431
rect 466430 1032062 467430 1032112
rect 467540 1032062 468540 1032112
rect 468661 1032062 469661 1032112
rect 469782 1032062 470782 1032112
rect 471339 1032062 472339 1032112
rect 472460 1032062 473460 1032112
rect 473581 1032062 474581 1032112
rect 474691 1032062 475691 1032112
rect 475812 1032062 476812 1032112
rect 476933 1032062 477933 1032112
rect 466430 1031892 467430 1031942
rect 467540 1031892 468540 1031942
rect 468661 1031892 469661 1031942
rect 469782 1031892 470782 1031942
rect 471339 1031892 472339 1031942
rect 472460 1031892 473460 1031942
rect 473581 1031892 474581 1031942
rect 474691 1031892 475691 1031942
rect 475812 1031892 476812 1031942
rect 476933 1031892 477933 1031942
rect 380040 1031605 380064 1031619
rect 428040 1031605 428064 1031619
rect 366035 1031595 380064 1031605
rect 366034 1031579 380064 1031595
rect 414034 1031579 415253 1031595
rect 426213 1031579 426228 1031595
rect 426258 1031579 428064 1031605
rect 466035 1031629 466170 1031633
rect 471044 1031629 471078 1031633
rect 478147 1031629 478286 1031663
rect 466035 1031605 478286 1031629
rect 480050 1031619 480064 1032463
rect 530213 1032409 530218 1032431
rect 518430 1032062 519253 1032112
rect 518430 1031892 519253 1031942
rect 532050 1031619 532064 1032463
rect 575104 1032409 582218 1032431
rect 570430 1032062 571430 1032112
rect 571540 1032062 572540 1032112
rect 572661 1032062 573661 1032112
rect 573782 1032062 574782 1032112
rect 575339 1032062 576339 1032112
rect 576460 1032062 577460 1032112
rect 577581 1032062 578581 1032112
rect 578691 1032062 579691 1032112
rect 579812 1032062 580812 1032112
rect 580933 1032062 581933 1032112
rect 570430 1031892 571430 1031942
rect 571540 1031892 572540 1031942
rect 572661 1031892 573661 1031942
rect 573782 1031892 574782 1031942
rect 575339 1031892 576339 1031942
rect 576460 1031892 577460 1031942
rect 577581 1031892 578581 1031942
rect 578691 1031892 579691 1031942
rect 579812 1031892 580812 1031942
rect 580933 1031892 581933 1031942
rect 480040 1031605 480064 1031619
rect 532040 1031605 532064 1031619
rect 466035 1031595 480064 1031605
rect 466034 1031579 480064 1031595
rect 518034 1031579 519253 1031595
rect 530213 1031579 530228 1031595
rect 530258 1031579 532064 1031605
rect 570035 1031629 570170 1031633
rect 575044 1031629 575078 1031633
rect 582147 1031629 582286 1031663
rect 570035 1031605 582286 1031629
rect 584050 1031619 584064 1032463
rect 584040 1031605 584064 1031619
rect 570035 1031595 584064 1031605
rect 570034 1031579 584064 1031595
rect 62035 1031541 74215 1031579
rect 74218 1031541 74228 1031579
rect 162035 1031541 174215 1031579
rect 174218 1031541 174228 1031579
rect 366035 1031541 378215 1031579
rect 378218 1031541 378228 1031579
rect 466035 1031541 478215 1031579
rect 478218 1031541 478228 1031579
rect 570035 1031541 582215 1031579
rect 582218 1031541 582228 1031579
rect 62657 1030211 62867 1030247
rect 74919 1030211 75032 1030247
rect 75481 1030211 75763 1030247
rect 123481 1030211 123763 1030247
rect 162657 1030211 162867 1030247
rect 174919 1030211 175032 1030247
rect 175481 1030211 175763 1030247
rect 227481 1030211 227763 1030247
rect 275481 1030211 275763 1030247
rect 327481 1030211 327763 1030247
rect 366657 1030211 366867 1030247
rect 378919 1030211 379032 1030247
rect 379481 1030211 379763 1030247
rect 427481 1030211 427763 1030247
rect 466657 1030211 466867 1030247
rect 478919 1030211 479032 1030247
rect 479481 1030211 479763 1030247
rect 531481 1030211 531763 1030247
rect 570657 1030211 570867 1030247
rect 582919 1030211 583032 1030247
rect 583481 1030211 583763 1030247
rect 62246 1029211 62324 1030211
rect 62446 1029211 62518 1030211
rect 62669 1029211 62697 1030211
rect 62734 1029211 62790 1030211
rect 62831 1029211 62867 1030211
rect 62881 1029211 62885 1030211
rect 63092 1029211 63152 1030211
rect 63352 1029211 63424 1030211
rect 63654 1029211 63710 1030211
rect 63726 1029211 63782 1030211
rect 64084 1029211 64144 1030211
rect 64344 1029211 64416 1030211
rect 64646 1029211 64702 1030211
rect 64718 1029211 64774 1030211
rect 65076 1029211 65136 1030211
rect 65336 1029211 65408 1030211
rect 65638 1029211 65694 1030211
rect 65710 1029211 65766 1030211
rect 66068 1029211 66128 1030211
rect 66328 1029211 66400 1030211
rect 66630 1029211 66686 1030211
rect 66702 1029211 66758 1030211
rect 67060 1029211 67120 1030211
rect 67320 1029211 67392 1030211
rect 67622 1029211 67678 1030211
rect 67694 1029211 67750 1030211
rect 68052 1029211 68112 1030211
rect 68312 1029211 68384 1030211
rect 68614 1029211 68670 1030211
rect 68686 1029211 68742 1030211
rect 69044 1029211 69104 1030211
rect 69304 1029211 69376 1030211
rect 69606 1029211 69662 1030211
rect 69678 1029211 69734 1030211
rect 70036 1029211 70096 1030211
rect 70296 1029211 70368 1030211
rect 70598 1029211 70654 1030211
rect 70670 1029211 70726 1030211
rect 71028 1029211 71088 1030211
rect 71288 1029211 71360 1030211
rect 71590 1029211 71646 1030211
rect 71662 1029211 71718 1030211
rect 72020 1029211 72080 1030211
rect 72280 1029211 72352 1030211
rect 72582 1029211 72638 1030211
rect 72654 1029211 72710 1030211
rect 73012 1029211 73072 1030211
rect 73272 1029211 73344 1030211
rect 73574 1029211 73630 1030211
rect 73646 1029211 73702 1030211
rect 74004 1029211 74064 1030211
rect 74264 1029211 74336 1030211
rect 74566 1029211 74622 1030211
rect 74638 1029211 74694 1030211
rect 74919 1029211 74959 1030211
rect 74996 1029211 75032 1030211
rect 75256 1029211 75328 1030211
rect 75481 1029211 75521 1030211
rect 75558 1029211 75614 1030211
rect 75630 1029211 75686 1030211
rect 75727 1029211 75763 1030211
rect 75777 1029211 75781 1030211
rect 75974 1029211 76034 1030211
rect 76070 1030194 76174 1030211
rect 110246 1030194 110324 1030211
rect 76070 1030160 76164 1030194
rect 76174 1030160 76208 1030194
rect 110256 1030160 110324 1030194
rect 76070 1030123 76174 1030160
rect 110246 1030123 110324 1030160
rect 76070 1030089 76164 1030123
rect 76174 1030089 76208 1030123
rect 110256 1030089 110324 1030123
rect 76070 1030049 76174 1030089
rect 110246 1030049 110324 1030089
rect 76070 1030015 76164 1030049
rect 76174 1030015 76208 1030049
rect 110256 1030015 110324 1030049
rect 76070 1029978 76174 1030015
rect 110246 1029978 110324 1030015
rect 76070 1029944 76164 1029978
rect 76174 1029944 76208 1029978
rect 110256 1029944 110324 1029978
rect 76070 1029904 76174 1029944
rect 110246 1029904 110324 1029944
rect 76070 1029870 76164 1029904
rect 76174 1029870 76208 1029904
rect 110256 1029870 110324 1029904
rect 76070 1029833 76174 1029870
rect 110246 1029833 110324 1029870
rect 76070 1029799 76164 1029833
rect 76174 1029799 76208 1029833
rect 110256 1029799 110324 1029833
rect 76070 1029759 76174 1029799
rect 110246 1029759 110324 1029799
rect 76070 1029725 76164 1029759
rect 76174 1029725 76208 1029759
rect 110256 1029725 110324 1029759
rect 76070 1029688 76174 1029725
rect 110246 1029688 110324 1029725
rect 76070 1029654 76164 1029688
rect 76174 1029654 76208 1029688
rect 110256 1029654 110324 1029688
rect 76070 1029614 76174 1029654
rect 110246 1029614 110324 1029654
rect 76070 1029580 76164 1029614
rect 76174 1029580 76208 1029614
rect 110256 1029580 110324 1029614
rect 76070 1029543 76174 1029580
rect 110246 1029543 110324 1029580
rect 76070 1029509 76164 1029543
rect 76174 1029509 76208 1029543
rect 110256 1029509 110324 1029543
rect 76070 1029469 76174 1029509
rect 110246 1029469 110324 1029509
rect 76070 1029435 76164 1029469
rect 76174 1029435 76208 1029469
rect 110256 1029435 110324 1029469
rect 76070 1029398 76174 1029435
rect 110246 1029398 110324 1029435
rect 76070 1029364 76164 1029398
rect 76174 1029364 76208 1029398
rect 110256 1029364 110324 1029398
rect 76070 1029304 76174 1029364
rect 110246 1029304 110324 1029364
rect 76070 1029270 76164 1029304
rect 76174 1029270 76208 1029304
rect 110256 1029270 110324 1029304
rect 76070 1029234 76174 1029270
rect 76070 1029211 76198 1029234
rect 110246 1029219 110324 1029270
rect 110256 1029211 110324 1029219
rect 110669 1029211 110693 1030211
rect 110734 1029211 110790 1030211
rect 122566 1029211 122622 1030211
rect 122638 1029211 122694 1030211
rect 123481 1029211 123521 1030211
rect 123558 1029211 123614 1030211
rect 123630 1029211 123686 1030211
rect 123727 1029211 123763 1030211
rect 123777 1029211 123781 1030211
rect 123974 1029211 124034 1030211
rect 124070 1030194 124174 1030211
rect 124070 1030160 124164 1030194
rect 124174 1030160 124208 1030194
rect 124070 1030123 124174 1030160
rect 124070 1030089 124164 1030123
rect 124174 1030089 124208 1030123
rect 124070 1030049 124174 1030089
rect 124070 1030015 124164 1030049
rect 124174 1030015 124208 1030049
rect 124070 1029978 124174 1030015
rect 124070 1029944 124164 1029978
rect 124174 1029944 124208 1029978
rect 124070 1029904 124174 1029944
rect 124070 1029870 124164 1029904
rect 124174 1029870 124208 1029904
rect 124070 1029833 124174 1029870
rect 124070 1029799 124164 1029833
rect 124174 1029799 124208 1029833
rect 124070 1029759 124174 1029799
rect 124070 1029725 124164 1029759
rect 124174 1029725 124208 1029759
rect 124070 1029688 124174 1029725
rect 124070 1029654 124164 1029688
rect 124174 1029654 124208 1029688
rect 124070 1029614 124174 1029654
rect 124070 1029580 124164 1029614
rect 124174 1029580 124208 1029614
rect 124070 1029543 124174 1029580
rect 124070 1029509 124164 1029543
rect 124174 1029509 124208 1029543
rect 124070 1029469 124174 1029509
rect 124070 1029435 124164 1029469
rect 124174 1029435 124208 1029469
rect 124070 1029398 124174 1029435
rect 124070 1029364 124164 1029398
rect 124174 1029364 124208 1029398
rect 124070 1029304 124174 1029364
rect 124070 1029270 124164 1029304
rect 124174 1029270 124208 1029304
rect 124070 1029234 124174 1029270
rect 124070 1029211 124198 1029234
rect 162246 1029211 162324 1030211
rect 162446 1029211 162518 1030211
rect 162669 1029211 162697 1030211
rect 162734 1029211 162790 1030211
rect 162831 1029211 162867 1030211
rect 162881 1029211 162885 1030211
rect 163092 1029211 163152 1030211
rect 163352 1029211 163424 1030211
rect 163654 1029211 163710 1030211
rect 163726 1029211 163782 1030211
rect 164084 1029211 164144 1030211
rect 164344 1029211 164416 1030211
rect 164646 1029211 164702 1030211
rect 164718 1029211 164774 1030211
rect 165076 1029211 165136 1030211
rect 165336 1029211 165408 1030211
rect 165638 1029211 165694 1030211
rect 165710 1029211 165766 1030211
rect 166068 1029211 166128 1030211
rect 166328 1029211 166400 1030211
rect 166630 1029211 166686 1030211
rect 166702 1029211 166758 1030211
rect 167060 1029211 167120 1030211
rect 167320 1029211 167392 1030211
rect 167622 1029211 167678 1030211
rect 167694 1029211 167750 1030211
rect 168052 1029211 168112 1030211
rect 168312 1029211 168384 1030211
rect 168614 1029211 168670 1030211
rect 168686 1029211 168742 1030211
rect 169044 1029211 169104 1030211
rect 169304 1029211 169376 1030211
rect 169606 1029211 169662 1030211
rect 169678 1029211 169734 1030211
rect 170036 1029211 170096 1030211
rect 170296 1029211 170368 1030211
rect 170598 1029211 170654 1030211
rect 170670 1029211 170726 1030211
rect 171028 1029211 171088 1030211
rect 171288 1029211 171360 1030211
rect 171590 1029211 171646 1030211
rect 171662 1029211 171718 1030211
rect 172020 1029211 172080 1030211
rect 172280 1029211 172352 1030211
rect 172582 1029211 172638 1030211
rect 172654 1029211 172710 1030211
rect 173012 1029211 173072 1030211
rect 173272 1029211 173344 1030211
rect 173574 1029211 173630 1030211
rect 173646 1029211 173702 1030211
rect 174004 1029211 174064 1030211
rect 174264 1029211 174336 1030211
rect 174566 1029211 174622 1030211
rect 174638 1029211 174694 1030211
rect 174919 1029211 174959 1030211
rect 174996 1029211 175032 1030211
rect 175256 1029211 175328 1030211
rect 175481 1029211 175521 1030211
rect 175558 1029211 175614 1030211
rect 175630 1029211 175686 1030211
rect 175727 1029211 175763 1030211
rect 175777 1029211 175781 1030211
rect 175974 1029211 176034 1030211
rect 176070 1030194 176174 1030211
rect 214246 1030194 214324 1030211
rect 176070 1030160 176164 1030194
rect 176174 1030160 176208 1030194
rect 214256 1030160 214324 1030194
rect 176070 1030123 176174 1030160
rect 214246 1030123 214324 1030160
rect 176070 1030089 176164 1030123
rect 176174 1030089 176208 1030123
rect 214256 1030089 214324 1030123
rect 176070 1030049 176174 1030089
rect 214246 1030049 214324 1030089
rect 176070 1030015 176164 1030049
rect 176174 1030015 176208 1030049
rect 214256 1030015 214324 1030049
rect 176070 1029978 176174 1030015
rect 214246 1029978 214324 1030015
rect 176070 1029944 176164 1029978
rect 176174 1029944 176208 1029978
rect 214256 1029944 214324 1029978
rect 176070 1029904 176174 1029944
rect 214246 1029904 214324 1029944
rect 176070 1029870 176164 1029904
rect 176174 1029870 176208 1029904
rect 214256 1029870 214324 1029904
rect 176070 1029833 176174 1029870
rect 214246 1029833 214324 1029870
rect 176070 1029799 176164 1029833
rect 176174 1029799 176208 1029833
rect 214256 1029799 214324 1029833
rect 176070 1029759 176174 1029799
rect 214246 1029759 214324 1029799
rect 176070 1029725 176164 1029759
rect 176174 1029725 176208 1029759
rect 214256 1029725 214324 1029759
rect 176070 1029688 176174 1029725
rect 214246 1029688 214324 1029725
rect 176070 1029654 176164 1029688
rect 176174 1029654 176208 1029688
rect 214256 1029654 214324 1029688
rect 176070 1029614 176174 1029654
rect 214246 1029614 214324 1029654
rect 176070 1029580 176164 1029614
rect 176174 1029580 176208 1029614
rect 214256 1029580 214324 1029614
rect 176070 1029543 176174 1029580
rect 214246 1029543 214324 1029580
rect 176070 1029509 176164 1029543
rect 176174 1029509 176208 1029543
rect 214256 1029509 214324 1029543
rect 176070 1029469 176174 1029509
rect 214246 1029469 214324 1029509
rect 176070 1029435 176164 1029469
rect 176174 1029435 176208 1029469
rect 214256 1029435 214324 1029469
rect 176070 1029398 176174 1029435
rect 214246 1029398 214324 1029435
rect 176070 1029364 176164 1029398
rect 176174 1029364 176208 1029398
rect 214256 1029364 214324 1029398
rect 176070 1029304 176174 1029364
rect 214246 1029304 214324 1029364
rect 176070 1029270 176164 1029304
rect 176174 1029270 176208 1029304
rect 214256 1029270 214324 1029304
rect 176070 1029234 176174 1029270
rect 176070 1029211 176198 1029234
rect 214246 1029219 214324 1029270
rect 214256 1029211 214324 1029219
rect 214669 1029211 214693 1030211
rect 214734 1029211 214790 1030211
rect 226566 1029211 226622 1030211
rect 226638 1029211 226694 1030211
rect 227481 1029211 227521 1030211
rect 227558 1029211 227614 1030211
rect 227630 1029211 227686 1030211
rect 227727 1029211 227763 1030211
rect 227777 1029211 227781 1030211
rect 227974 1029211 228034 1030211
rect 228070 1030194 228174 1030211
rect 228070 1030160 228164 1030194
rect 228174 1030160 228208 1030194
rect 228070 1030123 228174 1030160
rect 228070 1030089 228164 1030123
rect 228174 1030089 228208 1030123
rect 228070 1030049 228174 1030089
rect 228070 1030015 228164 1030049
rect 228174 1030015 228208 1030049
rect 228070 1029978 228174 1030015
rect 228070 1029944 228164 1029978
rect 228174 1029944 228208 1029978
rect 228070 1029904 228174 1029944
rect 228070 1029870 228164 1029904
rect 228174 1029870 228208 1029904
rect 228070 1029833 228174 1029870
rect 228070 1029799 228164 1029833
rect 228174 1029799 228208 1029833
rect 228070 1029759 228174 1029799
rect 228070 1029725 228164 1029759
rect 228174 1029725 228208 1029759
rect 228070 1029688 228174 1029725
rect 228070 1029654 228164 1029688
rect 228174 1029654 228208 1029688
rect 228070 1029614 228174 1029654
rect 228070 1029580 228164 1029614
rect 228174 1029580 228208 1029614
rect 228070 1029543 228174 1029580
rect 228070 1029509 228164 1029543
rect 228174 1029509 228208 1029543
rect 228070 1029469 228174 1029509
rect 228070 1029435 228164 1029469
rect 228174 1029435 228208 1029469
rect 228070 1029398 228174 1029435
rect 228070 1029364 228164 1029398
rect 228174 1029364 228208 1029398
rect 228070 1029304 228174 1029364
rect 228070 1029270 228164 1029304
rect 228174 1029270 228208 1029304
rect 228070 1029234 228174 1029270
rect 228070 1029211 228198 1029234
rect 274566 1029211 274622 1030211
rect 274638 1029211 274694 1030211
rect 275481 1029211 275521 1030211
rect 275558 1029211 275614 1030211
rect 275630 1029211 275686 1030211
rect 275727 1029211 275763 1030211
rect 275777 1029211 275781 1030211
rect 275974 1029211 276034 1030211
rect 276070 1030194 276174 1030211
rect 314246 1030194 314324 1030211
rect 276070 1030160 276164 1030194
rect 276174 1030160 276208 1030194
rect 314256 1030160 314324 1030194
rect 276070 1030123 276174 1030160
rect 314246 1030123 314324 1030160
rect 276070 1030089 276164 1030123
rect 276174 1030089 276208 1030123
rect 314256 1030089 314324 1030123
rect 276070 1030049 276174 1030089
rect 314246 1030049 314324 1030089
rect 276070 1030015 276164 1030049
rect 276174 1030015 276208 1030049
rect 314256 1030015 314324 1030049
rect 276070 1029978 276174 1030015
rect 314246 1029978 314324 1030015
rect 276070 1029944 276164 1029978
rect 276174 1029944 276208 1029978
rect 314256 1029944 314324 1029978
rect 276070 1029904 276174 1029944
rect 314246 1029904 314324 1029944
rect 276070 1029870 276164 1029904
rect 276174 1029870 276208 1029904
rect 314256 1029870 314324 1029904
rect 276070 1029833 276174 1029870
rect 314246 1029833 314324 1029870
rect 276070 1029799 276164 1029833
rect 276174 1029799 276208 1029833
rect 314256 1029799 314324 1029833
rect 276070 1029759 276174 1029799
rect 314246 1029759 314324 1029799
rect 276070 1029725 276164 1029759
rect 276174 1029725 276208 1029759
rect 314256 1029725 314324 1029759
rect 276070 1029688 276174 1029725
rect 314246 1029688 314324 1029725
rect 276070 1029654 276164 1029688
rect 276174 1029654 276208 1029688
rect 314256 1029654 314324 1029688
rect 276070 1029614 276174 1029654
rect 314246 1029614 314324 1029654
rect 276070 1029580 276164 1029614
rect 276174 1029580 276208 1029614
rect 314256 1029580 314324 1029614
rect 276070 1029543 276174 1029580
rect 314246 1029543 314324 1029580
rect 276070 1029509 276164 1029543
rect 276174 1029509 276208 1029543
rect 314256 1029509 314324 1029543
rect 276070 1029469 276174 1029509
rect 314246 1029469 314324 1029509
rect 276070 1029435 276164 1029469
rect 276174 1029435 276208 1029469
rect 314256 1029435 314324 1029469
rect 276070 1029398 276174 1029435
rect 314246 1029398 314324 1029435
rect 276070 1029364 276164 1029398
rect 276174 1029364 276208 1029398
rect 314256 1029364 314324 1029398
rect 276070 1029304 276174 1029364
rect 314246 1029304 314324 1029364
rect 276070 1029270 276164 1029304
rect 276174 1029270 276208 1029304
rect 314256 1029270 314324 1029304
rect 276070 1029234 276174 1029270
rect 276070 1029211 276198 1029234
rect 314246 1029219 314324 1029270
rect 314256 1029211 314324 1029219
rect 314669 1029211 314693 1030211
rect 314734 1029211 314790 1030211
rect 326566 1029211 326622 1030211
rect 326638 1029211 326694 1030211
rect 327481 1029211 327521 1030211
rect 327558 1029211 327614 1030211
rect 327630 1029211 327686 1030211
rect 327727 1029211 327763 1030211
rect 327777 1029211 327781 1030211
rect 327974 1029211 328034 1030211
rect 328070 1030194 328174 1030211
rect 328070 1030160 328164 1030194
rect 328174 1030160 328208 1030194
rect 328070 1030123 328174 1030160
rect 328070 1030089 328164 1030123
rect 328174 1030089 328208 1030123
rect 328070 1030049 328174 1030089
rect 328070 1030015 328164 1030049
rect 328174 1030015 328208 1030049
rect 328070 1029978 328174 1030015
rect 328070 1029944 328164 1029978
rect 328174 1029944 328208 1029978
rect 328070 1029904 328174 1029944
rect 328070 1029870 328164 1029904
rect 328174 1029870 328208 1029904
rect 328070 1029833 328174 1029870
rect 328070 1029799 328164 1029833
rect 328174 1029799 328208 1029833
rect 328070 1029759 328174 1029799
rect 328070 1029725 328164 1029759
rect 328174 1029725 328208 1029759
rect 328070 1029688 328174 1029725
rect 328070 1029654 328164 1029688
rect 328174 1029654 328208 1029688
rect 328070 1029614 328174 1029654
rect 328070 1029580 328164 1029614
rect 328174 1029580 328208 1029614
rect 328070 1029543 328174 1029580
rect 328070 1029509 328164 1029543
rect 328174 1029509 328208 1029543
rect 328070 1029469 328174 1029509
rect 328070 1029435 328164 1029469
rect 328174 1029435 328208 1029469
rect 328070 1029398 328174 1029435
rect 328070 1029364 328164 1029398
rect 328174 1029364 328208 1029398
rect 328070 1029304 328174 1029364
rect 328070 1029270 328164 1029304
rect 328174 1029270 328208 1029304
rect 328070 1029234 328174 1029270
rect 328070 1029211 328198 1029234
rect 366246 1029211 366324 1030211
rect 366446 1029211 366518 1030211
rect 366669 1029211 366697 1030211
rect 366734 1029211 366790 1030211
rect 366831 1029211 366867 1030211
rect 366881 1029211 366885 1030211
rect 367092 1029211 367152 1030211
rect 367352 1029211 367424 1030211
rect 367654 1029211 367710 1030211
rect 367726 1029211 367782 1030211
rect 368084 1029211 368144 1030211
rect 368344 1029211 368416 1030211
rect 368646 1029211 368702 1030211
rect 368718 1029211 368774 1030211
rect 369076 1029211 369136 1030211
rect 369336 1029211 369408 1030211
rect 369638 1029211 369694 1030211
rect 369710 1029211 369766 1030211
rect 370068 1029211 370128 1030211
rect 370328 1029211 370400 1030211
rect 370630 1029211 370686 1030211
rect 370702 1029211 370758 1030211
rect 371060 1029211 371120 1030211
rect 371320 1029211 371392 1030211
rect 371622 1029211 371678 1030211
rect 371694 1029211 371750 1030211
rect 372052 1029211 372112 1030211
rect 372312 1029211 372384 1030211
rect 372614 1029211 372670 1030211
rect 372686 1029211 372742 1030211
rect 373044 1029211 373104 1030211
rect 373304 1029211 373376 1030211
rect 373606 1029211 373662 1030211
rect 373678 1029211 373734 1030211
rect 374036 1029211 374096 1030211
rect 374296 1029211 374368 1030211
rect 374598 1029211 374654 1030211
rect 374670 1029211 374726 1030211
rect 375028 1029211 375088 1030211
rect 375288 1029211 375360 1030211
rect 375590 1029211 375646 1030211
rect 375662 1029211 375718 1030211
rect 376020 1029211 376080 1030211
rect 376280 1029211 376352 1030211
rect 376582 1029211 376638 1030211
rect 376654 1029211 376710 1030211
rect 377012 1029211 377072 1030211
rect 377272 1029211 377344 1030211
rect 377574 1029211 377630 1030211
rect 377646 1029211 377702 1030211
rect 378004 1029211 378064 1030211
rect 378264 1029211 378336 1030211
rect 378566 1029211 378622 1030211
rect 378638 1029211 378694 1030211
rect 378919 1029211 378959 1030211
rect 378996 1029211 379032 1030211
rect 379256 1029211 379328 1030211
rect 379481 1029211 379521 1030211
rect 379558 1029211 379614 1030211
rect 379630 1029211 379686 1030211
rect 379727 1029211 379763 1030211
rect 379777 1029211 379781 1030211
rect 379974 1029211 380034 1030211
rect 380070 1030194 380174 1030211
rect 414246 1030194 414324 1030211
rect 380070 1030160 380164 1030194
rect 380174 1030160 380208 1030194
rect 414256 1030160 414324 1030194
rect 380070 1030123 380174 1030160
rect 414246 1030123 414324 1030160
rect 380070 1030089 380164 1030123
rect 380174 1030089 380208 1030123
rect 414256 1030089 414324 1030123
rect 380070 1030049 380174 1030089
rect 414246 1030049 414324 1030089
rect 380070 1030015 380164 1030049
rect 380174 1030015 380208 1030049
rect 414256 1030015 414324 1030049
rect 380070 1029978 380174 1030015
rect 414246 1029978 414324 1030015
rect 380070 1029944 380164 1029978
rect 380174 1029944 380208 1029978
rect 414256 1029944 414324 1029978
rect 380070 1029904 380174 1029944
rect 414246 1029904 414324 1029944
rect 380070 1029870 380164 1029904
rect 380174 1029870 380208 1029904
rect 414256 1029870 414324 1029904
rect 380070 1029833 380174 1029870
rect 414246 1029833 414324 1029870
rect 380070 1029799 380164 1029833
rect 380174 1029799 380208 1029833
rect 414256 1029799 414324 1029833
rect 380070 1029759 380174 1029799
rect 414246 1029759 414324 1029799
rect 380070 1029725 380164 1029759
rect 380174 1029725 380208 1029759
rect 414256 1029725 414324 1029759
rect 380070 1029688 380174 1029725
rect 414246 1029688 414324 1029725
rect 380070 1029654 380164 1029688
rect 380174 1029654 380208 1029688
rect 414256 1029654 414324 1029688
rect 380070 1029614 380174 1029654
rect 414246 1029614 414324 1029654
rect 380070 1029580 380164 1029614
rect 380174 1029580 380208 1029614
rect 414256 1029580 414324 1029614
rect 380070 1029543 380174 1029580
rect 414246 1029543 414324 1029580
rect 380070 1029509 380164 1029543
rect 380174 1029509 380208 1029543
rect 414256 1029509 414324 1029543
rect 380070 1029469 380174 1029509
rect 414246 1029469 414324 1029509
rect 380070 1029435 380164 1029469
rect 380174 1029435 380208 1029469
rect 414256 1029435 414324 1029469
rect 380070 1029398 380174 1029435
rect 414246 1029398 414324 1029435
rect 380070 1029364 380164 1029398
rect 380174 1029364 380208 1029398
rect 414256 1029364 414324 1029398
rect 380070 1029304 380174 1029364
rect 414246 1029304 414324 1029364
rect 380070 1029270 380164 1029304
rect 380174 1029270 380208 1029304
rect 414256 1029270 414324 1029304
rect 380070 1029234 380174 1029270
rect 380070 1029211 380198 1029234
rect 414246 1029219 414324 1029270
rect 414256 1029211 414324 1029219
rect 414669 1029211 414693 1030211
rect 414734 1029211 414790 1030211
rect 426566 1029211 426622 1030211
rect 426638 1029211 426694 1030211
rect 427481 1029211 427521 1030211
rect 427558 1029211 427614 1030211
rect 427630 1029211 427686 1030211
rect 427727 1029211 427763 1030211
rect 427777 1029211 427781 1030211
rect 427974 1029211 428034 1030211
rect 428070 1030194 428174 1030211
rect 428070 1030160 428164 1030194
rect 428174 1030160 428208 1030194
rect 428070 1030123 428174 1030160
rect 428070 1030089 428164 1030123
rect 428174 1030089 428208 1030123
rect 428070 1030049 428174 1030089
rect 428070 1030015 428164 1030049
rect 428174 1030015 428208 1030049
rect 428070 1029978 428174 1030015
rect 428070 1029944 428164 1029978
rect 428174 1029944 428208 1029978
rect 428070 1029904 428174 1029944
rect 428070 1029870 428164 1029904
rect 428174 1029870 428208 1029904
rect 428070 1029833 428174 1029870
rect 428070 1029799 428164 1029833
rect 428174 1029799 428208 1029833
rect 428070 1029759 428174 1029799
rect 428070 1029725 428164 1029759
rect 428174 1029725 428208 1029759
rect 428070 1029688 428174 1029725
rect 428070 1029654 428164 1029688
rect 428174 1029654 428208 1029688
rect 428070 1029614 428174 1029654
rect 428070 1029580 428164 1029614
rect 428174 1029580 428208 1029614
rect 428070 1029543 428174 1029580
rect 428070 1029509 428164 1029543
rect 428174 1029509 428208 1029543
rect 428070 1029469 428174 1029509
rect 428070 1029435 428164 1029469
rect 428174 1029435 428208 1029469
rect 428070 1029398 428174 1029435
rect 428070 1029364 428164 1029398
rect 428174 1029364 428208 1029398
rect 428070 1029304 428174 1029364
rect 428070 1029270 428164 1029304
rect 428174 1029270 428208 1029304
rect 428070 1029234 428174 1029270
rect 428070 1029211 428198 1029234
rect 466246 1029211 466324 1030211
rect 466446 1029211 466518 1030211
rect 466669 1029211 466697 1030211
rect 466734 1029211 466790 1030211
rect 466831 1029211 466867 1030211
rect 466881 1029211 466885 1030211
rect 467092 1029211 467152 1030211
rect 467352 1029211 467424 1030211
rect 467654 1029211 467710 1030211
rect 467726 1029211 467782 1030211
rect 468084 1029211 468144 1030211
rect 468344 1029211 468416 1030211
rect 468646 1029211 468702 1030211
rect 468718 1029211 468774 1030211
rect 469076 1029211 469136 1030211
rect 469336 1029211 469408 1030211
rect 469638 1029211 469694 1030211
rect 469710 1029211 469766 1030211
rect 470068 1029211 470128 1030211
rect 470328 1029211 470400 1030211
rect 470630 1029211 470686 1030211
rect 470702 1029211 470758 1030211
rect 471060 1029211 471120 1030211
rect 471320 1029211 471392 1030211
rect 471622 1029211 471678 1030211
rect 471694 1029211 471750 1030211
rect 472052 1029211 472112 1030211
rect 472312 1029211 472384 1030211
rect 472614 1029211 472670 1030211
rect 472686 1029211 472742 1030211
rect 473044 1029211 473104 1030211
rect 473304 1029211 473376 1030211
rect 473606 1029211 473662 1030211
rect 473678 1029211 473734 1030211
rect 474036 1029211 474096 1030211
rect 474296 1029211 474368 1030211
rect 474598 1029211 474654 1030211
rect 474670 1029211 474726 1030211
rect 475028 1029211 475088 1030211
rect 475288 1029211 475360 1030211
rect 475590 1029211 475646 1030211
rect 475662 1029211 475718 1030211
rect 476020 1029211 476080 1030211
rect 476280 1029211 476352 1030211
rect 476582 1029211 476638 1030211
rect 476654 1029211 476710 1030211
rect 477012 1029211 477072 1030211
rect 477272 1029211 477344 1030211
rect 477574 1029211 477630 1030211
rect 477646 1029211 477702 1030211
rect 478004 1029211 478064 1030211
rect 478264 1029211 478336 1030211
rect 478566 1029211 478622 1030211
rect 478638 1029211 478694 1030211
rect 478919 1029211 478959 1030211
rect 478996 1029211 479032 1030211
rect 479256 1029211 479328 1030211
rect 479481 1029211 479521 1030211
rect 479558 1029211 479614 1030211
rect 479630 1029211 479686 1030211
rect 479727 1029211 479763 1030211
rect 479777 1029211 479781 1030211
rect 479974 1029211 480034 1030211
rect 480070 1030194 480174 1030211
rect 518246 1030194 518324 1030211
rect 480070 1030160 480164 1030194
rect 480174 1030160 480208 1030194
rect 518256 1030160 518324 1030194
rect 480070 1030123 480174 1030160
rect 518246 1030123 518324 1030160
rect 480070 1030089 480164 1030123
rect 480174 1030089 480208 1030123
rect 518256 1030089 518324 1030123
rect 480070 1030049 480174 1030089
rect 518246 1030049 518324 1030089
rect 480070 1030015 480164 1030049
rect 480174 1030015 480208 1030049
rect 518256 1030015 518324 1030049
rect 480070 1029978 480174 1030015
rect 518246 1029978 518324 1030015
rect 480070 1029944 480164 1029978
rect 480174 1029944 480208 1029978
rect 518256 1029944 518324 1029978
rect 480070 1029904 480174 1029944
rect 518246 1029904 518324 1029944
rect 480070 1029870 480164 1029904
rect 480174 1029870 480208 1029904
rect 518256 1029870 518324 1029904
rect 480070 1029833 480174 1029870
rect 518246 1029833 518324 1029870
rect 480070 1029799 480164 1029833
rect 480174 1029799 480208 1029833
rect 518256 1029799 518324 1029833
rect 480070 1029759 480174 1029799
rect 518246 1029759 518324 1029799
rect 480070 1029725 480164 1029759
rect 480174 1029725 480208 1029759
rect 518256 1029725 518324 1029759
rect 480070 1029688 480174 1029725
rect 518246 1029688 518324 1029725
rect 480070 1029654 480164 1029688
rect 480174 1029654 480208 1029688
rect 518256 1029654 518324 1029688
rect 480070 1029614 480174 1029654
rect 518246 1029614 518324 1029654
rect 480070 1029580 480164 1029614
rect 480174 1029580 480208 1029614
rect 518256 1029580 518324 1029614
rect 480070 1029543 480174 1029580
rect 518246 1029543 518324 1029580
rect 480070 1029509 480164 1029543
rect 480174 1029509 480208 1029543
rect 518256 1029509 518324 1029543
rect 480070 1029469 480174 1029509
rect 518246 1029469 518324 1029509
rect 480070 1029435 480164 1029469
rect 480174 1029435 480208 1029469
rect 518256 1029435 518324 1029469
rect 480070 1029398 480174 1029435
rect 518246 1029398 518324 1029435
rect 480070 1029364 480164 1029398
rect 480174 1029364 480208 1029398
rect 518256 1029364 518324 1029398
rect 480070 1029304 480174 1029364
rect 518246 1029304 518324 1029364
rect 480070 1029270 480164 1029304
rect 480174 1029270 480208 1029304
rect 518256 1029270 518324 1029304
rect 480070 1029234 480174 1029270
rect 480070 1029211 480198 1029234
rect 518246 1029219 518324 1029270
rect 518256 1029211 518324 1029219
rect 518669 1029211 518693 1030211
rect 518734 1029211 518790 1030211
rect 530566 1029211 530622 1030211
rect 530638 1029211 530694 1030211
rect 531481 1029211 531521 1030211
rect 531558 1029211 531614 1030211
rect 531630 1029211 531686 1030211
rect 531727 1029211 531763 1030211
rect 531777 1029211 531781 1030211
rect 531974 1029211 532034 1030211
rect 532070 1030194 532174 1030211
rect 532070 1030160 532164 1030194
rect 532174 1030160 532208 1030194
rect 532070 1030123 532174 1030160
rect 532070 1030089 532164 1030123
rect 532174 1030089 532208 1030123
rect 532070 1030049 532174 1030089
rect 532070 1030015 532164 1030049
rect 532174 1030015 532208 1030049
rect 532070 1029978 532174 1030015
rect 532070 1029944 532164 1029978
rect 532174 1029944 532208 1029978
rect 532070 1029904 532174 1029944
rect 532070 1029870 532164 1029904
rect 532174 1029870 532208 1029904
rect 532070 1029833 532174 1029870
rect 532070 1029799 532164 1029833
rect 532174 1029799 532208 1029833
rect 532070 1029759 532174 1029799
rect 532070 1029725 532164 1029759
rect 532174 1029725 532208 1029759
rect 532070 1029688 532174 1029725
rect 532070 1029654 532164 1029688
rect 532174 1029654 532208 1029688
rect 532070 1029614 532174 1029654
rect 532070 1029580 532164 1029614
rect 532174 1029580 532208 1029614
rect 532070 1029543 532174 1029580
rect 532070 1029509 532164 1029543
rect 532174 1029509 532208 1029543
rect 532070 1029469 532174 1029509
rect 532070 1029435 532164 1029469
rect 532174 1029435 532208 1029469
rect 532070 1029398 532174 1029435
rect 532070 1029364 532164 1029398
rect 532174 1029364 532208 1029398
rect 532070 1029304 532174 1029364
rect 532070 1029270 532164 1029304
rect 532174 1029270 532208 1029304
rect 532070 1029234 532174 1029270
rect 532070 1029211 532198 1029234
rect 570246 1029211 570324 1030211
rect 570446 1029211 570518 1030211
rect 570669 1029211 570697 1030211
rect 570734 1029211 570790 1030211
rect 570831 1029211 570867 1030211
rect 570881 1029211 570885 1030211
rect 571092 1029211 571152 1030211
rect 571352 1029211 571424 1030211
rect 571654 1029211 571710 1030211
rect 571726 1029211 571782 1030211
rect 572084 1029211 572144 1030211
rect 572344 1029211 572416 1030211
rect 572646 1029211 572702 1030211
rect 572718 1029211 572774 1030211
rect 573076 1029211 573136 1030211
rect 573336 1029211 573408 1030211
rect 573638 1029211 573694 1030211
rect 573710 1029211 573766 1030211
rect 574068 1029211 574128 1030211
rect 574328 1029211 574400 1030211
rect 574630 1029211 574686 1030211
rect 574702 1029211 574758 1030211
rect 575060 1029211 575120 1030211
rect 575320 1029211 575392 1030211
rect 575622 1029211 575678 1030211
rect 575694 1029211 575750 1030211
rect 576052 1029211 576112 1030211
rect 576312 1029211 576384 1030211
rect 576614 1029211 576670 1030211
rect 576686 1029211 576742 1030211
rect 577044 1029211 577104 1030211
rect 577304 1029211 577376 1030211
rect 577606 1029211 577662 1030211
rect 577678 1029211 577734 1030211
rect 578036 1029211 578096 1030211
rect 578296 1029211 578368 1030211
rect 578598 1029211 578654 1030211
rect 578670 1029211 578726 1030211
rect 579028 1029211 579088 1030211
rect 579288 1029211 579360 1030211
rect 579590 1029211 579646 1030211
rect 579662 1029211 579718 1030211
rect 580020 1029211 580080 1030211
rect 580280 1029211 580352 1030211
rect 580582 1029211 580638 1030211
rect 580654 1029211 580710 1030211
rect 581012 1029211 581072 1030211
rect 581272 1029211 581344 1030211
rect 581574 1029211 581630 1030211
rect 581646 1029211 581702 1030211
rect 582004 1029211 582064 1030211
rect 582264 1029211 582336 1030211
rect 582566 1029211 582622 1030211
rect 582638 1029211 582694 1030211
rect 582919 1029211 582959 1030211
rect 582996 1029211 583032 1030211
rect 583256 1029211 583328 1030211
rect 583481 1029211 583521 1030211
rect 583558 1029211 583614 1030211
rect 583630 1029211 583686 1030211
rect 583727 1029211 583763 1030211
rect 583777 1029211 583781 1030211
rect 583974 1029211 584034 1030211
rect 584070 1030194 584174 1030211
rect 584070 1030160 584164 1030194
rect 584174 1030160 584208 1030194
rect 584070 1030123 584174 1030160
rect 584070 1030089 584164 1030123
rect 584174 1030089 584208 1030123
rect 584070 1030049 584174 1030089
rect 584070 1030015 584164 1030049
rect 584174 1030015 584208 1030049
rect 584070 1029978 584174 1030015
rect 584070 1029944 584164 1029978
rect 584174 1029944 584208 1029978
rect 584070 1029904 584174 1029944
rect 584070 1029870 584164 1029904
rect 584174 1029870 584208 1029904
rect 584070 1029833 584174 1029870
rect 584070 1029799 584164 1029833
rect 584174 1029799 584208 1029833
rect 584070 1029759 584174 1029799
rect 584070 1029725 584164 1029759
rect 584174 1029725 584208 1029759
rect 584070 1029688 584174 1029725
rect 584070 1029654 584164 1029688
rect 584174 1029654 584208 1029688
rect 584070 1029614 584174 1029654
rect 584070 1029580 584164 1029614
rect 584174 1029580 584208 1029614
rect 584070 1029543 584174 1029580
rect 584070 1029509 584164 1029543
rect 584174 1029509 584208 1029543
rect 584070 1029469 584174 1029509
rect 584070 1029435 584164 1029469
rect 584174 1029435 584208 1029469
rect 584070 1029398 584174 1029435
rect 584070 1029364 584164 1029398
rect 584174 1029364 584208 1029398
rect 584070 1029304 584174 1029364
rect 584070 1029270 584164 1029304
rect 584174 1029270 584208 1029304
rect 584070 1029234 584174 1029270
rect 584070 1029211 584198 1029234
rect 62657 1029175 62867 1029211
rect 74919 1029175 75032 1029211
rect 75481 1029175 75763 1029211
rect 123481 1029175 123763 1029211
rect 162657 1029175 162867 1029211
rect 174919 1029175 175032 1029211
rect 175481 1029175 175763 1029211
rect 227481 1029175 227763 1029211
rect 275481 1029175 275763 1029211
rect 327481 1029175 327763 1029211
rect 366657 1029175 366867 1029211
rect 378919 1029175 379032 1029211
rect 379481 1029175 379763 1029211
rect 427481 1029175 427763 1029211
rect 466657 1029175 466867 1029211
rect 478919 1029175 479032 1029211
rect 479481 1029175 479763 1029211
rect 531481 1029175 531763 1029211
rect 570657 1029175 570867 1029211
rect 582919 1029175 583032 1029211
rect 583481 1029175 583763 1029211
rect 62212 1028638 62256 1028644
rect 62212 1028610 62222 1028638
rect 62246 1028610 62256 1028638
rect 62657 1028610 62867 1028646
rect 74919 1028610 75032 1028646
rect 75481 1028610 75763 1028646
rect 76164 1028610 76174 1028634
rect 123481 1028610 123763 1028646
rect 162212 1028638 162256 1028644
rect 124164 1028610 124174 1028634
rect 162212 1028610 162222 1028638
rect 162246 1028610 162256 1028638
rect 162657 1028610 162867 1028646
rect 174919 1028610 175032 1028646
rect 175481 1028610 175763 1028646
rect 176164 1028610 176174 1028634
rect 227481 1028610 227763 1028646
rect 228164 1028610 228174 1028634
rect 275481 1028610 275763 1028646
rect 276164 1028610 276174 1028634
rect 327481 1028610 327763 1028646
rect 366212 1028638 366256 1028644
rect 328164 1028610 328174 1028634
rect 366212 1028610 366222 1028638
rect 366246 1028610 366256 1028638
rect 366657 1028610 366867 1028646
rect 378919 1028610 379032 1028646
rect 379481 1028610 379763 1028646
rect 380164 1028610 380174 1028634
rect 427481 1028610 427763 1028646
rect 466212 1028638 466256 1028644
rect 428164 1028610 428174 1028634
rect 466212 1028610 466222 1028638
rect 466246 1028610 466256 1028638
rect 466657 1028610 466867 1028646
rect 478919 1028610 479032 1028646
rect 479481 1028610 479763 1028646
rect 480164 1028610 480174 1028634
rect 531481 1028610 531763 1028646
rect 570212 1028638 570256 1028644
rect 532164 1028610 532174 1028634
rect 570212 1028610 570222 1028638
rect 570246 1028610 570256 1028638
rect 570657 1028610 570867 1028646
rect 582919 1028610 583032 1028646
rect 583481 1028610 583763 1028646
rect 584164 1028610 584174 1028634
rect 62246 1027610 62350 1028610
rect 62446 1027610 62518 1028610
rect 62692 1027610 62697 1028610
rect 62734 1027610 62790 1028610
rect 62831 1027610 62832 1028610
rect 63092 1027610 63152 1028610
rect 63352 1027610 63424 1028610
rect 63654 1027610 63710 1028610
rect 63726 1027610 63782 1028610
rect 64084 1027610 64144 1028610
rect 64344 1027610 64416 1028610
rect 64646 1027610 64702 1028610
rect 64718 1027610 64774 1028610
rect 65076 1027610 65136 1028610
rect 65336 1027610 65408 1028610
rect 65638 1027610 65694 1028610
rect 65710 1027610 65766 1028610
rect 66068 1027610 66128 1028610
rect 66328 1027610 66400 1028610
rect 66630 1027610 66686 1028610
rect 66702 1027610 66758 1028610
rect 67060 1027610 67120 1028610
rect 67320 1027610 67392 1028610
rect 67622 1027610 67678 1028610
rect 67694 1027610 67750 1028610
rect 68052 1027610 68112 1028610
rect 68312 1027610 68384 1028610
rect 68614 1027610 68670 1028610
rect 68686 1027610 68742 1028610
rect 69044 1027610 69104 1028610
rect 69304 1027610 69376 1028610
rect 69606 1027610 69662 1028610
rect 69678 1027610 69734 1028610
rect 70036 1027610 70096 1028610
rect 70296 1027610 70368 1028610
rect 70598 1027610 70654 1028610
rect 70670 1027610 70726 1028610
rect 71028 1027610 71088 1028610
rect 71288 1027610 71360 1028610
rect 71590 1027610 71646 1028610
rect 71662 1027610 71718 1028610
rect 72020 1027610 72080 1028610
rect 72280 1027610 72352 1028610
rect 72582 1027610 72638 1028610
rect 72654 1027610 72710 1028610
rect 73012 1027610 73072 1028610
rect 73272 1027610 73344 1028610
rect 73574 1027610 73630 1028610
rect 73646 1027610 73702 1028610
rect 74004 1027610 74064 1028610
rect 74264 1027610 74336 1028610
rect 74566 1027610 74622 1028610
rect 74638 1027610 74694 1028610
rect 74919 1027610 74959 1028610
rect 74996 1027610 75032 1028610
rect 75256 1027610 75328 1028610
rect 75481 1027610 75521 1028610
rect 75558 1027610 75614 1028610
rect 75630 1027610 75686 1028610
rect 75727 1027610 75763 1028610
rect 75777 1027610 75781 1028610
rect 75974 1027610 76034 1028610
rect 76070 1028588 76164 1028610
rect 76174 1028588 76198 1028610
rect 110256 1028604 110350 1028610
rect 76070 1028554 76174 1028588
rect 110246 1028556 110350 1028604
rect 76070 1028520 76164 1028554
rect 76174 1028520 76198 1028554
rect 110256 1028522 110350 1028556
rect 76070 1028480 76174 1028520
rect 110246 1028480 110350 1028522
rect 76070 1028446 76164 1028480
rect 76174 1028446 76208 1028480
rect 110256 1028446 110350 1028480
rect 76070 1028403 76174 1028446
rect 110246 1028403 110350 1028446
rect 76070 1028369 76164 1028403
rect 76174 1028369 76208 1028403
rect 110256 1028369 110350 1028403
rect 76070 1028309 76174 1028369
rect 110246 1028309 110350 1028369
rect 76070 1028275 76164 1028309
rect 76174 1028275 76208 1028309
rect 110256 1028275 110350 1028309
rect 76070 1028238 76174 1028275
rect 110246 1028238 110350 1028275
rect 76070 1028204 76164 1028238
rect 76174 1028204 76208 1028238
rect 110256 1028204 110350 1028238
rect 76070 1028164 76174 1028204
rect 110246 1028164 110350 1028204
rect 76070 1028130 76164 1028164
rect 76174 1028130 76208 1028164
rect 110256 1028130 110350 1028164
rect 76070 1028093 76174 1028130
rect 110246 1028093 110350 1028130
rect 76070 1028059 76164 1028093
rect 76174 1028059 76208 1028093
rect 110256 1028059 110350 1028093
rect 76070 1028019 76174 1028059
rect 110246 1028019 110350 1028059
rect 76070 1027985 76164 1028019
rect 76174 1027985 76208 1028019
rect 110256 1027985 110350 1028019
rect 76070 1027948 76174 1027985
rect 110246 1027948 110350 1027985
rect 76070 1027914 76164 1027948
rect 76174 1027914 76208 1027948
rect 110256 1027914 110350 1027948
rect 76070 1027874 76174 1027914
rect 110246 1027874 110350 1027914
rect 76070 1027840 76164 1027874
rect 76174 1027840 76208 1027874
rect 110256 1027840 110350 1027874
rect 76070 1027803 76174 1027840
rect 110246 1027803 110350 1027840
rect 76070 1027769 76164 1027803
rect 76174 1027769 76208 1027803
rect 110256 1027769 110350 1027803
rect 76070 1027729 76174 1027769
rect 110246 1027729 110350 1027769
rect 76070 1027695 76164 1027729
rect 76174 1027695 76208 1027729
rect 110256 1027695 110350 1027729
rect 76070 1027658 76174 1027695
rect 110246 1027658 110350 1027695
rect 76070 1027624 76164 1027658
rect 76174 1027624 76208 1027658
rect 110256 1027624 110350 1027658
rect 76070 1027610 76174 1027624
rect 110246 1027610 110350 1027624
rect 110692 1027610 110693 1028610
rect 110734 1027610 110790 1028610
rect 110831 1027610 110832 1028610
rect 122566 1027610 122622 1028610
rect 122638 1027610 122694 1028610
rect 123481 1027610 123521 1028610
rect 123558 1027610 123614 1028610
rect 123630 1027610 123686 1028610
rect 123727 1027610 123763 1028610
rect 123777 1027610 123781 1028610
rect 123974 1027610 124034 1028610
rect 124070 1028588 124164 1028610
rect 124174 1028588 124198 1028610
rect 124070 1028554 124174 1028588
rect 124070 1028520 124164 1028554
rect 124174 1028520 124198 1028554
rect 124070 1028480 124174 1028520
rect 124070 1028446 124164 1028480
rect 124174 1028446 124208 1028480
rect 124070 1028403 124174 1028446
rect 124070 1028369 124164 1028403
rect 124174 1028369 124208 1028403
rect 124070 1028309 124174 1028369
rect 124070 1028275 124164 1028309
rect 124174 1028275 124208 1028309
rect 124070 1028238 124174 1028275
rect 124070 1028204 124164 1028238
rect 124174 1028204 124208 1028238
rect 124070 1028164 124174 1028204
rect 124070 1028130 124164 1028164
rect 124174 1028130 124208 1028164
rect 124070 1028093 124174 1028130
rect 124070 1028059 124164 1028093
rect 124174 1028059 124208 1028093
rect 124070 1028019 124174 1028059
rect 124070 1027985 124164 1028019
rect 124174 1027985 124208 1028019
rect 124070 1027948 124174 1027985
rect 124070 1027914 124164 1027948
rect 124174 1027914 124208 1027948
rect 124070 1027874 124174 1027914
rect 124070 1027840 124164 1027874
rect 124174 1027840 124208 1027874
rect 124070 1027803 124174 1027840
rect 124070 1027769 124164 1027803
rect 124174 1027769 124208 1027803
rect 124070 1027729 124174 1027769
rect 124070 1027695 124164 1027729
rect 124174 1027695 124208 1027729
rect 124070 1027658 124174 1027695
rect 124070 1027624 124164 1027658
rect 124174 1027624 124208 1027658
rect 124070 1027610 124174 1027624
rect 162246 1027610 162350 1028610
rect 162446 1027610 162518 1028610
rect 162692 1027610 162697 1028610
rect 162734 1027610 162790 1028610
rect 162831 1027610 162832 1028610
rect 163092 1027610 163152 1028610
rect 163352 1027610 163424 1028610
rect 163654 1027610 163710 1028610
rect 163726 1027610 163782 1028610
rect 164084 1027610 164144 1028610
rect 164344 1027610 164416 1028610
rect 164646 1027610 164702 1028610
rect 164718 1027610 164774 1028610
rect 165076 1027610 165136 1028610
rect 165336 1027610 165408 1028610
rect 165638 1027610 165694 1028610
rect 165710 1027610 165766 1028610
rect 166068 1027610 166128 1028610
rect 166328 1027610 166400 1028610
rect 166630 1027610 166686 1028610
rect 166702 1027610 166758 1028610
rect 167060 1027610 167120 1028610
rect 167320 1027610 167392 1028610
rect 167622 1027610 167678 1028610
rect 167694 1027610 167750 1028610
rect 168052 1027610 168112 1028610
rect 168312 1027610 168384 1028610
rect 168614 1027610 168670 1028610
rect 168686 1027610 168742 1028610
rect 169044 1027610 169104 1028610
rect 169304 1027610 169376 1028610
rect 169606 1027610 169662 1028610
rect 169678 1027610 169734 1028610
rect 170036 1027610 170096 1028610
rect 170296 1027610 170368 1028610
rect 170598 1027610 170654 1028610
rect 170670 1027610 170726 1028610
rect 171028 1027610 171088 1028610
rect 171288 1027610 171360 1028610
rect 171590 1027610 171646 1028610
rect 171662 1027610 171718 1028610
rect 172020 1027610 172080 1028610
rect 172280 1027610 172352 1028610
rect 172582 1027610 172638 1028610
rect 172654 1027610 172710 1028610
rect 173012 1027610 173072 1028610
rect 173272 1027610 173344 1028610
rect 173574 1027610 173630 1028610
rect 173646 1027610 173702 1028610
rect 174004 1027610 174064 1028610
rect 174264 1027610 174336 1028610
rect 174566 1027610 174622 1028610
rect 174638 1027610 174694 1028610
rect 174919 1027610 174959 1028610
rect 174996 1027610 175032 1028610
rect 175256 1027610 175328 1028610
rect 175481 1027610 175521 1028610
rect 175558 1027610 175614 1028610
rect 175630 1027610 175686 1028610
rect 175727 1027610 175763 1028610
rect 175777 1027610 175781 1028610
rect 175974 1027610 176034 1028610
rect 176070 1028588 176164 1028610
rect 176174 1028588 176198 1028610
rect 214256 1028604 214350 1028610
rect 176070 1028554 176174 1028588
rect 214246 1028556 214350 1028604
rect 176070 1028520 176164 1028554
rect 176174 1028520 176198 1028554
rect 214256 1028522 214350 1028556
rect 176070 1028480 176174 1028520
rect 214246 1028480 214350 1028522
rect 176070 1028446 176164 1028480
rect 176174 1028446 176208 1028480
rect 214256 1028446 214350 1028480
rect 176070 1028403 176174 1028446
rect 214246 1028403 214350 1028446
rect 176070 1028369 176164 1028403
rect 176174 1028369 176208 1028403
rect 214256 1028369 214350 1028403
rect 176070 1028309 176174 1028369
rect 214246 1028309 214350 1028369
rect 176070 1028275 176164 1028309
rect 176174 1028275 176208 1028309
rect 214256 1028275 214350 1028309
rect 176070 1028238 176174 1028275
rect 214246 1028238 214350 1028275
rect 176070 1028204 176164 1028238
rect 176174 1028204 176208 1028238
rect 214256 1028204 214350 1028238
rect 176070 1028164 176174 1028204
rect 214246 1028164 214350 1028204
rect 176070 1028130 176164 1028164
rect 176174 1028130 176208 1028164
rect 214256 1028130 214350 1028164
rect 176070 1028093 176174 1028130
rect 214246 1028093 214350 1028130
rect 176070 1028059 176164 1028093
rect 176174 1028059 176208 1028093
rect 214256 1028059 214350 1028093
rect 176070 1028019 176174 1028059
rect 214246 1028019 214350 1028059
rect 176070 1027985 176164 1028019
rect 176174 1027985 176208 1028019
rect 214256 1027985 214350 1028019
rect 176070 1027948 176174 1027985
rect 214246 1027948 214350 1027985
rect 176070 1027914 176164 1027948
rect 176174 1027914 176208 1027948
rect 214256 1027914 214350 1027948
rect 176070 1027874 176174 1027914
rect 214246 1027874 214350 1027914
rect 176070 1027840 176164 1027874
rect 176174 1027840 176208 1027874
rect 214256 1027840 214350 1027874
rect 176070 1027803 176174 1027840
rect 214246 1027803 214350 1027840
rect 176070 1027769 176164 1027803
rect 176174 1027769 176208 1027803
rect 214256 1027769 214350 1027803
rect 176070 1027729 176174 1027769
rect 214246 1027729 214350 1027769
rect 176070 1027695 176164 1027729
rect 176174 1027695 176208 1027729
rect 214256 1027695 214350 1027729
rect 176070 1027658 176174 1027695
rect 214246 1027658 214350 1027695
rect 176070 1027624 176164 1027658
rect 176174 1027624 176208 1027658
rect 214256 1027624 214350 1027658
rect 176070 1027610 176174 1027624
rect 214246 1027610 214350 1027624
rect 214692 1027610 214693 1028610
rect 214734 1027610 214790 1028610
rect 214831 1027610 214832 1028610
rect 226566 1027610 226622 1028610
rect 226638 1027610 226694 1028610
rect 227481 1027610 227521 1028610
rect 227558 1027610 227614 1028610
rect 227630 1027610 227686 1028610
rect 227727 1027610 227763 1028610
rect 227777 1027610 227781 1028610
rect 227974 1027610 228034 1028610
rect 228070 1028588 228164 1028610
rect 228174 1028588 228198 1028610
rect 228070 1028554 228174 1028588
rect 228070 1028520 228164 1028554
rect 228174 1028520 228198 1028554
rect 228070 1028480 228174 1028520
rect 228070 1028446 228164 1028480
rect 228174 1028446 228208 1028480
rect 228070 1028403 228174 1028446
rect 228070 1028369 228164 1028403
rect 228174 1028369 228208 1028403
rect 228070 1028309 228174 1028369
rect 228070 1028275 228164 1028309
rect 228174 1028275 228208 1028309
rect 228070 1028238 228174 1028275
rect 228070 1028204 228164 1028238
rect 228174 1028204 228208 1028238
rect 228070 1028164 228174 1028204
rect 228070 1028130 228164 1028164
rect 228174 1028130 228208 1028164
rect 228070 1028093 228174 1028130
rect 228070 1028059 228164 1028093
rect 228174 1028059 228208 1028093
rect 228070 1028019 228174 1028059
rect 228070 1027985 228164 1028019
rect 228174 1027985 228208 1028019
rect 228070 1027948 228174 1027985
rect 228070 1027914 228164 1027948
rect 228174 1027914 228208 1027948
rect 228070 1027874 228174 1027914
rect 228070 1027840 228164 1027874
rect 228174 1027840 228208 1027874
rect 228070 1027803 228174 1027840
rect 228070 1027769 228164 1027803
rect 228174 1027769 228208 1027803
rect 228070 1027729 228174 1027769
rect 228070 1027695 228164 1027729
rect 228174 1027695 228208 1027729
rect 228070 1027658 228174 1027695
rect 228070 1027624 228164 1027658
rect 228174 1027624 228208 1027658
rect 228070 1027610 228174 1027624
rect 274566 1027610 274622 1028610
rect 274638 1027610 274694 1028610
rect 275481 1027610 275521 1028610
rect 275558 1027610 275614 1028610
rect 275630 1027610 275686 1028610
rect 275727 1027610 275763 1028610
rect 275777 1027610 275781 1028610
rect 275974 1027610 276034 1028610
rect 276070 1028588 276164 1028610
rect 276174 1028588 276198 1028610
rect 314256 1028604 314350 1028610
rect 276070 1028554 276174 1028588
rect 314246 1028556 314350 1028604
rect 276070 1028520 276164 1028554
rect 276174 1028520 276198 1028554
rect 314256 1028522 314350 1028556
rect 276070 1028480 276174 1028520
rect 314246 1028480 314350 1028522
rect 276070 1028446 276164 1028480
rect 276174 1028446 276208 1028480
rect 314256 1028446 314350 1028480
rect 276070 1028403 276174 1028446
rect 314246 1028403 314350 1028446
rect 276070 1028369 276164 1028403
rect 276174 1028369 276208 1028403
rect 314256 1028369 314350 1028403
rect 276070 1028309 276174 1028369
rect 314246 1028309 314350 1028369
rect 276070 1028275 276164 1028309
rect 276174 1028275 276208 1028309
rect 314256 1028275 314350 1028309
rect 276070 1028238 276174 1028275
rect 314246 1028238 314350 1028275
rect 276070 1028204 276164 1028238
rect 276174 1028204 276208 1028238
rect 314256 1028204 314350 1028238
rect 276070 1028164 276174 1028204
rect 314246 1028164 314350 1028204
rect 276070 1028130 276164 1028164
rect 276174 1028130 276208 1028164
rect 314256 1028130 314350 1028164
rect 276070 1028093 276174 1028130
rect 314246 1028093 314350 1028130
rect 276070 1028059 276164 1028093
rect 276174 1028059 276208 1028093
rect 314256 1028059 314350 1028093
rect 276070 1028019 276174 1028059
rect 314246 1028019 314350 1028059
rect 276070 1027985 276164 1028019
rect 276174 1027985 276208 1028019
rect 314256 1027985 314350 1028019
rect 276070 1027948 276174 1027985
rect 314246 1027948 314350 1027985
rect 276070 1027914 276164 1027948
rect 276174 1027914 276208 1027948
rect 314256 1027914 314350 1027948
rect 276070 1027874 276174 1027914
rect 314246 1027874 314350 1027914
rect 276070 1027840 276164 1027874
rect 276174 1027840 276208 1027874
rect 314256 1027840 314350 1027874
rect 276070 1027803 276174 1027840
rect 314246 1027803 314350 1027840
rect 276070 1027769 276164 1027803
rect 276174 1027769 276208 1027803
rect 314256 1027769 314350 1027803
rect 276070 1027729 276174 1027769
rect 314246 1027729 314350 1027769
rect 276070 1027695 276164 1027729
rect 276174 1027695 276208 1027729
rect 314256 1027695 314350 1027729
rect 276070 1027658 276174 1027695
rect 314246 1027658 314350 1027695
rect 276070 1027624 276164 1027658
rect 276174 1027624 276208 1027658
rect 314256 1027624 314350 1027658
rect 276070 1027610 276174 1027624
rect 314246 1027610 314350 1027624
rect 314692 1027610 314693 1028610
rect 314734 1027610 314790 1028610
rect 314831 1027610 314832 1028610
rect 326566 1027610 326622 1028610
rect 326638 1027610 326694 1028610
rect 327481 1027610 327521 1028610
rect 327558 1027610 327614 1028610
rect 327630 1027610 327686 1028610
rect 327727 1027610 327763 1028610
rect 327777 1027610 327781 1028610
rect 327974 1027610 328034 1028610
rect 328070 1028588 328164 1028610
rect 328174 1028588 328198 1028610
rect 328070 1028554 328174 1028588
rect 328070 1028520 328164 1028554
rect 328174 1028520 328198 1028554
rect 328070 1028480 328174 1028520
rect 328070 1028446 328164 1028480
rect 328174 1028446 328208 1028480
rect 328070 1028403 328174 1028446
rect 328070 1028369 328164 1028403
rect 328174 1028369 328208 1028403
rect 328070 1028309 328174 1028369
rect 328070 1028275 328164 1028309
rect 328174 1028275 328208 1028309
rect 328070 1028238 328174 1028275
rect 328070 1028204 328164 1028238
rect 328174 1028204 328208 1028238
rect 328070 1028164 328174 1028204
rect 328070 1028130 328164 1028164
rect 328174 1028130 328208 1028164
rect 328070 1028093 328174 1028130
rect 328070 1028059 328164 1028093
rect 328174 1028059 328208 1028093
rect 328070 1028019 328174 1028059
rect 328070 1027985 328164 1028019
rect 328174 1027985 328208 1028019
rect 328070 1027948 328174 1027985
rect 328070 1027914 328164 1027948
rect 328174 1027914 328208 1027948
rect 328070 1027874 328174 1027914
rect 328070 1027840 328164 1027874
rect 328174 1027840 328208 1027874
rect 328070 1027803 328174 1027840
rect 328070 1027769 328164 1027803
rect 328174 1027769 328208 1027803
rect 328070 1027729 328174 1027769
rect 328070 1027695 328164 1027729
rect 328174 1027695 328208 1027729
rect 328070 1027658 328174 1027695
rect 328070 1027624 328164 1027658
rect 328174 1027624 328208 1027658
rect 328070 1027610 328174 1027624
rect 366246 1027610 366350 1028610
rect 366446 1027610 366518 1028610
rect 366692 1027610 366697 1028610
rect 366734 1027610 366790 1028610
rect 366831 1027610 366832 1028610
rect 367092 1027610 367152 1028610
rect 367352 1027610 367424 1028610
rect 367654 1027610 367710 1028610
rect 367726 1027610 367782 1028610
rect 368084 1027610 368144 1028610
rect 368344 1027610 368416 1028610
rect 368646 1027610 368702 1028610
rect 368718 1027610 368774 1028610
rect 369076 1027610 369136 1028610
rect 369336 1027610 369408 1028610
rect 369638 1027610 369694 1028610
rect 369710 1027610 369766 1028610
rect 370068 1027610 370128 1028610
rect 370328 1027610 370400 1028610
rect 370630 1027610 370686 1028610
rect 370702 1027610 370758 1028610
rect 371060 1027610 371120 1028610
rect 371320 1027610 371392 1028610
rect 371622 1027610 371678 1028610
rect 371694 1027610 371750 1028610
rect 372052 1027610 372112 1028610
rect 372312 1027610 372384 1028610
rect 372614 1027610 372670 1028610
rect 372686 1027610 372742 1028610
rect 373044 1027610 373104 1028610
rect 373304 1027610 373376 1028610
rect 373606 1027610 373662 1028610
rect 373678 1027610 373734 1028610
rect 374036 1027610 374096 1028610
rect 374296 1027610 374368 1028610
rect 374598 1027610 374654 1028610
rect 374670 1027610 374726 1028610
rect 375028 1027610 375088 1028610
rect 375288 1027610 375360 1028610
rect 375590 1027610 375646 1028610
rect 375662 1027610 375718 1028610
rect 376020 1027610 376080 1028610
rect 376280 1027610 376352 1028610
rect 376582 1027610 376638 1028610
rect 376654 1027610 376710 1028610
rect 377012 1027610 377072 1028610
rect 377272 1027610 377344 1028610
rect 377574 1027610 377630 1028610
rect 377646 1027610 377702 1028610
rect 378004 1027610 378064 1028610
rect 378264 1027610 378336 1028610
rect 378566 1027610 378622 1028610
rect 378638 1027610 378694 1028610
rect 378919 1027610 378959 1028610
rect 378996 1027610 379032 1028610
rect 379256 1027610 379328 1028610
rect 379481 1027610 379521 1028610
rect 379558 1027610 379614 1028610
rect 379630 1027610 379686 1028610
rect 379727 1027610 379763 1028610
rect 379777 1027610 379781 1028610
rect 379974 1027610 380034 1028610
rect 380070 1028588 380164 1028610
rect 380174 1028588 380198 1028610
rect 414256 1028604 414350 1028610
rect 380070 1028554 380174 1028588
rect 414246 1028556 414350 1028604
rect 380070 1028520 380164 1028554
rect 380174 1028520 380198 1028554
rect 414256 1028522 414350 1028556
rect 380070 1028480 380174 1028520
rect 414246 1028480 414350 1028522
rect 380070 1028446 380164 1028480
rect 380174 1028446 380208 1028480
rect 414256 1028446 414350 1028480
rect 380070 1028403 380174 1028446
rect 414246 1028403 414350 1028446
rect 380070 1028369 380164 1028403
rect 380174 1028369 380208 1028403
rect 414256 1028369 414350 1028403
rect 380070 1028309 380174 1028369
rect 414246 1028309 414350 1028369
rect 380070 1028275 380164 1028309
rect 380174 1028275 380208 1028309
rect 414256 1028275 414350 1028309
rect 380070 1028238 380174 1028275
rect 414246 1028238 414350 1028275
rect 380070 1028204 380164 1028238
rect 380174 1028204 380208 1028238
rect 414256 1028204 414350 1028238
rect 380070 1028164 380174 1028204
rect 414246 1028164 414350 1028204
rect 380070 1028130 380164 1028164
rect 380174 1028130 380208 1028164
rect 414256 1028130 414350 1028164
rect 380070 1028093 380174 1028130
rect 414246 1028093 414350 1028130
rect 380070 1028059 380164 1028093
rect 380174 1028059 380208 1028093
rect 414256 1028059 414350 1028093
rect 380070 1028019 380174 1028059
rect 414246 1028019 414350 1028059
rect 380070 1027985 380164 1028019
rect 380174 1027985 380208 1028019
rect 414256 1027985 414350 1028019
rect 380070 1027948 380174 1027985
rect 414246 1027948 414350 1027985
rect 380070 1027914 380164 1027948
rect 380174 1027914 380208 1027948
rect 414256 1027914 414350 1027948
rect 380070 1027874 380174 1027914
rect 414246 1027874 414350 1027914
rect 380070 1027840 380164 1027874
rect 380174 1027840 380208 1027874
rect 414256 1027840 414350 1027874
rect 380070 1027803 380174 1027840
rect 414246 1027803 414350 1027840
rect 380070 1027769 380164 1027803
rect 380174 1027769 380208 1027803
rect 414256 1027769 414350 1027803
rect 380070 1027729 380174 1027769
rect 414246 1027729 414350 1027769
rect 380070 1027695 380164 1027729
rect 380174 1027695 380208 1027729
rect 414256 1027695 414350 1027729
rect 380070 1027658 380174 1027695
rect 414246 1027658 414350 1027695
rect 380070 1027624 380164 1027658
rect 380174 1027624 380208 1027658
rect 414256 1027624 414350 1027658
rect 380070 1027610 380174 1027624
rect 414246 1027610 414350 1027624
rect 414692 1027610 414693 1028610
rect 414734 1027610 414790 1028610
rect 414831 1027610 414832 1028610
rect 426566 1027610 426622 1028610
rect 426638 1027610 426694 1028610
rect 427481 1027610 427521 1028610
rect 427558 1027610 427614 1028610
rect 427630 1027610 427686 1028610
rect 427727 1027610 427763 1028610
rect 427777 1027610 427781 1028610
rect 427974 1027610 428034 1028610
rect 428070 1028588 428164 1028610
rect 428174 1028588 428198 1028610
rect 428070 1028554 428174 1028588
rect 428070 1028520 428164 1028554
rect 428174 1028520 428198 1028554
rect 428070 1028480 428174 1028520
rect 428070 1028446 428164 1028480
rect 428174 1028446 428208 1028480
rect 428070 1028403 428174 1028446
rect 428070 1028369 428164 1028403
rect 428174 1028369 428208 1028403
rect 428070 1028309 428174 1028369
rect 428070 1028275 428164 1028309
rect 428174 1028275 428208 1028309
rect 428070 1028238 428174 1028275
rect 428070 1028204 428164 1028238
rect 428174 1028204 428208 1028238
rect 428070 1028164 428174 1028204
rect 428070 1028130 428164 1028164
rect 428174 1028130 428208 1028164
rect 428070 1028093 428174 1028130
rect 428070 1028059 428164 1028093
rect 428174 1028059 428208 1028093
rect 428070 1028019 428174 1028059
rect 428070 1027985 428164 1028019
rect 428174 1027985 428208 1028019
rect 428070 1027948 428174 1027985
rect 428070 1027914 428164 1027948
rect 428174 1027914 428208 1027948
rect 428070 1027874 428174 1027914
rect 428070 1027840 428164 1027874
rect 428174 1027840 428208 1027874
rect 428070 1027803 428174 1027840
rect 428070 1027769 428164 1027803
rect 428174 1027769 428208 1027803
rect 428070 1027729 428174 1027769
rect 428070 1027695 428164 1027729
rect 428174 1027695 428208 1027729
rect 428070 1027658 428174 1027695
rect 428070 1027624 428164 1027658
rect 428174 1027624 428208 1027658
rect 428070 1027610 428174 1027624
rect 466246 1027610 466350 1028610
rect 466446 1027610 466518 1028610
rect 466692 1027610 466697 1028610
rect 466734 1027610 466790 1028610
rect 466831 1027610 466832 1028610
rect 467092 1027610 467152 1028610
rect 467352 1027610 467424 1028610
rect 467654 1027610 467710 1028610
rect 467726 1027610 467782 1028610
rect 468084 1027610 468144 1028610
rect 468344 1027610 468416 1028610
rect 468646 1027610 468702 1028610
rect 468718 1027610 468774 1028610
rect 469076 1027610 469136 1028610
rect 469336 1027610 469408 1028610
rect 469638 1027610 469694 1028610
rect 469710 1027610 469766 1028610
rect 470068 1027610 470128 1028610
rect 470328 1027610 470400 1028610
rect 470630 1027610 470686 1028610
rect 470702 1027610 470758 1028610
rect 471060 1027610 471120 1028610
rect 471320 1027610 471392 1028610
rect 471622 1027610 471678 1028610
rect 471694 1027610 471750 1028610
rect 472052 1027610 472112 1028610
rect 472312 1027610 472384 1028610
rect 472614 1027610 472670 1028610
rect 472686 1027610 472742 1028610
rect 473044 1027610 473104 1028610
rect 473304 1027610 473376 1028610
rect 473606 1027610 473662 1028610
rect 473678 1027610 473734 1028610
rect 474036 1027610 474096 1028610
rect 474296 1027610 474368 1028610
rect 474598 1027610 474654 1028610
rect 474670 1027610 474726 1028610
rect 475028 1027610 475088 1028610
rect 475288 1027610 475360 1028610
rect 475590 1027610 475646 1028610
rect 475662 1027610 475718 1028610
rect 476020 1027610 476080 1028610
rect 476280 1027610 476352 1028610
rect 476582 1027610 476638 1028610
rect 476654 1027610 476710 1028610
rect 477012 1027610 477072 1028610
rect 477272 1027610 477344 1028610
rect 477574 1027610 477630 1028610
rect 477646 1027610 477702 1028610
rect 478004 1027610 478064 1028610
rect 478264 1027610 478336 1028610
rect 478566 1027610 478622 1028610
rect 478638 1027610 478694 1028610
rect 478919 1027610 478959 1028610
rect 478996 1027610 479032 1028610
rect 479256 1027610 479328 1028610
rect 479481 1027610 479521 1028610
rect 479558 1027610 479614 1028610
rect 479630 1027610 479686 1028610
rect 479727 1027610 479763 1028610
rect 479777 1027610 479781 1028610
rect 479974 1027610 480034 1028610
rect 480070 1028588 480164 1028610
rect 480174 1028588 480198 1028610
rect 518256 1028604 518350 1028610
rect 480070 1028554 480174 1028588
rect 518246 1028556 518350 1028604
rect 480070 1028520 480164 1028554
rect 480174 1028520 480198 1028554
rect 518256 1028522 518350 1028556
rect 480070 1028480 480174 1028520
rect 518246 1028480 518350 1028522
rect 480070 1028446 480164 1028480
rect 480174 1028446 480208 1028480
rect 518256 1028446 518350 1028480
rect 480070 1028403 480174 1028446
rect 518246 1028403 518350 1028446
rect 480070 1028369 480164 1028403
rect 480174 1028369 480208 1028403
rect 518256 1028369 518350 1028403
rect 480070 1028309 480174 1028369
rect 518246 1028309 518350 1028369
rect 480070 1028275 480164 1028309
rect 480174 1028275 480208 1028309
rect 518256 1028275 518350 1028309
rect 480070 1028238 480174 1028275
rect 518246 1028238 518350 1028275
rect 480070 1028204 480164 1028238
rect 480174 1028204 480208 1028238
rect 518256 1028204 518350 1028238
rect 480070 1028164 480174 1028204
rect 518246 1028164 518350 1028204
rect 480070 1028130 480164 1028164
rect 480174 1028130 480208 1028164
rect 518256 1028130 518350 1028164
rect 480070 1028093 480174 1028130
rect 518246 1028093 518350 1028130
rect 480070 1028059 480164 1028093
rect 480174 1028059 480208 1028093
rect 518256 1028059 518350 1028093
rect 480070 1028019 480174 1028059
rect 518246 1028019 518350 1028059
rect 480070 1027985 480164 1028019
rect 480174 1027985 480208 1028019
rect 518256 1027985 518350 1028019
rect 480070 1027948 480174 1027985
rect 518246 1027948 518350 1027985
rect 480070 1027914 480164 1027948
rect 480174 1027914 480208 1027948
rect 518256 1027914 518350 1027948
rect 480070 1027874 480174 1027914
rect 518246 1027874 518350 1027914
rect 480070 1027840 480164 1027874
rect 480174 1027840 480208 1027874
rect 518256 1027840 518350 1027874
rect 480070 1027803 480174 1027840
rect 518246 1027803 518350 1027840
rect 480070 1027769 480164 1027803
rect 480174 1027769 480208 1027803
rect 518256 1027769 518350 1027803
rect 480070 1027729 480174 1027769
rect 518246 1027729 518350 1027769
rect 480070 1027695 480164 1027729
rect 480174 1027695 480208 1027729
rect 518256 1027695 518350 1027729
rect 480070 1027658 480174 1027695
rect 518246 1027658 518350 1027695
rect 480070 1027624 480164 1027658
rect 480174 1027624 480208 1027658
rect 518256 1027624 518350 1027658
rect 480070 1027610 480174 1027624
rect 518246 1027610 518350 1027624
rect 518692 1027610 518693 1028610
rect 518734 1027610 518790 1028610
rect 518831 1027610 518832 1028610
rect 530566 1027610 530622 1028610
rect 530638 1027610 530694 1028610
rect 531481 1027610 531521 1028610
rect 531558 1027610 531614 1028610
rect 531630 1027610 531686 1028610
rect 531727 1027610 531763 1028610
rect 531777 1027610 531781 1028610
rect 531974 1027610 532034 1028610
rect 532070 1028588 532164 1028610
rect 532174 1028588 532198 1028610
rect 532070 1028554 532174 1028588
rect 532070 1028520 532164 1028554
rect 532174 1028520 532198 1028554
rect 532070 1028480 532174 1028520
rect 532070 1028446 532164 1028480
rect 532174 1028446 532208 1028480
rect 532070 1028403 532174 1028446
rect 532070 1028369 532164 1028403
rect 532174 1028369 532208 1028403
rect 532070 1028309 532174 1028369
rect 532070 1028275 532164 1028309
rect 532174 1028275 532208 1028309
rect 532070 1028238 532174 1028275
rect 532070 1028204 532164 1028238
rect 532174 1028204 532208 1028238
rect 532070 1028164 532174 1028204
rect 532070 1028130 532164 1028164
rect 532174 1028130 532208 1028164
rect 532070 1028093 532174 1028130
rect 532070 1028059 532164 1028093
rect 532174 1028059 532208 1028093
rect 532070 1028019 532174 1028059
rect 532070 1027985 532164 1028019
rect 532174 1027985 532208 1028019
rect 532070 1027948 532174 1027985
rect 532070 1027914 532164 1027948
rect 532174 1027914 532208 1027948
rect 532070 1027874 532174 1027914
rect 532070 1027840 532164 1027874
rect 532174 1027840 532208 1027874
rect 532070 1027803 532174 1027840
rect 532070 1027769 532164 1027803
rect 532174 1027769 532208 1027803
rect 532070 1027729 532174 1027769
rect 532070 1027695 532164 1027729
rect 532174 1027695 532208 1027729
rect 532070 1027658 532174 1027695
rect 532070 1027624 532164 1027658
rect 532174 1027624 532208 1027658
rect 532070 1027610 532174 1027624
rect 570246 1027610 570350 1028610
rect 570446 1027610 570518 1028610
rect 570692 1027610 570697 1028610
rect 570734 1027610 570790 1028610
rect 570831 1027610 570832 1028610
rect 571092 1027610 571152 1028610
rect 571352 1027610 571424 1028610
rect 571654 1027610 571710 1028610
rect 571726 1027610 571782 1028610
rect 572084 1027610 572144 1028610
rect 572344 1027610 572416 1028610
rect 572646 1027610 572702 1028610
rect 572718 1027610 572774 1028610
rect 573076 1027610 573136 1028610
rect 573336 1027610 573408 1028610
rect 573638 1027610 573694 1028610
rect 573710 1027610 573766 1028610
rect 574068 1027610 574128 1028610
rect 574328 1027610 574400 1028610
rect 574630 1027610 574686 1028610
rect 574702 1027610 574758 1028610
rect 575060 1027610 575120 1028610
rect 575320 1027610 575392 1028610
rect 575622 1027610 575678 1028610
rect 575694 1027610 575750 1028610
rect 576052 1027610 576112 1028610
rect 576312 1027610 576384 1028610
rect 576614 1027610 576670 1028610
rect 576686 1027610 576742 1028610
rect 577044 1027610 577104 1028610
rect 577304 1027610 577376 1028610
rect 577606 1027610 577662 1028610
rect 577678 1027610 577734 1028610
rect 578036 1027610 578096 1028610
rect 578296 1027610 578368 1028610
rect 578598 1027610 578654 1028610
rect 578670 1027610 578726 1028610
rect 579028 1027610 579088 1028610
rect 579288 1027610 579360 1028610
rect 579590 1027610 579646 1028610
rect 579662 1027610 579718 1028610
rect 580020 1027610 580080 1028610
rect 580280 1027610 580352 1028610
rect 580582 1027610 580638 1028610
rect 580654 1027610 580710 1028610
rect 581012 1027610 581072 1028610
rect 581272 1027610 581344 1028610
rect 581574 1027610 581630 1028610
rect 581646 1027610 581702 1028610
rect 582004 1027610 582064 1028610
rect 582264 1027610 582336 1028610
rect 582566 1027610 582622 1028610
rect 582638 1027610 582694 1028610
rect 582919 1027610 582959 1028610
rect 582996 1027610 583032 1028610
rect 583256 1027610 583328 1028610
rect 583481 1027610 583521 1028610
rect 583558 1027610 583614 1028610
rect 583630 1027610 583686 1028610
rect 583727 1027610 583763 1028610
rect 583777 1027610 583781 1028610
rect 583974 1027610 584034 1028610
rect 584070 1028588 584164 1028610
rect 584174 1028588 584198 1028610
rect 584070 1028554 584174 1028588
rect 584070 1028520 584164 1028554
rect 584174 1028520 584198 1028554
rect 584070 1028480 584174 1028520
rect 584070 1028446 584164 1028480
rect 584174 1028446 584208 1028480
rect 584070 1028403 584174 1028446
rect 584070 1028369 584164 1028403
rect 584174 1028369 584208 1028403
rect 584070 1028309 584174 1028369
rect 584070 1028275 584164 1028309
rect 584174 1028275 584208 1028309
rect 584070 1028238 584174 1028275
rect 584070 1028204 584164 1028238
rect 584174 1028204 584208 1028238
rect 584070 1028164 584174 1028204
rect 584070 1028130 584164 1028164
rect 584174 1028130 584208 1028164
rect 584070 1028093 584174 1028130
rect 584070 1028059 584164 1028093
rect 584174 1028059 584208 1028093
rect 584070 1028019 584174 1028059
rect 584070 1027985 584164 1028019
rect 584174 1027985 584208 1028019
rect 584070 1027948 584174 1027985
rect 584070 1027914 584164 1027948
rect 584174 1027914 584208 1027948
rect 584070 1027874 584174 1027914
rect 584070 1027840 584164 1027874
rect 584174 1027840 584208 1027874
rect 584070 1027803 584174 1027840
rect 584070 1027769 584164 1027803
rect 584174 1027769 584208 1027803
rect 584070 1027729 584174 1027769
rect 584070 1027695 584164 1027729
rect 584174 1027695 584208 1027729
rect 584070 1027658 584174 1027695
rect 584070 1027624 584164 1027658
rect 584174 1027624 584208 1027658
rect 584070 1027610 584174 1027624
rect 62657 1027574 62867 1027610
rect 74919 1027574 75032 1027610
rect 75481 1027574 75763 1027610
rect 123481 1027574 123763 1027610
rect 162657 1027574 162867 1027610
rect 174919 1027574 175032 1027610
rect 175481 1027574 175763 1027610
rect 227481 1027574 227763 1027610
rect 275481 1027574 275763 1027610
rect 327481 1027574 327763 1027610
rect 366657 1027574 366867 1027610
rect 378919 1027574 379032 1027610
rect 379481 1027574 379763 1027610
rect 427481 1027574 427763 1027610
rect 466657 1027574 466867 1027610
rect 478919 1027574 479032 1027610
rect 479481 1027574 479763 1027610
rect 531481 1027574 531763 1027610
rect 570657 1027574 570867 1027610
rect 582919 1027574 583032 1027610
rect 583481 1027574 583763 1027610
rect 62069 1025107 62085 1025173
rect 64093 1025107 64109 1025173
rect 110069 1025107 110085 1025173
rect 162069 1025107 162085 1025173
rect 164093 1025107 164109 1025173
rect 214069 1025107 214085 1025173
rect 262069 1025107 262080 1025173
rect 314069 1025107 314085 1025173
rect 366069 1025107 366085 1025173
rect 368093 1025107 368109 1025173
rect 414069 1025107 414085 1025173
rect 466069 1025107 466085 1025173
rect 468093 1025107 468109 1025173
rect 518069 1025107 518085 1025173
rect 570069 1025107 570085 1025173
rect 572093 1025107 572109 1025173
rect 70260 1025041 70276 1025057
rect 70158 1024735 70276 1025041
rect 70260 1024719 70276 1024735
rect 72448 1025041 72464 1025057
rect 170260 1025041 170276 1025057
rect 72448 1024735 72566 1025041
rect 170158 1024735 170276 1025041
rect 72448 1024719 72464 1024735
rect 170260 1024719 170276 1024735
rect 172448 1025041 172464 1025057
rect 374260 1025041 374276 1025057
rect 172448 1024735 172566 1025041
rect 374158 1024735 374276 1025041
rect 172448 1024719 172464 1024735
rect 374260 1024719 374276 1024735
rect 376448 1025041 376464 1025057
rect 474260 1025041 474276 1025057
rect 376448 1024735 376566 1025041
rect 474158 1024735 474276 1025041
rect 376448 1024719 376464 1024735
rect 474260 1024719 474276 1024735
rect 476448 1025041 476464 1025057
rect 578260 1025041 578276 1025057
rect 476448 1024735 476566 1025041
rect 578158 1024735 578276 1025041
rect 476448 1024719 476464 1024735
rect 578260 1024719 578276 1024735
rect 580448 1025041 580464 1025057
rect 580448 1024735 580566 1025041
rect 580448 1024719 580464 1024735
rect 61692 1022853 61716 1023645
rect 71531 1023541 71535 1023701
rect 71677 1023541 71681 1023701
rect 72873 1023541 72877 1023701
rect 73019 1023539 73023 1023699
rect 109692 1022853 109716 1023645
rect 161692 1022853 161716 1023645
rect 171531 1023541 171535 1023701
rect 171677 1023541 171681 1023701
rect 172873 1023541 172877 1023701
rect 173019 1023539 173023 1023699
rect 213692 1022853 213716 1023645
rect 261692 1022853 261716 1023645
rect 313692 1022853 313716 1023645
rect 365692 1022853 365716 1023645
rect 375531 1023541 375535 1023701
rect 375677 1023541 375681 1023701
rect 376873 1023541 376877 1023701
rect 377019 1023539 377023 1023699
rect 413692 1022853 413716 1023645
rect 465692 1022853 465716 1023645
rect 475531 1023541 475535 1023701
rect 475677 1023541 475681 1023701
rect 476873 1023541 476877 1023701
rect 477019 1023539 477023 1023699
rect 517692 1022853 517716 1023645
rect 569692 1022853 569716 1023645
rect 579531 1023541 579535 1023701
rect 579677 1023541 579681 1023701
rect 580873 1023541 580877 1023701
rect 581019 1023539 581023 1023699
rect 61561 1022756 61716 1022853
rect 109561 1022756 109716 1022853
rect 161561 1022756 161716 1022853
rect 213561 1022756 213716 1022853
rect 261561 1022756 261716 1022853
rect 313561 1022756 313716 1022853
rect 365561 1022756 365716 1022853
rect 413561 1022756 413716 1022853
rect 465561 1022756 465716 1022853
rect 517561 1022756 517716 1022853
rect 569561 1022756 569716 1022853
rect 61561 1018210 61668 1022756
rect 62356 1020922 62406 1021922
rect 62617 1020922 62673 1021922
rect 62689 1020922 62745 1021922
rect 63047 1021842 63247 1021922
rect 63262 1021852 63296 1021876
rect 63307 1021852 63379 1021922
rect 63262 1021842 63379 1021852
rect 63034 1021818 63379 1021842
rect 63047 1021774 63247 1021818
rect 63262 1021808 63286 1021818
rect 63262 1021784 63296 1021808
rect 63307 1021784 63379 1021818
rect 63262 1021774 63379 1021784
rect 63034 1021750 63379 1021774
rect 63047 1021706 63247 1021750
rect 63262 1021740 63286 1021750
rect 63262 1021716 63296 1021740
rect 63307 1021716 63379 1021750
rect 63262 1021706 63379 1021716
rect 63034 1021682 63379 1021706
rect 63047 1021638 63247 1021682
rect 63262 1021672 63286 1021682
rect 63262 1021648 63296 1021672
rect 63307 1021648 63379 1021682
rect 63262 1021638 63379 1021648
rect 63034 1021614 63379 1021638
rect 63047 1021570 63247 1021614
rect 63262 1021604 63286 1021614
rect 63262 1021580 63296 1021604
rect 63307 1021580 63379 1021614
rect 63262 1021570 63379 1021580
rect 63034 1021546 63379 1021570
rect 63047 1021502 63247 1021546
rect 63262 1021536 63286 1021546
rect 63262 1021512 63296 1021536
rect 63307 1021512 63379 1021546
rect 63262 1021502 63379 1021512
rect 63034 1021478 63379 1021502
rect 63047 1021434 63247 1021478
rect 63262 1021468 63286 1021478
rect 63262 1021444 63296 1021468
rect 63307 1021444 63379 1021478
rect 63262 1021434 63379 1021444
rect 63034 1021410 63379 1021434
rect 63047 1021366 63247 1021410
rect 63262 1021400 63286 1021410
rect 63262 1021376 63296 1021400
rect 63307 1021376 63379 1021410
rect 63262 1021366 63379 1021376
rect 63034 1021342 63379 1021366
rect 63047 1021298 63247 1021342
rect 63262 1021332 63286 1021342
rect 63262 1021308 63296 1021332
rect 63307 1021308 63379 1021342
rect 63262 1021298 63379 1021308
rect 63034 1021274 63379 1021298
rect 63047 1021230 63247 1021274
rect 63262 1021264 63286 1021274
rect 63262 1021240 63296 1021264
rect 63307 1021240 63379 1021274
rect 63262 1021230 63379 1021240
rect 63034 1021206 63379 1021230
rect 63047 1021162 63247 1021206
rect 63262 1021196 63286 1021206
rect 63262 1021172 63296 1021196
rect 63307 1021172 63379 1021206
rect 63262 1021162 63379 1021172
rect 63034 1021138 63379 1021162
rect 63047 1021094 63247 1021138
rect 63262 1021128 63286 1021138
rect 63262 1021104 63296 1021128
rect 63307 1021104 63379 1021138
rect 63262 1021094 63379 1021104
rect 63034 1021070 63379 1021094
rect 63047 1021026 63247 1021070
rect 63262 1021060 63286 1021070
rect 63262 1021036 63296 1021060
rect 63307 1021036 63379 1021070
rect 63262 1021026 63379 1021036
rect 63034 1021002 63379 1021026
rect 63047 1020958 63247 1021002
rect 63262 1020992 63286 1021002
rect 63262 1020968 63296 1020992
rect 63307 1020968 63379 1021002
rect 63262 1020958 63379 1020968
rect 63034 1020934 63379 1020958
rect 63047 1020922 63247 1020934
rect 63058 1020910 63082 1020922
rect 63262 1020910 63286 1020934
rect 63307 1020922 63379 1020934
rect 63609 1020922 63665 1021922
rect 63681 1020922 63737 1021922
rect 64039 1021842 64239 1021922
rect 64254 1021852 64288 1021876
rect 64299 1021852 64371 1021922
rect 64254 1021842 64371 1021852
rect 64026 1021818 64371 1021842
rect 64039 1021774 64239 1021818
rect 64254 1021808 64278 1021818
rect 64254 1021784 64288 1021808
rect 64299 1021784 64371 1021818
rect 64254 1021774 64371 1021784
rect 64026 1021750 64371 1021774
rect 64039 1021706 64239 1021750
rect 64254 1021740 64278 1021750
rect 64254 1021716 64288 1021740
rect 64299 1021716 64371 1021750
rect 64254 1021706 64371 1021716
rect 64026 1021682 64371 1021706
rect 64039 1021638 64239 1021682
rect 64254 1021672 64278 1021682
rect 64254 1021648 64288 1021672
rect 64299 1021648 64371 1021682
rect 64254 1021638 64371 1021648
rect 64026 1021614 64371 1021638
rect 64039 1021570 64239 1021614
rect 64254 1021604 64278 1021614
rect 64254 1021580 64288 1021604
rect 64299 1021580 64371 1021614
rect 64254 1021570 64371 1021580
rect 64026 1021546 64371 1021570
rect 64039 1021502 64239 1021546
rect 64254 1021536 64278 1021546
rect 64254 1021512 64288 1021536
rect 64299 1021512 64371 1021546
rect 64254 1021502 64371 1021512
rect 64026 1021478 64371 1021502
rect 64039 1021434 64239 1021478
rect 64254 1021468 64278 1021478
rect 64254 1021444 64288 1021468
rect 64299 1021444 64371 1021478
rect 64254 1021434 64371 1021444
rect 64026 1021410 64371 1021434
rect 64039 1021366 64239 1021410
rect 64254 1021400 64278 1021410
rect 64254 1021376 64288 1021400
rect 64299 1021376 64371 1021410
rect 64254 1021366 64371 1021376
rect 64026 1021342 64371 1021366
rect 64039 1021298 64239 1021342
rect 64254 1021332 64278 1021342
rect 64254 1021308 64288 1021332
rect 64299 1021308 64371 1021342
rect 64254 1021298 64371 1021308
rect 64026 1021274 64371 1021298
rect 64039 1021230 64239 1021274
rect 64254 1021264 64278 1021274
rect 64254 1021240 64288 1021264
rect 64299 1021240 64371 1021274
rect 64254 1021230 64371 1021240
rect 64026 1021206 64371 1021230
rect 64039 1021162 64239 1021206
rect 64254 1021196 64278 1021206
rect 64254 1021172 64288 1021196
rect 64299 1021172 64371 1021206
rect 64254 1021162 64371 1021172
rect 64026 1021138 64371 1021162
rect 64039 1021094 64239 1021138
rect 64254 1021128 64278 1021138
rect 64254 1021104 64288 1021128
rect 64299 1021104 64371 1021138
rect 64254 1021094 64371 1021104
rect 64026 1021070 64371 1021094
rect 64039 1021026 64239 1021070
rect 64254 1021060 64278 1021070
rect 64254 1021036 64288 1021060
rect 64299 1021036 64371 1021070
rect 64254 1021026 64371 1021036
rect 64026 1021002 64371 1021026
rect 64039 1020958 64239 1021002
rect 64254 1020992 64278 1021002
rect 64254 1020968 64288 1020992
rect 64299 1020968 64371 1021002
rect 64254 1020958 64371 1020968
rect 64026 1020934 64371 1020958
rect 64039 1020922 64239 1020934
rect 64050 1020910 64074 1020922
rect 64254 1020910 64278 1020934
rect 64299 1020922 64371 1020934
rect 64601 1020922 64657 1021922
rect 64673 1020922 64729 1021922
rect 65031 1021842 65231 1021922
rect 65246 1021852 65280 1021876
rect 65291 1021852 65363 1021922
rect 65246 1021842 65363 1021852
rect 65018 1021818 65363 1021842
rect 65031 1021774 65231 1021818
rect 65246 1021808 65270 1021818
rect 65246 1021784 65280 1021808
rect 65291 1021784 65363 1021818
rect 65246 1021774 65363 1021784
rect 65018 1021750 65363 1021774
rect 65031 1021706 65231 1021750
rect 65246 1021740 65270 1021750
rect 65246 1021716 65280 1021740
rect 65291 1021716 65363 1021750
rect 65246 1021706 65363 1021716
rect 65018 1021682 65363 1021706
rect 65031 1021638 65231 1021682
rect 65246 1021672 65270 1021682
rect 65246 1021648 65280 1021672
rect 65291 1021648 65363 1021682
rect 65246 1021638 65363 1021648
rect 65018 1021614 65363 1021638
rect 65031 1021570 65231 1021614
rect 65246 1021604 65270 1021614
rect 65246 1021580 65280 1021604
rect 65291 1021580 65363 1021614
rect 65246 1021570 65363 1021580
rect 65018 1021546 65363 1021570
rect 65031 1021502 65231 1021546
rect 65246 1021536 65270 1021546
rect 65246 1021512 65280 1021536
rect 65291 1021512 65363 1021546
rect 65246 1021502 65363 1021512
rect 65018 1021478 65363 1021502
rect 65031 1021434 65231 1021478
rect 65246 1021468 65270 1021478
rect 65246 1021444 65280 1021468
rect 65291 1021444 65363 1021478
rect 65246 1021434 65363 1021444
rect 65018 1021410 65363 1021434
rect 65031 1021366 65231 1021410
rect 65246 1021400 65270 1021410
rect 65246 1021376 65280 1021400
rect 65291 1021376 65363 1021410
rect 65246 1021366 65363 1021376
rect 65018 1021342 65363 1021366
rect 65031 1021298 65231 1021342
rect 65246 1021332 65270 1021342
rect 65246 1021308 65280 1021332
rect 65291 1021308 65363 1021342
rect 65246 1021298 65363 1021308
rect 65018 1021274 65363 1021298
rect 65031 1021230 65231 1021274
rect 65246 1021264 65270 1021274
rect 65246 1021240 65280 1021264
rect 65291 1021240 65363 1021274
rect 65246 1021230 65363 1021240
rect 65018 1021206 65363 1021230
rect 65031 1021162 65231 1021206
rect 65246 1021196 65270 1021206
rect 65246 1021172 65280 1021196
rect 65291 1021172 65363 1021206
rect 65246 1021162 65363 1021172
rect 65018 1021138 65363 1021162
rect 65031 1021094 65231 1021138
rect 65246 1021128 65270 1021138
rect 65246 1021104 65280 1021128
rect 65291 1021104 65363 1021138
rect 65246 1021094 65363 1021104
rect 65018 1021070 65363 1021094
rect 65031 1021026 65231 1021070
rect 65246 1021060 65270 1021070
rect 65246 1021036 65280 1021060
rect 65291 1021036 65363 1021070
rect 65246 1021026 65363 1021036
rect 65018 1021002 65363 1021026
rect 65031 1020958 65231 1021002
rect 65246 1020992 65270 1021002
rect 65246 1020968 65280 1020992
rect 65291 1020968 65363 1021002
rect 65246 1020958 65363 1020968
rect 65018 1020934 65363 1020958
rect 65031 1020922 65231 1020934
rect 65042 1020910 65066 1020922
rect 65246 1020910 65270 1020934
rect 65291 1020922 65363 1020934
rect 65593 1020922 65649 1021922
rect 65665 1020922 65721 1021922
rect 66023 1021842 66223 1021922
rect 66238 1021852 66272 1021876
rect 66283 1021852 66355 1021922
rect 66238 1021842 66355 1021852
rect 66010 1021818 66355 1021842
rect 66023 1021774 66223 1021818
rect 66238 1021808 66262 1021818
rect 66238 1021784 66272 1021808
rect 66283 1021784 66355 1021818
rect 66238 1021774 66355 1021784
rect 66010 1021750 66355 1021774
rect 66023 1021706 66223 1021750
rect 66238 1021740 66262 1021750
rect 66238 1021716 66272 1021740
rect 66283 1021716 66355 1021750
rect 66238 1021706 66355 1021716
rect 66010 1021682 66355 1021706
rect 66023 1021638 66223 1021682
rect 66238 1021672 66262 1021682
rect 66238 1021648 66272 1021672
rect 66283 1021648 66355 1021682
rect 66238 1021638 66355 1021648
rect 66010 1021614 66355 1021638
rect 66023 1021570 66223 1021614
rect 66238 1021604 66262 1021614
rect 66238 1021580 66272 1021604
rect 66283 1021580 66355 1021614
rect 66238 1021570 66355 1021580
rect 66010 1021546 66355 1021570
rect 66023 1021502 66223 1021546
rect 66238 1021536 66262 1021546
rect 66238 1021512 66272 1021536
rect 66283 1021512 66355 1021546
rect 66238 1021502 66355 1021512
rect 66010 1021478 66355 1021502
rect 66023 1021434 66223 1021478
rect 66238 1021468 66262 1021478
rect 66238 1021444 66272 1021468
rect 66283 1021444 66355 1021478
rect 66238 1021434 66355 1021444
rect 66010 1021410 66355 1021434
rect 66023 1021366 66223 1021410
rect 66238 1021400 66262 1021410
rect 66238 1021376 66272 1021400
rect 66283 1021376 66355 1021410
rect 66238 1021366 66355 1021376
rect 66010 1021342 66355 1021366
rect 66023 1021298 66223 1021342
rect 66238 1021332 66262 1021342
rect 66238 1021308 66272 1021332
rect 66283 1021308 66355 1021342
rect 66238 1021298 66355 1021308
rect 66010 1021274 66355 1021298
rect 66023 1021230 66223 1021274
rect 66238 1021264 66262 1021274
rect 66238 1021240 66272 1021264
rect 66283 1021240 66355 1021274
rect 66238 1021230 66355 1021240
rect 66010 1021206 66355 1021230
rect 66023 1021162 66223 1021206
rect 66238 1021196 66262 1021206
rect 66238 1021172 66272 1021196
rect 66283 1021172 66355 1021206
rect 66238 1021162 66355 1021172
rect 66010 1021138 66355 1021162
rect 66023 1021094 66223 1021138
rect 66238 1021128 66262 1021138
rect 66238 1021104 66272 1021128
rect 66283 1021104 66355 1021138
rect 66238 1021094 66355 1021104
rect 66010 1021070 66355 1021094
rect 66023 1021026 66223 1021070
rect 66238 1021060 66262 1021070
rect 66238 1021036 66272 1021060
rect 66283 1021036 66355 1021070
rect 66238 1021026 66355 1021036
rect 66010 1021002 66355 1021026
rect 66023 1020958 66223 1021002
rect 66238 1020992 66262 1021002
rect 66238 1020968 66272 1020992
rect 66283 1020968 66355 1021002
rect 66238 1020958 66355 1020968
rect 66010 1020934 66355 1020958
rect 66023 1020922 66223 1020934
rect 66034 1020910 66058 1020922
rect 66238 1020910 66262 1020934
rect 66283 1020922 66355 1020934
rect 66585 1020922 66641 1021922
rect 66657 1020922 66713 1021922
rect 67015 1021842 67215 1021922
rect 67230 1021852 67264 1021876
rect 67275 1021852 67347 1021922
rect 67230 1021842 67347 1021852
rect 67002 1021818 67347 1021842
rect 67015 1021774 67215 1021818
rect 67230 1021808 67254 1021818
rect 67230 1021784 67264 1021808
rect 67275 1021784 67347 1021818
rect 67230 1021774 67347 1021784
rect 67002 1021750 67347 1021774
rect 67015 1021706 67215 1021750
rect 67230 1021740 67254 1021750
rect 67230 1021716 67264 1021740
rect 67275 1021716 67347 1021750
rect 67230 1021706 67347 1021716
rect 67002 1021682 67347 1021706
rect 67015 1021638 67215 1021682
rect 67230 1021672 67254 1021682
rect 67230 1021648 67264 1021672
rect 67275 1021648 67347 1021682
rect 67230 1021638 67347 1021648
rect 67002 1021614 67347 1021638
rect 67015 1021570 67215 1021614
rect 67230 1021604 67254 1021614
rect 67230 1021580 67264 1021604
rect 67275 1021580 67347 1021614
rect 67230 1021570 67347 1021580
rect 67002 1021546 67347 1021570
rect 67015 1021502 67215 1021546
rect 67230 1021536 67254 1021546
rect 67230 1021512 67264 1021536
rect 67275 1021512 67347 1021546
rect 67230 1021502 67347 1021512
rect 67002 1021478 67347 1021502
rect 67015 1021434 67215 1021478
rect 67230 1021468 67254 1021478
rect 67230 1021444 67264 1021468
rect 67275 1021444 67347 1021478
rect 67230 1021434 67347 1021444
rect 67002 1021410 67347 1021434
rect 67015 1021366 67215 1021410
rect 67230 1021400 67254 1021410
rect 67230 1021376 67264 1021400
rect 67275 1021376 67347 1021410
rect 67230 1021366 67347 1021376
rect 67002 1021342 67347 1021366
rect 67015 1021298 67215 1021342
rect 67230 1021332 67254 1021342
rect 67230 1021308 67264 1021332
rect 67275 1021308 67347 1021342
rect 67230 1021298 67347 1021308
rect 67002 1021274 67347 1021298
rect 67015 1021230 67215 1021274
rect 67230 1021264 67254 1021274
rect 67230 1021240 67264 1021264
rect 67275 1021240 67347 1021274
rect 67230 1021230 67347 1021240
rect 67002 1021206 67347 1021230
rect 67015 1021162 67215 1021206
rect 67230 1021196 67254 1021206
rect 67230 1021172 67264 1021196
rect 67275 1021172 67347 1021206
rect 67230 1021162 67347 1021172
rect 67002 1021138 67347 1021162
rect 67015 1021094 67215 1021138
rect 67230 1021128 67254 1021138
rect 67230 1021104 67264 1021128
rect 67275 1021104 67347 1021138
rect 67230 1021094 67347 1021104
rect 67002 1021070 67347 1021094
rect 67015 1021026 67215 1021070
rect 67230 1021060 67254 1021070
rect 67230 1021036 67264 1021060
rect 67275 1021036 67347 1021070
rect 67230 1021026 67347 1021036
rect 67002 1021002 67347 1021026
rect 67015 1020958 67215 1021002
rect 67230 1020992 67254 1021002
rect 67230 1020968 67264 1020992
rect 67275 1020968 67347 1021002
rect 67230 1020958 67347 1020968
rect 67002 1020934 67347 1020958
rect 67015 1020922 67215 1020934
rect 67026 1020910 67050 1020922
rect 67230 1020910 67254 1020934
rect 67275 1020922 67347 1020934
rect 67577 1020922 67633 1021922
rect 67649 1020922 67705 1021922
rect 68007 1021842 68207 1021922
rect 68222 1021852 68256 1021876
rect 68267 1021852 68339 1021922
rect 68222 1021842 68339 1021852
rect 67994 1021818 68339 1021842
rect 68007 1021774 68207 1021818
rect 68222 1021808 68246 1021818
rect 68222 1021784 68256 1021808
rect 68267 1021784 68339 1021818
rect 68222 1021774 68339 1021784
rect 67994 1021750 68339 1021774
rect 68007 1021706 68207 1021750
rect 68222 1021740 68246 1021750
rect 68222 1021716 68256 1021740
rect 68267 1021716 68339 1021750
rect 68222 1021706 68339 1021716
rect 67994 1021682 68339 1021706
rect 68007 1021638 68207 1021682
rect 68222 1021672 68246 1021682
rect 68222 1021648 68256 1021672
rect 68267 1021648 68339 1021682
rect 68222 1021638 68339 1021648
rect 67994 1021614 68339 1021638
rect 68007 1021570 68207 1021614
rect 68222 1021604 68246 1021614
rect 68222 1021580 68256 1021604
rect 68267 1021580 68339 1021614
rect 68222 1021570 68339 1021580
rect 67994 1021546 68339 1021570
rect 68007 1021502 68207 1021546
rect 68222 1021536 68246 1021546
rect 68222 1021512 68256 1021536
rect 68267 1021512 68339 1021546
rect 68222 1021502 68339 1021512
rect 67994 1021478 68339 1021502
rect 68007 1021434 68207 1021478
rect 68222 1021468 68246 1021478
rect 68222 1021444 68256 1021468
rect 68267 1021444 68339 1021478
rect 68222 1021434 68339 1021444
rect 67994 1021410 68339 1021434
rect 68007 1021366 68207 1021410
rect 68222 1021400 68246 1021410
rect 68222 1021376 68256 1021400
rect 68267 1021376 68339 1021410
rect 68222 1021366 68339 1021376
rect 67994 1021342 68339 1021366
rect 68007 1021298 68207 1021342
rect 68222 1021332 68246 1021342
rect 68222 1021308 68256 1021332
rect 68267 1021308 68339 1021342
rect 68222 1021298 68339 1021308
rect 67994 1021274 68339 1021298
rect 68007 1021230 68207 1021274
rect 68222 1021264 68246 1021274
rect 68222 1021240 68256 1021264
rect 68267 1021240 68339 1021274
rect 68222 1021230 68339 1021240
rect 67994 1021206 68339 1021230
rect 68007 1021162 68207 1021206
rect 68222 1021196 68246 1021206
rect 68222 1021172 68256 1021196
rect 68267 1021172 68339 1021206
rect 68222 1021162 68339 1021172
rect 67994 1021138 68339 1021162
rect 68007 1021094 68207 1021138
rect 68222 1021128 68246 1021138
rect 68222 1021104 68256 1021128
rect 68267 1021104 68339 1021138
rect 68222 1021094 68339 1021104
rect 67994 1021070 68339 1021094
rect 68007 1021026 68207 1021070
rect 68222 1021060 68246 1021070
rect 68222 1021036 68256 1021060
rect 68267 1021036 68339 1021070
rect 68222 1021026 68339 1021036
rect 67994 1021002 68339 1021026
rect 68007 1020958 68207 1021002
rect 68222 1020992 68246 1021002
rect 68222 1020968 68256 1020992
rect 68267 1020968 68339 1021002
rect 68222 1020958 68339 1020968
rect 67994 1020934 68339 1020958
rect 68007 1020922 68207 1020934
rect 68018 1020910 68042 1020922
rect 68222 1020910 68246 1020934
rect 68267 1020922 68339 1020934
rect 68569 1020922 68625 1021922
rect 68641 1020922 68697 1021922
rect 68999 1021842 69199 1021922
rect 69214 1021852 69248 1021876
rect 69259 1021852 69331 1021922
rect 69214 1021842 69331 1021852
rect 68986 1021818 69331 1021842
rect 68999 1021774 69199 1021818
rect 69214 1021808 69238 1021818
rect 69214 1021784 69248 1021808
rect 69259 1021784 69331 1021818
rect 69214 1021774 69331 1021784
rect 68986 1021750 69331 1021774
rect 68999 1021706 69199 1021750
rect 69214 1021740 69238 1021750
rect 69214 1021716 69248 1021740
rect 69259 1021716 69331 1021750
rect 69214 1021706 69331 1021716
rect 68986 1021682 69331 1021706
rect 68999 1021638 69199 1021682
rect 69214 1021672 69238 1021682
rect 69214 1021648 69248 1021672
rect 69259 1021648 69331 1021682
rect 69214 1021638 69331 1021648
rect 68986 1021614 69331 1021638
rect 68999 1021570 69199 1021614
rect 69214 1021604 69238 1021614
rect 69214 1021580 69248 1021604
rect 69259 1021580 69331 1021614
rect 69214 1021570 69331 1021580
rect 68986 1021546 69331 1021570
rect 68999 1021502 69199 1021546
rect 69214 1021536 69238 1021546
rect 69214 1021512 69248 1021536
rect 69259 1021512 69331 1021546
rect 69214 1021502 69331 1021512
rect 68986 1021478 69331 1021502
rect 68999 1021434 69199 1021478
rect 69214 1021468 69238 1021478
rect 69214 1021444 69248 1021468
rect 69259 1021444 69331 1021478
rect 69214 1021434 69331 1021444
rect 68986 1021410 69331 1021434
rect 68999 1021366 69199 1021410
rect 69214 1021400 69238 1021410
rect 69214 1021376 69248 1021400
rect 69259 1021376 69331 1021410
rect 69214 1021366 69331 1021376
rect 68986 1021342 69331 1021366
rect 68999 1021298 69199 1021342
rect 69214 1021332 69238 1021342
rect 69214 1021308 69248 1021332
rect 69259 1021308 69331 1021342
rect 69214 1021298 69331 1021308
rect 68986 1021274 69331 1021298
rect 68999 1021230 69199 1021274
rect 69214 1021264 69238 1021274
rect 69214 1021240 69248 1021264
rect 69259 1021240 69331 1021274
rect 69214 1021230 69331 1021240
rect 68986 1021206 69331 1021230
rect 68999 1021162 69199 1021206
rect 69214 1021196 69238 1021206
rect 69214 1021172 69248 1021196
rect 69259 1021172 69331 1021206
rect 69214 1021162 69331 1021172
rect 68986 1021138 69331 1021162
rect 68999 1021094 69199 1021138
rect 69214 1021128 69238 1021138
rect 69214 1021104 69248 1021128
rect 69259 1021104 69331 1021138
rect 69214 1021094 69331 1021104
rect 68986 1021070 69331 1021094
rect 68999 1021026 69199 1021070
rect 69214 1021060 69238 1021070
rect 69214 1021036 69248 1021060
rect 69259 1021036 69331 1021070
rect 69214 1021026 69331 1021036
rect 68986 1021002 69331 1021026
rect 68999 1020958 69199 1021002
rect 69214 1020992 69238 1021002
rect 69214 1020968 69248 1020992
rect 69259 1020968 69331 1021002
rect 69214 1020958 69331 1020968
rect 68986 1020934 69331 1020958
rect 68999 1020922 69199 1020934
rect 69010 1020910 69034 1020922
rect 69214 1020910 69238 1020934
rect 69259 1020922 69331 1020934
rect 69561 1020922 69617 1021922
rect 69633 1020922 69689 1021922
rect 69991 1021842 70191 1021922
rect 70206 1021852 70240 1021876
rect 70251 1021852 70323 1021922
rect 70206 1021842 70323 1021852
rect 69978 1021818 70323 1021842
rect 69991 1021774 70191 1021818
rect 70206 1021808 70230 1021818
rect 70206 1021784 70240 1021808
rect 70251 1021784 70323 1021818
rect 70206 1021774 70323 1021784
rect 69978 1021750 70323 1021774
rect 69991 1021706 70191 1021750
rect 70206 1021740 70230 1021750
rect 70206 1021716 70240 1021740
rect 70251 1021716 70323 1021750
rect 70206 1021706 70323 1021716
rect 69978 1021682 70323 1021706
rect 69991 1021638 70191 1021682
rect 70206 1021672 70230 1021682
rect 70206 1021648 70240 1021672
rect 70251 1021648 70323 1021682
rect 70206 1021638 70323 1021648
rect 69978 1021614 70323 1021638
rect 69991 1021570 70191 1021614
rect 70206 1021604 70230 1021614
rect 70206 1021580 70240 1021604
rect 70251 1021580 70323 1021614
rect 70206 1021570 70323 1021580
rect 69978 1021546 70323 1021570
rect 69991 1021502 70191 1021546
rect 70206 1021536 70230 1021546
rect 70206 1021512 70240 1021536
rect 70251 1021512 70323 1021546
rect 70206 1021502 70323 1021512
rect 69978 1021478 70323 1021502
rect 69991 1021434 70191 1021478
rect 70206 1021468 70230 1021478
rect 70206 1021444 70240 1021468
rect 70251 1021444 70323 1021478
rect 70206 1021434 70323 1021444
rect 69978 1021410 70323 1021434
rect 69991 1021366 70191 1021410
rect 70206 1021400 70230 1021410
rect 70206 1021376 70240 1021400
rect 70251 1021376 70323 1021410
rect 70206 1021366 70323 1021376
rect 69978 1021342 70323 1021366
rect 69991 1021298 70191 1021342
rect 70206 1021332 70230 1021342
rect 70206 1021308 70240 1021332
rect 70251 1021308 70323 1021342
rect 70206 1021298 70323 1021308
rect 69978 1021274 70323 1021298
rect 69991 1021230 70191 1021274
rect 70206 1021264 70230 1021274
rect 70206 1021240 70240 1021264
rect 70251 1021240 70323 1021274
rect 70206 1021230 70323 1021240
rect 69978 1021206 70323 1021230
rect 69991 1021162 70191 1021206
rect 70206 1021196 70230 1021206
rect 70206 1021172 70240 1021196
rect 70251 1021172 70323 1021206
rect 70206 1021162 70323 1021172
rect 69978 1021138 70323 1021162
rect 69991 1021094 70191 1021138
rect 70206 1021128 70230 1021138
rect 70206 1021104 70240 1021128
rect 70251 1021104 70323 1021138
rect 70206 1021094 70323 1021104
rect 69978 1021070 70323 1021094
rect 69991 1021026 70191 1021070
rect 70206 1021060 70230 1021070
rect 70206 1021036 70240 1021060
rect 70251 1021036 70323 1021070
rect 70206 1021026 70323 1021036
rect 69978 1021002 70323 1021026
rect 69991 1020958 70191 1021002
rect 70206 1020992 70230 1021002
rect 70206 1020968 70240 1020992
rect 70251 1020968 70323 1021002
rect 70206 1020958 70323 1020968
rect 69978 1020934 70323 1020958
rect 69991 1020922 70191 1020934
rect 70002 1020910 70026 1020922
rect 70206 1020910 70230 1020934
rect 70251 1020922 70323 1020934
rect 70553 1020922 70609 1021922
rect 70625 1020922 70681 1021922
rect 70983 1021842 71183 1021922
rect 71198 1021852 71232 1021876
rect 71243 1021852 71315 1021922
rect 71198 1021842 71315 1021852
rect 70970 1021818 71315 1021842
rect 70983 1021774 71183 1021818
rect 71198 1021808 71222 1021818
rect 71198 1021784 71232 1021808
rect 71243 1021784 71315 1021818
rect 71198 1021774 71315 1021784
rect 70970 1021750 71315 1021774
rect 70983 1021706 71183 1021750
rect 71198 1021740 71222 1021750
rect 71198 1021716 71232 1021740
rect 71243 1021716 71315 1021750
rect 71198 1021706 71315 1021716
rect 70970 1021682 71315 1021706
rect 70983 1021638 71183 1021682
rect 71198 1021672 71222 1021682
rect 71198 1021648 71232 1021672
rect 71243 1021648 71315 1021682
rect 71198 1021638 71315 1021648
rect 70970 1021614 71315 1021638
rect 70983 1021570 71183 1021614
rect 71198 1021604 71222 1021614
rect 71198 1021580 71232 1021604
rect 71243 1021580 71315 1021614
rect 71198 1021570 71315 1021580
rect 70970 1021546 71315 1021570
rect 70983 1021502 71183 1021546
rect 71198 1021536 71222 1021546
rect 71198 1021512 71232 1021536
rect 71243 1021512 71315 1021546
rect 71198 1021502 71315 1021512
rect 70970 1021478 71315 1021502
rect 70983 1021434 71183 1021478
rect 71198 1021468 71222 1021478
rect 71198 1021444 71232 1021468
rect 71243 1021444 71315 1021478
rect 71198 1021434 71315 1021444
rect 70970 1021410 71315 1021434
rect 70983 1021366 71183 1021410
rect 71198 1021400 71222 1021410
rect 71198 1021376 71232 1021400
rect 71243 1021376 71315 1021410
rect 71198 1021366 71315 1021376
rect 70970 1021342 71315 1021366
rect 70983 1021298 71183 1021342
rect 71198 1021332 71222 1021342
rect 71198 1021308 71232 1021332
rect 71243 1021308 71315 1021342
rect 71198 1021298 71315 1021308
rect 70970 1021274 71315 1021298
rect 70983 1021230 71183 1021274
rect 71198 1021264 71222 1021274
rect 71198 1021240 71232 1021264
rect 71243 1021240 71315 1021274
rect 71198 1021230 71315 1021240
rect 70970 1021206 71315 1021230
rect 70983 1021162 71183 1021206
rect 71198 1021196 71222 1021206
rect 71198 1021172 71232 1021196
rect 71243 1021172 71315 1021206
rect 71198 1021162 71315 1021172
rect 70970 1021138 71315 1021162
rect 70983 1021094 71183 1021138
rect 71198 1021128 71222 1021138
rect 71198 1021104 71232 1021128
rect 71243 1021104 71315 1021138
rect 71198 1021094 71315 1021104
rect 70970 1021070 71315 1021094
rect 70983 1021026 71183 1021070
rect 71198 1021060 71222 1021070
rect 71198 1021036 71232 1021060
rect 71243 1021036 71315 1021070
rect 71198 1021026 71315 1021036
rect 70970 1021002 71315 1021026
rect 70983 1020958 71183 1021002
rect 71198 1020992 71222 1021002
rect 71198 1020968 71232 1020992
rect 71243 1020968 71315 1021002
rect 71198 1020958 71315 1020968
rect 70970 1020934 71315 1020958
rect 70983 1020922 71183 1020934
rect 70994 1020910 71018 1020922
rect 71198 1020910 71222 1020934
rect 71243 1020922 71315 1020934
rect 71545 1020922 71601 1021922
rect 71617 1020922 71673 1021922
rect 71975 1021842 72175 1021922
rect 72190 1021852 72224 1021876
rect 72235 1021852 72307 1021922
rect 72190 1021842 72307 1021852
rect 71962 1021818 72307 1021842
rect 71975 1021774 72175 1021818
rect 72190 1021808 72214 1021818
rect 72190 1021784 72224 1021808
rect 72235 1021784 72307 1021818
rect 72190 1021774 72307 1021784
rect 71962 1021750 72307 1021774
rect 71975 1021706 72175 1021750
rect 72190 1021740 72214 1021750
rect 72190 1021716 72224 1021740
rect 72235 1021716 72307 1021750
rect 72190 1021706 72307 1021716
rect 71962 1021682 72307 1021706
rect 71975 1021638 72175 1021682
rect 72190 1021672 72214 1021682
rect 72190 1021648 72224 1021672
rect 72235 1021648 72307 1021682
rect 72190 1021638 72307 1021648
rect 71962 1021614 72307 1021638
rect 71975 1021570 72175 1021614
rect 72190 1021604 72214 1021614
rect 72190 1021580 72224 1021604
rect 72235 1021580 72307 1021614
rect 72190 1021570 72307 1021580
rect 71962 1021546 72307 1021570
rect 71975 1021502 72175 1021546
rect 72190 1021536 72214 1021546
rect 72190 1021512 72224 1021536
rect 72235 1021512 72307 1021546
rect 72190 1021502 72307 1021512
rect 71962 1021478 72307 1021502
rect 71975 1021434 72175 1021478
rect 72190 1021468 72214 1021478
rect 72190 1021444 72224 1021468
rect 72235 1021444 72307 1021478
rect 72190 1021434 72307 1021444
rect 71962 1021410 72307 1021434
rect 71975 1021366 72175 1021410
rect 72190 1021400 72214 1021410
rect 72190 1021376 72224 1021400
rect 72235 1021376 72307 1021410
rect 72190 1021366 72307 1021376
rect 71962 1021342 72307 1021366
rect 71975 1021298 72175 1021342
rect 72190 1021332 72214 1021342
rect 72190 1021308 72224 1021332
rect 72235 1021308 72307 1021342
rect 72190 1021298 72307 1021308
rect 71962 1021274 72307 1021298
rect 71975 1021230 72175 1021274
rect 72190 1021264 72214 1021274
rect 72190 1021240 72224 1021264
rect 72235 1021240 72307 1021274
rect 72190 1021230 72307 1021240
rect 71962 1021206 72307 1021230
rect 71975 1021162 72175 1021206
rect 72190 1021196 72214 1021206
rect 72190 1021172 72224 1021196
rect 72235 1021172 72307 1021206
rect 72190 1021162 72307 1021172
rect 71962 1021138 72307 1021162
rect 71975 1021094 72175 1021138
rect 72190 1021128 72214 1021138
rect 72190 1021104 72224 1021128
rect 72235 1021104 72307 1021138
rect 72190 1021094 72307 1021104
rect 71962 1021070 72307 1021094
rect 71975 1021026 72175 1021070
rect 72190 1021060 72214 1021070
rect 72190 1021036 72224 1021060
rect 72235 1021036 72307 1021070
rect 72190 1021026 72307 1021036
rect 71962 1021002 72307 1021026
rect 71975 1020958 72175 1021002
rect 72190 1020992 72214 1021002
rect 72190 1020968 72224 1020992
rect 72235 1020968 72307 1021002
rect 72190 1020958 72307 1020968
rect 71962 1020934 72307 1020958
rect 71975 1020922 72175 1020934
rect 71986 1020910 72010 1020922
rect 72190 1020910 72214 1020934
rect 72235 1020922 72307 1020934
rect 72537 1020922 72593 1021922
rect 72609 1020922 72665 1021922
rect 72967 1021842 73167 1021922
rect 73182 1021852 73216 1021876
rect 73227 1021852 73299 1021922
rect 73182 1021842 73299 1021852
rect 72954 1021818 73299 1021842
rect 72967 1021774 73167 1021818
rect 73182 1021808 73206 1021818
rect 73182 1021784 73216 1021808
rect 73227 1021784 73299 1021818
rect 73182 1021774 73299 1021784
rect 72954 1021750 73299 1021774
rect 72967 1021706 73167 1021750
rect 73182 1021740 73206 1021750
rect 73182 1021716 73216 1021740
rect 73227 1021716 73299 1021750
rect 73182 1021706 73299 1021716
rect 72954 1021682 73299 1021706
rect 72967 1021638 73167 1021682
rect 73182 1021672 73206 1021682
rect 73182 1021648 73216 1021672
rect 73227 1021648 73299 1021682
rect 73182 1021638 73299 1021648
rect 72954 1021614 73299 1021638
rect 72967 1021570 73167 1021614
rect 73182 1021604 73206 1021614
rect 73182 1021580 73216 1021604
rect 73227 1021580 73299 1021614
rect 73182 1021570 73299 1021580
rect 72954 1021546 73299 1021570
rect 72967 1021502 73167 1021546
rect 73182 1021536 73206 1021546
rect 73182 1021512 73216 1021536
rect 73227 1021512 73299 1021546
rect 73182 1021502 73299 1021512
rect 72954 1021478 73299 1021502
rect 72967 1021434 73167 1021478
rect 73182 1021468 73206 1021478
rect 73182 1021444 73216 1021468
rect 73227 1021444 73299 1021478
rect 73182 1021434 73299 1021444
rect 72954 1021410 73299 1021434
rect 72967 1021366 73167 1021410
rect 73182 1021400 73206 1021410
rect 73182 1021376 73216 1021400
rect 73227 1021376 73299 1021410
rect 73182 1021366 73299 1021376
rect 72954 1021342 73299 1021366
rect 72967 1021298 73167 1021342
rect 73182 1021332 73206 1021342
rect 73182 1021308 73216 1021332
rect 73227 1021308 73299 1021342
rect 73182 1021298 73299 1021308
rect 72954 1021274 73299 1021298
rect 72967 1021230 73167 1021274
rect 73182 1021264 73206 1021274
rect 73182 1021240 73216 1021264
rect 73227 1021240 73299 1021274
rect 73182 1021230 73299 1021240
rect 72954 1021206 73299 1021230
rect 72967 1021162 73167 1021206
rect 73182 1021196 73206 1021206
rect 73182 1021172 73216 1021196
rect 73227 1021172 73299 1021206
rect 73182 1021162 73299 1021172
rect 72954 1021138 73299 1021162
rect 72967 1021094 73167 1021138
rect 73182 1021128 73206 1021138
rect 73182 1021104 73216 1021128
rect 73227 1021104 73299 1021138
rect 73182 1021094 73299 1021104
rect 72954 1021070 73299 1021094
rect 72967 1021026 73167 1021070
rect 73182 1021060 73206 1021070
rect 73182 1021036 73216 1021060
rect 73227 1021036 73299 1021070
rect 73182 1021026 73299 1021036
rect 72954 1021002 73299 1021026
rect 72967 1020958 73167 1021002
rect 73182 1020992 73206 1021002
rect 73182 1020968 73216 1020992
rect 73227 1020968 73299 1021002
rect 73182 1020958 73299 1020968
rect 72954 1020934 73299 1020958
rect 72967 1020922 73167 1020934
rect 72978 1020910 73002 1020922
rect 73182 1020910 73206 1020934
rect 73227 1020922 73299 1020934
rect 73529 1020922 73585 1021922
rect 73601 1020922 73657 1021922
rect 73959 1021842 74159 1021922
rect 74174 1021852 74208 1021876
rect 74219 1021852 74291 1021922
rect 74174 1021842 74291 1021852
rect 73946 1021818 74291 1021842
rect 73959 1021774 74159 1021818
rect 74174 1021808 74198 1021818
rect 74174 1021784 74208 1021808
rect 74219 1021784 74291 1021818
rect 74174 1021774 74291 1021784
rect 73946 1021750 74291 1021774
rect 73959 1021706 74159 1021750
rect 74174 1021740 74198 1021750
rect 74174 1021716 74208 1021740
rect 74219 1021716 74291 1021750
rect 74174 1021706 74291 1021716
rect 73946 1021682 74291 1021706
rect 73959 1021638 74159 1021682
rect 74174 1021672 74198 1021682
rect 74174 1021648 74208 1021672
rect 74219 1021648 74291 1021682
rect 74174 1021638 74291 1021648
rect 73946 1021614 74291 1021638
rect 73959 1021570 74159 1021614
rect 74174 1021604 74198 1021614
rect 74174 1021580 74208 1021604
rect 74219 1021580 74291 1021614
rect 74174 1021570 74291 1021580
rect 73946 1021546 74291 1021570
rect 73959 1021502 74159 1021546
rect 74174 1021536 74198 1021546
rect 74174 1021512 74208 1021536
rect 74219 1021512 74291 1021546
rect 74174 1021502 74291 1021512
rect 73946 1021478 74291 1021502
rect 73959 1021434 74159 1021478
rect 74174 1021468 74198 1021478
rect 74174 1021444 74208 1021468
rect 74219 1021444 74291 1021478
rect 74174 1021434 74291 1021444
rect 73946 1021410 74291 1021434
rect 73959 1021366 74159 1021410
rect 74174 1021400 74198 1021410
rect 74174 1021376 74208 1021400
rect 74219 1021376 74291 1021410
rect 74174 1021366 74291 1021376
rect 73946 1021342 74291 1021366
rect 73959 1021298 74159 1021342
rect 74174 1021332 74198 1021342
rect 74174 1021308 74208 1021332
rect 74219 1021308 74291 1021342
rect 74174 1021298 74291 1021308
rect 73946 1021274 74291 1021298
rect 73959 1021230 74159 1021274
rect 74174 1021264 74198 1021274
rect 74174 1021240 74208 1021264
rect 74219 1021240 74291 1021274
rect 74174 1021230 74291 1021240
rect 73946 1021206 74291 1021230
rect 73959 1021162 74159 1021206
rect 74174 1021196 74198 1021206
rect 74174 1021172 74208 1021196
rect 74219 1021172 74291 1021206
rect 74174 1021162 74291 1021172
rect 73946 1021138 74291 1021162
rect 73959 1021094 74159 1021138
rect 74174 1021128 74198 1021138
rect 74174 1021104 74208 1021128
rect 74219 1021104 74291 1021138
rect 74174 1021094 74291 1021104
rect 73946 1021070 74291 1021094
rect 73959 1021026 74159 1021070
rect 74174 1021060 74198 1021070
rect 74174 1021036 74208 1021060
rect 74219 1021036 74291 1021070
rect 74174 1021026 74291 1021036
rect 73946 1021002 74291 1021026
rect 73959 1020958 74159 1021002
rect 74174 1020992 74198 1021002
rect 74174 1020968 74208 1020992
rect 74219 1020968 74291 1021002
rect 74174 1020958 74291 1020968
rect 73946 1020934 74291 1020958
rect 73959 1020922 74159 1020934
rect 73970 1020910 73994 1020922
rect 74174 1020910 74198 1020934
rect 74219 1020922 74291 1020934
rect 74521 1020922 74577 1021922
rect 74593 1020922 74649 1021922
rect 74951 1021842 75151 1021922
rect 75166 1021852 75200 1021876
rect 75211 1021852 75283 1021922
rect 75166 1021842 75283 1021852
rect 74938 1021818 75283 1021842
rect 74951 1021774 75151 1021818
rect 75166 1021808 75190 1021818
rect 75166 1021784 75200 1021808
rect 75211 1021784 75283 1021818
rect 75166 1021774 75283 1021784
rect 74938 1021750 75283 1021774
rect 74951 1021706 75151 1021750
rect 75166 1021740 75190 1021750
rect 75166 1021716 75200 1021740
rect 75211 1021716 75283 1021750
rect 75166 1021706 75283 1021716
rect 74938 1021682 75283 1021706
rect 74951 1021638 75151 1021682
rect 75166 1021672 75190 1021682
rect 75166 1021648 75200 1021672
rect 75211 1021648 75283 1021682
rect 75166 1021638 75283 1021648
rect 74938 1021614 75283 1021638
rect 74951 1021570 75151 1021614
rect 75166 1021604 75190 1021614
rect 75166 1021580 75200 1021604
rect 75211 1021580 75283 1021614
rect 75166 1021570 75283 1021580
rect 74938 1021546 75283 1021570
rect 74951 1021502 75151 1021546
rect 75166 1021536 75190 1021546
rect 75166 1021512 75200 1021536
rect 75211 1021512 75283 1021546
rect 75166 1021502 75283 1021512
rect 74938 1021478 75283 1021502
rect 74951 1021434 75151 1021478
rect 75166 1021468 75190 1021478
rect 75166 1021444 75200 1021468
rect 75211 1021444 75283 1021478
rect 75166 1021434 75283 1021444
rect 74938 1021410 75283 1021434
rect 74951 1021366 75151 1021410
rect 75166 1021400 75190 1021410
rect 75166 1021376 75200 1021400
rect 75211 1021376 75283 1021410
rect 75166 1021366 75283 1021376
rect 74938 1021342 75283 1021366
rect 74951 1021298 75151 1021342
rect 75166 1021332 75190 1021342
rect 75166 1021308 75200 1021332
rect 75211 1021308 75283 1021342
rect 75166 1021298 75283 1021308
rect 74938 1021274 75283 1021298
rect 74951 1021230 75151 1021274
rect 75166 1021264 75190 1021274
rect 75166 1021240 75200 1021264
rect 75211 1021240 75283 1021274
rect 75166 1021230 75283 1021240
rect 74938 1021206 75283 1021230
rect 74951 1021162 75151 1021206
rect 75166 1021196 75190 1021206
rect 75166 1021172 75200 1021196
rect 75211 1021172 75283 1021206
rect 75166 1021162 75283 1021172
rect 74938 1021138 75283 1021162
rect 74951 1021094 75151 1021138
rect 75166 1021128 75190 1021138
rect 75166 1021104 75200 1021128
rect 75211 1021104 75283 1021138
rect 75166 1021094 75283 1021104
rect 74938 1021070 75283 1021094
rect 74951 1021026 75151 1021070
rect 75166 1021060 75190 1021070
rect 75166 1021036 75200 1021060
rect 75211 1021036 75283 1021070
rect 75166 1021026 75283 1021036
rect 74938 1021002 75283 1021026
rect 74951 1020958 75151 1021002
rect 75166 1020992 75190 1021002
rect 75166 1020968 75200 1020992
rect 75211 1020968 75283 1021002
rect 75166 1020958 75283 1020968
rect 74938 1020934 75283 1020958
rect 74951 1020922 75151 1020934
rect 74962 1020910 74986 1020922
rect 75166 1020910 75190 1020934
rect 75211 1020922 75283 1020934
rect 75472 1020922 75544 1021922
rect 75610 1020922 75627 1021922
rect 75797 1020922 75830 1021922
rect 75953 1021730 76025 1021760
rect 75953 1021692 75987 1021722
rect 63058 1020322 63092 1020334
rect 62356 1019322 62406 1020322
rect 62617 1019322 62673 1020322
rect 62689 1019322 62745 1020322
rect 63047 1020300 63247 1020322
rect 63262 1020310 63296 1020334
rect 64050 1020322 64084 1020334
rect 63307 1020310 63379 1020322
rect 63262 1020300 63379 1020310
rect 63034 1020276 63379 1020300
rect 63047 1020232 63247 1020276
rect 63262 1020266 63286 1020276
rect 63262 1020242 63296 1020266
rect 63307 1020242 63379 1020276
rect 63262 1020232 63379 1020242
rect 63034 1020208 63379 1020232
rect 63047 1020164 63247 1020208
rect 63262 1020198 63286 1020208
rect 63262 1020174 63296 1020198
rect 63307 1020174 63379 1020208
rect 63262 1020164 63379 1020174
rect 63034 1020140 63379 1020164
rect 63047 1020096 63247 1020140
rect 63262 1020130 63286 1020140
rect 63262 1020106 63296 1020130
rect 63307 1020106 63379 1020140
rect 63262 1020096 63379 1020106
rect 63034 1020072 63379 1020096
rect 63047 1020028 63247 1020072
rect 63262 1020062 63286 1020072
rect 63262 1020038 63296 1020062
rect 63307 1020038 63379 1020072
rect 63262 1020028 63379 1020038
rect 63034 1020004 63379 1020028
rect 63047 1019960 63247 1020004
rect 63262 1019994 63286 1020004
rect 63262 1019970 63296 1019994
rect 63307 1019970 63379 1020004
rect 63262 1019960 63379 1019970
rect 63034 1019936 63379 1019960
rect 63047 1019892 63247 1019936
rect 63262 1019926 63286 1019936
rect 63262 1019902 63296 1019926
rect 63307 1019902 63379 1019936
rect 63262 1019892 63379 1019902
rect 63034 1019868 63379 1019892
rect 63047 1019824 63247 1019868
rect 63262 1019858 63286 1019868
rect 63262 1019834 63296 1019858
rect 63307 1019834 63379 1019868
rect 63262 1019824 63379 1019834
rect 63034 1019800 63379 1019824
rect 63047 1019756 63247 1019800
rect 63262 1019790 63286 1019800
rect 63262 1019766 63296 1019790
rect 63307 1019766 63379 1019800
rect 63262 1019756 63379 1019766
rect 63034 1019732 63379 1019756
rect 63047 1019688 63247 1019732
rect 63262 1019722 63286 1019732
rect 63262 1019698 63296 1019722
rect 63307 1019698 63379 1019732
rect 63262 1019688 63379 1019698
rect 63034 1019664 63379 1019688
rect 63047 1019620 63247 1019664
rect 63262 1019654 63286 1019664
rect 63262 1019630 63296 1019654
rect 63307 1019630 63379 1019664
rect 63262 1019620 63379 1019630
rect 63034 1019596 63379 1019620
rect 63047 1019552 63247 1019596
rect 63262 1019586 63286 1019596
rect 63262 1019562 63296 1019586
rect 63307 1019562 63379 1019596
rect 63262 1019552 63379 1019562
rect 63034 1019528 63379 1019552
rect 63047 1019484 63247 1019528
rect 63262 1019518 63286 1019528
rect 63262 1019494 63296 1019518
rect 63307 1019494 63379 1019528
rect 63262 1019484 63379 1019494
rect 63034 1019460 63379 1019484
rect 63047 1019416 63247 1019460
rect 63262 1019450 63286 1019460
rect 63262 1019426 63296 1019450
rect 63307 1019426 63379 1019460
rect 63262 1019416 63379 1019426
rect 63034 1019392 63379 1019416
rect 63047 1019322 63247 1019392
rect 63262 1019368 63286 1019392
rect 63307 1019322 63379 1019392
rect 63609 1019322 63665 1020322
rect 63681 1019322 63737 1020322
rect 64039 1020300 64239 1020322
rect 64254 1020310 64288 1020334
rect 65042 1020322 65076 1020334
rect 64299 1020310 64371 1020322
rect 64254 1020300 64371 1020310
rect 64026 1020276 64371 1020300
rect 64039 1020232 64239 1020276
rect 64254 1020266 64278 1020276
rect 64254 1020242 64288 1020266
rect 64299 1020242 64371 1020276
rect 64254 1020232 64371 1020242
rect 64026 1020208 64371 1020232
rect 64039 1020164 64239 1020208
rect 64254 1020198 64278 1020208
rect 64254 1020174 64288 1020198
rect 64299 1020174 64371 1020208
rect 64254 1020164 64371 1020174
rect 64026 1020140 64371 1020164
rect 64039 1020096 64239 1020140
rect 64254 1020130 64278 1020140
rect 64254 1020106 64288 1020130
rect 64299 1020106 64371 1020140
rect 64254 1020096 64371 1020106
rect 64026 1020072 64371 1020096
rect 64039 1020028 64239 1020072
rect 64254 1020062 64278 1020072
rect 64254 1020038 64288 1020062
rect 64299 1020038 64371 1020072
rect 64254 1020028 64371 1020038
rect 64026 1020004 64371 1020028
rect 64039 1019960 64239 1020004
rect 64254 1019994 64278 1020004
rect 64254 1019970 64288 1019994
rect 64299 1019970 64371 1020004
rect 64254 1019960 64371 1019970
rect 64026 1019936 64371 1019960
rect 64039 1019892 64239 1019936
rect 64254 1019926 64278 1019936
rect 64254 1019902 64288 1019926
rect 64299 1019902 64371 1019936
rect 64254 1019892 64371 1019902
rect 64026 1019868 64371 1019892
rect 64039 1019824 64239 1019868
rect 64254 1019858 64278 1019868
rect 64254 1019834 64288 1019858
rect 64299 1019834 64371 1019868
rect 64254 1019824 64371 1019834
rect 64026 1019800 64371 1019824
rect 64039 1019756 64239 1019800
rect 64254 1019790 64278 1019800
rect 64254 1019766 64288 1019790
rect 64299 1019766 64371 1019800
rect 64254 1019756 64371 1019766
rect 64026 1019732 64371 1019756
rect 64039 1019688 64239 1019732
rect 64254 1019722 64278 1019732
rect 64254 1019698 64288 1019722
rect 64299 1019698 64371 1019732
rect 64254 1019688 64371 1019698
rect 64026 1019664 64371 1019688
rect 64039 1019620 64239 1019664
rect 64254 1019654 64278 1019664
rect 64254 1019630 64288 1019654
rect 64299 1019630 64371 1019664
rect 64254 1019620 64371 1019630
rect 64026 1019596 64371 1019620
rect 64039 1019552 64239 1019596
rect 64254 1019586 64278 1019596
rect 64254 1019562 64288 1019586
rect 64299 1019562 64371 1019596
rect 64254 1019552 64371 1019562
rect 64026 1019528 64371 1019552
rect 64039 1019484 64239 1019528
rect 64254 1019518 64278 1019528
rect 64254 1019494 64288 1019518
rect 64299 1019494 64371 1019528
rect 64254 1019484 64371 1019494
rect 64026 1019460 64371 1019484
rect 64039 1019416 64239 1019460
rect 64254 1019450 64278 1019460
rect 64254 1019426 64288 1019450
rect 64299 1019426 64371 1019460
rect 64254 1019416 64371 1019426
rect 64026 1019392 64371 1019416
rect 64039 1019322 64239 1019392
rect 64254 1019368 64278 1019392
rect 64299 1019322 64371 1019392
rect 64601 1019322 64657 1020322
rect 64673 1019322 64729 1020322
rect 65031 1020300 65231 1020322
rect 65246 1020310 65280 1020334
rect 66034 1020322 66068 1020334
rect 65291 1020310 65363 1020322
rect 65246 1020300 65363 1020310
rect 65018 1020276 65363 1020300
rect 65031 1020232 65231 1020276
rect 65246 1020266 65270 1020276
rect 65246 1020242 65280 1020266
rect 65291 1020242 65363 1020276
rect 65246 1020232 65363 1020242
rect 65018 1020208 65363 1020232
rect 65031 1020164 65231 1020208
rect 65246 1020198 65270 1020208
rect 65246 1020174 65280 1020198
rect 65291 1020174 65363 1020208
rect 65246 1020164 65363 1020174
rect 65018 1020140 65363 1020164
rect 65031 1020096 65231 1020140
rect 65246 1020130 65270 1020140
rect 65246 1020106 65280 1020130
rect 65291 1020106 65363 1020140
rect 65246 1020096 65363 1020106
rect 65018 1020072 65363 1020096
rect 65031 1020028 65231 1020072
rect 65246 1020062 65270 1020072
rect 65246 1020038 65280 1020062
rect 65291 1020038 65363 1020072
rect 65246 1020028 65363 1020038
rect 65018 1020004 65363 1020028
rect 65031 1019960 65231 1020004
rect 65246 1019994 65270 1020004
rect 65246 1019970 65280 1019994
rect 65291 1019970 65363 1020004
rect 65246 1019960 65363 1019970
rect 65018 1019936 65363 1019960
rect 65031 1019892 65231 1019936
rect 65246 1019926 65270 1019936
rect 65246 1019902 65280 1019926
rect 65291 1019902 65363 1019936
rect 65246 1019892 65363 1019902
rect 65018 1019868 65363 1019892
rect 65031 1019824 65231 1019868
rect 65246 1019858 65270 1019868
rect 65246 1019834 65280 1019858
rect 65291 1019834 65363 1019868
rect 65246 1019824 65363 1019834
rect 65018 1019800 65363 1019824
rect 65031 1019756 65231 1019800
rect 65246 1019790 65270 1019800
rect 65246 1019766 65280 1019790
rect 65291 1019766 65363 1019800
rect 65246 1019756 65363 1019766
rect 65018 1019732 65363 1019756
rect 65031 1019688 65231 1019732
rect 65246 1019722 65270 1019732
rect 65246 1019698 65280 1019722
rect 65291 1019698 65363 1019732
rect 65246 1019688 65363 1019698
rect 65018 1019664 65363 1019688
rect 65031 1019620 65231 1019664
rect 65246 1019654 65270 1019664
rect 65246 1019630 65280 1019654
rect 65291 1019630 65363 1019664
rect 65246 1019620 65363 1019630
rect 65018 1019596 65363 1019620
rect 65031 1019552 65231 1019596
rect 65246 1019586 65270 1019596
rect 65246 1019562 65280 1019586
rect 65291 1019562 65363 1019596
rect 65246 1019552 65363 1019562
rect 65018 1019528 65363 1019552
rect 65031 1019484 65231 1019528
rect 65246 1019518 65270 1019528
rect 65246 1019494 65280 1019518
rect 65291 1019494 65363 1019528
rect 65246 1019484 65363 1019494
rect 65018 1019460 65363 1019484
rect 65031 1019416 65231 1019460
rect 65246 1019450 65270 1019460
rect 65246 1019426 65280 1019450
rect 65291 1019426 65363 1019460
rect 65246 1019416 65363 1019426
rect 65018 1019392 65363 1019416
rect 65031 1019322 65231 1019392
rect 65246 1019368 65270 1019392
rect 65291 1019322 65363 1019392
rect 65593 1019322 65649 1020322
rect 65665 1019322 65721 1020322
rect 66023 1020300 66223 1020322
rect 66238 1020310 66272 1020334
rect 67026 1020322 67060 1020334
rect 66283 1020310 66355 1020322
rect 66238 1020300 66355 1020310
rect 66010 1020276 66355 1020300
rect 66023 1020232 66223 1020276
rect 66238 1020266 66262 1020276
rect 66238 1020242 66272 1020266
rect 66283 1020242 66355 1020276
rect 66238 1020232 66355 1020242
rect 66010 1020208 66355 1020232
rect 66023 1020164 66223 1020208
rect 66238 1020198 66262 1020208
rect 66238 1020174 66272 1020198
rect 66283 1020174 66355 1020208
rect 66238 1020164 66355 1020174
rect 66010 1020140 66355 1020164
rect 66023 1020096 66223 1020140
rect 66238 1020130 66262 1020140
rect 66238 1020106 66272 1020130
rect 66283 1020106 66355 1020140
rect 66238 1020096 66355 1020106
rect 66010 1020072 66355 1020096
rect 66023 1020028 66223 1020072
rect 66238 1020062 66262 1020072
rect 66238 1020038 66272 1020062
rect 66283 1020038 66355 1020072
rect 66238 1020028 66355 1020038
rect 66010 1020004 66355 1020028
rect 66023 1019960 66223 1020004
rect 66238 1019994 66262 1020004
rect 66238 1019970 66272 1019994
rect 66283 1019970 66355 1020004
rect 66238 1019960 66355 1019970
rect 66010 1019936 66355 1019960
rect 66023 1019892 66223 1019936
rect 66238 1019926 66262 1019936
rect 66238 1019902 66272 1019926
rect 66283 1019902 66355 1019936
rect 66238 1019892 66355 1019902
rect 66010 1019868 66355 1019892
rect 66023 1019824 66223 1019868
rect 66238 1019858 66262 1019868
rect 66238 1019834 66272 1019858
rect 66283 1019834 66355 1019868
rect 66238 1019824 66355 1019834
rect 66010 1019800 66355 1019824
rect 66023 1019756 66223 1019800
rect 66238 1019790 66262 1019800
rect 66238 1019766 66272 1019790
rect 66283 1019766 66355 1019800
rect 66238 1019756 66355 1019766
rect 66010 1019732 66355 1019756
rect 66023 1019688 66223 1019732
rect 66238 1019722 66262 1019732
rect 66238 1019698 66272 1019722
rect 66283 1019698 66355 1019732
rect 66238 1019688 66355 1019698
rect 66010 1019664 66355 1019688
rect 66023 1019620 66223 1019664
rect 66238 1019654 66262 1019664
rect 66238 1019630 66272 1019654
rect 66283 1019630 66355 1019664
rect 66238 1019620 66355 1019630
rect 66010 1019596 66355 1019620
rect 66023 1019552 66223 1019596
rect 66238 1019586 66262 1019596
rect 66238 1019562 66272 1019586
rect 66283 1019562 66355 1019596
rect 66238 1019552 66355 1019562
rect 66010 1019528 66355 1019552
rect 66023 1019484 66223 1019528
rect 66238 1019518 66262 1019528
rect 66238 1019494 66272 1019518
rect 66283 1019494 66355 1019528
rect 66238 1019484 66355 1019494
rect 66010 1019460 66355 1019484
rect 66023 1019416 66223 1019460
rect 66238 1019450 66262 1019460
rect 66238 1019426 66272 1019450
rect 66283 1019426 66355 1019460
rect 66238 1019416 66355 1019426
rect 66010 1019392 66355 1019416
rect 66023 1019322 66223 1019392
rect 66238 1019368 66262 1019392
rect 66283 1019322 66355 1019392
rect 66585 1019322 66641 1020322
rect 66657 1019322 66713 1020322
rect 67015 1020300 67215 1020322
rect 67230 1020310 67264 1020334
rect 68018 1020322 68052 1020334
rect 67275 1020310 67347 1020322
rect 67230 1020300 67347 1020310
rect 67002 1020276 67347 1020300
rect 67015 1020232 67215 1020276
rect 67230 1020266 67254 1020276
rect 67230 1020242 67264 1020266
rect 67275 1020242 67347 1020276
rect 67230 1020232 67347 1020242
rect 67002 1020208 67347 1020232
rect 67015 1020164 67215 1020208
rect 67230 1020198 67254 1020208
rect 67230 1020174 67264 1020198
rect 67275 1020174 67347 1020208
rect 67230 1020164 67347 1020174
rect 67002 1020140 67347 1020164
rect 67015 1020096 67215 1020140
rect 67230 1020130 67254 1020140
rect 67230 1020106 67264 1020130
rect 67275 1020106 67347 1020140
rect 67230 1020096 67347 1020106
rect 67002 1020072 67347 1020096
rect 67015 1020028 67215 1020072
rect 67230 1020062 67254 1020072
rect 67230 1020038 67264 1020062
rect 67275 1020038 67347 1020072
rect 67230 1020028 67347 1020038
rect 67002 1020004 67347 1020028
rect 67015 1019960 67215 1020004
rect 67230 1019994 67254 1020004
rect 67230 1019970 67264 1019994
rect 67275 1019970 67347 1020004
rect 67230 1019960 67347 1019970
rect 67002 1019936 67347 1019960
rect 67015 1019892 67215 1019936
rect 67230 1019926 67254 1019936
rect 67230 1019902 67264 1019926
rect 67275 1019902 67347 1019936
rect 67230 1019892 67347 1019902
rect 67002 1019868 67347 1019892
rect 67015 1019824 67215 1019868
rect 67230 1019858 67254 1019868
rect 67230 1019834 67264 1019858
rect 67275 1019834 67347 1019868
rect 67230 1019824 67347 1019834
rect 67002 1019800 67347 1019824
rect 67015 1019756 67215 1019800
rect 67230 1019790 67254 1019800
rect 67230 1019766 67264 1019790
rect 67275 1019766 67347 1019800
rect 67230 1019756 67347 1019766
rect 67002 1019732 67347 1019756
rect 67015 1019688 67215 1019732
rect 67230 1019722 67254 1019732
rect 67230 1019698 67264 1019722
rect 67275 1019698 67347 1019732
rect 67230 1019688 67347 1019698
rect 67002 1019664 67347 1019688
rect 67015 1019620 67215 1019664
rect 67230 1019654 67254 1019664
rect 67230 1019630 67264 1019654
rect 67275 1019630 67347 1019664
rect 67230 1019620 67347 1019630
rect 67002 1019596 67347 1019620
rect 67015 1019552 67215 1019596
rect 67230 1019586 67254 1019596
rect 67230 1019562 67264 1019586
rect 67275 1019562 67347 1019596
rect 67230 1019552 67347 1019562
rect 67002 1019528 67347 1019552
rect 67015 1019484 67215 1019528
rect 67230 1019518 67254 1019528
rect 67230 1019494 67264 1019518
rect 67275 1019494 67347 1019528
rect 67230 1019484 67347 1019494
rect 67002 1019460 67347 1019484
rect 67015 1019416 67215 1019460
rect 67230 1019450 67254 1019460
rect 67230 1019426 67264 1019450
rect 67275 1019426 67347 1019460
rect 67230 1019416 67347 1019426
rect 67002 1019392 67347 1019416
rect 67015 1019322 67215 1019392
rect 67230 1019368 67254 1019392
rect 67275 1019322 67347 1019392
rect 67577 1019322 67633 1020322
rect 67649 1019322 67705 1020322
rect 68007 1020300 68207 1020322
rect 68222 1020310 68256 1020334
rect 69010 1020322 69044 1020334
rect 68267 1020310 68339 1020322
rect 68222 1020300 68339 1020310
rect 67994 1020276 68339 1020300
rect 68007 1020232 68207 1020276
rect 68222 1020266 68246 1020276
rect 68222 1020242 68256 1020266
rect 68267 1020242 68339 1020276
rect 68222 1020232 68339 1020242
rect 67994 1020208 68339 1020232
rect 68007 1020164 68207 1020208
rect 68222 1020198 68246 1020208
rect 68222 1020174 68256 1020198
rect 68267 1020174 68339 1020208
rect 68222 1020164 68339 1020174
rect 67994 1020140 68339 1020164
rect 68007 1020096 68207 1020140
rect 68222 1020130 68246 1020140
rect 68222 1020106 68256 1020130
rect 68267 1020106 68339 1020140
rect 68222 1020096 68339 1020106
rect 67994 1020072 68339 1020096
rect 68007 1020028 68207 1020072
rect 68222 1020062 68246 1020072
rect 68222 1020038 68256 1020062
rect 68267 1020038 68339 1020072
rect 68222 1020028 68339 1020038
rect 67994 1020004 68339 1020028
rect 68007 1019960 68207 1020004
rect 68222 1019994 68246 1020004
rect 68222 1019970 68256 1019994
rect 68267 1019970 68339 1020004
rect 68222 1019960 68339 1019970
rect 67994 1019936 68339 1019960
rect 68007 1019892 68207 1019936
rect 68222 1019926 68246 1019936
rect 68222 1019902 68256 1019926
rect 68267 1019902 68339 1019936
rect 68222 1019892 68339 1019902
rect 67994 1019868 68339 1019892
rect 68007 1019824 68207 1019868
rect 68222 1019858 68246 1019868
rect 68222 1019834 68256 1019858
rect 68267 1019834 68339 1019868
rect 68222 1019824 68339 1019834
rect 67994 1019800 68339 1019824
rect 68007 1019756 68207 1019800
rect 68222 1019790 68246 1019800
rect 68222 1019766 68256 1019790
rect 68267 1019766 68339 1019800
rect 68222 1019756 68339 1019766
rect 67994 1019732 68339 1019756
rect 68007 1019688 68207 1019732
rect 68222 1019722 68246 1019732
rect 68222 1019698 68256 1019722
rect 68267 1019698 68339 1019732
rect 68222 1019688 68339 1019698
rect 67994 1019664 68339 1019688
rect 68007 1019620 68207 1019664
rect 68222 1019654 68246 1019664
rect 68222 1019630 68256 1019654
rect 68267 1019630 68339 1019664
rect 68222 1019620 68339 1019630
rect 67994 1019596 68339 1019620
rect 68007 1019552 68207 1019596
rect 68222 1019586 68246 1019596
rect 68222 1019562 68256 1019586
rect 68267 1019562 68339 1019596
rect 68222 1019552 68339 1019562
rect 67994 1019528 68339 1019552
rect 68007 1019484 68207 1019528
rect 68222 1019518 68246 1019528
rect 68222 1019494 68256 1019518
rect 68267 1019494 68339 1019528
rect 68222 1019484 68339 1019494
rect 67994 1019460 68339 1019484
rect 68007 1019416 68207 1019460
rect 68222 1019450 68246 1019460
rect 68222 1019426 68256 1019450
rect 68267 1019426 68339 1019460
rect 68222 1019416 68339 1019426
rect 67994 1019392 68339 1019416
rect 68007 1019322 68207 1019392
rect 68222 1019368 68246 1019392
rect 68267 1019322 68339 1019392
rect 68569 1019322 68625 1020322
rect 68641 1019322 68697 1020322
rect 68999 1020300 69199 1020322
rect 69214 1020310 69248 1020334
rect 70002 1020322 70036 1020334
rect 69259 1020310 69331 1020322
rect 69214 1020300 69331 1020310
rect 68986 1020276 69331 1020300
rect 68999 1020232 69199 1020276
rect 69214 1020266 69238 1020276
rect 69214 1020242 69248 1020266
rect 69259 1020242 69331 1020276
rect 69214 1020232 69331 1020242
rect 68986 1020208 69331 1020232
rect 68999 1020164 69199 1020208
rect 69214 1020198 69238 1020208
rect 69214 1020174 69248 1020198
rect 69259 1020174 69331 1020208
rect 69214 1020164 69331 1020174
rect 68986 1020140 69331 1020164
rect 68999 1020096 69199 1020140
rect 69214 1020130 69238 1020140
rect 69214 1020106 69248 1020130
rect 69259 1020106 69331 1020140
rect 69214 1020096 69331 1020106
rect 68986 1020072 69331 1020096
rect 68999 1020028 69199 1020072
rect 69214 1020062 69238 1020072
rect 69214 1020038 69248 1020062
rect 69259 1020038 69331 1020072
rect 69214 1020028 69331 1020038
rect 68986 1020004 69331 1020028
rect 68999 1019960 69199 1020004
rect 69214 1019994 69238 1020004
rect 69214 1019970 69248 1019994
rect 69259 1019970 69331 1020004
rect 69214 1019960 69331 1019970
rect 68986 1019936 69331 1019960
rect 68999 1019892 69199 1019936
rect 69214 1019926 69238 1019936
rect 69214 1019902 69248 1019926
rect 69259 1019902 69331 1019936
rect 69214 1019892 69331 1019902
rect 68986 1019868 69331 1019892
rect 68999 1019824 69199 1019868
rect 69214 1019858 69238 1019868
rect 69214 1019834 69248 1019858
rect 69259 1019834 69331 1019868
rect 69214 1019824 69331 1019834
rect 68986 1019800 69331 1019824
rect 68999 1019756 69199 1019800
rect 69214 1019790 69238 1019800
rect 69214 1019766 69248 1019790
rect 69259 1019766 69331 1019800
rect 69214 1019756 69331 1019766
rect 68986 1019732 69331 1019756
rect 68999 1019688 69199 1019732
rect 69214 1019722 69238 1019732
rect 69214 1019698 69248 1019722
rect 69259 1019698 69331 1019732
rect 69214 1019688 69331 1019698
rect 68986 1019664 69331 1019688
rect 68999 1019620 69199 1019664
rect 69214 1019654 69238 1019664
rect 69214 1019630 69248 1019654
rect 69259 1019630 69331 1019664
rect 69214 1019620 69331 1019630
rect 68986 1019596 69331 1019620
rect 68999 1019552 69199 1019596
rect 69214 1019586 69238 1019596
rect 69214 1019562 69248 1019586
rect 69259 1019562 69331 1019596
rect 69214 1019552 69331 1019562
rect 68986 1019528 69331 1019552
rect 68999 1019484 69199 1019528
rect 69214 1019518 69238 1019528
rect 69214 1019494 69248 1019518
rect 69259 1019494 69331 1019528
rect 69214 1019484 69331 1019494
rect 68986 1019460 69331 1019484
rect 68999 1019416 69199 1019460
rect 69214 1019450 69238 1019460
rect 69214 1019426 69248 1019450
rect 69259 1019426 69331 1019460
rect 69214 1019416 69331 1019426
rect 68986 1019392 69331 1019416
rect 68999 1019322 69199 1019392
rect 69214 1019368 69238 1019392
rect 69259 1019322 69331 1019392
rect 69561 1019322 69617 1020322
rect 69633 1019322 69689 1020322
rect 69991 1020300 70191 1020322
rect 70206 1020310 70240 1020334
rect 70994 1020322 71028 1020334
rect 70251 1020310 70323 1020322
rect 70206 1020300 70323 1020310
rect 69978 1020276 70323 1020300
rect 69991 1020232 70191 1020276
rect 70206 1020266 70230 1020276
rect 70206 1020242 70240 1020266
rect 70251 1020242 70323 1020276
rect 70206 1020232 70323 1020242
rect 69978 1020208 70323 1020232
rect 69991 1020164 70191 1020208
rect 70206 1020198 70230 1020208
rect 70206 1020174 70240 1020198
rect 70251 1020174 70323 1020208
rect 70206 1020164 70323 1020174
rect 69978 1020140 70323 1020164
rect 69991 1020096 70191 1020140
rect 70206 1020130 70230 1020140
rect 70206 1020106 70240 1020130
rect 70251 1020106 70323 1020140
rect 70206 1020096 70323 1020106
rect 69978 1020072 70323 1020096
rect 69991 1020028 70191 1020072
rect 70206 1020062 70230 1020072
rect 70206 1020038 70240 1020062
rect 70251 1020038 70323 1020072
rect 70206 1020028 70323 1020038
rect 69978 1020004 70323 1020028
rect 69991 1019960 70191 1020004
rect 70206 1019994 70230 1020004
rect 70206 1019970 70240 1019994
rect 70251 1019970 70323 1020004
rect 70206 1019960 70323 1019970
rect 69978 1019936 70323 1019960
rect 69991 1019892 70191 1019936
rect 70206 1019926 70230 1019936
rect 70206 1019902 70240 1019926
rect 70251 1019902 70323 1019936
rect 70206 1019892 70323 1019902
rect 69978 1019868 70323 1019892
rect 69991 1019824 70191 1019868
rect 70206 1019858 70230 1019868
rect 70206 1019834 70240 1019858
rect 70251 1019834 70323 1019868
rect 70206 1019824 70323 1019834
rect 69978 1019800 70323 1019824
rect 69991 1019756 70191 1019800
rect 70206 1019790 70230 1019800
rect 70206 1019766 70240 1019790
rect 70251 1019766 70323 1019800
rect 70206 1019756 70323 1019766
rect 69978 1019732 70323 1019756
rect 69991 1019688 70191 1019732
rect 70206 1019722 70230 1019732
rect 70206 1019698 70240 1019722
rect 70251 1019698 70323 1019732
rect 70206 1019688 70323 1019698
rect 69978 1019664 70323 1019688
rect 69991 1019620 70191 1019664
rect 70206 1019654 70230 1019664
rect 70206 1019630 70240 1019654
rect 70251 1019630 70323 1019664
rect 70206 1019620 70323 1019630
rect 69978 1019596 70323 1019620
rect 69991 1019552 70191 1019596
rect 70206 1019586 70230 1019596
rect 70206 1019562 70240 1019586
rect 70251 1019562 70323 1019596
rect 70206 1019552 70323 1019562
rect 69978 1019528 70323 1019552
rect 69991 1019484 70191 1019528
rect 70206 1019518 70230 1019528
rect 70206 1019494 70240 1019518
rect 70251 1019494 70323 1019528
rect 70206 1019484 70323 1019494
rect 69978 1019460 70323 1019484
rect 69991 1019416 70191 1019460
rect 70206 1019450 70230 1019460
rect 70206 1019426 70240 1019450
rect 70251 1019426 70323 1019460
rect 70206 1019416 70323 1019426
rect 69978 1019392 70323 1019416
rect 69991 1019322 70191 1019392
rect 70206 1019368 70230 1019392
rect 70251 1019322 70323 1019392
rect 70553 1019322 70609 1020322
rect 70625 1019322 70681 1020322
rect 70983 1020300 71183 1020322
rect 71198 1020310 71232 1020334
rect 71986 1020322 72020 1020334
rect 71243 1020310 71315 1020322
rect 71198 1020300 71315 1020310
rect 70970 1020276 71315 1020300
rect 70983 1020232 71183 1020276
rect 71198 1020266 71222 1020276
rect 71198 1020242 71232 1020266
rect 71243 1020242 71315 1020276
rect 71198 1020232 71315 1020242
rect 70970 1020208 71315 1020232
rect 70983 1020164 71183 1020208
rect 71198 1020198 71222 1020208
rect 71198 1020174 71232 1020198
rect 71243 1020174 71315 1020208
rect 71198 1020164 71315 1020174
rect 70970 1020140 71315 1020164
rect 70983 1020096 71183 1020140
rect 71198 1020130 71222 1020140
rect 71198 1020106 71232 1020130
rect 71243 1020106 71315 1020140
rect 71198 1020096 71315 1020106
rect 70970 1020072 71315 1020096
rect 70983 1020028 71183 1020072
rect 71198 1020062 71222 1020072
rect 71198 1020038 71232 1020062
rect 71243 1020038 71315 1020072
rect 71198 1020028 71315 1020038
rect 70970 1020004 71315 1020028
rect 70983 1019960 71183 1020004
rect 71198 1019994 71222 1020004
rect 71198 1019970 71232 1019994
rect 71243 1019970 71315 1020004
rect 71198 1019960 71315 1019970
rect 70970 1019936 71315 1019960
rect 70983 1019892 71183 1019936
rect 71198 1019926 71222 1019936
rect 71198 1019902 71232 1019926
rect 71243 1019902 71315 1019936
rect 71198 1019892 71315 1019902
rect 70970 1019868 71315 1019892
rect 70983 1019824 71183 1019868
rect 71198 1019858 71222 1019868
rect 71198 1019834 71232 1019858
rect 71243 1019834 71315 1019868
rect 71198 1019824 71315 1019834
rect 70970 1019800 71315 1019824
rect 70983 1019756 71183 1019800
rect 71198 1019790 71222 1019800
rect 71198 1019766 71232 1019790
rect 71243 1019766 71315 1019800
rect 71198 1019756 71315 1019766
rect 70970 1019732 71315 1019756
rect 70983 1019688 71183 1019732
rect 71198 1019722 71222 1019732
rect 71198 1019698 71232 1019722
rect 71243 1019698 71315 1019732
rect 71198 1019688 71315 1019698
rect 70970 1019664 71315 1019688
rect 70983 1019620 71183 1019664
rect 71198 1019654 71222 1019664
rect 71198 1019630 71232 1019654
rect 71243 1019630 71315 1019664
rect 71198 1019620 71315 1019630
rect 70970 1019596 71315 1019620
rect 70983 1019552 71183 1019596
rect 71198 1019586 71222 1019596
rect 71198 1019562 71232 1019586
rect 71243 1019562 71315 1019596
rect 71198 1019552 71315 1019562
rect 70970 1019528 71315 1019552
rect 70983 1019484 71183 1019528
rect 71198 1019518 71222 1019528
rect 71198 1019494 71232 1019518
rect 71243 1019494 71315 1019528
rect 71198 1019484 71315 1019494
rect 70970 1019460 71315 1019484
rect 70983 1019416 71183 1019460
rect 71198 1019450 71222 1019460
rect 71198 1019426 71232 1019450
rect 71243 1019426 71315 1019460
rect 71198 1019416 71315 1019426
rect 70970 1019392 71315 1019416
rect 70983 1019322 71183 1019392
rect 71198 1019368 71222 1019392
rect 71243 1019322 71315 1019392
rect 71545 1019322 71601 1020322
rect 71617 1019322 71673 1020322
rect 71975 1020300 72175 1020322
rect 72190 1020310 72224 1020334
rect 72978 1020322 73012 1020334
rect 72235 1020310 72307 1020322
rect 72190 1020300 72307 1020310
rect 71962 1020276 72307 1020300
rect 71975 1020232 72175 1020276
rect 72190 1020266 72214 1020276
rect 72190 1020242 72224 1020266
rect 72235 1020242 72307 1020276
rect 72190 1020232 72307 1020242
rect 71962 1020208 72307 1020232
rect 71975 1020164 72175 1020208
rect 72190 1020198 72214 1020208
rect 72190 1020174 72224 1020198
rect 72235 1020174 72307 1020208
rect 72190 1020164 72307 1020174
rect 71962 1020140 72307 1020164
rect 71975 1020096 72175 1020140
rect 72190 1020130 72214 1020140
rect 72190 1020106 72224 1020130
rect 72235 1020106 72307 1020140
rect 72190 1020096 72307 1020106
rect 71962 1020072 72307 1020096
rect 71975 1020028 72175 1020072
rect 72190 1020062 72214 1020072
rect 72190 1020038 72224 1020062
rect 72235 1020038 72307 1020072
rect 72190 1020028 72307 1020038
rect 71962 1020004 72307 1020028
rect 71975 1019960 72175 1020004
rect 72190 1019994 72214 1020004
rect 72190 1019970 72224 1019994
rect 72235 1019970 72307 1020004
rect 72190 1019960 72307 1019970
rect 71962 1019936 72307 1019960
rect 71975 1019892 72175 1019936
rect 72190 1019926 72214 1019936
rect 72190 1019902 72224 1019926
rect 72235 1019902 72307 1019936
rect 72190 1019892 72307 1019902
rect 71962 1019868 72307 1019892
rect 71975 1019824 72175 1019868
rect 72190 1019858 72214 1019868
rect 72190 1019834 72224 1019858
rect 72235 1019834 72307 1019868
rect 72190 1019824 72307 1019834
rect 71962 1019800 72307 1019824
rect 71975 1019756 72175 1019800
rect 72190 1019790 72214 1019800
rect 72190 1019766 72224 1019790
rect 72235 1019766 72307 1019800
rect 72190 1019756 72307 1019766
rect 71962 1019732 72307 1019756
rect 71975 1019688 72175 1019732
rect 72190 1019722 72214 1019732
rect 72190 1019698 72224 1019722
rect 72235 1019698 72307 1019732
rect 72190 1019688 72307 1019698
rect 71962 1019664 72307 1019688
rect 71975 1019620 72175 1019664
rect 72190 1019654 72214 1019664
rect 72190 1019630 72224 1019654
rect 72235 1019630 72307 1019664
rect 72190 1019620 72307 1019630
rect 71962 1019596 72307 1019620
rect 71975 1019552 72175 1019596
rect 72190 1019586 72214 1019596
rect 72190 1019562 72224 1019586
rect 72235 1019562 72307 1019596
rect 72190 1019552 72307 1019562
rect 71962 1019528 72307 1019552
rect 71975 1019484 72175 1019528
rect 72190 1019518 72214 1019528
rect 72190 1019494 72224 1019518
rect 72235 1019494 72307 1019528
rect 72190 1019484 72307 1019494
rect 71962 1019460 72307 1019484
rect 71975 1019416 72175 1019460
rect 72190 1019450 72214 1019460
rect 72190 1019426 72224 1019450
rect 72235 1019426 72307 1019460
rect 72190 1019416 72307 1019426
rect 71962 1019392 72307 1019416
rect 71975 1019322 72175 1019392
rect 72190 1019368 72214 1019392
rect 72235 1019322 72307 1019392
rect 72537 1019322 72593 1020322
rect 72609 1019322 72665 1020322
rect 72967 1020300 73167 1020322
rect 73182 1020310 73216 1020334
rect 73970 1020322 74004 1020334
rect 73227 1020310 73299 1020322
rect 73182 1020300 73299 1020310
rect 72954 1020276 73299 1020300
rect 72967 1020232 73167 1020276
rect 73182 1020266 73206 1020276
rect 73182 1020242 73216 1020266
rect 73227 1020242 73299 1020276
rect 73182 1020232 73299 1020242
rect 72954 1020208 73299 1020232
rect 72967 1020164 73167 1020208
rect 73182 1020198 73206 1020208
rect 73182 1020174 73216 1020198
rect 73227 1020174 73299 1020208
rect 73182 1020164 73299 1020174
rect 72954 1020140 73299 1020164
rect 72967 1020096 73167 1020140
rect 73182 1020130 73206 1020140
rect 73182 1020106 73216 1020130
rect 73227 1020106 73299 1020140
rect 73182 1020096 73299 1020106
rect 72954 1020072 73299 1020096
rect 72967 1020028 73167 1020072
rect 73182 1020062 73206 1020072
rect 73182 1020038 73216 1020062
rect 73227 1020038 73299 1020072
rect 73182 1020028 73299 1020038
rect 72954 1020004 73299 1020028
rect 72967 1019960 73167 1020004
rect 73182 1019994 73206 1020004
rect 73182 1019970 73216 1019994
rect 73227 1019970 73299 1020004
rect 73182 1019960 73299 1019970
rect 72954 1019936 73299 1019960
rect 72967 1019892 73167 1019936
rect 73182 1019926 73206 1019936
rect 73182 1019902 73216 1019926
rect 73227 1019902 73299 1019936
rect 73182 1019892 73299 1019902
rect 72954 1019868 73299 1019892
rect 72967 1019824 73167 1019868
rect 73182 1019858 73206 1019868
rect 73182 1019834 73216 1019858
rect 73227 1019834 73299 1019868
rect 73182 1019824 73299 1019834
rect 72954 1019800 73299 1019824
rect 72967 1019756 73167 1019800
rect 73182 1019790 73206 1019800
rect 73182 1019766 73216 1019790
rect 73227 1019766 73299 1019800
rect 73182 1019756 73299 1019766
rect 72954 1019732 73299 1019756
rect 72967 1019688 73167 1019732
rect 73182 1019722 73206 1019732
rect 73182 1019698 73216 1019722
rect 73227 1019698 73299 1019732
rect 73182 1019688 73299 1019698
rect 72954 1019664 73299 1019688
rect 72967 1019620 73167 1019664
rect 73182 1019654 73206 1019664
rect 73182 1019630 73216 1019654
rect 73227 1019630 73299 1019664
rect 73182 1019620 73299 1019630
rect 72954 1019596 73299 1019620
rect 72967 1019552 73167 1019596
rect 73182 1019586 73206 1019596
rect 73182 1019562 73216 1019586
rect 73227 1019562 73299 1019596
rect 73182 1019552 73299 1019562
rect 72954 1019528 73299 1019552
rect 72967 1019484 73167 1019528
rect 73182 1019518 73206 1019528
rect 73182 1019494 73216 1019518
rect 73227 1019494 73299 1019528
rect 73182 1019484 73299 1019494
rect 72954 1019460 73299 1019484
rect 72967 1019416 73167 1019460
rect 73182 1019450 73206 1019460
rect 73182 1019426 73216 1019450
rect 73227 1019426 73299 1019460
rect 73182 1019416 73299 1019426
rect 72954 1019392 73299 1019416
rect 72967 1019322 73167 1019392
rect 73182 1019368 73206 1019392
rect 73227 1019322 73299 1019392
rect 73529 1019322 73585 1020322
rect 73601 1019322 73657 1020322
rect 73959 1020300 74159 1020322
rect 74174 1020310 74208 1020334
rect 74962 1020322 74996 1020334
rect 74219 1020310 74291 1020322
rect 74174 1020300 74291 1020310
rect 73946 1020276 74291 1020300
rect 73959 1020232 74159 1020276
rect 74174 1020266 74198 1020276
rect 74174 1020242 74208 1020266
rect 74219 1020242 74291 1020276
rect 74174 1020232 74291 1020242
rect 73946 1020208 74291 1020232
rect 73959 1020164 74159 1020208
rect 74174 1020198 74198 1020208
rect 74174 1020174 74208 1020198
rect 74219 1020174 74291 1020208
rect 74174 1020164 74291 1020174
rect 73946 1020140 74291 1020164
rect 73959 1020096 74159 1020140
rect 74174 1020130 74198 1020140
rect 74174 1020106 74208 1020130
rect 74219 1020106 74291 1020140
rect 74174 1020096 74291 1020106
rect 73946 1020072 74291 1020096
rect 73959 1020028 74159 1020072
rect 74174 1020062 74198 1020072
rect 74174 1020038 74208 1020062
rect 74219 1020038 74291 1020072
rect 74174 1020028 74291 1020038
rect 73946 1020004 74291 1020028
rect 73959 1019960 74159 1020004
rect 74174 1019994 74198 1020004
rect 74174 1019970 74208 1019994
rect 74219 1019970 74291 1020004
rect 74174 1019960 74291 1019970
rect 73946 1019936 74291 1019960
rect 73959 1019892 74159 1019936
rect 74174 1019926 74198 1019936
rect 74174 1019902 74208 1019926
rect 74219 1019902 74291 1019936
rect 74174 1019892 74291 1019902
rect 73946 1019868 74291 1019892
rect 73959 1019824 74159 1019868
rect 74174 1019858 74198 1019868
rect 74174 1019834 74208 1019858
rect 74219 1019834 74291 1019868
rect 74174 1019824 74291 1019834
rect 73946 1019800 74291 1019824
rect 73959 1019756 74159 1019800
rect 74174 1019790 74198 1019800
rect 74174 1019766 74208 1019790
rect 74219 1019766 74291 1019800
rect 74174 1019756 74291 1019766
rect 73946 1019732 74291 1019756
rect 73959 1019688 74159 1019732
rect 74174 1019722 74198 1019732
rect 74174 1019698 74208 1019722
rect 74219 1019698 74291 1019732
rect 74174 1019688 74291 1019698
rect 73946 1019664 74291 1019688
rect 73959 1019620 74159 1019664
rect 74174 1019654 74198 1019664
rect 74174 1019630 74208 1019654
rect 74219 1019630 74291 1019664
rect 74174 1019620 74291 1019630
rect 73946 1019596 74291 1019620
rect 73959 1019552 74159 1019596
rect 74174 1019586 74198 1019596
rect 74174 1019562 74208 1019586
rect 74219 1019562 74291 1019596
rect 74174 1019552 74291 1019562
rect 73946 1019528 74291 1019552
rect 73959 1019484 74159 1019528
rect 74174 1019518 74198 1019528
rect 74174 1019494 74208 1019518
rect 74219 1019494 74291 1019528
rect 74174 1019484 74291 1019494
rect 73946 1019460 74291 1019484
rect 73959 1019416 74159 1019460
rect 74174 1019450 74198 1019460
rect 74174 1019426 74208 1019450
rect 74219 1019426 74291 1019460
rect 74174 1019416 74291 1019426
rect 73946 1019392 74291 1019416
rect 73959 1019322 74159 1019392
rect 74174 1019368 74198 1019392
rect 74219 1019322 74291 1019392
rect 74521 1019322 74577 1020322
rect 74593 1019322 74649 1020322
rect 74951 1020300 75151 1020322
rect 75166 1020310 75200 1020334
rect 75211 1020310 75283 1020322
rect 75166 1020300 75283 1020310
rect 74938 1020276 75283 1020300
rect 74951 1020232 75151 1020276
rect 75166 1020266 75190 1020276
rect 75166 1020242 75200 1020266
rect 75211 1020242 75283 1020276
rect 75166 1020232 75283 1020242
rect 74938 1020208 75283 1020232
rect 74951 1020164 75151 1020208
rect 75166 1020198 75190 1020208
rect 75166 1020174 75200 1020198
rect 75211 1020174 75283 1020208
rect 75166 1020164 75283 1020174
rect 74938 1020140 75283 1020164
rect 74951 1020096 75151 1020140
rect 75166 1020130 75190 1020140
rect 75166 1020106 75200 1020130
rect 75211 1020106 75283 1020140
rect 75166 1020096 75283 1020106
rect 74938 1020072 75283 1020096
rect 74951 1020028 75151 1020072
rect 75166 1020062 75190 1020072
rect 75166 1020038 75200 1020062
rect 75211 1020038 75283 1020072
rect 75166 1020028 75283 1020038
rect 74938 1020004 75283 1020028
rect 74951 1019960 75151 1020004
rect 75166 1019994 75190 1020004
rect 75166 1019970 75200 1019994
rect 75211 1019970 75283 1020004
rect 75166 1019960 75283 1019970
rect 74938 1019936 75283 1019960
rect 74951 1019892 75151 1019936
rect 75166 1019926 75190 1019936
rect 75166 1019902 75200 1019926
rect 75211 1019902 75283 1019936
rect 75166 1019892 75283 1019902
rect 74938 1019868 75283 1019892
rect 74951 1019824 75151 1019868
rect 75166 1019858 75190 1019868
rect 75166 1019834 75200 1019858
rect 75211 1019834 75283 1019868
rect 75166 1019824 75283 1019834
rect 74938 1019800 75283 1019824
rect 74951 1019756 75151 1019800
rect 75166 1019790 75190 1019800
rect 75166 1019766 75200 1019790
rect 75211 1019766 75283 1019800
rect 75166 1019756 75283 1019766
rect 74938 1019732 75283 1019756
rect 74951 1019688 75151 1019732
rect 75166 1019722 75190 1019732
rect 75166 1019698 75200 1019722
rect 75211 1019698 75283 1019732
rect 75166 1019688 75283 1019698
rect 74938 1019664 75283 1019688
rect 74951 1019620 75151 1019664
rect 75166 1019654 75190 1019664
rect 75166 1019630 75200 1019654
rect 75211 1019630 75283 1019664
rect 75166 1019620 75283 1019630
rect 74938 1019596 75283 1019620
rect 74951 1019552 75151 1019596
rect 75166 1019586 75190 1019596
rect 75166 1019562 75200 1019586
rect 75211 1019562 75283 1019596
rect 75166 1019552 75283 1019562
rect 74938 1019528 75283 1019552
rect 74951 1019484 75151 1019528
rect 75166 1019518 75190 1019528
rect 75166 1019494 75200 1019518
rect 75211 1019494 75283 1019528
rect 75166 1019484 75283 1019494
rect 74938 1019460 75283 1019484
rect 74951 1019416 75151 1019460
rect 75166 1019450 75190 1019460
rect 75166 1019426 75200 1019450
rect 75211 1019426 75283 1019460
rect 75166 1019416 75283 1019426
rect 74938 1019392 75283 1019416
rect 74951 1019322 75151 1019392
rect 75166 1019368 75190 1019392
rect 75211 1019322 75283 1019392
rect 75472 1019322 75544 1020322
rect 75610 1019322 75627 1020322
rect 75797 1019322 75830 1020322
rect 109561 1018210 109668 1022756
rect 110356 1020922 110406 1021922
rect 110617 1020922 110673 1021922
rect 110689 1020922 110745 1021922
rect 111107 1020922 111247 1021922
rect 122521 1020922 122577 1021922
rect 122593 1020922 122649 1021922
rect 123011 1020922 123151 1021922
rect 123473 1020922 123544 1021922
rect 123610 1020922 123627 1021922
rect 123797 1020922 123830 1021922
rect 123953 1021730 124025 1021760
rect 123953 1021692 123987 1021722
rect 110356 1019322 110406 1020322
rect 110617 1019322 110673 1020322
rect 110689 1019322 110745 1020322
rect 111107 1019322 111247 1020322
rect 122521 1019322 122577 1020322
rect 122593 1019322 122649 1020322
rect 123011 1019322 123151 1020322
rect 123473 1019322 123544 1020322
rect 123610 1019322 123627 1020322
rect 123797 1019322 123830 1020322
rect 161561 1018210 161668 1022756
rect 162356 1020922 162406 1021922
rect 162617 1020922 162673 1021922
rect 162689 1020922 162745 1021922
rect 163047 1021842 163247 1021922
rect 163262 1021852 163296 1021876
rect 163307 1021852 163379 1021922
rect 163262 1021842 163379 1021852
rect 163034 1021818 163379 1021842
rect 163047 1021774 163247 1021818
rect 163262 1021808 163286 1021818
rect 163262 1021784 163296 1021808
rect 163307 1021784 163379 1021818
rect 163262 1021774 163379 1021784
rect 163034 1021750 163379 1021774
rect 163047 1021706 163247 1021750
rect 163262 1021740 163286 1021750
rect 163262 1021716 163296 1021740
rect 163307 1021716 163379 1021750
rect 163262 1021706 163379 1021716
rect 163034 1021682 163379 1021706
rect 163047 1021638 163247 1021682
rect 163262 1021672 163286 1021682
rect 163262 1021648 163296 1021672
rect 163307 1021648 163379 1021682
rect 163262 1021638 163379 1021648
rect 163034 1021614 163379 1021638
rect 163047 1021570 163247 1021614
rect 163262 1021604 163286 1021614
rect 163262 1021580 163296 1021604
rect 163307 1021580 163379 1021614
rect 163262 1021570 163379 1021580
rect 163034 1021546 163379 1021570
rect 163047 1021502 163247 1021546
rect 163262 1021536 163286 1021546
rect 163262 1021512 163296 1021536
rect 163307 1021512 163379 1021546
rect 163262 1021502 163379 1021512
rect 163034 1021478 163379 1021502
rect 163047 1021434 163247 1021478
rect 163262 1021468 163286 1021478
rect 163262 1021444 163296 1021468
rect 163307 1021444 163379 1021478
rect 163262 1021434 163379 1021444
rect 163034 1021410 163379 1021434
rect 163047 1021366 163247 1021410
rect 163262 1021400 163286 1021410
rect 163262 1021376 163296 1021400
rect 163307 1021376 163379 1021410
rect 163262 1021366 163379 1021376
rect 163034 1021342 163379 1021366
rect 163047 1021298 163247 1021342
rect 163262 1021332 163286 1021342
rect 163262 1021308 163296 1021332
rect 163307 1021308 163379 1021342
rect 163262 1021298 163379 1021308
rect 163034 1021274 163379 1021298
rect 163047 1021230 163247 1021274
rect 163262 1021264 163286 1021274
rect 163262 1021240 163296 1021264
rect 163307 1021240 163379 1021274
rect 163262 1021230 163379 1021240
rect 163034 1021206 163379 1021230
rect 163047 1021162 163247 1021206
rect 163262 1021196 163286 1021206
rect 163262 1021172 163296 1021196
rect 163307 1021172 163379 1021206
rect 163262 1021162 163379 1021172
rect 163034 1021138 163379 1021162
rect 163047 1021094 163247 1021138
rect 163262 1021128 163286 1021138
rect 163262 1021104 163296 1021128
rect 163307 1021104 163379 1021138
rect 163262 1021094 163379 1021104
rect 163034 1021070 163379 1021094
rect 163047 1021026 163247 1021070
rect 163262 1021060 163286 1021070
rect 163262 1021036 163296 1021060
rect 163307 1021036 163379 1021070
rect 163262 1021026 163379 1021036
rect 163034 1021002 163379 1021026
rect 163047 1020958 163247 1021002
rect 163262 1020992 163286 1021002
rect 163262 1020968 163296 1020992
rect 163307 1020968 163379 1021002
rect 163262 1020958 163379 1020968
rect 163034 1020934 163379 1020958
rect 163047 1020922 163247 1020934
rect 163058 1020910 163082 1020922
rect 163262 1020910 163286 1020934
rect 163307 1020922 163379 1020934
rect 163609 1020922 163665 1021922
rect 163681 1020922 163737 1021922
rect 164039 1021842 164239 1021922
rect 164254 1021852 164288 1021876
rect 164299 1021852 164371 1021922
rect 164254 1021842 164371 1021852
rect 164026 1021818 164371 1021842
rect 164039 1021774 164239 1021818
rect 164254 1021808 164278 1021818
rect 164254 1021784 164288 1021808
rect 164299 1021784 164371 1021818
rect 164254 1021774 164371 1021784
rect 164026 1021750 164371 1021774
rect 164039 1021706 164239 1021750
rect 164254 1021740 164278 1021750
rect 164254 1021716 164288 1021740
rect 164299 1021716 164371 1021750
rect 164254 1021706 164371 1021716
rect 164026 1021682 164371 1021706
rect 164039 1021638 164239 1021682
rect 164254 1021672 164278 1021682
rect 164254 1021648 164288 1021672
rect 164299 1021648 164371 1021682
rect 164254 1021638 164371 1021648
rect 164026 1021614 164371 1021638
rect 164039 1021570 164239 1021614
rect 164254 1021604 164278 1021614
rect 164254 1021580 164288 1021604
rect 164299 1021580 164371 1021614
rect 164254 1021570 164371 1021580
rect 164026 1021546 164371 1021570
rect 164039 1021502 164239 1021546
rect 164254 1021536 164278 1021546
rect 164254 1021512 164288 1021536
rect 164299 1021512 164371 1021546
rect 164254 1021502 164371 1021512
rect 164026 1021478 164371 1021502
rect 164039 1021434 164239 1021478
rect 164254 1021468 164278 1021478
rect 164254 1021444 164288 1021468
rect 164299 1021444 164371 1021478
rect 164254 1021434 164371 1021444
rect 164026 1021410 164371 1021434
rect 164039 1021366 164239 1021410
rect 164254 1021400 164278 1021410
rect 164254 1021376 164288 1021400
rect 164299 1021376 164371 1021410
rect 164254 1021366 164371 1021376
rect 164026 1021342 164371 1021366
rect 164039 1021298 164239 1021342
rect 164254 1021332 164278 1021342
rect 164254 1021308 164288 1021332
rect 164299 1021308 164371 1021342
rect 164254 1021298 164371 1021308
rect 164026 1021274 164371 1021298
rect 164039 1021230 164239 1021274
rect 164254 1021264 164278 1021274
rect 164254 1021240 164288 1021264
rect 164299 1021240 164371 1021274
rect 164254 1021230 164371 1021240
rect 164026 1021206 164371 1021230
rect 164039 1021162 164239 1021206
rect 164254 1021196 164278 1021206
rect 164254 1021172 164288 1021196
rect 164299 1021172 164371 1021206
rect 164254 1021162 164371 1021172
rect 164026 1021138 164371 1021162
rect 164039 1021094 164239 1021138
rect 164254 1021128 164278 1021138
rect 164254 1021104 164288 1021128
rect 164299 1021104 164371 1021138
rect 164254 1021094 164371 1021104
rect 164026 1021070 164371 1021094
rect 164039 1021026 164239 1021070
rect 164254 1021060 164278 1021070
rect 164254 1021036 164288 1021060
rect 164299 1021036 164371 1021070
rect 164254 1021026 164371 1021036
rect 164026 1021002 164371 1021026
rect 164039 1020958 164239 1021002
rect 164254 1020992 164278 1021002
rect 164254 1020968 164288 1020992
rect 164299 1020968 164371 1021002
rect 164254 1020958 164371 1020968
rect 164026 1020934 164371 1020958
rect 164039 1020922 164239 1020934
rect 164050 1020910 164074 1020922
rect 164254 1020910 164278 1020934
rect 164299 1020922 164371 1020934
rect 164601 1020922 164657 1021922
rect 164673 1020922 164729 1021922
rect 165031 1021842 165231 1021922
rect 165246 1021852 165280 1021876
rect 165291 1021852 165363 1021922
rect 165246 1021842 165363 1021852
rect 165018 1021818 165363 1021842
rect 165031 1021774 165231 1021818
rect 165246 1021808 165270 1021818
rect 165246 1021784 165280 1021808
rect 165291 1021784 165363 1021818
rect 165246 1021774 165363 1021784
rect 165018 1021750 165363 1021774
rect 165031 1021706 165231 1021750
rect 165246 1021740 165270 1021750
rect 165246 1021716 165280 1021740
rect 165291 1021716 165363 1021750
rect 165246 1021706 165363 1021716
rect 165018 1021682 165363 1021706
rect 165031 1021638 165231 1021682
rect 165246 1021672 165270 1021682
rect 165246 1021648 165280 1021672
rect 165291 1021648 165363 1021682
rect 165246 1021638 165363 1021648
rect 165018 1021614 165363 1021638
rect 165031 1021570 165231 1021614
rect 165246 1021604 165270 1021614
rect 165246 1021580 165280 1021604
rect 165291 1021580 165363 1021614
rect 165246 1021570 165363 1021580
rect 165018 1021546 165363 1021570
rect 165031 1021502 165231 1021546
rect 165246 1021536 165270 1021546
rect 165246 1021512 165280 1021536
rect 165291 1021512 165363 1021546
rect 165246 1021502 165363 1021512
rect 165018 1021478 165363 1021502
rect 165031 1021434 165231 1021478
rect 165246 1021468 165270 1021478
rect 165246 1021444 165280 1021468
rect 165291 1021444 165363 1021478
rect 165246 1021434 165363 1021444
rect 165018 1021410 165363 1021434
rect 165031 1021366 165231 1021410
rect 165246 1021400 165270 1021410
rect 165246 1021376 165280 1021400
rect 165291 1021376 165363 1021410
rect 165246 1021366 165363 1021376
rect 165018 1021342 165363 1021366
rect 165031 1021298 165231 1021342
rect 165246 1021332 165270 1021342
rect 165246 1021308 165280 1021332
rect 165291 1021308 165363 1021342
rect 165246 1021298 165363 1021308
rect 165018 1021274 165363 1021298
rect 165031 1021230 165231 1021274
rect 165246 1021264 165270 1021274
rect 165246 1021240 165280 1021264
rect 165291 1021240 165363 1021274
rect 165246 1021230 165363 1021240
rect 165018 1021206 165363 1021230
rect 165031 1021162 165231 1021206
rect 165246 1021196 165270 1021206
rect 165246 1021172 165280 1021196
rect 165291 1021172 165363 1021206
rect 165246 1021162 165363 1021172
rect 165018 1021138 165363 1021162
rect 165031 1021094 165231 1021138
rect 165246 1021128 165270 1021138
rect 165246 1021104 165280 1021128
rect 165291 1021104 165363 1021138
rect 165246 1021094 165363 1021104
rect 165018 1021070 165363 1021094
rect 165031 1021026 165231 1021070
rect 165246 1021060 165270 1021070
rect 165246 1021036 165280 1021060
rect 165291 1021036 165363 1021070
rect 165246 1021026 165363 1021036
rect 165018 1021002 165363 1021026
rect 165031 1020958 165231 1021002
rect 165246 1020992 165270 1021002
rect 165246 1020968 165280 1020992
rect 165291 1020968 165363 1021002
rect 165246 1020958 165363 1020968
rect 165018 1020934 165363 1020958
rect 165031 1020922 165231 1020934
rect 165042 1020910 165066 1020922
rect 165246 1020910 165270 1020934
rect 165291 1020922 165363 1020934
rect 165593 1020922 165649 1021922
rect 165665 1020922 165721 1021922
rect 166023 1021842 166223 1021922
rect 166238 1021852 166272 1021876
rect 166283 1021852 166355 1021922
rect 166238 1021842 166355 1021852
rect 166010 1021818 166355 1021842
rect 166023 1021774 166223 1021818
rect 166238 1021808 166262 1021818
rect 166238 1021784 166272 1021808
rect 166283 1021784 166355 1021818
rect 166238 1021774 166355 1021784
rect 166010 1021750 166355 1021774
rect 166023 1021706 166223 1021750
rect 166238 1021740 166262 1021750
rect 166238 1021716 166272 1021740
rect 166283 1021716 166355 1021750
rect 166238 1021706 166355 1021716
rect 166010 1021682 166355 1021706
rect 166023 1021638 166223 1021682
rect 166238 1021672 166262 1021682
rect 166238 1021648 166272 1021672
rect 166283 1021648 166355 1021682
rect 166238 1021638 166355 1021648
rect 166010 1021614 166355 1021638
rect 166023 1021570 166223 1021614
rect 166238 1021604 166262 1021614
rect 166238 1021580 166272 1021604
rect 166283 1021580 166355 1021614
rect 166238 1021570 166355 1021580
rect 166010 1021546 166355 1021570
rect 166023 1021502 166223 1021546
rect 166238 1021536 166262 1021546
rect 166238 1021512 166272 1021536
rect 166283 1021512 166355 1021546
rect 166238 1021502 166355 1021512
rect 166010 1021478 166355 1021502
rect 166023 1021434 166223 1021478
rect 166238 1021468 166262 1021478
rect 166238 1021444 166272 1021468
rect 166283 1021444 166355 1021478
rect 166238 1021434 166355 1021444
rect 166010 1021410 166355 1021434
rect 166023 1021366 166223 1021410
rect 166238 1021400 166262 1021410
rect 166238 1021376 166272 1021400
rect 166283 1021376 166355 1021410
rect 166238 1021366 166355 1021376
rect 166010 1021342 166355 1021366
rect 166023 1021298 166223 1021342
rect 166238 1021332 166262 1021342
rect 166238 1021308 166272 1021332
rect 166283 1021308 166355 1021342
rect 166238 1021298 166355 1021308
rect 166010 1021274 166355 1021298
rect 166023 1021230 166223 1021274
rect 166238 1021264 166262 1021274
rect 166238 1021240 166272 1021264
rect 166283 1021240 166355 1021274
rect 166238 1021230 166355 1021240
rect 166010 1021206 166355 1021230
rect 166023 1021162 166223 1021206
rect 166238 1021196 166262 1021206
rect 166238 1021172 166272 1021196
rect 166283 1021172 166355 1021206
rect 166238 1021162 166355 1021172
rect 166010 1021138 166355 1021162
rect 166023 1021094 166223 1021138
rect 166238 1021128 166262 1021138
rect 166238 1021104 166272 1021128
rect 166283 1021104 166355 1021138
rect 166238 1021094 166355 1021104
rect 166010 1021070 166355 1021094
rect 166023 1021026 166223 1021070
rect 166238 1021060 166262 1021070
rect 166238 1021036 166272 1021060
rect 166283 1021036 166355 1021070
rect 166238 1021026 166355 1021036
rect 166010 1021002 166355 1021026
rect 166023 1020958 166223 1021002
rect 166238 1020992 166262 1021002
rect 166238 1020968 166272 1020992
rect 166283 1020968 166355 1021002
rect 166238 1020958 166355 1020968
rect 166010 1020934 166355 1020958
rect 166023 1020922 166223 1020934
rect 166034 1020910 166058 1020922
rect 166238 1020910 166262 1020934
rect 166283 1020922 166355 1020934
rect 166585 1020922 166641 1021922
rect 166657 1020922 166713 1021922
rect 167015 1021842 167215 1021922
rect 167230 1021852 167264 1021876
rect 167275 1021852 167347 1021922
rect 167230 1021842 167347 1021852
rect 167002 1021818 167347 1021842
rect 167015 1021774 167215 1021818
rect 167230 1021808 167254 1021818
rect 167230 1021784 167264 1021808
rect 167275 1021784 167347 1021818
rect 167230 1021774 167347 1021784
rect 167002 1021750 167347 1021774
rect 167015 1021706 167215 1021750
rect 167230 1021740 167254 1021750
rect 167230 1021716 167264 1021740
rect 167275 1021716 167347 1021750
rect 167230 1021706 167347 1021716
rect 167002 1021682 167347 1021706
rect 167015 1021638 167215 1021682
rect 167230 1021672 167254 1021682
rect 167230 1021648 167264 1021672
rect 167275 1021648 167347 1021682
rect 167230 1021638 167347 1021648
rect 167002 1021614 167347 1021638
rect 167015 1021570 167215 1021614
rect 167230 1021604 167254 1021614
rect 167230 1021580 167264 1021604
rect 167275 1021580 167347 1021614
rect 167230 1021570 167347 1021580
rect 167002 1021546 167347 1021570
rect 167015 1021502 167215 1021546
rect 167230 1021536 167254 1021546
rect 167230 1021512 167264 1021536
rect 167275 1021512 167347 1021546
rect 167230 1021502 167347 1021512
rect 167002 1021478 167347 1021502
rect 167015 1021434 167215 1021478
rect 167230 1021468 167254 1021478
rect 167230 1021444 167264 1021468
rect 167275 1021444 167347 1021478
rect 167230 1021434 167347 1021444
rect 167002 1021410 167347 1021434
rect 167015 1021366 167215 1021410
rect 167230 1021400 167254 1021410
rect 167230 1021376 167264 1021400
rect 167275 1021376 167347 1021410
rect 167230 1021366 167347 1021376
rect 167002 1021342 167347 1021366
rect 167015 1021298 167215 1021342
rect 167230 1021332 167254 1021342
rect 167230 1021308 167264 1021332
rect 167275 1021308 167347 1021342
rect 167230 1021298 167347 1021308
rect 167002 1021274 167347 1021298
rect 167015 1021230 167215 1021274
rect 167230 1021264 167254 1021274
rect 167230 1021240 167264 1021264
rect 167275 1021240 167347 1021274
rect 167230 1021230 167347 1021240
rect 167002 1021206 167347 1021230
rect 167015 1021162 167215 1021206
rect 167230 1021196 167254 1021206
rect 167230 1021172 167264 1021196
rect 167275 1021172 167347 1021206
rect 167230 1021162 167347 1021172
rect 167002 1021138 167347 1021162
rect 167015 1021094 167215 1021138
rect 167230 1021128 167254 1021138
rect 167230 1021104 167264 1021128
rect 167275 1021104 167347 1021138
rect 167230 1021094 167347 1021104
rect 167002 1021070 167347 1021094
rect 167015 1021026 167215 1021070
rect 167230 1021060 167254 1021070
rect 167230 1021036 167264 1021060
rect 167275 1021036 167347 1021070
rect 167230 1021026 167347 1021036
rect 167002 1021002 167347 1021026
rect 167015 1020958 167215 1021002
rect 167230 1020992 167254 1021002
rect 167230 1020968 167264 1020992
rect 167275 1020968 167347 1021002
rect 167230 1020958 167347 1020968
rect 167002 1020934 167347 1020958
rect 167015 1020922 167215 1020934
rect 167026 1020910 167050 1020922
rect 167230 1020910 167254 1020934
rect 167275 1020922 167347 1020934
rect 167577 1020922 167633 1021922
rect 167649 1020922 167705 1021922
rect 168007 1021842 168207 1021922
rect 168222 1021852 168256 1021876
rect 168267 1021852 168339 1021922
rect 168222 1021842 168339 1021852
rect 167994 1021818 168339 1021842
rect 168007 1021774 168207 1021818
rect 168222 1021808 168246 1021818
rect 168222 1021784 168256 1021808
rect 168267 1021784 168339 1021818
rect 168222 1021774 168339 1021784
rect 167994 1021750 168339 1021774
rect 168007 1021706 168207 1021750
rect 168222 1021740 168246 1021750
rect 168222 1021716 168256 1021740
rect 168267 1021716 168339 1021750
rect 168222 1021706 168339 1021716
rect 167994 1021682 168339 1021706
rect 168007 1021638 168207 1021682
rect 168222 1021672 168246 1021682
rect 168222 1021648 168256 1021672
rect 168267 1021648 168339 1021682
rect 168222 1021638 168339 1021648
rect 167994 1021614 168339 1021638
rect 168007 1021570 168207 1021614
rect 168222 1021604 168246 1021614
rect 168222 1021580 168256 1021604
rect 168267 1021580 168339 1021614
rect 168222 1021570 168339 1021580
rect 167994 1021546 168339 1021570
rect 168007 1021502 168207 1021546
rect 168222 1021536 168246 1021546
rect 168222 1021512 168256 1021536
rect 168267 1021512 168339 1021546
rect 168222 1021502 168339 1021512
rect 167994 1021478 168339 1021502
rect 168007 1021434 168207 1021478
rect 168222 1021468 168246 1021478
rect 168222 1021444 168256 1021468
rect 168267 1021444 168339 1021478
rect 168222 1021434 168339 1021444
rect 167994 1021410 168339 1021434
rect 168007 1021366 168207 1021410
rect 168222 1021400 168246 1021410
rect 168222 1021376 168256 1021400
rect 168267 1021376 168339 1021410
rect 168222 1021366 168339 1021376
rect 167994 1021342 168339 1021366
rect 168007 1021298 168207 1021342
rect 168222 1021332 168246 1021342
rect 168222 1021308 168256 1021332
rect 168267 1021308 168339 1021342
rect 168222 1021298 168339 1021308
rect 167994 1021274 168339 1021298
rect 168007 1021230 168207 1021274
rect 168222 1021264 168246 1021274
rect 168222 1021240 168256 1021264
rect 168267 1021240 168339 1021274
rect 168222 1021230 168339 1021240
rect 167994 1021206 168339 1021230
rect 168007 1021162 168207 1021206
rect 168222 1021196 168246 1021206
rect 168222 1021172 168256 1021196
rect 168267 1021172 168339 1021206
rect 168222 1021162 168339 1021172
rect 167994 1021138 168339 1021162
rect 168007 1021094 168207 1021138
rect 168222 1021128 168246 1021138
rect 168222 1021104 168256 1021128
rect 168267 1021104 168339 1021138
rect 168222 1021094 168339 1021104
rect 167994 1021070 168339 1021094
rect 168007 1021026 168207 1021070
rect 168222 1021060 168246 1021070
rect 168222 1021036 168256 1021060
rect 168267 1021036 168339 1021070
rect 168222 1021026 168339 1021036
rect 167994 1021002 168339 1021026
rect 168007 1020958 168207 1021002
rect 168222 1020992 168246 1021002
rect 168222 1020968 168256 1020992
rect 168267 1020968 168339 1021002
rect 168222 1020958 168339 1020968
rect 167994 1020934 168339 1020958
rect 168007 1020922 168207 1020934
rect 168018 1020910 168042 1020922
rect 168222 1020910 168246 1020934
rect 168267 1020922 168339 1020934
rect 168569 1020922 168625 1021922
rect 168641 1020922 168697 1021922
rect 168999 1021842 169199 1021922
rect 169214 1021852 169248 1021876
rect 169259 1021852 169331 1021922
rect 169214 1021842 169331 1021852
rect 168986 1021818 169331 1021842
rect 168999 1021774 169199 1021818
rect 169214 1021808 169238 1021818
rect 169214 1021784 169248 1021808
rect 169259 1021784 169331 1021818
rect 169214 1021774 169331 1021784
rect 168986 1021750 169331 1021774
rect 168999 1021706 169199 1021750
rect 169214 1021740 169238 1021750
rect 169214 1021716 169248 1021740
rect 169259 1021716 169331 1021750
rect 169214 1021706 169331 1021716
rect 168986 1021682 169331 1021706
rect 168999 1021638 169199 1021682
rect 169214 1021672 169238 1021682
rect 169214 1021648 169248 1021672
rect 169259 1021648 169331 1021682
rect 169214 1021638 169331 1021648
rect 168986 1021614 169331 1021638
rect 168999 1021570 169199 1021614
rect 169214 1021604 169238 1021614
rect 169214 1021580 169248 1021604
rect 169259 1021580 169331 1021614
rect 169214 1021570 169331 1021580
rect 168986 1021546 169331 1021570
rect 168999 1021502 169199 1021546
rect 169214 1021536 169238 1021546
rect 169214 1021512 169248 1021536
rect 169259 1021512 169331 1021546
rect 169214 1021502 169331 1021512
rect 168986 1021478 169331 1021502
rect 168999 1021434 169199 1021478
rect 169214 1021468 169238 1021478
rect 169214 1021444 169248 1021468
rect 169259 1021444 169331 1021478
rect 169214 1021434 169331 1021444
rect 168986 1021410 169331 1021434
rect 168999 1021366 169199 1021410
rect 169214 1021400 169238 1021410
rect 169214 1021376 169248 1021400
rect 169259 1021376 169331 1021410
rect 169214 1021366 169331 1021376
rect 168986 1021342 169331 1021366
rect 168999 1021298 169199 1021342
rect 169214 1021332 169238 1021342
rect 169214 1021308 169248 1021332
rect 169259 1021308 169331 1021342
rect 169214 1021298 169331 1021308
rect 168986 1021274 169331 1021298
rect 168999 1021230 169199 1021274
rect 169214 1021264 169238 1021274
rect 169214 1021240 169248 1021264
rect 169259 1021240 169331 1021274
rect 169214 1021230 169331 1021240
rect 168986 1021206 169331 1021230
rect 168999 1021162 169199 1021206
rect 169214 1021196 169238 1021206
rect 169214 1021172 169248 1021196
rect 169259 1021172 169331 1021206
rect 169214 1021162 169331 1021172
rect 168986 1021138 169331 1021162
rect 168999 1021094 169199 1021138
rect 169214 1021128 169238 1021138
rect 169214 1021104 169248 1021128
rect 169259 1021104 169331 1021138
rect 169214 1021094 169331 1021104
rect 168986 1021070 169331 1021094
rect 168999 1021026 169199 1021070
rect 169214 1021060 169238 1021070
rect 169214 1021036 169248 1021060
rect 169259 1021036 169331 1021070
rect 169214 1021026 169331 1021036
rect 168986 1021002 169331 1021026
rect 168999 1020958 169199 1021002
rect 169214 1020992 169238 1021002
rect 169214 1020968 169248 1020992
rect 169259 1020968 169331 1021002
rect 169214 1020958 169331 1020968
rect 168986 1020934 169331 1020958
rect 168999 1020922 169199 1020934
rect 169010 1020910 169034 1020922
rect 169214 1020910 169238 1020934
rect 169259 1020922 169331 1020934
rect 169561 1020922 169617 1021922
rect 169633 1020922 169689 1021922
rect 169991 1021842 170191 1021922
rect 170206 1021852 170240 1021876
rect 170251 1021852 170323 1021922
rect 170206 1021842 170323 1021852
rect 169978 1021818 170323 1021842
rect 169991 1021774 170191 1021818
rect 170206 1021808 170230 1021818
rect 170206 1021784 170240 1021808
rect 170251 1021784 170323 1021818
rect 170206 1021774 170323 1021784
rect 169978 1021750 170323 1021774
rect 169991 1021706 170191 1021750
rect 170206 1021740 170230 1021750
rect 170206 1021716 170240 1021740
rect 170251 1021716 170323 1021750
rect 170206 1021706 170323 1021716
rect 169978 1021682 170323 1021706
rect 169991 1021638 170191 1021682
rect 170206 1021672 170230 1021682
rect 170206 1021648 170240 1021672
rect 170251 1021648 170323 1021682
rect 170206 1021638 170323 1021648
rect 169978 1021614 170323 1021638
rect 169991 1021570 170191 1021614
rect 170206 1021604 170230 1021614
rect 170206 1021580 170240 1021604
rect 170251 1021580 170323 1021614
rect 170206 1021570 170323 1021580
rect 169978 1021546 170323 1021570
rect 169991 1021502 170191 1021546
rect 170206 1021536 170230 1021546
rect 170206 1021512 170240 1021536
rect 170251 1021512 170323 1021546
rect 170206 1021502 170323 1021512
rect 169978 1021478 170323 1021502
rect 169991 1021434 170191 1021478
rect 170206 1021468 170230 1021478
rect 170206 1021444 170240 1021468
rect 170251 1021444 170323 1021478
rect 170206 1021434 170323 1021444
rect 169978 1021410 170323 1021434
rect 169991 1021366 170191 1021410
rect 170206 1021400 170230 1021410
rect 170206 1021376 170240 1021400
rect 170251 1021376 170323 1021410
rect 170206 1021366 170323 1021376
rect 169978 1021342 170323 1021366
rect 169991 1021298 170191 1021342
rect 170206 1021332 170230 1021342
rect 170206 1021308 170240 1021332
rect 170251 1021308 170323 1021342
rect 170206 1021298 170323 1021308
rect 169978 1021274 170323 1021298
rect 169991 1021230 170191 1021274
rect 170206 1021264 170230 1021274
rect 170206 1021240 170240 1021264
rect 170251 1021240 170323 1021274
rect 170206 1021230 170323 1021240
rect 169978 1021206 170323 1021230
rect 169991 1021162 170191 1021206
rect 170206 1021196 170230 1021206
rect 170206 1021172 170240 1021196
rect 170251 1021172 170323 1021206
rect 170206 1021162 170323 1021172
rect 169978 1021138 170323 1021162
rect 169991 1021094 170191 1021138
rect 170206 1021128 170230 1021138
rect 170206 1021104 170240 1021128
rect 170251 1021104 170323 1021138
rect 170206 1021094 170323 1021104
rect 169978 1021070 170323 1021094
rect 169991 1021026 170191 1021070
rect 170206 1021060 170230 1021070
rect 170206 1021036 170240 1021060
rect 170251 1021036 170323 1021070
rect 170206 1021026 170323 1021036
rect 169978 1021002 170323 1021026
rect 169991 1020958 170191 1021002
rect 170206 1020992 170230 1021002
rect 170206 1020968 170240 1020992
rect 170251 1020968 170323 1021002
rect 170206 1020958 170323 1020968
rect 169978 1020934 170323 1020958
rect 169991 1020922 170191 1020934
rect 170002 1020910 170026 1020922
rect 170206 1020910 170230 1020934
rect 170251 1020922 170323 1020934
rect 170553 1020922 170609 1021922
rect 170625 1020922 170681 1021922
rect 170983 1021842 171183 1021922
rect 171198 1021852 171232 1021876
rect 171243 1021852 171315 1021922
rect 171198 1021842 171315 1021852
rect 170970 1021818 171315 1021842
rect 170983 1021774 171183 1021818
rect 171198 1021808 171222 1021818
rect 171198 1021784 171232 1021808
rect 171243 1021784 171315 1021818
rect 171198 1021774 171315 1021784
rect 170970 1021750 171315 1021774
rect 170983 1021706 171183 1021750
rect 171198 1021740 171222 1021750
rect 171198 1021716 171232 1021740
rect 171243 1021716 171315 1021750
rect 171198 1021706 171315 1021716
rect 170970 1021682 171315 1021706
rect 170983 1021638 171183 1021682
rect 171198 1021672 171222 1021682
rect 171198 1021648 171232 1021672
rect 171243 1021648 171315 1021682
rect 171198 1021638 171315 1021648
rect 170970 1021614 171315 1021638
rect 170983 1021570 171183 1021614
rect 171198 1021604 171222 1021614
rect 171198 1021580 171232 1021604
rect 171243 1021580 171315 1021614
rect 171198 1021570 171315 1021580
rect 170970 1021546 171315 1021570
rect 170983 1021502 171183 1021546
rect 171198 1021536 171222 1021546
rect 171198 1021512 171232 1021536
rect 171243 1021512 171315 1021546
rect 171198 1021502 171315 1021512
rect 170970 1021478 171315 1021502
rect 170983 1021434 171183 1021478
rect 171198 1021468 171222 1021478
rect 171198 1021444 171232 1021468
rect 171243 1021444 171315 1021478
rect 171198 1021434 171315 1021444
rect 170970 1021410 171315 1021434
rect 170983 1021366 171183 1021410
rect 171198 1021400 171222 1021410
rect 171198 1021376 171232 1021400
rect 171243 1021376 171315 1021410
rect 171198 1021366 171315 1021376
rect 170970 1021342 171315 1021366
rect 170983 1021298 171183 1021342
rect 171198 1021332 171222 1021342
rect 171198 1021308 171232 1021332
rect 171243 1021308 171315 1021342
rect 171198 1021298 171315 1021308
rect 170970 1021274 171315 1021298
rect 170983 1021230 171183 1021274
rect 171198 1021264 171222 1021274
rect 171198 1021240 171232 1021264
rect 171243 1021240 171315 1021274
rect 171198 1021230 171315 1021240
rect 170970 1021206 171315 1021230
rect 170983 1021162 171183 1021206
rect 171198 1021196 171222 1021206
rect 171198 1021172 171232 1021196
rect 171243 1021172 171315 1021206
rect 171198 1021162 171315 1021172
rect 170970 1021138 171315 1021162
rect 170983 1021094 171183 1021138
rect 171198 1021128 171222 1021138
rect 171198 1021104 171232 1021128
rect 171243 1021104 171315 1021138
rect 171198 1021094 171315 1021104
rect 170970 1021070 171315 1021094
rect 170983 1021026 171183 1021070
rect 171198 1021060 171222 1021070
rect 171198 1021036 171232 1021060
rect 171243 1021036 171315 1021070
rect 171198 1021026 171315 1021036
rect 170970 1021002 171315 1021026
rect 170983 1020958 171183 1021002
rect 171198 1020992 171222 1021002
rect 171198 1020968 171232 1020992
rect 171243 1020968 171315 1021002
rect 171198 1020958 171315 1020968
rect 170970 1020934 171315 1020958
rect 170983 1020922 171183 1020934
rect 170994 1020910 171018 1020922
rect 171198 1020910 171222 1020934
rect 171243 1020922 171315 1020934
rect 171545 1020922 171601 1021922
rect 171617 1020922 171673 1021922
rect 171975 1021842 172175 1021922
rect 172190 1021852 172224 1021876
rect 172235 1021852 172307 1021922
rect 172190 1021842 172307 1021852
rect 171962 1021818 172307 1021842
rect 171975 1021774 172175 1021818
rect 172190 1021808 172214 1021818
rect 172190 1021784 172224 1021808
rect 172235 1021784 172307 1021818
rect 172190 1021774 172307 1021784
rect 171962 1021750 172307 1021774
rect 171975 1021706 172175 1021750
rect 172190 1021740 172214 1021750
rect 172190 1021716 172224 1021740
rect 172235 1021716 172307 1021750
rect 172190 1021706 172307 1021716
rect 171962 1021682 172307 1021706
rect 171975 1021638 172175 1021682
rect 172190 1021672 172214 1021682
rect 172190 1021648 172224 1021672
rect 172235 1021648 172307 1021682
rect 172190 1021638 172307 1021648
rect 171962 1021614 172307 1021638
rect 171975 1021570 172175 1021614
rect 172190 1021604 172214 1021614
rect 172190 1021580 172224 1021604
rect 172235 1021580 172307 1021614
rect 172190 1021570 172307 1021580
rect 171962 1021546 172307 1021570
rect 171975 1021502 172175 1021546
rect 172190 1021536 172214 1021546
rect 172190 1021512 172224 1021536
rect 172235 1021512 172307 1021546
rect 172190 1021502 172307 1021512
rect 171962 1021478 172307 1021502
rect 171975 1021434 172175 1021478
rect 172190 1021468 172214 1021478
rect 172190 1021444 172224 1021468
rect 172235 1021444 172307 1021478
rect 172190 1021434 172307 1021444
rect 171962 1021410 172307 1021434
rect 171975 1021366 172175 1021410
rect 172190 1021400 172214 1021410
rect 172190 1021376 172224 1021400
rect 172235 1021376 172307 1021410
rect 172190 1021366 172307 1021376
rect 171962 1021342 172307 1021366
rect 171975 1021298 172175 1021342
rect 172190 1021332 172214 1021342
rect 172190 1021308 172224 1021332
rect 172235 1021308 172307 1021342
rect 172190 1021298 172307 1021308
rect 171962 1021274 172307 1021298
rect 171975 1021230 172175 1021274
rect 172190 1021264 172214 1021274
rect 172190 1021240 172224 1021264
rect 172235 1021240 172307 1021274
rect 172190 1021230 172307 1021240
rect 171962 1021206 172307 1021230
rect 171975 1021162 172175 1021206
rect 172190 1021196 172214 1021206
rect 172190 1021172 172224 1021196
rect 172235 1021172 172307 1021206
rect 172190 1021162 172307 1021172
rect 171962 1021138 172307 1021162
rect 171975 1021094 172175 1021138
rect 172190 1021128 172214 1021138
rect 172190 1021104 172224 1021128
rect 172235 1021104 172307 1021138
rect 172190 1021094 172307 1021104
rect 171962 1021070 172307 1021094
rect 171975 1021026 172175 1021070
rect 172190 1021060 172214 1021070
rect 172190 1021036 172224 1021060
rect 172235 1021036 172307 1021070
rect 172190 1021026 172307 1021036
rect 171962 1021002 172307 1021026
rect 171975 1020958 172175 1021002
rect 172190 1020992 172214 1021002
rect 172190 1020968 172224 1020992
rect 172235 1020968 172307 1021002
rect 172190 1020958 172307 1020968
rect 171962 1020934 172307 1020958
rect 171975 1020922 172175 1020934
rect 171986 1020910 172010 1020922
rect 172190 1020910 172214 1020934
rect 172235 1020922 172307 1020934
rect 172537 1020922 172593 1021922
rect 172609 1020922 172665 1021922
rect 172967 1021842 173167 1021922
rect 173182 1021852 173216 1021876
rect 173227 1021852 173299 1021922
rect 173182 1021842 173299 1021852
rect 172954 1021818 173299 1021842
rect 172967 1021774 173167 1021818
rect 173182 1021808 173206 1021818
rect 173182 1021784 173216 1021808
rect 173227 1021784 173299 1021818
rect 173182 1021774 173299 1021784
rect 172954 1021750 173299 1021774
rect 172967 1021706 173167 1021750
rect 173182 1021740 173206 1021750
rect 173182 1021716 173216 1021740
rect 173227 1021716 173299 1021750
rect 173182 1021706 173299 1021716
rect 172954 1021682 173299 1021706
rect 172967 1021638 173167 1021682
rect 173182 1021672 173206 1021682
rect 173182 1021648 173216 1021672
rect 173227 1021648 173299 1021682
rect 173182 1021638 173299 1021648
rect 172954 1021614 173299 1021638
rect 172967 1021570 173167 1021614
rect 173182 1021604 173206 1021614
rect 173182 1021580 173216 1021604
rect 173227 1021580 173299 1021614
rect 173182 1021570 173299 1021580
rect 172954 1021546 173299 1021570
rect 172967 1021502 173167 1021546
rect 173182 1021536 173206 1021546
rect 173182 1021512 173216 1021536
rect 173227 1021512 173299 1021546
rect 173182 1021502 173299 1021512
rect 172954 1021478 173299 1021502
rect 172967 1021434 173167 1021478
rect 173182 1021468 173206 1021478
rect 173182 1021444 173216 1021468
rect 173227 1021444 173299 1021478
rect 173182 1021434 173299 1021444
rect 172954 1021410 173299 1021434
rect 172967 1021366 173167 1021410
rect 173182 1021400 173206 1021410
rect 173182 1021376 173216 1021400
rect 173227 1021376 173299 1021410
rect 173182 1021366 173299 1021376
rect 172954 1021342 173299 1021366
rect 172967 1021298 173167 1021342
rect 173182 1021332 173206 1021342
rect 173182 1021308 173216 1021332
rect 173227 1021308 173299 1021342
rect 173182 1021298 173299 1021308
rect 172954 1021274 173299 1021298
rect 172967 1021230 173167 1021274
rect 173182 1021264 173206 1021274
rect 173182 1021240 173216 1021264
rect 173227 1021240 173299 1021274
rect 173182 1021230 173299 1021240
rect 172954 1021206 173299 1021230
rect 172967 1021162 173167 1021206
rect 173182 1021196 173206 1021206
rect 173182 1021172 173216 1021196
rect 173227 1021172 173299 1021206
rect 173182 1021162 173299 1021172
rect 172954 1021138 173299 1021162
rect 172967 1021094 173167 1021138
rect 173182 1021128 173206 1021138
rect 173182 1021104 173216 1021128
rect 173227 1021104 173299 1021138
rect 173182 1021094 173299 1021104
rect 172954 1021070 173299 1021094
rect 172967 1021026 173167 1021070
rect 173182 1021060 173206 1021070
rect 173182 1021036 173216 1021060
rect 173227 1021036 173299 1021070
rect 173182 1021026 173299 1021036
rect 172954 1021002 173299 1021026
rect 172967 1020958 173167 1021002
rect 173182 1020992 173206 1021002
rect 173182 1020968 173216 1020992
rect 173227 1020968 173299 1021002
rect 173182 1020958 173299 1020968
rect 172954 1020934 173299 1020958
rect 172967 1020922 173167 1020934
rect 172978 1020910 173002 1020922
rect 173182 1020910 173206 1020934
rect 173227 1020922 173299 1020934
rect 173529 1020922 173585 1021922
rect 173601 1020922 173657 1021922
rect 173959 1021842 174159 1021922
rect 174174 1021852 174208 1021876
rect 174219 1021852 174291 1021922
rect 174174 1021842 174291 1021852
rect 173946 1021818 174291 1021842
rect 173959 1021774 174159 1021818
rect 174174 1021808 174198 1021818
rect 174174 1021784 174208 1021808
rect 174219 1021784 174291 1021818
rect 174174 1021774 174291 1021784
rect 173946 1021750 174291 1021774
rect 173959 1021706 174159 1021750
rect 174174 1021740 174198 1021750
rect 174174 1021716 174208 1021740
rect 174219 1021716 174291 1021750
rect 174174 1021706 174291 1021716
rect 173946 1021682 174291 1021706
rect 173959 1021638 174159 1021682
rect 174174 1021672 174198 1021682
rect 174174 1021648 174208 1021672
rect 174219 1021648 174291 1021682
rect 174174 1021638 174291 1021648
rect 173946 1021614 174291 1021638
rect 173959 1021570 174159 1021614
rect 174174 1021604 174198 1021614
rect 174174 1021580 174208 1021604
rect 174219 1021580 174291 1021614
rect 174174 1021570 174291 1021580
rect 173946 1021546 174291 1021570
rect 173959 1021502 174159 1021546
rect 174174 1021536 174198 1021546
rect 174174 1021512 174208 1021536
rect 174219 1021512 174291 1021546
rect 174174 1021502 174291 1021512
rect 173946 1021478 174291 1021502
rect 173959 1021434 174159 1021478
rect 174174 1021468 174198 1021478
rect 174174 1021444 174208 1021468
rect 174219 1021444 174291 1021478
rect 174174 1021434 174291 1021444
rect 173946 1021410 174291 1021434
rect 173959 1021366 174159 1021410
rect 174174 1021400 174198 1021410
rect 174174 1021376 174208 1021400
rect 174219 1021376 174291 1021410
rect 174174 1021366 174291 1021376
rect 173946 1021342 174291 1021366
rect 173959 1021298 174159 1021342
rect 174174 1021332 174198 1021342
rect 174174 1021308 174208 1021332
rect 174219 1021308 174291 1021342
rect 174174 1021298 174291 1021308
rect 173946 1021274 174291 1021298
rect 173959 1021230 174159 1021274
rect 174174 1021264 174198 1021274
rect 174174 1021240 174208 1021264
rect 174219 1021240 174291 1021274
rect 174174 1021230 174291 1021240
rect 173946 1021206 174291 1021230
rect 173959 1021162 174159 1021206
rect 174174 1021196 174198 1021206
rect 174174 1021172 174208 1021196
rect 174219 1021172 174291 1021206
rect 174174 1021162 174291 1021172
rect 173946 1021138 174291 1021162
rect 173959 1021094 174159 1021138
rect 174174 1021128 174198 1021138
rect 174174 1021104 174208 1021128
rect 174219 1021104 174291 1021138
rect 174174 1021094 174291 1021104
rect 173946 1021070 174291 1021094
rect 173959 1021026 174159 1021070
rect 174174 1021060 174198 1021070
rect 174174 1021036 174208 1021060
rect 174219 1021036 174291 1021070
rect 174174 1021026 174291 1021036
rect 173946 1021002 174291 1021026
rect 173959 1020958 174159 1021002
rect 174174 1020992 174198 1021002
rect 174174 1020968 174208 1020992
rect 174219 1020968 174291 1021002
rect 174174 1020958 174291 1020968
rect 173946 1020934 174291 1020958
rect 173959 1020922 174159 1020934
rect 173970 1020910 173994 1020922
rect 174174 1020910 174198 1020934
rect 174219 1020922 174291 1020934
rect 174521 1020922 174577 1021922
rect 174593 1020922 174649 1021922
rect 174951 1021842 175151 1021922
rect 175166 1021852 175200 1021876
rect 175211 1021852 175283 1021922
rect 175166 1021842 175283 1021852
rect 174938 1021818 175283 1021842
rect 174951 1021774 175151 1021818
rect 175166 1021808 175190 1021818
rect 175166 1021784 175200 1021808
rect 175211 1021784 175283 1021818
rect 175166 1021774 175283 1021784
rect 174938 1021750 175283 1021774
rect 174951 1021706 175151 1021750
rect 175166 1021740 175190 1021750
rect 175166 1021716 175200 1021740
rect 175211 1021716 175283 1021750
rect 175166 1021706 175283 1021716
rect 174938 1021682 175283 1021706
rect 174951 1021638 175151 1021682
rect 175166 1021672 175190 1021682
rect 175166 1021648 175200 1021672
rect 175211 1021648 175283 1021682
rect 175166 1021638 175283 1021648
rect 174938 1021614 175283 1021638
rect 174951 1021570 175151 1021614
rect 175166 1021604 175190 1021614
rect 175166 1021580 175200 1021604
rect 175211 1021580 175283 1021614
rect 175166 1021570 175283 1021580
rect 174938 1021546 175283 1021570
rect 174951 1021502 175151 1021546
rect 175166 1021536 175190 1021546
rect 175166 1021512 175200 1021536
rect 175211 1021512 175283 1021546
rect 175166 1021502 175283 1021512
rect 174938 1021478 175283 1021502
rect 174951 1021434 175151 1021478
rect 175166 1021468 175190 1021478
rect 175166 1021444 175200 1021468
rect 175211 1021444 175283 1021478
rect 175166 1021434 175283 1021444
rect 174938 1021410 175283 1021434
rect 174951 1021366 175151 1021410
rect 175166 1021400 175190 1021410
rect 175166 1021376 175200 1021400
rect 175211 1021376 175283 1021410
rect 175166 1021366 175283 1021376
rect 174938 1021342 175283 1021366
rect 174951 1021298 175151 1021342
rect 175166 1021332 175190 1021342
rect 175166 1021308 175200 1021332
rect 175211 1021308 175283 1021342
rect 175166 1021298 175283 1021308
rect 174938 1021274 175283 1021298
rect 174951 1021230 175151 1021274
rect 175166 1021264 175190 1021274
rect 175166 1021240 175200 1021264
rect 175211 1021240 175283 1021274
rect 175166 1021230 175283 1021240
rect 174938 1021206 175283 1021230
rect 174951 1021162 175151 1021206
rect 175166 1021196 175190 1021206
rect 175166 1021172 175200 1021196
rect 175211 1021172 175283 1021206
rect 175166 1021162 175283 1021172
rect 174938 1021138 175283 1021162
rect 174951 1021094 175151 1021138
rect 175166 1021128 175190 1021138
rect 175166 1021104 175200 1021128
rect 175211 1021104 175283 1021138
rect 175166 1021094 175283 1021104
rect 174938 1021070 175283 1021094
rect 174951 1021026 175151 1021070
rect 175166 1021060 175190 1021070
rect 175166 1021036 175200 1021060
rect 175211 1021036 175283 1021070
rect 175166 1021026 175283 1021036
rect 174938 1021002 175283 1021026
rect 174951 1020958 175151 1021002
rect 175166 1020992 175190 1021002
rect 175166 1020968 175200 1020992
rect 175211 1020968 175283 1021002
rect 175166 1020958 175283 1020968
rect 174938 1020934 175283 1020958
rect 174951 1020922 175151 1020934
rect 174962 1020910 174986 1020922
rect 175166 1020910 175190 1020934
rect 175211 1020922 175283 1020934
rect 175472 1020922 175544 1021922
rect 175610 1020922 175627 1021922
rect 175797 1020922 175830 1021922
rect 175953 1021730 176025 1021760
rect 175953 1021692 175987 1021722
rect 163058 1020322 163092 1020334
rect 162356 1019322 162406 1020322
rect 162617 1019322 162673 1020322
rect 162689 1019322 162745 1020322
rect 163047 1020300 163247 1020322
rect 163262 1020310 163296 1020334
rect 164050 1020322 164084 1020334
rect 163307 1020310 163379 1020322
rect 163262 1020300 163379 1020310
rect 163034 1020276 163379 1020300
rect 163047 1020232 163247 1020276
rect 163262 1020266 163286 1020276
rect 163262 1020242 163296 1020266
rect 163307 1020242 163379 1020276
rect 163262 1020232 163379 1020242
rect 163034 1020208 163379 1020232
rect 163047 1020164 163247 1020208
rect 163262 1020198 163286 1020208
rect 163262 1020174 163296 1020198
rect 163307 1020174 163379 1020208
rect 163262 1020164 163379 1020174
rect 163034 1020140 163379 1020164
rect 163047 1020096 163247 1020140
rect 163262 1020130 163286 1020140
rect 163262 1020106 163296 1020130
rect 163307 1020106 163379 1020140
rect 163262 1020096 163379 1020106
rect 163034 1020072 163379 1020096
rect 163047 1020028 163247 1020072
rect 163262 1020062 163286 1020072
rect 163262 1020038 163296 1020062
rect 163307 1020038 163379 1020072
rect 163262 1020028 163379 1020038
rect 163034 1020004 163379 1020028
rect 163047 1019960 163247 1020004
rect 163262 1019994 163286 1020004
rect 163262 1019970 163296 1019994
rect 163307 1019970 163379 1020004
rect 163262 1019960 163379 1019970
rect 163034 1019936 163379 1019960
rect 163047 1019892 163247 1019936
rect 163262 1019926 163286 1019936
rect 163262 1019902 163296 1019926
rect 163307 1019902 163379 1019936
rect 163262 1019892 163379 1019902
rect 163034 1019868 163379 1019892
rect 163047 1019824 163247 1019868
rect 163262 1019858 163286 1019868
rect 163262 1019834 163296 1019858
rect 163307 1019834 163379 1019868
rect 163262 1019824 163379 1019834
rect 163034 1019800 163379 1019824
rect 163047 1019756 163247 1019800
rect 163262 1019790 163286 1019800
rect 163262 1019766 163296 1019790
rect 163307 1019766 163379 1019800
rect 163262 1019756 163379 1019766
rect 163034 1019732 163379 1019756
rect 163047 1019688 163247 1019732
rect 163262 1019722 163286 1019732
rect 163262 1019698 163296 1019722
rect 163307 1019698 163379 1019732
rect 163262 1019688 163379 1019698
rect 163034 1019664 163379 1019688
rect 163047 1019620 163247 1019664
rect 163262 1019654 163286 1019664
rect 163262 1019630 163296 1019654
rect 163307 1019630 163379 1019664
rect 163262 1019620 163379 1019630
rect 163034 1019596 163379 1019620
rect 163047 1019552 163247 1019596
rect 163262 1019586 163286 1019596
rect 163262 1019562 163296 1019586
rect 163307 1019562 163379 1019596
rect 163262 1019552 163379 1019562
rect 163034 1019528 163379 1019552
rect 163047 1019484 163247 1019528
rect 163262 1019518 163286 1019528
rect 163262 1019494 163296 1019518
rect 163307 1019494 163379 1019528
rect 163262 1019484 163379 1019494
rect 163034 1019460 163379 1019484
rect 163047 1019416 163247 1019460
rect 163262 1019450 163286 1019460
rect 163262 1019426 163296 1019450
rect 163307 1019426 163379 1019460
rect 163262 1019416 163379 1019426
rect 163034 1019392 163379 1019416
rect 163047 1019322 163247 1019392
rect 163262 1019368 163286 1019392
rect 163307 1019322 163379 1019392
rect 163609 1019322 163665 1020322
rect 163681 1019322 163737 1020322
rect 164039 1020300 164239 1020322
rect 164254 1020310 164288 1020334
rect 165042 1020322 165076 1020334
rect 164299 1020310 164371 1020322
rect 164254 1020300 164371 1020310
rect 164026 1020276 164371 1020300
rect 164039 1020232 164239 1020276
rect 164254 1020266 164278 1020276
rect 164254 1020242 164288 1020266
rect 164299 1020242 164371 1020276
rect 164254 1020232 164371 1020242
rect 164026 1020208 164371 1020232
rect 164039 1020164 164239 1020208
rect 164254 1020198 164278 1020208
rect 164254 1020174 164288 1020198
rect 164299 1020174 164371 1020208
rect 164254 1020164 164371 1020174
rect 164026 1020140 164371 1020164
rect 164039 1020096 164239 1020140
rect 164254 1020130 164278 1020140
rect 164254 1020106 164288 1020130
rect 164299 1020106 164371 1020140
rect 164254 1020096 164371 1020106
rect 164026 1020072 164371 1020096
rect 164039 1020028 164239 1020072
rect 164254 1020062 164278 1020072
rect 164254 1020038 164288 1020062
rect 164299 1020038 164371 1020072
rect 164254 1020028 164371 1020038
rect 164026 1020004 164371 1020028
rect 164039 1019960 164239 1020004
rect 164254 1019994 164278 1020004
rect 164254 1019970 164288 1019994
rect 164299 1019970 164371 1020004
rect 164254 1019960 164371 1019970
rect 164026 1019936 164371 1019960
rect 164039 1019892 164239 1019936
rect 164254 1019926 164278 1019936
rect 164254 1019902 164288 1019926
rect 164299 1019902 164371 1019936
rect 164254 1019892 164371 1019902
rect 164026 1019868 164371 1019892
rect 164039 1019824 164239 1019868
rect 164254 1019858 164278 1019868
rect 164254 1019834 164288 1019858
rect 164299 1019834 164371 1019868
rect 164254 1019824 164371 1019834
rect 164026 1019800 164371 1019824
rect 164039 1019756 164239 1019800
rect 164254 1019790 164278 1019800
rect 164254 1019766 164288 1019790
rect 164299 1019766 164371 1019800
rect 164254 1019756 164371 1019766
rect 164026 1019732 164371 1019756
rect 164039 1019688 164239 1019732
rect 164254 1019722 164278 1019732
rect 164254 1019698 164288 1019722
rect 164299 1019698 164371 1019732
rect 164254 1019688 164371 1019698
rect 164026 1019664 164371 1019688
rect 164039 1019620 164239 1019664
rect 164254 1019654 164278 1019664
rect 164254 1019630 164288 1019654
rect 164299 1019630 164371 1019664
rect 164254 1019620 164371 1019630
rect 164026 1019596 164371 1019620
rect 164039 1019552 164239 1019596
rect 164254 1019586 164278 1019596
rect 164254 1019562 164288 1019586
rect 164299 1019562 164371 1019596
rect 164254 1019552 164371 1019562
rect 164026 1019528 164371 1019552
rect 164039 1019484 164239 1019528
rect 164254 1019518 164278 1019528
rect 164254 1019494 164288 1019518
rect 164299 1019494 164371 1019528
rect 164254 1019484 164371 1019494
rect 164026 1019460 164371 1019484
rect 164039 1019416 164239 1019460
rect 164254 1019450 164278 1019460
rect 164254 1019426 164288 1019450
rect 164299 1019426 164371 1019460
rect 164254 1019416 164371 1019426
rect 164026 1019392 164371 1019416
rect 164039 1019322 164239 1019392
rect 164254 1019368 164278 1019392
rect 164299 1019322 164371 1019392
rect 164601 1019322 164657 1020322
rect 164673 1019322 164729 1020322
rect 165031 1020300 165231 1020322
rect 165246 1020310 165280 1020334
rect 166034 1020322 166068 1020334
rect 165291 1020310 165363 1020322
rect 165246 1020300 165363 1020310
rect 165018 1020276 165363 1020300
rect 165031 1020232 165231 1020276
rect 165246 1020266 165270 1020276
rect 165246 1020242 165280 1020266
rect 165291 1020242 165363 1020276
rect 165246 1020232 165363 1020242
rect 165018 1020208 165363 1020232
rect 165031 1020164 165231 1020208
rect 165246 1020198 165270 1020208
rect 165246 1020174 165280 1020198
rect 165291 1020174 165363 1020208
rect 165246 1020164 165363 1020174
rect 165018 1020140 165363 1020164
rect 165031 1020096 165231 1020140
rect 165246 1020130 165270 1020140
rect 165246 1020106 165280 1020130
rect 165291 1020106 165363 1020140
rect 165246 1020096 165363 1020106
rect 165018 1020072 165363 1020096
rect 165031 1020028 165231 1020072
rect 165246 1020062 165270 1020072
rect 165246 1020038 165280 1020062
rect 165291 1020038 165363 1020072
rect 165246 1020028 165363 1020038
rect 165018 1020004 165363 1020028
rect 165031 1019960 165231 1020004
rect 165246 1019994 165270 1020004
rect 165246 1019970 165280 1019994
rect 165291 1019970 165363 1020004
rect 165246 1019960 165363 1019970
rect 165018 1019936 165363 1019960
rect 165031 1019892 165231 1019936
rect 165246 1019926 165270 1019936
rect 165246 1019902 165280 1019926
rect 165291 1019902 165363 1019936
rect 165246 1019892 165363 1019902
rect 165018 1019868 165363 1019892
rect 165031 1019824 165231 1019868
rect 165246 1019858 165270 1019868
rect 165246 1019834 165280 1019858
rect 165291 1019834 165363 1019868
rect 165246 1019824 165363 1019834
rect 165018 1019800 165363 1019824
rect 165031 1019756 165231 1019800
rect 165246 1019790 165270 1019800
rect 165246 1019766 165280 1019790
rect 165291 1019766 165363 1019800
rect 165246 1019756 165363 1019766
rect 165018 1019732 165363 1019756
rect 165031 1019688 165231 1019732
rect 165246 1019722 165270 1019732
rect 165246 1019698 165280 1019722
rect 165291 1019698 165363 1019732
rect 165246 1019688 165363 1019698
rect 165018 1019664 165363 1019688
rect 165031 1019620 165231 1019664
rect 165246 1019654 165270 1019664
rect 165246 1019630 165280 1019654
rect 165291 1019630 165363 1019664
rect 165246 1019620 165363 1019630
rect 165018 1019596 165363 1019620
rect 165031 1019552 165231 1019596
rect 165246 1019586 165270 1019596
rect 165246 1019562 165280 1019586
rect 165291 1019562 165363 1019596
rect 165246 1019552 165363 1019562
rect 165018 1019528 165363 1019552
rect 165031 1019484 165231 1019528
rect 165246 1019518 165270 1019528
rect 165246 1019494 165280 1019518
rect 165291 1019494 165363 1019528
rect 165246 1019484 165363 1019494
rect 165018 1019460 165363 1019484
rect 165031 1019416 165231 1019460
rect 165246 1019450 165270 1019460
rect 165246 1019426 165280 1019450
rect 165291 1019426 165363 1019460
rect 165246 1019416 165363 1019426
rect 165018 1019392 165363 1019416
rect 165031 1019322 165231 1019392
rect 165246 1019368 165270 1019392
rect 165291 1019322 165363 1019392
rect 165593 1019322 165649 1020322
rect 165665 1019322 165721 1020322
rect 166023 1020300 166223 1020322
rect 166238 1020310 166272 1020334
rect 167026 1020322 167060 1020334
rect 166283 1020310 166355 1020322
rect 166238 1020300 166355 1020310
rect 166010 1020276 166355 1020300
rect 166023 1020232 166223 1020276
rect 166238 1020266 166262 1020276
rect 166238 1020242 166272 1020266
rect 166283 1020242 166355 1020276
rect 166238 1020232 166355 1020242
rect 166010 1020208 166355 1020232
rect 166023 1020164 166223 1020208
rect 166238 1020198 166262 1020208
rect 166238 1020174 166272 1020198
rect 166283 1020174 166355 1020208
rect 166238 1020164 166355 1020174
rect 166010 1020140 166355 1020164
rect 166023 1020096 166223 1020140
rect 166238 1020130 166262 1020140
rect 166238 1020106 166272 1020130
rect 166283 1020106 166355 1020140
rect 166238 1020096 166355 1020106
rect 166010 1020072 166355 1020096
rect 166023 1020028 166223 1020072
rect 166238 1020062 166262 1020072
rect 166238 1020038 166272 1020062
rect 166283 1020038 166355 1020072
rect 166238 1020028 166355 1020038
rect 166010 1020004 166355 1020028
rect 166023 1019960 166223 1020004
rect 166238 1019994 166262 1020004
rect 166238 1019970 166272 1019994
rect 166283 1019970 166355 1020004
rect 166238 1019960 166355 1019970
rect 166010 1019936 166355 1019960
rect 166023 1019892 166223 1019936
rect 166238 1019926 166262 1019936
rect 166238 1019902 166272 1019926
rect 166283 1019902 166355 1019936
rect 166238 1019892 166355 1019902
rect 166010 1019868 166355 1019892
rect 166023 1019824 166223 1019868
rect 166238 1019858 166262 1019868
rect 166238 1019834 166272 1019858
rect 166283 1019834 166355 1019868
rect 166238 1019824 166355 1019834
rect 166010 1019800 166355 1019824
rect 166023 1019756 166223 1019800
rect 166238 1019790 166262 1019800
rect 166238 1019766 166272 1019790
rect 166283 1019766 166355 1019800
rect 166238 1019756 166355 1019766
rect 166010 1019732 166355 1019756
rect 166023 1019688 166223 1019732
rect 166238 1019722 166262 1019732
rect 166238 1019698 166272 1019722
rect 166283 1019698 166355 1019732
rect 166238 1019688 166355 1019698
rect 166010 1019664 166355 1019688
rect 166023 1019620 166223 1019664
rect 166238 1019654 166262 1019664
rect 166238 1019630 166272 1019654
rect 166283 1019630 166355 1019664
rect 166238 1019620 166355 1019630
rect 166010 1019596 166355 1019620
rect 166023 1019552 166223 1019596
rect 166238 1019586 166262 1019596
rect 166238 1019562 166272 1019586
rect 166283 1019562 166355 1019596
rect 166238 1019552 166355 1019562
rect 166010 1019528 166355 1019552
rect 166023 1019484 166223 1019528
rect 166238 1019518 166262 1019528
rect 166238 1019494 166272 1019518
rect 166283 1019494 166355 1019528
rect 166238 1019484 166355 1019494
rect 166010 1019460 166355 1019484
rect 166023 1019416 166223 1019460
rect 166238 1019450 166262 1019460
rect 166238 1019426 166272 1019450
rect 166283 1019426 166355 1019460
rect 166238 1019416 166355 1019426
rect 166010 1019392 166355 1019416
rect 166023 1019322 166223 1019392
rect 166238 1019368 166262 1019392
rect 166283 1019322 166355 1019392
rect 166585 1019322 166641 1020322
rect 166657 1019322 166713 1020322
rect 167015 1020300 167215 1020322
rect 167230 1020310 167264 1020334
rect 168018 1020322 168052 1020334
rect 167275 1020310 167347 1020322
rect 167230 1020300 167347 1020310
rect 167002 1020276 167347 1020300
rect 167015 1020232 167215 1020276
rect 167230 1020266 167254 1020276
rect 167230 1020242 167264 1020266
rect 167275 1020242 167347 1020276
rect 167230 1020232 167347 1020242
rect 167002 1020208 167347 1020232
rect 167015 1020164 167215 1020208
rect 167230 1020198 167254 1020208
rect 167230 1020174 167264 1020198
rect 167275 1020174 167347 1020208
rect 167230 1020164 167347 1020174
rect 167002 1020140 167347 1020164
rect 167015 1020096 167215 1020140
rect 167230 1020130 167254 1020140
rect 167230 1020106 167264 1020130
rect 167275 1020106 167347 1020140
rect 167230 1020096 167347 1020106
rect 167002 1020072 167347 1020096
rect 167015 1020028 167215 1020072
rect 167230 1020062 167254 1020072
rect 167230 1020038 167264 1020062
rect 167275 1020038 167347 1020072
rect 167230 1020028 167347 1020038
rect 167002 1020004 167347 1020028
rect 167015 1019960 167215 1020004
rect 167230 1019994 167254 1020004
rect 167230 1019970 167264 1019994
rect 167275 1019970 167347 1020004
rect 167230 1019960 167347 1019970
rect 167002 1019936 167347 1019960
rect 167015 1019892 167215 1019936
rect 167230 1019926 167254 1019936
rect 167230 1019902 167264 1019926
rect 167275 1019902 167347 1019936
rect 167230 1019892 167347 1019902
rect 167002 1019868 167347 1019892
rect 167015 1019824 167215 1019868
rect 167230 1019858 167254 1019868
rect 167230 1019834 167264 1019858
rect 167275 1019834 167347 1019868
rect 167230 1019824 167347 1019834
rect 167002 1019800 167347 1019824
rect 167015 1019756 167215 1019800
rect 167230 1019790 167254 1019800
rect 167230 1019766 167264 1019790
rect 167275 1019766 167347 1019800
rect 167230 1019756 167347 1019766
rect 167002 1019732 167347 1019756
rect 167015 1019688 167215 1019732
rect 167230 1019722 167254 1019732
rect 167230 1019698 167264 1019722
rect 167275 1019698 167347 1019732
rect 167230 1019688 167347 1019698
rect 167002 1019664 167347 1019688
rect 167015 1019620 167215 1019664
rect 167230 1019654 167254 1019664
rect 167230 1019630 167264 1019654
rect 167275 1019630 167347 1019664
rect 167230 1019620 167347 1019630
rect 167002 1019596 167347 1019620
rect 167015 1019552 167215 1019596
rect 167230 1019586 167254 1019596
rect 167230 1019562 167264 1019586
rect 167275 1019562 167347 1019596
rect 167230 1019552 167347 1019562
rect 167002 1019528 167347 1019552
rect 167015 1019484 167215 1019528
rect 167230 1019518 167254 1019528
rect 167230 1019494 167264 1019518
rect 167275 1019494 167347 1019528
rect 167230 1019484 167347 1019494
rect 167002 1019460 167347 1019484
rect 167015 1019416 167215 1019460
rect 167230 1019450 167254 1019460
rect 167230 1019426 167264 1019450
rect 167275 1019426 167347 1019460
rect 167230 1019416 167347 1019426
rect 167002 1019392 167347 1019416
rect 167015 1019322 167215 1019392
rect 167230 1019368 167254 1019392
rect 167275 1019322 167347 1019392
rect 167577 1019322 167633 1020322
rect 167649 1019322 167705 1020322
rect 168007 1020300 168207 1020322
rect 168222 1020310 168256 1020334
rect 169010 1020322 169044 1020334
rect 168267 1020310 168339 1020322
rect 168222 1020300 168339 1020310
rect 167994 1020276 168339 1020300
rect 168007 1020232 168207 1020276
rect 168222 1020266 168246 1020276
rect 168222 1020242 168256 1020266
rect 168267 1020242 168339 1020276
rect 168222 1020232 168339 1020242
rect 167994 1020208 168339 1020232
rect 168007 1020164 168207 1020208
rect 168222 1020198 168246 1020208
rect 168222 1020174 168256 1020198
rect 168267 1020174 168339 1020208
rect 168222 1020164 168339 1020174
rect 167994 1020140 168339 1020164
rect 168007 1020096 168207 1020140
rect 168222 1020130 168246 1020140
rect 168222 1020106 168256 1020130
rect 168267 1020106 168339 1020140
rect 168222 1020096 168339 1020106
rect 167994 1020072 168339 1020096
rect 168007 1020028 168207 1020072
rect 168222 1020062 168246 1020072
rect 168222 1020038 168256 1020062
rect 168267 1020038 168339 1020072
rect 168222 1020028 168339 1020038
rect 167994 1020004 168339 1020028
rect 168007 1019960 168207 1020004
rect 168222 1019994 168246 1020004
rect 168222 1019970 168256 1019994
rect 168267 1019970 168339 1020004
rect 168222 1019960 168339 1019970
rect 167994 1019936 168339 1019960
rect 168007 1019892 168207 1019936
rect 168222 1019926 168246 1019936
rect 168222 1019902 168256 1019926
rect 168267 1019902 168339 1019936
rect 168222 1019892 168339 1019902
rect 167994 1019868 168339 1019892
rect 168007 1019824 168207 1019868
rect 168222 1019858 168246 1019868
rect 168222 1019834 168256 1019858
rect 168267 1019834 168339 1019868
rect 168222 1019824 168339 1019834
rect 167994 1019800 168339 1019824
rect 168007 1019756 168207 1019800
rect 168222 1019790 168246 1019800
rect 168222 1019766 168256 1019790
rect 168267 1019766 168339 1019800
rect 168222 1019756 168339 1019766
rect 167994 1019732 168339 1019756
rect 168007 1019688 168207 1019732
rect 168222 1019722 168246 1019732
rect 168222 1019698 168256 1019722
rect 168267 1019698 168339 1019732
rect 168222 1019688 168339 1019698
rect 167994 1019664 168339 1019688
rect 168007 1019620 168207 1019664
rect 168222 1019654 168246 1019664
rect 168222 1019630 168256 1019654
rect 168267 1019630 168339 1019664
rect 168222 1019620 168339 1019630
rect 167994 1019596 168339 1019620
rect 168007 1019552 168207 1019596
rect 168222 1019586 168246 1019596
rect 168222 1019562 168256 1019586
rect 168267 1019562 168339 1019596
rect 168222 1019552 168339 1019562
rect 167994 1019528 168339 1019552
rect 168007 1019484 168207 1019528
rect 168222 1019518 168246 1019528
rect 168222 1019494 168256 1019518
rect 168267 1019494 168339 1019528
rect 168222 1019484 168339 1019494
rect 167994 1019460 168339 1019484
rect 168007 1019416 168207 1019460
rect 168222 1019450 168246 1019460
rect 168222 1019426 168256 1019450
rect 168267 1019426 168339 1019460
rect 168222 1019416 168339 1019426
rect 167994 1019392 168339 1019416
rect 168007 1019322 168207 1019392
rect 168222 1019368 168246 1019392
rect 168267 1019322 168339 1019392
rect 168569 1019322 168625 1020322
rect 168641 1019322 168697 1020322
rect 168999 1020300 169199 1020322
rect 169214 1020310 169248 1020334
rect 170002 1020322 170036 1020334
rect 169259 1020310 169331 1020322
rect 169214 1020300 169331 1020310
rect 168986 1020276 169331 1020300
rect 168999 1020232 169199 1020276
rect 169214 1020266 169238 1020276
rect 169214 1020242 169248 1020266
rect 169259 1020242 169331 1020276
rect 169214 1020232 169331 1020242
rect 168986 1020208 169331 1020232
rect 168999 1020164 169199 1020208
rect 169214 1020198 169238 1020208
rect 169214 1020174 169248 1020198
rect 169259 1020174 169331 1020208
rect 169214 1020164 169331 1020174
rect 168986 1020140 169331 1020164
rect 168999 1020096 169199 1020140
rect 169214 1020130 169238 1020140
rect 169214 1020106 169248 1020130
rect 169259 1020106 169331 1020140
rect 169214 1020096 169331 1020106
rect 168986 1020072 169331 1020096
rect 168999 1020028 169199 1020072
rect 169214 1020062 169238 1020072
rect 169214 1020038 169248 1020062
rect 169259 1020038 169331 1020072
rect 169214 1020028 169331 1020038
rect 168986 1020004 169331 1020028
rect 168999 1019960 169199 1020004
rect 169214 1019994 169238 1020004
rect 169214 1019970 169248 1019994
rect 169259 1019970 169331 1020004
rect 169214 1019960 169331 1019970
rect 168986 1019936 169331 1019960
rect 168999 1019892 169199 1019936
rect 169214 1019926 169238 1019936
rect 169214 1019902 169248 1019926
rect 169259 1019902 169331 1019936
rect 169214 1019892 169331 1019902
rect 168986 1019868 169331 1019892
rect 168999 1019824 169199 1019868
rect 169214 1019858 169238 1019868
rect 169214 1019834 169248 1019858
rect 169259 1019834 169331 1019868
rect 169214 1019824 169331 1019834
rect 168986 1019800 169331 1019824
rect 168999 1019756 169199 1019800
rect 169214 1019790 169238 1019800
rect 169214 1019766 169248 1019790
rect 169259 1019766 169331 1019800
rect 169214 1019756 169331 1019766
rect 168986 1019732 169331 1019756
rect 168999 1019688 169199 1019732
rect 169214 1019722 169238 1019732
rect 169214 1019698 169248 1019722
rect 169259 1019698 169331 1019732
rect 169214 1019688 169331 1019698
rect 168986 1019664 169331 1019688
rect 168999 1019620 169199 1019664
rect 169214 1019654 169238 1019664
rect 169214 1019630 169248 1019654
rect 169259 1019630 169331 1019664
rect 169214 1019620 169331 1019630
rect 168986 1019596 169331 1019620
rect 168999 1019552 169199 1019596
rect 169214 1019586 169238 1019596
rect 169214 1019562 169248 1019586
rect 169259 1019562 169331 1019596
rect 169214 1019552 169331 1019562
rect 168986 1019528 169331 1019552
rect 168999 1019484 169199 1019528
rect 169214 1019518 169238 1019528
rect 169214 1019494 169248 1019518
rect 169259 1019494 169331 1019528
rect 169214 1019484 169331 1019494
rect 168986 1019460 169331 1019484
rect 168999 1019416 169199 1019460
rect 169214 1019450 169238 1019460
rect 169214 1019426 169248 1019450
rect 169259 1019426 169331 1019460
rect 169214 1019416 169331 1019426
rect 168986 1019392 169331 1019416
rect 168999 1019322 169199 1019392
rect 169214 1019368 169238 1019392
rect 169259 1019322 169331 1019392
rect 169561 1019322 169617 1020322
rect 169633 1019322 169689 1020322
rect 169991 1020300 170191 1020322
rect 170206 1020310 170240 1020334
rect 170994 1020322 171028 1020334
rect 170251 1020310 170323 1020322
rect 170206 1020300 170323 1020310
rect 169978 1020276 170323 1020300
rect 169991 1020232 170191 1020276
rect 170206 1020266 170230 1020276
rect 170206 1020242 170240 1020266
rect 170251 1020242 170323 1020276
rect 170206 1020232 170323 1020242
rect 169978 1020208 170323 1020232
rect 169991 1020164 170191 1020208
rect 170206 1020198 170230 1020208
rect 170206 1020174 170240 1020198
rect 170251 1020174 170323 1020208
rect 170206 1020164 170323 1020174
rect 169978 1020140 170323 1020164
rect 169991 1020096 170191 1020140
rect 170206 1020130 170230 1020140
rect 170206 1020106 170240 1020130
rect 170251 1020106 170323 1020140
rect 170206 1020096 170323 1020106
rect 169978 1020072 170323 1020096
rect 169991 1020028 170191 1020072
rect 170206 1020062 170230 1020072
rect 170206 1020038 170240 1020062
rect 170251 1020038 170323 1020072
rect 170206 1020028 170323 1020038
rect 169978 1020004 170323 1020028
rect 169991 1019960 170191 1020004
rect 170206 1019994 170230 1020004
rect 170206 1019970 170240 1019994
rect 170251 1019970 170323 1020004
rect 170206 1019960 170323 1019970
rect 169978 1019936 170323 1019960
rect 169991 1019892 170191 1019936
rect 170206 1019926 170230 1019936
rect 170206 1019902 170240 1019926
rect 170251 1019902 170323 1019936
rect 170206 1019892 170323 1019902
rect 169978 1019868 170323 1019892
rect 169991 1019824 170191 1019868
rect 170206 1019858 170230 1019868
rect 170206 1019834 170240 1019858
rect 170251 1019834 170323 1019868
rect 170206 1019824 170323 1019834
rect 169978 1019800 170323 1019824
rect 169991 1019756 170191 1019800
rect 170206 1019790 170230 1019800
rect 170206 1019766 170240 1019790
rect 170251 1019766 170323 1019800
rect 170206 1019756 170323 1019766
rect 169978 1019732 170323 1019756
rect 169991 1019688 170191 1019732
rect 170206 1019722 170230 1019732
rect 170206 1019698 170240 1019722
rect 170251 1019698 170323 1019732
rect 170206 1019688 170323 1019698
rect 169978 1019664 170323 1019688
rect 169991 1019620 170191 1019664
rect 170206 1019654 170230 1019664
rect 170206 1019630 170240 1019654
rect 170251 1019630 170323 1019664
rect 170206 1019620 170323 1019630
rect 169978 1019596 170323 1019620
rect 169991 1019552 170191 1019596
rect 170206 1019586 170230 1019596
rect 170206 1019562 170240 1019586
rect 170251 1019562 170323 1019596
rect 170206 1019552 170323 1019562
rect 169978 1019528 170323 1019552
rect 169991 1019484 170191 1019528
rect 170206 1019518 170230 1019528
rect 170206 1019494 170240 1019518
rect 170251 1019494 170323 1019528
rect 170206 1019484 170323 1019494
rect 169978 1019460 170323 1019484
rect 169991 1019416 170191 1019460
rect 170206 1019450 170230 1019460
rect 170206 1019426 170240 1019450
rect 170251 1019426 170323 1019460
rect 170206 1019416 170323 1019426
rect 169978 1019392 170323 1019416
rect 169991 1019322 170191 1019392
rect 170206 1019368 170230 1019392
rect 170251 1019322 170323 1019392
rect 170553 1019322 170609 1020322
rect 170625 1019322 170681 1020322
rect 170983 1020300 171183 1020322
rect 171198 1020310 171232 1020334
rect 171986 1020322 172020 1020334
rect 171243 1020310 171315 1020322
rect 171198 1020300 171315 1020310
rect 170970 1020276 171315 1020300
rect 170983 1020232 171183 1020276
rect 171198 1020266 171222 1020276
rect 171198 1020242 171232 1020266
rect 171243 1020242 171315 1020276
rect 171198 1020232 171315 1020242
rect 170970 1020208 171315 1020232
rect 170983 1020164 171183 1020208
rect 171198 1020198 171222 1020208
rect 171198 1020174 171232 1020198
rect 171243 1020174 171315 1020208
rect 171198 1020164 171315 1020174
rect 170970 1020140 171315 1020164
rect 170983 1020096 171183 1020140
rect 171198 1020130 171222 1020140
rect 171198 1020106 171232 1020130
rect 171243 1020106 171315 1020140
rect 171198 1020096 171315 1020106
rect 170970 1020072 171315 1020096
rect 170983 1020028 171183 1020072
rect 171198 1020062 171222 1020072
rect 171198 1020038 171232 1020062
rect 171243 1020038 171315 1020072
rect 171198 1020028 171315 1020038
rect 170970 1020004 171315 1020028
rect 170983 1019960 171183 1020004
rect 171198 1019994 171222 1020004
rect 171198 1019970 171232 1019994
rect 171243 1019970 171315 1020004
rect 171198 1019960 171315 1019970
rect 170970 1019936 171315 1019960
rect 170983 1019892 171183 1019936
rect 171198 1019926 171222 1019936
rect 171198 1019902 171232 1019926
rect 171243 1019902 171315 1019936
rect 171198 1019892 171315 1019902
rect 170970 1019868 171315 1019892
rect 170983 1019824 171183 1019868
rect 171198 1019858 171222 1019868
rect 171198 1019834 171232 1019858
rect 171243 1019834 171315 1019868
rect 171198 1019824 171315 1019834
rect 170970 1019800 171315 1019824
rect 170983 1019756 171183 1019800
rect 171198 1019790 171222 1019800
rect 171198 1019766 171232 1019790
rect 171243 1019766 171315 1019800
rect 171198 1019756 171315 1019766
rect 170970 1019732 171315 1019756
rect 170983 1019688 171183 1019732
rect 171198 1019722 171222 1019732
rect 171198 1019698 171232 1019722
rect 171243 1019698 171315 1019732
rect 171198 1019688 171315 1019698
rect 170970 1019664 171315 1019688
rect 170983 1019620 171183 1019664
rect 171198 1019654 171222 1019664
rect 171198 1019630 171232 1019654
rect 171243 1019630 171315 1019664
rect 171198 1019620 171315 1019630
rect 170970 1019596 171315 1019620
rect 170983 1019552 171183 1019596
rect 171198 1019586 171222 1019596
rect 171198 1019562 171232 1019586
rect 171243 1019562 171315 1019596
rect 171198 1019552 171315 1019562
rect 170970 1019528 171315 1019552
rect 170983 1019484 171183 1019528
rect 171198 1019518 171222 1019528
rect 171198 1019494 171232 1019518
rect 171243 1019494 171315 1019528
rect 171198 1019484 171315 1019494
rect 170970 1019460 171315 1019484
rect 170983 1019416 171183 1019460
rect 171198 1019450 171222 1019460
rect 171198 1019426 171232 1019450
rect 171243 1019426 171315 1019460
rect 171198 1019416 171315 1019426
rect 170970 1019392 171315 1019416
rect 170983 1019322 171183 1019392
rect 171198 1019368 171222 1019392
rect 171243 1019322 171315 1019392
rect 171545 1019322 171601 1020322
rect 171617 1019322 171673 1020322
rect 171975 1020300 172175 1020322
rect 172190 1020310 172224 1020334
rect 172978 1020322 173012 1020334
rect 172235 1020310 172307 1020322
rect 172190 1020300 172307 1020310
rect 171962 1020276 172307 1020300
rect 171975 1020232 172175 1020276
rect 172190 1020266 172214 1020276
rect 172190 1020242 172224 1020266
rect 172235 1020242 172307 1020276
rect 172190 1020232 172307 1020242
rect 171962 1020208 172307 1020232
rect 171975 1020164 172175 1020208
rect 172190 1020198 172214 1020208
rect 172190 1020174 172224 1020198
rect 172235 1020174 172307 1020208
rect 172190 1020164 172307 1020174
rect 171962 1020140 172307 1020164
rect 171975 1020096 172175 1020140
rect 172190 1020130 172214 1020140
rect 172190 1020106 172224 1020130
rect 172235 1020106 172307 1020140
rect 172190 1020096 172307 1020106
rect 171962 1020072 172307 1020096
rect 171975 1020028 172175 1020072
rect 172190 1020062 172214 1020072
rect 172190 1020038 172224 1020062
rect 172235 1020038 172307 1020072
rect 172190 1020028 172307 1020038
rect 171962 1020004 172307 1020028
rect 171975 1019960 172175 1020004
rect 172190 1019994 172214 1020004
rect 172190 1019970 172224 1019994
rect 172235 1019970 172307 1020004
rect 172190 1019960 172307 1019970
rect 171962 1019936 172307 1019960
rect 171975 1019892 172175 1019936
rect 172190 1019926 172214 1019936
rect 172190 1019902 172224 1019926
rect 172235 1019902 172307 1019936
rect 172190 1019892 172307 1019902
rect 171962 1019868 172307 1019892
rect 171975 1019824 172175 1019868
rect 172190 1019858 172214 1019868
rect 172190 1019834 172224 1019858
rect 172235 1019834 172307 1019868
rect 172190 1019824 172307 1019834
rect 171962 1019800 172307 1019824
rect 171975 1019756 172175 1019800
rect 172190 1019790 172214 1019800
rect 172190 1019766 172224 1019790
rect 172235 1019766 172307 1019800
rect 172190 1019756 172307 1019766
rect 171962 1019732 172307 1019756
rect 171975 1019688 172175 1019732
rect 172190 1019722 172214 1019732
rect 172190 1019698 172224 1019722
rect 172235 1019698 172307 1019732
rect 172190 1019688 172307 1019698
rect 171962 1019664 172307 1019688
rect 171975 1019620 172175 1019664
rect 172190 1019654 172214 1019664
rect 172190 1019630 172224 1019654
rect 172235 1019630 172307 1019664
rect 172190 1019620 172307 1019630
rect 171962 1019596 172307 1019620
rect 171975 1019552 172175 1019596
rect 172190 1019586 172214 1019596
rect 172190 1019562 172224 1019586
rect 172235 1019562 172307 1019596
rect 172190 1019552 172307 1019562
rect 171962 1019528 172307 1019552
rect 171975 1019484 172175 1019528
rect 172190 1019518 172214 1019528
rect 172190 1019494 172224 1019518
rect 172235 1019494 172307 1019528
rect 172190 1019484 172307 1019494
rect 171962 1019460 172307 1019484
rect 171975 1019416 172175 1019460
rect 172190 1019450 172214 1019460
rect 172190 1019426 172224 1019450
rect 172235 1019426 172307 1019460
rect 172190 1019416 172307 1019426
rect 171962 1019392 172307 1019416
rect 171975 1019322 172175 1019392
rect 172190 1019368 172214 1019392
rect 172235 1019322 172307 1019392
rect 172537 1019322 172593 1020322
rect 172609 1019322 172665 1020322
rect 172967 1020300 173167 1020322
rect 173182 1020310 173216 1020334
rect 173970 1020322 174004 1020334
rect 173227 1020310 173299 1020322
rect 173182 1020300 173299 1020310
rect 172954 1020276 173299 1020300
rect 172967 1020232 173167 1020276
rect 173182 1020266 173206 1020276
rect 173182 1020242 173216 1020266
rect 173227 1020242 173299 1020276
rect 173182 1020232 173299 1020242
rect 172954 1020208 173299 1020232
rect 172967 1020164 173167 1020208
rect 173182 1020198 173206 1020208
rect 173182 1020174 173216 1020198
rect 173227 1020174 173299 1020208
rect 173182 1020164 173299 1020174
rect 172954 1020140 173299 1020164
rect 172967 1020096 173167 1020140
rect 173182 1020130 173206 1020140
rect 173182 1020106 173216 1020130
rect 173227 1020106 173299 1020140
rect 173182 1020096 173299 1020106
rect 172954 1020072 173299 1020096
rect 172967 1020028 173167 1020072
rect 173182 1020062 173206 1020072
rect 173182 1020038 173216 1020062
rect 173227 1020038 173299 1020072
rect 173182 1020028 173299 1020038
rect 172954 1020004 173299 1020028
rect 172967 1019960 173167 1020004
rect 173182 1019994 173206 1020004
rect 173182 1019970 173216 1019994
rect 173227 1019970 173299 1020004
rect 173182 1019960 173299 1019970
rect 172954 1019936 173299 1019960
rect 172967 1019892 173167 1019936
rect 173182 1019926 173206 1019936
rect 173182 1019902 173216 1019926
rect 173227 1019902 173299 1019936
rect 173182 1019892 173299 1019902
rect 172954 1019868 173299 1019892
rect 172967 1019824 173167 1019868
rect 173182 1019858 173206 1019868
rect 173182 1019834 173216 1019858
rect 173227 1019834 173299 1019868
rect 173182 1019824 173299 1019834
rect 172954 1019800 173299 1019824
rect 172967 1019756 173167 1019800
rect 173182 1019790 173206 1019800
rect 173182 1019766 173216 1019790
rect 173227 1019766 173299 1019800
rect 173182 1019756 173299 1019766
rect 172954 1019732 173299 1019756
rect 172967 1019688 173167 1019732
rect 173182 1019722 173206 1019732
rect 173182 1019698 173216 1019722
rect 173227 1019698 173299 1019732
rect 173182 1019688 173299 1019698
rect 172954 1019664 173299 1019688
rect 172967 1019620 173167 1019664
rect 173182 1019654 173206 1019664
rect 173182 1019630 173216 1019654
rect 173227 1019630 173299 1019664
rect 173182 1019620 173299 1019630
rect 172954 1019596 173299 1019620
rect 172967 1019552 173167 1019596
rect 173182 1019586 173206 1019596
rect 173182 1019562 173216 1019586
rect 173227 1019562 173299 1019596
rect 173182 1019552 173299 1019562
rect 172954 1019528 173299 1019552
rect 172967 1019484 173167 1019528
rect 173182 1019518 173206 1019528
rect 173182 1019494 173216 1019518
rect 173227 1019494 173299 1019528
rect 173182 1019484 173299 1019494
rect 172954 1019460 173299 1019484
rect 172967 1019416 173167 1019460
rect 173182 1019450 173206 1019460
rect 173182 1019426 173216 1019450
rect 173227 1019426 173299 1019460
rect 173182 1019416 173299 1019426
rect 172954 1019392 173299 1019416
rect 172967 1019322 173167 1019392
rect 173182 1019368 173206 1019392
rect 173227 1019322 173299 1019392
rect 173529 1019322 173585 1020322
rect 173601 1019322 173657 1020322
rect 173959 1020300 174159 1020322
rect 174174 1020310 174208 1020334
rect 174962 1020322 174996 1020334
rect 174219 1020310 174291 1020322
rect 174174 1020300 174291 1020310
rect 173946 1020276 174291 1020300
rect 173959 1020232 174159 1020276
rect 174174 1020266 174198 1020276
rect 174174 1020242 174208 1020266
rect 174219 1020242 174291 1020276
rect 174174 1020232 174291 1020242
rect 173946 1020208 174291 1020232
rect 173959 1020164 174159 1020208
rect 174174 1020198 174198 1020208
rect 174174 1020174 174208 1020198
rect 174219 1020174 174291 1020208
rect 174174 1020164 174291 1020174
rect 173946 1020140 174291 1020164
rect 173959 1020096 174159 1020140
rect 174174 1020130 174198 1020140
rect 174174 1020106 174208 1020130
rect 174219 1020106 174291 1020140
rect 174174 1020096 174291 1020106
rect 173946 1020072 174291 1020096
rect 173959 1020028 174159 1020072
rect 174174 1020062 174198 1020072
rect 174174 1020038 174208 1020062
rect 174219 1020038 174291 1020072
rect 174174 1020028 174291 1020038
rect 173946 1020004 174291 1020028
rect 173959 1019960 174159 1020004
rect 174174 1019994 174198 1020004
rect 174174 1019970 174208 1019994
rect 174219 1019970 174291 1020004
rect 174174 1019960 174291 1019970
rect 173946 1019936 174291 1019960
rect 173959 1019892 174159 1019936
rect 174174 1019926 174198 1019936
rect 174174 1019902 174208 1019926
rect 174219 1019902 174291 1019936
rect 174174 1019892 174291 1019902
rect 173946 1019868 174291 1019892
rect 173959 1019824 174159 1019868
rect 174174 1019858 174198 1019868
rect 174174 1019834 174208 1019858
rect 174219 1019834 174291 1019868
rect 174174 1019824 174291 1019834
rect 173946 1019800 174291 1019824
rect 173959 1019756 174159 1019800
rect 174174 1019790 174198 1019800
rect 174174 1019766 174208 1019790
rect 174219 1019766 174291 1019800
rect 174174 1019756 174291 1019766
rect 173946 1019732 174291 1019756
rect 173959 1019688 174159 1019732
rect 174174 1019722 174198 1019732
rect 174174 1019698 174208 1019722
rect 174219 1019698 174291 1019732
rect 174174 1019688 174291 1019698
rect 173946 1019664 174291 1019688
rect 173959 1019620 174159 1019664
rect 174174 1019654 174198 1019664
rect 174174 1019630 174208 1019654
rect 174219 1019630 174291 1019664
rect 174174 1019620 174291 1019630
rect 173946 1019596 174291 1019620
rect 173959 1019552 174159 1019596
rect 174174 1019586 174198 1019596
rect 174174 1019562 174208 1019586
rect 174219 1019562 174291 1019596
rect 174174 1019552 174291 1019562
rect 173946 1019528 174291 1019552
rect 173959 1019484 174159 1019528
rect 174174 1019518 174198 1019528
rect 174174 1019494 174208 1019518
rect 174219 1019494 174291 1019528
rect 174174 1019484 174291 1019494
rect 173946 1019460 174291 1019484
rect 173959 1019416 174159 1019460
rect 174174 1019450 174198 1019460
rect 174174 1019426 174208 1019450
rect 174219 1019426 174291 1019460
rect 174174 1019416 174291 1019426
rect 173946 1019392 174291 1019416
rect 173959 1019322 174159 1019392
rect 174174 1019368 174198 1019392
rect 174219 1019322 174291 1019392
rect 174521 1019322 174577 1020322
rect 174593 1019322 174649 1020322
rect 174951 1020300 175151 1020322
rect 175166 1020310 175200 1020334
rect 175211 1020310 175283 1020322
rect 175166 1020300 175283 1020310
rect 174938 1020276 175283 1020300
rect 174951 1020232 175151 1020276
rect 175166 1020266 175190 1020276
rect 175166 1020242 175200 1020266
rect 175211 1020242 175283 1020276
rect 175166 1020232 175283 1020242
rect 174938 1020208 175283 1020232
rect 174951 1020164 175151 1020208
rect 175166 1020198 175190 1020208
rect 175166 1020174 175200 1020198
rect 175211 1020174 175283 1020208
rect 175166 1020164 175283 1020174
rect 174938 1020140 175283 1020164
rect 174951 1020096 175151 1020140
rect 175166 1020130 175190 1020140
rect 175166 1020106 175200 1020130
rect 175211 1020106 175283 1020140
rect 175166 1020096 175283 1020106
rect 174938 1020072 175283 1020096
rect 174951 1020028 175151 1020072
rect 175166 1020062 175190 1020072
rect 175166 1020038 175200 1020062
rect 175211 1020038 175283 1020072
rect 175166 1020028 175283 1020038
rect 174938 1020004 175283 1020028
rect 174951 1019960 175151 1020004
rect 175166 1019994 175190 1020004
rect 175166 1019970 175200 1019994
rect 175211 1019970 175283 1020004
rect 175166 1019960 175283 1019970
rect 174938 1019936 175283 1019960
rect 174951 1019892 175151 1019936
rect 175166 1019926 175190 1019936
rect 175166 1019902 175200 1019926
rect 175211 1019902 175283 1019936
rect 175166 1019892 175283 1019902
rect 174938 1019868 175283 1019892
rect 174951 1019824 175151 1019868
rect 175166 1019858 175190 1019868
rect 175166 1019834 175200 1019858
rect 175211 1019834 175283 1019868
rect 175166 1019824 175283 1019834
rect 174938 1019800 175283 1019824
rect 174951 1019756 175151 1019800
rect 175166 1019790 175190 1019800
rect 175166 1019766 175200 1019790
rect 175211 1019766 175283 1019800
rect 175166 1019756 175283 1019766
rect 174938 1019732 175283 1019756
rect 174951 1019688 175151 1019732
rect 175166 1019722 175190 1019732
rect 175166 1019698 175200 1019722
rect 175211 1019698 175283 1019732
rect 175166 1019688 175283 1019698
rect 174938 1019664 175283 1019688
rect 174951 1019620 175151 1019664
rect 175166 1019654 175190 1019664
rect 175166 1019630 175200 1019654
rect 175211 1019630 175283 1019664
rect 175166 1019620 175283 1019630
rect 174938 1019596 175283 1019620
rect 174951 1019552 175151 1019596
rect 175166 1019586 175190 1019596
rect 175166 1019562 175200 1019586
rect 175211 1019562 175283 1019596
rect 175166 1019552 175283 1019562
rect 174938 1019528 175283 1019552
rect 174951 1019484 175151 1019528
rect 175166 1019518 175190 1019528
rect 175166 1019494 175200 1019518
rect 175211 1019494 175283 1019528
rect 175166 1019484 175283 1019494
rect 174938 1019460 175283 1019484
rect 174951 1019416 175151 1019460
rect 175166 1019450 175190 1019460
rect 175166 1019426 175200 1019450
rect 175211 1019426 175283 1019460
rect 175166 1019416 175283 1019426
rect 174938 1019392 175283 1019416
rect 174951 1019322 175151 1019392
rect 175166 1019368 175190 1019392
rect 175211 1019322 175283 1019392
rect 175472 1019322 175544 1020322
rect 175610 1019322 175627 1020322
rect 175797 1019322 175830 1020322
rect 213561 1018210 213668 1022756
rect 214356 1020922 214406 1021922
rect 214617 1020922 214673 1021922
rect 214689 1020922 214745 1021922
rect 215107 1020922 215247 1021922
rect 226521 1020922 226577 1021922
rect 226593 1020922 226649 1021922
rect 227011 1020922 227151 1021922
rect 227473 1020922 227544 1021922
rect 227610 1020922 227627 1021922
rect 227797 1020922 227830 1021922
rect 227953 1021730 228025 1021760
rect 227953 1021692 227987 1021722
rect 214356 1019322 214406 1020322
rect 214617 1019322 214673 1020322
rect 214689 1019322 214745 1020322
rect 215107 1019322 215247 1020322
rect 226521 1019322 226577 1020322
rect 226593 1019322 226649 1020322
rect 227011 1019322 227151 1020322
rect 227473 1019322 227544 1020322
rect 227610 1019322 227627 1020322
rect 227797 1019322 227830 1020322
rect 261561 1018210 261668 1022756
rect 274521 1020922 274577 1021922
rect 274593 1020922 274649 1021922
rect 275011 1020922 275151 1021922
rect 275473 1020922 275544 1021922
rect 275610 1020922 275627 1021922
rect 275797 1020922 275830 1021922
rect 275953 1021730 276025 1021760
rect 275953 1021692 275987 1021722
rect 274521 1019322 274577 1020322
rect 274593 1019322 274649 1020322
rect 275011 1019322 275151 1020322
rect 275473 1019322 275544 1020322
rect 275610 1019322 275627 1020322
rect 275797 1019322 275830 1020322
rect 313561 1018210 313668 1022756
rect 314356 1020922 314406 1021922
rect 314617 1020922 314673 1021922
rect 314689 1020922 314745 1021922
rect 315107 1020922 315247 1021922
rect 326521 1020922 326577 1021922
rect 326593 1020922 326649 1021922
rect 327011 1020922 327151 1021922
rect 327473 1020922 327544 1021922
rect 327610 1020922 327627 1021922
rect 327797 1020922 327830 1021922
rect 327953 1021730 328025 1021760
rect 327953 1021692 327987 1021722
rect 314356 1019322 314406 1020322
rect 314617 1019322 314673 1020322
rect 314689 1019322 314745 1020322
rect 315107 1019322 315247 1020322
rect 326521 1019322 326577 1020322
rect 326593 1019322 326649 1020322
rect 327011 1019322 327151 1020322
rect 327473 1019322 327544 1020322
rect 327610 1019322 327627 1020322
rect 327797 1019322 327830 1020322
rect 365561 1018210 365668 1022756
rect 366356 1020922 366406 1021922
rect 366617 1020922 366673 1021922
rect 366689 1020922 366745 1021922
rect 367047 1021842 367247 1021922
rect 367262 1021852 367296 1021876
rect 367307 1021852 367379 1021922
rect 367262 1021842 367379 1021852
rect 367034 1021818 367379 1021842
rect 367047 1021774 367247 1021818
rect 367262 1021808 367286 1021818
rect 367262 1021784 367296 1021808
rect 367307 1021784 367379 1021818
rect 367262 1021774 367379 1021784
rect 367034 1021750 367379 1021774
rect 367047 1021706 367247 1021750
rect 367262 1021740 367286 1021750
rect 367262 1021716 367296 1021740
rect 367307 1021716 367379 1021750
rect 367262 1021706 367379 1021716
rect 367034 1021682 367379 1021706
rect 367047 1021638 367247 1021682
rect 367262 1021672 367286 1021682
rect 367262 1021648 367296 1021672
rect 367307 1021648 367379 1021682
rect 367262 1021638 367379 1021648
rect 367034 1021614 367379 1021638
rect 367047 1021570 367247 1021614
rect 367262 1021604 367286 1021614
rect 367262 1021580 367296 1021604
rect 367307 1021580 367379 1021614
rect 367262 1021570 367379 1021580
rect 367034 1021546 367379 1021570
rect 367047 1021502 367247 1021546
rect 367262 1021536 367286 1021546
rect 367262 1021512 367296 1021536
rect 367307 1021512 367379 1021546
rect 367262 1021502 367379 1021512
rect 367034 1021478 367379 1021502
rect 367047 1021434 367247 1021478
rect 367262 1021468 367286 1021478
rect 367262 1021444 367296 1021468
rect 367307 1021444 367379 1021478
rect 367262 1021434 367379 1021444
rect 367034 1021410 367379 1021434
rect 367047 1021366 367247 1021410
rect 367262 1021400 367286 1021410
rect 367262 1021376 367296 1021400
rect 367307 1021376 367379 1021410
rect 367262 1021366 367379 1021376
rect 367034 1021342 367379 1021366
rect 367047 1021298 367247 1021342
rect 367262 1021332 367286 1021342
rect 367262 1021308 367296 1021332
rect 367307 1021308 367379 1021342
rect 367262 1021298 367379 1021308
rect 367034 1021274 367379 1021298
rect 367047 1021230 367247 1021274
rect 367262 1021264 367286 1021274
rect 367262 1021240 367296 1021264
rect 367307 1021240 367379 1021274
rect 367262 1021230 367379 1021240
rect 367034 1021206 367379 1021230
rect 367047 1021162 367247 1021206
rect 367262 1021196 367286 1021206
rect 367262 1021172 367296 1021196
rect 367307 1021172 367379 1021206
rect 367262 1021162 367379 1021172
rect 367034 1021138 367379 1021162
rect 367047 1021094 367247 1021138
rect 367262 1021128 367286 1021138
rect 367262 1021104 367296 1021128
rect 367307 1021104 367379 1021138
rect 367262 1021094 367379 1021104
rect 367034 1021070 367379 1021094
rect 367047 1021026 367247 1021070
rect 367262 1021060 367286 1021070
rect 367262 1021036 367296 1021060
rect 367307 1021036 367379 1021070
rect 367262 1021026 367379 1021036
rect 367034 1021002 367379 1021026
rect 367047 1020958 367247 1021002
rect 367262 1020992 367286 1021002
rect 367262 1020968 367296 1020992
rect 367307 1020968 367379 1021002
rect 367262 1020958 367379 1020968
rect 367034 1020934 367379 1020958
rect 367047 1020922 367247 1020934
rect 367058 1020910 367082 1020922
rect 367262 1020910 367286 1020934
rect 367307 1020922 367379 1020934
rect 367609 1020922 367665 1021922
rect 367681 1020922 367737 1021922
rect 368039 1021842 368239 1021922
rect 368254 1021852 368288 1021876
rect 368299 1021852 368371 1021922
rect 368254 1021842 368371 1021852
rect 368026 1021818 368371 1021842
rect 368039 1021774 368239 1021818
rect 368254 1021808 368278 1021818
rect 368254 1021784 368288 1021808
rect 368299 1021784 368371 1021818
rect 368254 1021774 368371 1021784
rect 368026 1021750 368371 1021774
rect 368039 1021706 368239 1021750
rect 368254 1021740 368278 1021750
rect 368254 1021716 368288 1021740
rect 368299 1021716 368371 1021750
rect 368254 1021706 368371 1021716
rect 368026 1021682 368371 1021706
rect 368039 1021638 368239 1021682
rect 368254 1021672 368278 1021682
rect 368254 1021648 368288 1021672
rect 368299 1021648 368371 1021682
rect 368254 1021638 368371 1021648
rect 368026 1021614 368371 1021638
rect 368039 1021570 368239 1021614
rect 368254 1021604 368278 1021614
rect 368254 1021580 368288 1021604
rect 368299 1021580 368371 1021614
rect 368254 1021570 368371 1021580
rect 368026 1021546 368371 1021570
rect 368039 1021502 368239 1021546
rect 368254 1021536 368278 1021546
rect 368254 1021512 368288 1021536
rect 368299 1021512 368371 1021546
rect 368254 1021502 368371 1021512
rect 368026 1021478 368371 1021502
rect 368039 1021434 368239 1021478
rect 368254 1021468 368278 1021478
rect 368254 1021444 368288 1021468
rect 368299 1021444 368371 1021478
rect 368254 1021434 368371 1021444
rect 368026 1021410 368371 1021434
rect 368039 1021366 368239 1021410
rect 368254 1021400 368278 1021410
rect 368254 1021376 368288 1021400
rect 368299 1021376 368371 1021410
rect 368254 1021366 368371 1021376
rect 368026 1021342 368371 1021366
rect 368039 1021298 368239 1021342
rect 368254 1021332 368278 1021342
rect 368254 1021308 368288 1021332
rect 368299 1021308 368371 1021342
rect 368254 1021298 368371 1021308
rect 368026 1021274 368371 1021298
rect 368039 1021230 368239 1021274
rect 368254 1021264 368278 1021274
rect 368254 1021240 368288 1021264
rect 368299 1021240 368371 1021274
rect 368254 1021230 368371 1021240
rect 368026 1021206 368371 1021230
rect 368039 1021162 368239 1021206
rect 368254 1021196 368278 1021206
rect 368254 1021172 368288 1021196
rect 368299 1021172 368371 1021206
rect 368254 1021162 368371 1021172
rect 368026 1021138 368371 1021162
rect 368039 1021094 368239 1021138
rect 368254 1021128 368278 1021138
rect 368254 1021104 368288 1021128
rect 368299 1021104 368371 1021138
rect 368254 1021094 368371 1021104
rect 368026 1021070 368371 1021094
rect 368039 1021026 368239 1021070
rect 368254 1021060 368278 1021070
rect 368254 1021036 368288 1021060
rect 368299 1021036 368371 1021070
rect 368254 1021026 368371 1021036
rect 368026 1021002 368371 1021026
rect 368039 1020958 368239 1021002
rect 368254 1020992 368278 1021002
rect 368254 1020968 368288 1020992
rect 368299 1020968 368371 1021002
rect 368254 1020958 368371 1020968
rect 368026 1020934 368371 1020958
rect 368039 1020922 368239 1020934
rect 368050 1020910 368074 1020922
rect 368254 1020910 368278 1020934
rect 368299 1020922 368371 1020934
rect 368601 1020922 368657 1021922
rect 368673 1020922 368729 1021922
rect 369031 1021842 369231 1021922
rect 369246 1021852 369280 1021876
rect 369291 1021852 369363 1021922
rect 369246 1021842 369363 1021852
rect 369018 1021818 369363 1021842
rect 369031 1021774 369231 1021818
rect 369246 1021808 369270 1021818
rect 369246 1021784 369280 1021808
rect 369291 1021784 369363 1021818
rect 369246 1021774 369363 1021784
rect 369018 1021750 369363 1021774
rect 369031 1021706 369231 1021750
rect 369246 1021740 369270 1021750
rect 369246 1021716 369280 1021740
rect 369291 1021716 369363 1021750
rect 369246 1021706 369363 1021716
rect 369018 1021682 369363 1021706
rect 369031 1021638 369231 1021682
rect 369246 1021672 369270 1021682
rect 369246 1021648 369280 1021672
rect 369291 1021648 369363 1021682
rect 369246 1021638 369363 1021648
rect 369018 1021614 369363 1021638
rect 369031 1021570 369231 1021614
rect 369246 1021604 369270 1021614
rect 369246 1021580 369280 1021604
rect 369291 1021580 369363 1021614
rect 369246 1021570 369363 1021580
rect 369018 1021546 369363 1021570
rect 369031 1021502 369231 1021546
rect 369246 1021536 369270 1021546
rect 369246 1021512 369280 1021536
rect 369291 1021512 369363 1021546
rect 369246 1021502 369363 1021512
rect 369018 1021478 369363 1021502
rect 369031 1021434 369231 1021478
rect 369246 1021468 369270 1021478
rect 369246 1021444 369280 1021468
rect 369291 1021444 369363 1021478
rect 369246 1021434 369363 1021444
rect 369018 1021410 369363 1021434
rect 369031 1021366 369231 1021410
rect 369246 1021400 369270 1021410
rect 369246 1021376 369280 1021400
rect 369291 1021376 369363 1021410
rect 369246 1021366 369363 1021376
rect 369018 1021342 369363 1021366
rect 369031 1021298 369231 1021342
rect 369246 1021332 369270 1021342
rect 369246 1021308 369280 1021332
rect 369291 1021308 369363 1021342
rect 369246 1021298 369363 1021308
rect 369018 1021274 369363 1021298
rect 369031 1021230 369231 1021274
rect 369246 1021264 369270 1021274
rect 369246 1021240 369280 1021264
rect 369291 1021240 369363 1021274
rect 369246 1021230 369363 1021240
rect 369018 1021206 369363 1021230
rect 369031 1021162 369231 1021206
rect 369246 1021196 369270 1021206
rect 369246 1021172 369280 1021196
rect 369291 1021172 369363 1021206
rect 369246 1021162 369363 1021172
rect 369018 1021138 369363 1021162
rect 369031 1021094 369231 1021138
rect 369246 1021128 369270 1021138
rect 369246 1021104 369280 1021128
rect 369291 1021104 369363 1021138
rect 369246 1021094 369363 1021104
rect 369018 1021070 369363 1021094
rect 369031 1021026 369231 1021070
rect 369246 1021060 369270 1021070
rect 369246 1021036 369280 1021060
rect 369291 1021036 369363 1021070
rect 369246 1021026 369363 1021036
rect 369018 1021002 369363 1021026
rect 369031 1020958 369231 1021002
rect 369246 1020992 369270 1021002
rect 369246 1020968 369280 1020992
rect 369291 1020968 369363 1021002
rect 369246 1020958 369363 1020968
rect 369018 1020934 369363 1020958
rect 369031 1020922 369231 1020934
rect 369042 1020910 369066 1020922
rect 369246 1020910 369270 1020934
rect 369291 1020922 369363 1020934
rect 369593 1020922 369649 1021922
rect 369665 1020922 369721 1021922
rect 370023 1021842 370223 1021922
rect 370238 1021852 370272 1021876
rect 370283 1021852 370355 1021922
rect 370238 1021842 370355 1021852
rect 370010 1021818 370355 1021842
rect 370023 1021774 370223 1021818
rect 370238 1021808 370262 1021818
rect 370238 1021784 370272 1021808
rect 370283 1021784 370355 1021818
rect 370238 1021774 370355 1021784
rect 370010 1021750 370355 1021774
rect 370023 1021706 370223 1021750
rect 370238 1021740 370262 1021750
rect 370238 1021716 370272 1021740
rect 370283 1021716 370355 1021750
rect 370238 1021706 370355 1021716
rect 370010 1021682 370355 1021706
rect 370023 1021638 370223 1021682
rect 370238 1021672 370262 1021682
rect 370238 1021648 370272 1021672
rect 370283 1021648 370355 1021682
rect 370238 1021638 370355 1021648
rect 370010 1021614 370355 1021638
rect 370023 1021570 370223 1021614
rect 370238 1021604 370262 1021614
rect 370238 1021580 370272 1021604
rect 370283 1021580 370355 1021614
rect 370238 1021570 370355 1021580
rect 370010 1021546 370355 1021570
rect 370023 1021502 370223 1021546
rect 370238 1021536 370262 1021546
rect 370238 1021512 370272 1021536
rect 370283 1021512 370355 1021546
rect 370238 1021502 370355 1021512
rect 370010 1021478 370355 1021502
rect 370023 1021434 370223 1021478
rect 370238 1021468 370262 1021478
rect 370238 1021444 370272 1021468
rect 370283 1021444 370355 1021478
rect 370238 1021434 370355 1021444
rect 370010 1021410 370355 1021434
rect 370023 1021366 370223 1021410
rect 370238 1021400 370262 1021410
rect 370238 1021376 370272 1021400
rect 370283 1021376 370355 1021410
rect 370238 1021366 370355 1021376
rect 370010 1021342 370355 1021366
rect 370023 1021298 370223 1021342
rect 370238 1021332 370262 1021342
rect 370238 1021308 370272 1021332
rect 370283 1021308 370355 1021342
rect 370238 1021298 370355 1021308
rect 370010 1021274 370355 1021298
rect 370023 1021230 370223 1021274
rect 370238 1021264 370262 1021274
rect 370238 1021240 370272 1021264
rect 370283 1021240 370355 1021274
rect 370238 1021230 370355 1021240
rect 370010 1021206 370355 1021230
rect 370023 1021162 370223 1021206
rect 370238 1021196 370262 1021206
rect 370238 1021172 370272 1021196
rect 370283 1021172 370355 1021206
rect 370238 1021162 370355 1021172
rect 370010 1021138 370355 1021162
rect 370023 1021094 370223 1021138
rect 370238 1021128 370262 1021138
rect 370238 1021104 370272 1021128
rect 370283 1021104 370355 1021138
rect 370238 1021094 370355 1021104
rect 370010 1021070 370355 1021094
rect 370023 1021026 370223 1021070
rect 370238 1021060 370262 1021070
rect 370238 1021036 370272 1021060
rect 370283 1021036 370355 1021070
rect 370238 1021026 370355 1021036
rect 370010 1021002 370355 1021026
rect 370023 1020958 370223 1021002
rect 370238 1020992 370262 1021002
rect 370238 1020968 370272 1020992
rect 370283 1020968 370355 1021002
rect 370238 1020958 370355 1020968
rect 370010 1020934 370355 1020958
rect 370023 1020922 370223 1020934
rect 370034 1020910 370058 1020922
rect 370238 1020910 370262 1020934
rect 370283 1020922 370355 1020934
rect 370585 1020922 370641 1021922
rect 370657 1020922 370713 1021922
rect 371015 1021842 371215 1021922
rect 371230 1021852 371264 1021876
rect 371275 1021852 371347 1021922
rect 371230 1021842 371347 1021852
rect 371002 1021818 371347 1021842
rect 371015 1021774 371215 1021818
rect 371230 1021808 371254 1021818
rect 371230 1021784 371264 1021808
rect 371275 1021784 371347 1021818
rect 371230 1021774 371347 1021784
rect 371002 1021750 371347 1021774
rect 371015 1021706 371215 1021750
rect 371230 1021740 371254 1021750
rect 371230 1021716 371264 1021740
rect 371275 1021716 371347 1021750
rect 371230 1021706 371347 1021716
rect 371002 1021682 371347 1021706
rect 371015 1021638 371215 1021682
rect 371230 1021672 371254 1021682
rect 371230 1021648 371264 1021672
rect 371275 1021648 371347 1021682
rect 371230 1021638 371347 1021648
rect 371002 1021614 371347 1021638
rect 371015 1021570 371215 1021614
rect 371230 1021604 371254 1021614
rect 371230 1021580 371264 1021604
rect 371275 1021580 371347 1021614
rect 371230 1021570 371347 1021580
rect 371002 1021546 371347 1021570
rect 371015 1021502 371215 1021546
rect 371230 1021536 371254 1021546
rect 371230 1021512 371264 1021536
rect 371275 1021512 371347 1021546
rect 371230 1021502 371347 1021512
rect 371002 1021478 371347 1021502
rect 371015 1021434 371215 1021478
rect 371230 1021468 371254 1021478
rect 371230 1021444 371264 1021468
rect 371275 1021444 371347 1021478
rect 371230 1021434 371347 1021444
rect 371002 1021410 371347 1021434
rect 371015 1021366 371215 1021410
rect 371230 1021400 371254 1021410
rect 371230 1021376 371264 1021400
rect 371275 1021376 371347 1021410
rect 371230 1021366 371347 1021376
rect 371002 1021342 371347 1021366
rect 371015 1021298 371215 1021342
rect 371230 1021332 371254 1021342
rect 371230 1021308 371264 1021332
rect 371275 1021308 371347 1021342
rect 371230 1021298 371347 1021308
rect 371002 1021274 371347 1021298
rect 371015 1021230 371215 1021274
rect 371230 1021264 371254 1021274
rect 371230 1021240 371264 1021264
rect 371275 1021240 371347 1021274
rect 371230 1021230 371347 1021240
rect 371002 1021206 371347 1021230
rect 371015 1021162 371215 1021206
rect 371230 1021196 371254 1021206
rect 371230 1021172 371264 1021196
rect 371275 1021172 371347 1021206
rect 371230 1021162 371347 1021172
rect 371002 1021138 371347 1021162
rect 371015 1021094 371215 1021138
rect 371230 1021128 371254 1021138
rect 371230 1021104 371264 1021128
rect 371275 1021104 371347 1021138
rect 371230 1021094 371347 1021104
rect 371002 1021070 371347 1021094
rect 371015 1021026 371215 1021070
rect 371230 1021060 371254 1021070
rect 371230 1021036 371264 1021060
rect 371275 1021036 371347 1021070
rect 371230 1021026 371347 1021036
rect 371002 1021002 371347 1021026
rect 371015 1020958 371215 1021002
rect 371230 1020992 371254 1021002
rect 371230 1020968 371264 1020992
rect 371275 1020968 371347 1021002
rect 371230 1020958 371347 1020968
rect 371002 1020934 371347 1020958
rect 371015 1020922 371215 1020934
rect 371026 1020910 371050 1020922
rect 371230 1020910 371254 1020934
rect 371275 1020922 371347 1020934
rect 371577 1020922 371633 1021922
rect 371649 1020922 371705 1021922
rect 372007 1021842 372207 1021922
rect 372222 1021852 372256 1021876
rect 372267 1021852 372339 1021922
rect 372222 1021842 372339 1021852
rect 371994 1021818 372339 1021842
rect 372007 1021774 372207 1021818
rect 372222 1021808 372246 1021818
rect 372222 1021784 372256 1021808
rect 372267 1021784 372339 1021818
rect 372222 1021774 372339 1021784
rect 371994 1021750 372339 1021774
rect 372007 1021706 372207 1021750
rect 372222 1021740 372246 1021750
rect 372222 1021716 372256 1021740
rect 372267 1021716 372339 1021750
rect 372222 1021706 372339 1021716
rect 371994 1021682 372339 1021706
rect 372007 1021638 372207 1021682
rect 372222 1021672 372246 1021682
rect 372222 1021648 372256 1021672
rect 372267 1021648 372339 1021682
rect 372222 1021638 372339 1021648
rect 371994 1021614 372339 1021638
rect 372007 1021570 372207 1021614
rect 372222 1021604 372246 1021614
rect 372222 1021580 372256 1021604
rect 372267 1021580 372339 1021614
rect 372222 1021570 372339 1021580
rect 371994 1021546 372339 1021570
rect 372007 1021502 372207 1021546
rect 372222 1021536 372246 1021546
rect 372222 1021512 372256 1021536
rect 372267 1021512 372339 1021546
rect 372222 1021502 372339 1021512
rect 371994 1021478 372339 1021502
rect 372007 1021434 372207 1021478
rect 372222 1021468 372246 1021478
rect 372222 1021444 372256 1021468
rect 372267 1021444 372339 1021478
rect 372222 1021434 372339 1021444
rect 371994 1021410 372339 1021434
rect 372007 1021366 372207 1021410
rect 372222 1021400 372246 1021410
rect 372222 1021376 372256 1021400
rect 372267 1021376 372339 1021410
rect 372222 1021366 372339 1021376
rect 371994 1021342 372339 1021366
rect 372007 1021298 372207 1021342
rect 372222 1021332 372246 1021342
rect 372222 1021308 372256 1021332
rect 372267 1021308 372339 1021342
rect 372222 1021298 372339 1021308
rect 371994 1021274 372339 1021298
rect 372007 1021230 372207 1021274
rect 372222 1021264 372246 1021274
rect 372222 1021240 372256 1021264
rect 372267 1021240 372339 1021274
rect 372222 1021230 372339 1021240
rect 371994 1021206 372339 1021230
rect 372007 1021162 372207 1021206
rect 372222 1021196 372246 1021206
rect 372222 1021172 372256 1021196
rect 372267 1021172 372339 1021206
rect 372222 1021162 372339 1021172
rect 371994 1021138 372339 1021162
rect 372007 1021094 372207 1021138
rect 372222 1021128 372246 1021138
rect 372222 1021104 372256 1021128
rect 372267 1021104 372339 1021138
rect 372222 1021094 372339 1021104
rect 371994 1021070 372339 1021094
rect 372007 1021026 372207 1021070
rect 372222 1021060 372246 1021070
rect 372222 1021036 372256 1021060
rect 372267 1021036 372339 1021070
rect 372222 1021026 372339 1021036
rect 371994 1021002 372339 1021026
rect 372007 1020958 372207 1021002
rect 372222 1020992 372246 1021002
rect 372222 1020968 372256 1020992
rect 372267 1020968 372339 1021002
rect 372222 1020958 372339 1020968
rect 371994 1020934 372339 1020958
rect 372007 1020922 372207 1020934
rect 372018 1020910 372042 1020922
rect 372222 1020910 372246 1020934
rect 372267 1020922 372339 1020934
rect 372569 1020922 372625 1021922
rect 372641 1020922 372697 1021922
rect 372999 1021842 373199 1021922
rect 373214 1021852 373248 1021876
rect 373259 1021852 373331 1021922
rect 373214 1021842 373331 1021852
rect 372986 1021818 373331 1021842
rect 372999 1021774 373199 1021818
rect 373214 1021808 373238 1021818
rect 373214 1021784 373248 1021808
rect 373259 1021784 373331 1021818
rect 373214 1021774 373331 1021784
rect 372986 1021750 373331 1021774
rect 372999 1021706 373199 1021750
rect 373214 1021740 373238 1021750
rect 373214 1021716 373248 1021740
rect 373259 1021716 373331 1021750
rect 373214 1021706 373331 1021716
rect 372986 1021682 373331 1021706
rect 372999 1021638 373199 1021682
rect 373214 1021672 373238 1021682
rect 373214 1021648 373248 1021672
rect 373259 1021648 373331 1021682
rect 373214 1021638 373331 1021648
rect 372986 1021614 373331 1021638
rect 372999 1021570 373199 1021614
rect 373214 1021604 373238 1021614
rect 373214 1021580 373248 1021604
rect 373259 1021580 373331 1021614
rect 373214 1021570 373331 1021580
rect 372986 1021546 373331 1021570
rect 372999 1021502 373199 1021546
rect 373214 1021536 373238 1021546
rect 373214 1021512 373248 1021536
rect 373259 1021512 373331 1021546
rect 373214 1021502 373331 1021512
rect 372986 1021478 373331 1021502
rect 372999 1021434 373199 1021478
rect 373214 1021468 373238 1021478
rect 373214 1021444 373248 1021468
rect 373259 1021444 373331 1021478
rect 373214 1021434 373331 1021444
rect 372986 1021410 373331 1021434
rect 372999 1021366 373199 1021410
rect 373214 1021400 373238 1021410
rect 373214 1021376 373248 1021400
rect 373259 1021376 373331 1021410
rect 373214 1021366 373331 1021376
rect 372986 1021342 373331 1021366
rect 372999 1021298 373199 1021342
rect 373214 1021332 373238 1021342
rect 373214 1021308 373248 1021332
rect 373259 1021308 373331 1021342
rect 373214 1021298 373331 1021308
rect 372986 1021274 373331 1021298
rect 372999 1021230 373199 1021274
rect 373214 1021264 373238 1021274
rect 373214 1021240 373248 1021264
rect 373259 1021240 373331 1021274
rect 373214 1021230 373331 1021240
rect 372986 1021206 373331 1021230
rect 372999 1021162 373199 1021206
rect 373214 1021196 373238 1021206
rect 373214 1021172 373248 1021196
rect 373259 1021172 373331 1021206
rect 373214 1021162 373331 1021172
rect 372986 1021138 373331 1021162
rect 372999 1021094 373199 1021138
rect 373214 1021128 373238 1021138
rect 373214 1021104 373248 1021128
rect 373259 1021104 373331 1021138
rect 373214 1021094 373331 1021104
rect 372986 1021070 373331 1021094
rect 372999 1021026 373199 1021070
rect 373214 1021060 373238 1021070
rect 373214 1021036 373248 1021060
rect 373259 1021036 373331 1021070
rect 373214 1021026 373331 1021036
rect 372986 1021002 373331 1021026
rect 372999 1020958 373199 1021002
rect 373214 1020992 373238 1021002
rect 373214 1020968 373248 1020992
rect 373259 1020968 373331 1021002
rect 373214 1020958 373331 1020968
rect 372986 1020934 373331 1020958
rect 372999 1020922 373199 1020934
rect 373010 1020910 373034 1020922
rect 373214 1020910 373238 1020934
rect 373259 1020922 373331 1020934
rect 373561 1020922 373617 1021922
rect 373633 1020922 373689 1021922
rect 373991 1021842 374191 1021922
rect 374206 1021852 374240 1021876
rect 374251 1021852 374323 1021922
rect 374206 1021842 374323 1021852
rect 373978 1021818 374323 1021842
rect 373991 1021774 374191 1021818
rect 374206 1021808 374230 1021818
rect 374206 1021784 374240 1021808
rect 374251 1021784 374323 1021818
rect 374206 1021774 374323 1021784
rect 373978 1021750 374323 1021774
rect 373991 1021706 374191 1021750
rect 374206 1021740 374230 1021750
rect 374206 1021716 374240 1021740
rect 374251 1021716 374323 1021750
rect 374206 1021706 374323 1021716
rect 373978 1021682 374323 1021706
rect 373991 1021638 374191 1021682
rect 374206 1021672 374230 1021682
rect 374206 1021648 374240 1021672
rect 374251 1021648 374323 1021682
rect 374206 1021638 374323 1021648
rect 373978 1021614 374323 1021638
rect 373991 1021570 374191 1021614
rect 374206 1021604 374230 1021614
rect 374206 1021580 374240 1021604
rect 374251 1021580 374323 1021614
rect 374206 1021570 374323 1021580
rect 373978 1021546 374323 1021570
rect 373991 1021502 374191 1021546
rect 374206 1021536 374230 1021546
rect 374206 1021512 374240 1021536
rect 374251 1021512 374323 1021546
rect 374206 1021502 374323 1021512
rect 373978 1021478 374323 1021502
rect 373991 1021434 374191 1021478
rect 374206 1021468 374230 1021478
rect 374206 1021444 374240 1021468
rect 374251 1021444 374323 1021478
rect 374206 1021434 374323 1021444
rect 373978 1021410 374323 1021434
rect 373991 1021366 374191 1021410
rect 374206 1021400 374230 1021410
rect 374206 1021376 374240 1021400
rect 374251 1021376 374323 1021410
rect 374206 1021366 374323 1021376
rect 373978 1021342 374323 1021366
rect 373991 1021298 374191 1021342
rect 374206 1021332 374230 1021342
rect 374206 1021308 374240 1021332
rect 374251 1021308 374323 1021342
rect 374206 1021298 374323 1021308
rect 373978 1021274 374323 1021298
rect 373991 1021230 374191 1021274
rect 374206 1021264 374230 1021274
rect 374206 1021240 374240 1021264
rect 374251 1021240 374323 1021274
rect 374206 1021230 374323 1021240
rect 373978 1021206 374323 1021230
rect 373991 1021162 374191 1021206
rect 374206 1021196 374230 1021206
rect 374206 1021172 374240 1021196
rect 374251 1021172 374323 1021206
rect 374206 1021162 374323 1021172
rect 373978 1021138 374323 1021162
rect 373991 1021094 374191 1021138
rect 374206 1021128 374230 1021138
rect 374206 1021104 374240 1021128
rect 374251 1021104 374323 1021138
rect 374206 1021094 374323 1021104
rect 373978 1021070 374323 1021094
rect 373991 1021026 374191 1021070
rect 374206 1021060 374230 1021070
rect 374206 1021036 374240 1021060
rect 374251 1021036 374323 1021070
rect 374206 1021026 374323 1021036
rect 373978 1021002 374323 1021026
rect 373991 1020958 374191 1021002
rect 374206 1020992 374230 1021002
rect 374206 1020968 374240 1020992
rect 374251 1020968 374323 1021002
rect 374206 1020958 374323 1020968
rect 373978 1020934 374323 1020958
rect 373991 1020922 374191 1020934
rect 374002 1020910 374026 1020922
rect 374206 1020910 374230 1020934
rect 374251 1020922 374323 1020934
rect 374553 1020922 374609 1021922
rect 374625 1020922 374681 1021922
rect 374983 1021842 375183 1021922
rect 375198 1021852 375232 1021876
rect 375243 1021852 375315 1021922
rect 375198 1021842 375315 1021852
rect 374970 1021818 375315 1021842
rect 374983 1021774 375183 1021818
rect 375198 1021808 375222 1021818
rect 375198 1021784 375232 1021808
rect 375243 1021784 375315 1021818
rect 375198 1021774 375315 1021784
rect 374970 1021750 375315 1021774
rect 374983 1021706 375183 1021750
rect 375198 1021740 375222 1021750
rect 375198 1021716 375232 1021740
rect 375243 1021716 375315 1021750
rect 375198 1021706 375315 1021716
rect 374970 1021682 375315 1021706
rect 374983 1021638 375183 1021682
rect 375198 1021672 375222 1021682
rect 375198 1021648 375232 1021672
rect 375243 1021648 375315 1021682
rect 375198 1021638 375315 1021648
rect 374970 1021614 375315 1021638
rect 374983 1021570 375183 1021614
rect 375198 1021604 375222 1021614
rect 375198 1021580 375232 1021604
rect 375243 1021580 375315 1021614
rect 375198 1021570 375315 1021580
rect 374970 1021546 375315 1021570
rect 374983 1021502 375183 1021546
rect 375198 1021536 375222 1021546
rect 375198 1021512 375232 1021536
rect 375243 1021512 375315 1021546
rect 375198 1021502 375315 1021512
rect 374970 1021478 375315 1021502
rect 374983 1021434 375183 1021478
rect 375198 1021468 375222 1021478
rect 375198 1021444 375232 1021468
rect 375243 1021444 375315 1021478
rect 375198 1021434 375315 1021444
rect 374970 1021410 375315 1021434
rect 374983 1021366 375183 1021410
rect 375198 1021400 375222 1021410
rect 375198 1021376 375232 1021400
rect 375243 1021376 375315 1021410
rect 375198 1021366 375315 1021376
rect 374970 1021342 375315 1021366
rect 374983 1021298 375183 1021342
rect 375198 1021332 375222 1021342
rect 375198 1021308 375232 1021332
rect 375243 1021308 375315 1021342
rect 375198 1021298 375315 1021308
rect 374970 1021274 375315 1021298
rect 374983 1021230 375183 1021274
rect 375198 1021264 375222 1021274
rect 375198 1021240 375232 1021264
rect 375243 1021240 375315 1021274
rect 375198 1021230 375315 1021240
rect 374970 1021206 375315 1021230
rect 374983 1021162 375183 1021206
rect 375198 1021196 375222 1021206
rect 375198 1021172 375232 1021196
rect 375243 1021172 375315 1021206
rect 375198 1021162 375315 1021172
rect 374970 1021138 375315 1021162
rect 374983 1021094 375183 1021138
rect 375198 1021128 375222 1021138
rect 375198 1021104 375232 1021128
rect 375243 1021104 375315 1021138
rect 375198 1021094 375315 1021104
rect 374970 1021070 375315 1021094
rect 374983 1021026 375183 1021070
rect 375198 1021060 375222 1021070
rect 375198 1021036 375232 1021060
rect 375243 1021036 375315 1021070
rect 375198 1021026 375315 1021036
rect 374970 1021002 375315 1021026
rect 374983 1020958 375183 1021002
rect 375198 1020992 375222 1021002
rect 375198 1020968 375232 1020992
rect 375243 1020968 375315 1021002
rect 375198 1020958 375315 1020968
rect 374970 1020934 375315 1020958
rect 374983 1020922 375183 1020934
rect 374994 1020910 375018 1020922
rect 375198 1020910 375222 1020934
rect 375243 1020922 375315 1020934
rect 375545 1020922 375601 1021922
rect 375617 1020922 375673 1021922
rect 375975 1021842 376175 1021922
rect 376190 1021852 376224 1021876
rect 376235 1021852 376307 1021922
rect 376190 1021842 376307 1021852
rect 375962 1021818 376307 1021842
rect 375975 1021774 376175 1021818
rect 376190 1021808 376214 1021818
rect 376190 1021784 376224 1021808
rect 376235 1021784 376307 1021818
rect 376190 1021774 376307 1021784
rect 375962 1021750 376307 1021774
rect 375975 1021706 376175 1021750
rect 376190 1021740 376214 1021750
rect 376190 1021716 376224 1021740
rect 376235 1021716 376307 1021750
rect 376190 1021706 376307 1021716
rect 375962 1021682 376307 1021706
rect 375975 1021638 376175 1021682
rect 376190 1021672 376214 1021682
rect 376190 1021648 376224 1021672
rect 376235 1021648 376307 1021682
rect 376190 1021638 376307 1021648
rect 375962 1021614 376307 1021638
rect 375975 1021570 376175 1021614
rect 376190 1021604 376214 1021614
rect 376190 1021580 376224 1021604
rect 376235 1021580 376307 1021614
rect 376190 1021570 376307 1021580
rect 375962 1021546 376307 1021570
rect 375975 1021502 376175 1021546
rect 376190 1021536 376214 1021546
rect 376190 1021512 376224 1021536
rect 376235 1021512 376307 1021546
rect 376190 1021502 376307 1021512
rect 375962 1021478 376307 1021502
rect 375975 1021434 376175 1021478
rect 376190 1021468 376214 1021478
rect 376190 1021444 376224 1021468
rect 376235 1021444 376307 1021478
rect 376190 1021434 376307 1021444
rect 375962 1021410 376307 1021434
rect 375975 1021366 376175 1021410
rect 376190 1021400 376214 1021410
rect 376190 1021376 376224 1021400
rect 376235 1021376 376307 1021410
rect 376190 1021366 376307 1021376
rect 375962 1021342 376307 1021366
rect 375975 1021298 376175 1021342
rect 376190 1021332 376214 1021342
rect 376190 1021308 376224 1021332
rect 376235 1021308 376307 1021342
rect 376190 1021298 376307 1021308
rect 375962 1021274 376307 1021298
rect 375975 1021230 376175 1021274
rect 376190 1021264 376214 1021274
rect 376190 1021240 376224 1021264
rect 376235 1021240 376307 1021274
rect 376190 1021230 376307 1021240
rect 375962 1021206 376307 1021230
rect 375975 1021162 376175 1021206
rect 376190 1021196 376214 1021206
rect 376190 1021172 376224 1021196
rect 376235 1021172 376307 1021206
rect 376190 1021162 376307 1021172
rect 375962 1021138 376307 1021162
rect 375975 1021094 376175 1021138
rect 376190 1021128 376214 1021138
rect 376190 1021104 376224 1021128
rect 376235 1021104 376307 1021138
rect 376190 1021094 376307 1021104
rect 375962 1021070 376307 1021094
rect 375975 1021026 376175 1021070
rect 376190 1021060 376214 1021070
rect 376190 1021036 376224 1021060
rect 376235 1021036 376307 1021070
rect 376190 1021026 376307 1021036
rect 375962 1021002 376307 1021026
rect 375975 1020958 376175 1021002
rect 376190 1020992 376214 1021002
rect 376190 1020968 376224 1020992
rect 376235 1020968 376307 1021002
rect 376190 1020958 376307 1020968
rect 375962 1020934 376307 1020958
rect 375975 1020922 376175 1020934
rect 375986 1020910 376010 1020922
rect 376190 1020910 376214 1020934
rect 376235 1020922 376307 1020934
rect 376537 1020922 376593 1021922
rect 376609 1020922 376665 1021922
rect 376967 1021842 377167 1021922
rect 377182 1021852 377216 1021876
rect 377227 1021852 377299 1021922
rect 377182 1021842 377299 1021852
rect 376954 1021818 377299 1021842
rect 376967 1021774 377167 1021818
rect 377182 1021808 377206 1021818
rect 377182 1021784 377216 1021808
rect 377227 1021784 377299 1021818
rect 377182 1021774 377299 1021784
rect 376954 1021750 377299 1021774
rect 376967 1021706 377167 1021750
rect 377182 1021740 377206 1021750
rect 377182 1021716 377216 1021740
rect 377227 1021716 377299 1021750
rect 377182 1021706 377299 1021716
rect 376954 1021682 377299 1021706
rect 376967 1021638 377167 1021682
rect 377182 1021672 377206 1021682
rect 377182 1021648 377216 1021672
rect 377227 1021648 377299 1021682
rect 377182 1021638 377299 1021648
rect 376954 1021614 377299 1021638
rect 376967 1021570 377167 1021614
rect 377182 1021604 377206 1021614
rect 377182 1021580 377216 1021604
rect 377227 1021580 377299 1021614
rect 377182 1021570 377299 1021580
rect 376954 1021546 377299 1021570
rect 376967 1021502 377167 1021546
rect 377182 1021536 377206 1021546
rect 377182 1021512 377216 1021536
rect 377227 1021512 377299 1021546
rect 377182 1021502 377299 1021512
rect 376954 1021478 377299 1021502
rect 376967 1021434 377167 1021478
rect 377182 1021468 377206 1021478
rect 377182 1021444 377216 1021468
rect 377227 1021444 377299 1021478
rect 377182 1021434 377299 1021444
rect 376954 1021410 377299 1021434
rect 376967 1021366 377167 1021410
rect 377182 1021400 377206 1021410
rect 377182 1021376 377216 1021400
rect 377227 1021376 377299 1021410
rect 377182 1021366 377299 1021376
rect 376954 1021342 377299 1021366
rect 376967 1021298 377167 1021342
rect 377182 1021332 377206 1021342
rect 377182 1021308 377216 1021332
rect 377227 1021308 377299 1021342
rect 377182 1021298 377299 1021308
rect 376954 1021274 377299 1021298
rect 376967 1021230 377167 1021274
rect 377182 1021264 377206 1021274
rect 377182 1021240 377216 1021264
rect 377227 1021240 377299 1021274
rect 377182 1021230 377299 1021240
rect 376954 1021206 377299 1021230
rect 376967 1021162 377167 1021206
rect 377182 1021196 377206 1021206
rect 377182 1021172 377216 1021196
rect 377227 1021172 377299 1021206
rect 377182 1021162 377299 1021172
rect 376954 1021138 377299 1021162
rect 376967 1021094 377167 1021138
rect 377182 1021128 377206 1021138
rect 377182 1021104 377216 1021128
rect 377227 1021104 377299 1021138
rect 377182 1021094 377299 1021104
rect 376954 1021070 377299 1021094
rect 376967 1021026 377167 1021070
rect 377182 1021060 377206 1021070
rect 377182 1021036 377216 1021060
rect 377227 1021036 377299 1021070
rect 377182 1021026 377299 1021036
rect 376954 1021002 377299 1021026
rect 376967 1020958 377167 1021002
rect 377182 1020992 377206 1021002
rect 377182 1020968 377216 1020992
rect 377227 1020968 377299 1021002
rect 377182 1020958 377299 1020968
rect 376954 1020934 377299 1020958
rect 376967 1020922 377167 1020934
rect 376978 1020910 377002 1020922
rect 377182 1020910 377206 1020934
rect 377227 1020922 377299 1020934
rect 377529 1020922 377585 1021922
rect 377601 1020922 377657 1021922
rect 377959 1021842 378159 1021922
rect 378174 1021852 378208 1021876
rect 378219 1021852 378291 1021922
rect 378174 1021842 378291 1021852
rect 377946 1021818 378291 1021842
rect 377959 1021774 378159 1021818
rect 378174 1021808 378198 1021818
rect 378174 1021784 378208 1021808
rect 378219 1021784 378291 1021818
rect 378174 1021774 378291 1021784
rect 377946 1021750 378291 1021774
rect 377959 1021706 378159 1021750
rect 378174 1021740 378198 1021750
rect 378174 1021716 378208 1021740
rect 378219 1021716 378291 1021750
rect 378174 1021706 378291 1021716
rect 377946 1021682 378291 1021706
rect 377959 1021638 378159 1021682
rect 378174 1021672 378198 1021682
rect 378174 1021648 378208 1021672
rect 378219 1021648 378291 1021682
rect 378174 1021638 378291 1021648
rect 377946 1021614 378291 1021638
rect 377959 1021570 378159 1021614
rect 378174 1021604 378198 1021614
rect 378174 1021580 378208 1021604
rect 378219 1021580 378291 1021614
rect 378174 1021570 378291 1021580
rect 377946 1021546 378291 1021570
rect 377959 1021502 378159 1021546
rect 378174 1021536 378198 1021546
rect 378174 1021512 378208 1021536
rect 378219 1021512 378291 1021546
rect 378174 1021502 378291 1021512
rect 377946 1021478 378291 1021502
rect 377959 1021434 378159 1021478
rect 378174 1021468 378198 1021478
rect 378174 1021444 378208 1021468
rect 378219 1021444 378291 1021478
rect 378174 1021434 378291 1021444
rect 377946 1021410 378291 1021434
rect 377959 1021366 378159 1021410
rect 378174 1021400 378198 1021410
rect 378174 1021376 378208 1021400
rect 378219 1021376 378291 1021410
rect 378174 1021366 378291 1021376
rect 377946 1021342 378291 1021366
rect 377959 1021298 378159 1021342
rect 378174 1021332 378198 1021342
rect 378174 1021308 378208 1021332
rect 378219 1021308 378291 1021342
rect 378174 1021298 378291 1021308
rect 377946 1021274 378291 1021298
rect 377959 1021230 378159 1021274
rect 378174 1021264 378198 1021274
rect 378174 1021240 378208 1021264
rect 378219 1021240 378291 1021274
rect 378174 1021230 378291 1021240
rect 377946 1021206 378291 1021230
rect 377959 1021162 378159 1021206
rect 378174 1021196 378198 1021206
rect 378174 1021172 378208 1021196
rect 378219 1021172 378291 1021206
rect 378174 1021162 378291 1021172
rect 377946 1021138 378291 1021162
rect 377959 1021094 378159 1021138
rect 378174 1021128 378198 1021138
rect 378174 1021104 378208 1021128
rect 378219 1021104 378291 1021138
rect 378174 1021094 378291 1021104
rect 377946 1021070 378291 1021094
rect 377959 1021026 378159 1021070
rect 378174 1021060 378198 1021070
rect 378174 1021036 378208 1021060
rect 378219 1021036 378291 1021070
rect 378174 1021026 378291 1021036
rect 377946 1021002 378291 1021026
rect 377959 1020958 378159 1021002
rect 378174 1020992 378198 1021002
rect 378174 1020968 378208 1020992
rect 378219 1020968 378291 1021002
rect 378174 1020958 378291 1020968
rect 377946 1020934 378291 1020958
rect 377959 1020922 378159 1020934
rect 377970 1020910 377994 1020922
rect 378174 1020910 378198 1020934
rect 378219 1020922 378291 1020934
rect 378521 1020922 378577 1021922
rect 378593 1020922 378649 1021922
rect 378951 1021842 379151 1021922
rect 379166 1021852 379200 1021876
rect 379211 1021852 379283 1021922
rect 379166 1021842 379283 1021852
rect 378938 1021818 379283 1021842
rect 378951 1021774 379151 1021818
rect 379166 1021808 379190 1021818
rect 379166 1021784 379200 1021808
rect 379211 1021784 379283 1021818
rect 379166 1021774 379283 1021784
rect 378938 1021750 379283 1021774
rect 378951 1021706 379151 1021750
rect 379166 1021740 379190 1021750
rect 379166 1021716 379200 1021740
rect 379211 1021716 379283 1021750
rect 379166 1021706 379283 1021716
rect 378938 1021682 379283 1021706
rect 378951 1021638 379151 1021682
rect 379166 1021672 379190 1021682
rect 379166 1021648 379200 1021672
rect 379211 1021648 379283 1021682
rect 379166 1021638 379283 1021648
rect 378938 1021614 379283 1021638
rect 378951 1021570 379151 1021614
rect 379166 1021604 379190 1021614
rect 379166 1021580 379200 1021604
rect 379211 1021580 379283 1021614
rect 379166 1021570 379283 1021580
rect 378938 1021546 379283 1021570
rect 378951 1021502 379151 1021546
rect 379166 1021536 379190 1021546
rect 379166 1021512 379200 1021536
rect 379211 1021512 379283 1021546
rect 379166 1021502 379283 1021512
rect 378938 1021478 379283 1021502
rect 378951 1021434 379151 1021478
rect 379166 1021468 379190 1021478
rect 379166 1021444 379200 1021468
rect 379211 1021444 379283 1021478
rect 379166 1021434 379283 1021444
rect 378938 1021410 379283 1021434
rect 378951 1021366 379151 1021410
rect 379166 1021400 379190 1021410
rect 379166 1021376 379200 1021400
rect 379211 1021376 379283 1021410
rect 379166 1021366 379283 1021376
rect 378938 1021342 379283 1021366
rect 378951 1021298 379151 1021342
rect 379166 1021332 379190 1021342
rect 379166 1021308 379200 1021332
rect 379211 1021308 379283 1021342
rect 379166 1021298 379283 1021308
rect 378938 1021274 379283 1021298
rect 378951 1021230 379151 1021274
rect 379166 1021264 379190 1021274
rect 379166 1021240 379200 1021264
rect 379211 1021240 379283 1021274
rect 379166 1021230 379283 1021240
rect 378938 1021206 379283 1021230
rect 378951 1021162 379151 1021206
rect 379166 1021196 379190 1021206
rect 379166 1021172 379200 1021196
rect 379211 1021172 379283 1021206
rect 379166 1021162 379283 1021172
rect 378938 1021138 379283 1021162
rect 378951 1021094 379151 1021138
rect 379166 1021128 379190 1021138
rect 379166 1021104 379200 1021128
rect 379211 1021104 379283 1021138
rect 379166 1021094 379283 1021104
rect 378938 1021070 379283 1021094
rect 378951 1021026 379151 1021070
rect 379166 1021060 379190 1021070
rect 379166 1021036 379200 1021060
rect 379211 1021036 379283 1021070
rect 379166 1021026 379283 1021036
rect 378938 1021002 379283 1021026
rect 378951 1020958 379151 1021002
rect 379166 1020992 379190 1021002
rect 379166 1020968 379200 1020992
rect 379211 1020968 379283 1021002
rect 379166 1020958 379283 1020968
rect 378938 1020934 379283 1020958
rect 378951 1020922 379151 1020934
rect 378962 1020910 378986 1020922
rect 379166 1020910 379190 1020934
rect 379211 1020922 379283 1020934
rect 379472 1020922 379544 1021922
rect 379610 1020922 379627 1021922
rect 379797 1020922 379830 1021922
rect 379953 1021730 380025 1021760
rect 379953 1021692 379987 1021722
rect 367058 1020322 367092 1020334
rect 366356 1019322 366406 1020322
rect 366617 1019322 366673 1020322
rect 366689 1019322 366745 1020322
rect 367047 1020300 367247 1020322
rect 367262 1020310 367296 1020334
rect 368050 1020322 368084 1020334
rect 367307 1020310 367379 1020322
rect 367262 1020300 367379 1020310
rect 367034 1020276 367379 1020300
rect 367047 1020232 367247 1020276
rect 367262 1020266 367286 1020276
rect 367262 1020242 367296 1020266
rect 367307 1020242 367379 1020276
rect 367262 1020232 367379 1020242
rect 367034 1020208 367379 1020232
rect 367047 1020164 367247 1020208
rect 367262 1020198 367286 1020208
rect 367262 1020174 367296 1020198
rect 367307 1020174 367379 1020208
rect 367262 1020164 367379 1020174
rect 367034 1020140 367379 1020164
rect 367047 1020096 367247 1020140
rect 367262 1020130 367286 1020140
rect 367262 1020106 367296 1020130
rect 367307 1020106 367379 1020140
rect 367262 1020096 367379 1020106
rect 367034 1020072 367379 1020096
rect 367047 1020028 367247 1020072
rect 367262 1020062 367286 1020072
rect 367262 1020038 367296 1020062
rect 367307 1020038 367379 1020072
rect 367262 1020028 367379 1020038
rect 367034 1020004 367379 1020028
rect 367047 1019960 367247 1020004
rect 367262 1019994 367286 1020004
rect 367262 1019970 367296 1019994
rect 367307 1019970 367379 1020004
rect 367262 1019960 367379 1019970
rect 367034 1019936 367379 1019960
rect 367047 1019892 367247 1019936
rect 367262 1019926 367286 1019936
rect 367262 1019902 367296 1019926
rect 367307 1019902 367379 1019936
rect 367262 1019892 367379 1019902
rect 367034 1019868 367379 1019892
rect 367047 1019824 367247 1019868
rect 367262 1019858 367286 1019868
rect 367262 1019834 367296 1019858
rect 367307 1019834 367379 1019868
rect 367262 1019824 367379 1019834
rect 367034 1019800 367379 1019824
rect 367047 1019756 367247 1019800
rect 367262 1019790 367286 1019800
rect 367262 1019766 367296 1019790
rect 367307 1019766 367379 1019800
rect 367262 1019756 367379 1019766
rect 367034 1019732 367379 1019756
rect 367047 1019688 367247 1019732
rect 367262 1019722 367286 1019732
rect 367262 1019698 367296 1019722
rect 367307 1019698 367379 1019732
rect 367262 1019688 367379 1019698
rect 367034 1019664 367379 1019688
rect 367047 1019620 367247 1019664
rect 367262 1019654 367286 1019664
rect 367262 1019630 367296 1019654
rect 367307 1019630 367379 1019664
rect 367262 1019620 367379 1019630
rect 367034 1019596 367379 1019620
rect 367047 1019552 367247 1019596
rect 367262 1019586 367286 1019596
rect 367262 1019562 367296 1019586
rect 367307 1019562 367379 1019596
rect 367262 1019552 367379 1019562
rect 367034 1019528 367379 1019552
rect 367047 1019484 367247 1019528
rect 367262 1019518 367286 1019528
rect 367262 1019494 367296 1019518
rect 367307 1019494 367379 1019528
rect 367262 1019484 367379 1019494
rect 367034 1019460 367379 1019484
rect 367047 1019416 367247 1019460
rect 367262 1019450 367286 1019460
rect 367262 1019426 367296 1019450
rect 367307 1019426 367379 1019460
rect 367262 1019416 367379 1019426
rect 367034 1019392 367379 1019416
rect 367047 1019322 367247 1019392
rect 367262 1019368 367286 1019392
rect 367307 1019322 367379 1019392
rect 367609 1019322 367665 1020322
rect 367681 1019322 367737 1020322
rect 368039 1020300 368239 1020322
rect 368254 1020310 368288 1020334
rect 369042 1020322 369076 1020334
rect 368299 1020310 368371 1020322
rect 368254 1020300 368371 1020310
rect 368026 1020276 368371 1020300
rect 368039 1020232 368239 1020276
rect 368254 1020266 368278 1020276
rect 368254 1020242 368288 1020266
rect 368299 1020242 368371 1020276
rect 368254 1020232 368371 1020242
rect 368026 1020208 368371 1020232
rect 368039 1020164 368239 1020208
rect 368254 1020198 368278 1020208
rect 368254 1020174 368288 1020198
rect 368299 1020174 368371 1020208
rect 368254 1020164 368371 1020174
rect 368026 1020140 368371 1020164
rect 368039 1020096 368239 1020140
rect 368254 1020130 368278 1020140
rect 368254 1020106 368288 1020130
rect 368299 1020106 368371 1020140
rect 368254 1020096 368371 1020106
rect 368026 1020072 368371 1020096
rect 368039 1020028 368239 1020072
rect 368254 1020062 368278 1020072
rect 368254 1020038 368288 1020062
rect 368299 1020038 368371 1020072
rect 368254 1020028 368371 1020038
rect 368026 1020004 368371 1020028
rect 368039 1019960 368239 1020004
rect 368254 1019994 368278 1020004
rect 368254 1019970 368288 1019994
rect 368299 1019970 368371 1020004
rect 368254 1019960 368371 1019970
rect 368026 1019936 368371 1019960
rect 368039 1019892 368239 1019936
rect 368254 1019926 368278 1019936
rect 368254 1019902 368288 1019926
rect 368299 1019902 368371 1019936
rect 368254 1019892 368371 1019902
rect 368026 1019868 368371 1019892
rect 368039 1019824 368239 1019868
rect 368254 1019858 368278 1019868
rect 368254 1019834 368288 1019858
rect 368299 1019834 368371 1019868
rect 368254 1019824 368371 1019834
rect 368026 1019800 368371 1019824
rect 368039 1019756 368239 1019800
rect 368254 1019790 368278 1019800
rect 368254 1019766 368288 1019790
rect 368299 1019766 368371 1019800
rect 368254 1019756 368371 1019766
rect 368026 1019732 368371 1019756
rect 368039 1019688 368239 1019732
rect 368254 1019722 368278 1019732
rect 368254 1019698 368288 1019722
rect 368299 1019698 368371 1019732
rect 368254 1019688 368371 1019698
rect 368026 1019664 368371 1019688
rect 368039 1019620 368239 1019664
rect 368254 1019654 368278 1019664
rect 368254 1019630 368288 1019654
rect 368299 1019630 368371 1019664
rect 368254 1019620 368371 1019630
rect 368026 1019596 368371 1019620
rect 368039 1019552 368239 1019596
rect 368254 1019586 368278 1019596
rect 368254 1019562 368288 1019586
rect 368299 1019562 368371 1019596
rect 368254 1019552 368371 1019562
rect 368026 1019528 368371 1019552
rect 368039 1019484 368239 1019528
rect 368254 1019518 368278 1019528
rect 368254 1019494 368288 1019518
rect 368299 1019494 368371 1019528
rect 368254 1019484 368371 1019494
rect 368026 1019460 368371 1019484
rect 368039 1019416 368239 1019460
rect 368254 1019450 368278 1019460
rect 368254 1019426 368288 1019450
rect 368299 1019426 368371 1019460
rect 368254 1019416 368371 1019426
rect 368026 1019392 368371 1019416
rect 368039 1019322 368239 1019392
rect 368254 1019368 368278 1019392
rect 368299 1019322 368371 1019392
rect 368601 1019322 368657 1020322
rect 368673 1019322 368729 1020322
rect 369031 1020300 369231 1020322
rect 369246 1020310 369280 1020334
rect 370034 1020322 370068 1020334
rect 369291 1020310 369363 1020322
rect 369246 1020300 369363 1020310
rect 369018 1020276 369363 1020300
rect 369031 1020232 369231 1020276
rect 369246 1020266 369270 1020276
rect 369246 1020242 369280 1020266
rect 369291 1020242 369363 1020276
rect 369246 1020232 369363 1020242
rect 369018 1020208 369363 1020232
rect 369031 1020164 369231 1020208
rect 369246 1020198 369270 1020208
rect 369246 1020174 369280 1020198
rect 369291 1020174 369363 1020208
rect 369246 1020164 369363 1020174
rect 369018 1020140 369363 1020164
rect 369031 1020096 369231 1020140
rect 369246 1020130 369270 1020140
rect 369246 1020106 369280 1020130
rect 369291 1020106 369363 1020140
rect 369246 1020096 369363 1020106
rect 369018 1020072 369363 1020096
rect 369031 1020028 369231 1020072
rect 369246 1020062 369270 1020072
rect 369246 1020038 369280 1020062
rect 369291 1020038 369363 1020072
rect 369246 1020028 369363 1020038
rect 369018 1020004 369363 1020028
rect 369031 1019960 369231 1020004
rect 369246 1019994 369270 1020004
rect 369246 1019970 369280 1019994
rect 369291 1019970 369363 1020004
rect 369246 1019960 369363 1019970
rect 369018 1019936 369363 1019960
rect 369031 1019892 369231 1019936
rect 369246 1019926 369270 1019936
rect 369246 1019902 369280 1019926
rect 369291 1019902 369363 1019936
rect 369246 1019892 369363 1019902
rect 369018 1019868 369363 1019892
rect 369031 1019824 369231 1019868
rect 369246 1019858 369270 1019868
rect 369246 1019834 369280 1019858
rect 369291 1019834 369363 1019868
rect 369246 1019824 369363 1019834
rect 369018 1019800 369363 1019824
rect 369031 1019756 369231 1019800
rect 369246 1019790 369270 1019800
rect 369246 1019766 369280 1019790
rect 369291 1019766 369363 1019800
rect 369246 1019756 369363 1019766
rect 369018 1019732 369363 1019756
rect 369031 1019688 369231 1019732
rect 369246 1019722 369270 1019732
rect 369246 1019698 369280 1019722
rect 369291 1019698 369363 1019732
rect 369246 1019688 369363 1019698
rect 369018 1019664 369363 1019688
rect 369031 1019620 369231 1019664
rect 369246 1019654 369270 1019664
rect 369246 1019630 369280 1019654
rect 369291 1019630 369363 1019664
rect 369246 1019620 369363 1019630
rect 369018 1019596 369363 1019620
rect 369031 1019552 369231 1019596
rect 369246 1019586 369270 1019596
rect 369246 1019562 369280 1019586
rect 369291 1019562 369363 1019596
rect 369246 1019552 369363 1019562
rect 369018 1019528 369363 1019552
rect 369031 1019484 369231 1019528
rect 369246 1019518 369270 1019528
rect 369246 1019494 369280 1019518
rect 369291 1019494 369363 1019528
rect 369246 1019484 369363 1019494
rect 369018 1019460 369363 1019484
rect 369031 1019416 369231 1019460
rect 369246 1019450 369270 1019460
rect 369246 1019426 369280 1019450
rect 369291 1019426 369363 1019460
rect 369246 1019416 369363 1019426
rect 369018 1019392 369363 1019416
rect 369031 1019322 369231 1019392
rect 369246 1019368 369270 1019392
rect 369291 1019322 369363 1019392
rect 369593 1019322 369649 1020322
rect 369665 1019322 369721 1020322
rect 370023 1020300 370223 1020322
rect 370238 1020310 370272 1020334
rect 371026 1020322 371060 1020334
rect 370283 1020310 370355 1020322
rect 370238 1020300 370355 1020310
rect 370010 1020276 370355 1020300
rect 370023 1020232 370223 1020276
rect 370238 1020266 370262 1020276
rect 370238 1020242 370272 1020266
rect 370283 1020242 370355 1020276
rect 370238 1020232 370355 1020242
rect 370010 1020208 370355 1020232
rect 370023 1020164 370223 1020208
rect 370238 1020198 370262 1020208
rect 370238 1020174 370272 1020198
rect 370283 1020174 370355 1020208
rect 370238 1020164 370355 1020174
rect 370010 1020140 370355 1020164
rect 370023 1020096 370223 1020140
rect 370238 1020130 370262 1020140
rect 370238 1020106 370272 1020130
rect 370283 1020106 370355 1020140
rect 370238 1020096 370355 1020106
rect 370010 1020072 370355 1020096
rect 370023 1020028 370223 1020072
rect 370238 1020062 370262 1020072
rect 370238 1020038 370272 1020062
rect 370283 1020038 370355 1020072
rect 370238 1020028 370355 1020038
rect 370010 1020004 370355 1020028
rect 370023 1019960 370223 1020004
rect 370238 1019994 370262 1020004
rect 370238 1019970 370272 1019994
rect 370283 1019970 370355 1020004
rect 370238 1019960 370355 1019970
rect 370010 1019936 370355 1019960
rect 370023 1019892 370223 1019936
rect 370238 1019926 370262 1019936
rect 370238 1019902 370272 1019926
rect 370283 1019902 370355 1019936
rect 370238 1019892 370355 1019902
rect 370010 1019868 370355 1019892
rect 370023 1019824 370223 1019868
rect 370238 1019858 370262 1019868
rect 370238 1019834 370272 1019858
rect 370283 1019834 370355 1019868
rect 370238 1019824 370355 1019834
rect 370010 1019800 370355 1019824
rect 370023 1019756 370223 1019800
rect 370238 1019790 370262 1019800
rect 370238 1019766 370272 1019790
rect 370283 1019766 370355 1019800
rect 370238 1019756 370355 1019766
rect 370010 1019732 370355 1019756
rect 370023 1019688 370223 1019732
rect 370238 1019722 370262 1019732
rect 370238 1019698 370272 1019722
rect 370283 1019698 370355 1019732
rect 370238 1019688 370355 1019698
rect 370010 1019664 370355 1019688
rect 370023 1019620 370223 1019664
rect 370238 1019654 370262 1019664
rect 370238 1019630 370272 1019654
rect 370283 1019630 370355 1019664
rect 370238 1019620 370355 1019630
rect 370010 1019596 370355 1019620
rect 370023 1019552 370223 1019596
rect 370238 1019586 370262 1019596
rect 370238 1019562 370272 1019586
rect 370283 1019562 370355 1019596
rect 370238 1019552 370355 1019562
rect 370010 1019528 370355 1019552
rect 370023 1019484 370223 1019528
rect 370238 1019518 370262 1019528
rect 370238 1019494 370272 1019518
rect 370283 1019494 370355 1019528
rect 370238 1019484 370355 1019494
rect 370010 1019460 370355 1019484
rect 370023 1019416 370223 1019460
rect 370238 1019450 370262 1019460
rect 370238 1019426 370272 1019450
rect 370283 1019426 370355 1019460
rect 370238 1019416 370355 1019426
rect 370010 1019392 370355 1019416
rect 370023 1019322 370223 1019392
rect 370238 1019368 370262 1019392
rect 370283 1019322 370355 1019392
rect 370585 1019322 370641 1020322
rect 370657 1019322 370713 1020322
rect 371015 1020300 371215 1020322
rect 371230 1020310 371264 1020334
rect 372018 1020322 372052 1020334
rect 371275 1020310 371347 1020322
rect 371230 1020300 371347 1020310
rect 371002 1020276 371347 1020300
rect 371015 1020232 371215 1020276
rect 371230 1020266 371254 1020276
rect 371230 1020242 371264 1020266
rect 371275 1020242 371347 1020276
rect 371230 1020232 371347 1020242
rect 371002 1020208 371347 1020232
rect 371015 1020164 371215 1020208
rect 371230 1020198 371254 1020208
rect 371230 1020174 371264 1020198
rect 371275 1020174 371347 1020208
rect 371230 1020164 371347 1020174
rect 371002 1020140 371347 1020164
rect 371015 1020096 371215 1020140
rect 371230 1020130 371254 1020140
rect 371230 1020106 371264 1020130
rect 371275 1020106 371347 1020140
rect 371230 1020096 371347 1020106
rect 371002 1020072 371347 1020096
rect 371015 1020028 371215 1020072
rect 371230 1020062 371254 1020072
rect 371230 1020038 371264 1020062
rect 371275 1020038 371347 1020072
rect 371230 1020028 371347 1020038
rect 371002 1020004 371347 1020028
rect 371015 1019960 371215 1020004
rect 371230 1019994 371254 1020004
rect 371230 1019970 371264 1019994
rect 371275 1019970 371347 1020004
rect 371230 1019960 371347 1019970
rect 371002 1019936 371347 1019960
rect 371015 1019892 371215 1019936
rect 371230 1019926 371254 1019936
rect 371230 1019902 371264 1019926
rect 371275 1019902 371347 1019936
rect 371230 1019892 371347 1019902
rect 371002 1019868 371347 1019892
rect 371015 1019824 371215 1019868
rect 371230 1019858 371254 1019868
rect 371230 1019834 371264 1019858
rect 371275 1019834 371347 1019868
rect 371230 1019824 371347 1019834
rect 371002 1019800 371347 1019824
rect 371015 1019756 371215 1019800
rect 371230 1019790 371254 1019800
rect 371230 1019766 371264 1019790
rect 371275 1019766 371347 1019800
rect 371230 1019756 371347 1019766
rect 371002 1019732 371347 1019756
rect 371015 1019688 371215 1019732
rect 371230 1019722 371254 1019732
rect 371230 1019698 371264 1019722
rect 371275 1019698 371347 1019732
rect 371230 1019688 371347 1019698
rect 371002 1019664 371347 1019688
rect 371015 1019620 371215 1019664
rect 371230 1019654 371254 1019664
rect 371230 1019630 371264 1019654
rect 371275 1019630 371347 1019664
rect 371230 1019620 371347 1019630
rect 371002 1019596 371347 1019620
rect 371015 1019552 371215 1019596
rect 371230 1019586 371254 1019596
rect 371230 1019562 371264 1019586
rect 371275 1019562 371347 1019596
rect 371230 1019552 371347 1019562
rect 371002 1019528 371347 1019552
rect 371015 1019484 371215 1019528
rect 371230 1019518 371254 1019528
rect 371230 1019494 371264 1019518
rect 371275 1019494 371347 1019528
rect 371230 1019484 371347 1019494
rect 371002 1019460 371347 1019484
rect 371015 1019416 371215 1019460
rect 371230 1019450 371254 1019460
rect 371230 1019426 371264 1019450
rect 371275 1019426 371347 1019460
rect 371230 1019416 371347 1019426
rect 371002 1019392 371347 1019416
rect 371015 1019322 371215 1019392
rect 371230 1019368 371254 1019392
rect 371275 1019322 371347 1019392
rect 371577 1019322 371633 1020322
rect 371649 1019322 371705 1020322
rect 372007 1020300 372207 1020322
rect 372222 1020310 372256 1020334
rect 373010 1020322 373044 1020334
rect 372267 1020310 372339 1020322
rect 372222 1020300 372339 1020310
rect 371994 1020276 372339 1020300
rect 372007 1020232 372207 1020276
rect 372222 1020266 372246 1020276
rect 372222 1020242 372256 1020266
rect 372267 1020242 372339 1020276
rect 372222 1020232 372339 1020242
rect 371994 1020208 372339 1020232
rect 372007 1020164 372207 1020208
rect 372222 1020198 372246 1020208
rect 372222 1020174 372256 1020198
rect 372267 1020174 372339 1020208
rect 372222 1020164 372339 1020174
rect 371994 1020140 372339 1020164
rect 372007 1020096 372207 1020140
rect 372222 1020130 372246 1020140
rect 372222 1020106 372256 1020130
rect 372267 1020106 372339 1020140
rect 372222 1020096 372339 1020106
rect 371994 1020072 372339 1020096
rect 372007 1020028 372207 1020072
rect 372222 1020062 372246 1020072
rect 372222 1020038 372256 1020062
rect 372267 1020038 372339 1020072
rect 372222 1020028 372339 1020038
rect 371994 1020004 372339 1020028
rect 372007 1019960 372207 1020004
rect 372222 1019994 372246 1020004
rect 372222 1019970 372256 1019994
rect 372267 1019970 372339 1020004
rect 372222 1019960 372339 1019970
rect 371994 1019936 372339 1019960
rect 372007 1019892 372207 1019936
rect 372222 1019926 372246 1019936
rect 372222 1019902 372256 1019926
rect 372267 1019902 372339 1019936
rect 372222 1019892 372339 1019902
rect 371994 1019868 372339 1019892
rect 372007 1019824 372207 1019868
rect 372222 1019858 372246 1019868
rect 372222 1019834 372256 1019858
rect 372267 1019834 372339 1019868
rect 372222 1019824 372339 1019834
rect 371994 1019800 372339 1019824
rect 372007 1019756 372207 1019800
rect 372222 1019790 372246 1019800
rect 372222 1019766 372256 1019790
rect 372267 1019766 372339 1019800
rect 372222 1019756 372339 1019766
rect 371994 1019732 372339 1019756
rect 372007 1019688 372207 1019732
rect 372222 1019722 372246 1019732
rect 372222 1019698 372256 1019722
rect 372267 1019698 372339 1019732
rect 372222 1019688 372339 1019698
rect 371994 1019664 372339 1019688
rect 372007 1019620 372207 1019664
rect 372222 1019654 372246 1019664
rect 372222 1019630 372256 1019654
rect 372267 1019630 372339 1019664
rect 372222 1019620 372339 1019630
rect 371994 1019596 372339 1019620
rect 372007 1019552 372207 1019596
rect 372222 1019586 372246 1019596
rect 372222 1019562 372256 1019586
rect 372267 1019562 372339 1019596
rect 372222 1019552 372339 1019562
rect 371994 1019528 372339 1019552
rect 372007 1019484 372207 1019528
rect 372222 1019518 372246 1019528
rect 372222 1019494 372256 1019518
rect 372267 1019494 372339 1019528
rect 372222 1019484 372339 1019494
rect 371994 1019460 372339 1019484
rect 372007 1019416 372207 1019460
rect 372222 1019450 372246 1019460
rect 372222 1019426 372256 1019450
rect 372267 1019426 372339 1019460
rect 372222 1019416 372339 1019426
rect 371994 1019392 372339 1019416
rect 372007 1019322 372207 1019392
rect 372222 1019368 372246 1019392
rect 372267 1019322 372339 1019392
rect 372569 1019322 372625 1020322
rect 372641 1019322 372697 1020322
rect 372999 1020300 373199 1020322
rect 373214 1020310 373248 1020334
rect 374002 1020322 374036 1020334
rect 373259 1020310 373331 1020322
rect 373214 1020300 373331 1020310
rect 372986 1020276 373331 1020300
rect 372999 1020232 373199 1020276
rect 373214 1020266 373238 1020276
rect 373214 1020242 373248 1020266
rect 373259 1020242 373331 1020276
rect 373214 1020232 373331 1020242
rect 372986 1020208 373331 1020232
rect 372999 1020164 373199 1020208
rect 373214 1020198 373238 1020208
rect 373214 1020174 373248 1020198
rect 373259 1020174 373331 1020208
rect 373214 1020164 373331 1020174
rect 372986 1020140 373331 1020164
rect 372999 1020096 373199 1020140
rect 373214 1020130 373238 1020140
rect 373214 1020106 373248 1020130
rect 373259 1020106 373331 1020140
rect 373214 1020096 373331 1020106
rect 372986 1020072 373331 1020096
rect 372999 1020028 373199 1020072
rect 373214 1020062 373238 1020072
rect 373214 1020038 373248 1020062
rect 373259 1020038 373331 1020072
rect 373214 1020028 373331 1020038
rect 372986 1020004 373331 1020028
rect 372999 1019960 373199 1020004
rect 373214 1019994 373238 1020004
rect 373214 1019970 373248 1019994
rect 373259 1019970 373331 1020004
rect 373214 1019960 373331 1019970
rect 372986 1019936 373331 1019960
rect 372999 1019892 373199 1019936
rect 373214 1019926 373238 1019936
rect 373214 1019902 373248 1019926
rect 373259 1019902 373331 1019936
rect 373214 1019892 373331 1019902
rect 372986 1019868 373331 1019892
rect 372999 1019824 373199 1019868
rect 373214 1019858 373238 1019868
rect 373214 1019834 373248 1019858
rect 373259 1019834 373331 1019868
rect 373214 1019824 373331 1019834
rect 372986 1019800 373331 1019824
rect 372999 1019756 373199 1019800
rect 373214 1019790 373238 1019800
rect 373214 1019766 373248 1019790
rect 373259 1019766 373331 1019800
rect 373214 1019756 373331 1019766
rect 372986 1019732 373331 1019756
rect 372999 1019688 373199 1019732
rect 373214 1019722 373238 1019732
rect 373214 1019698 373248 1019722
rect 373259 1019698 373331 1019732
rect 373214 1019688 373331 1019698
rect 372986 1019664 373331 1019688
rect 372999 1019620 373199 1019664
rect 373214 1019654 373238 1019664
rect 373214 1019630 373248 1019654
rect 373259 1019630 373331 1019664
rect 373214 1019620 373331 1019630
rect 372986 1019596 373331 1019620
rect 372999 1019552 373199 1019596
rect 373214 1019586 373238 1019596
rect 373214 1019562 373248 1019586
rect 373259 1019562 373331 1019596
rect 373214 1019552 373331 1019562
rect 372986 1019528 373331 1019552
rect 372999 1019484 373199 1019528
rect 373214 1019518 373238 1019528
rect 373214 1019494 373248 1019518
rect 373259 1019494 373331 1019528
rect 373214 1019484 373331 1019494
rect 372986 1019460 373331 1019484
rect 372999 1019416 373199 1019460
rect 373214 1019450 373238 1019460
rect 373214 1019426 373248 1019450
rect 373259 1019426 373331 1019460
rect 373214 1019416 373331 1019426
rect 372986 1019392 373331 1019416
rect 372999 1019322 373199 1019392
rect 373214 1019368 373238 1019392
rect 373259 1019322 373331 1019392
rect 373561 1019322 373617 1020322
rect 373633 1019322 373689 1020322
rect 373991 1020300 374191 1020322
rect 374206 1020310 374240 1020334
rect 374994 1020322 375028 1020334
rect 374251 1020310 374323 1020322
rect 374206 1020300 374323 1020310
rect 373978 1020276 374323 1020300
rect 373991 1020232 374191 1020276
rect 374206 1020266 374230 1020276
rect 374206 1020242 374240 1020266
rect 374251 1020242 374323 1020276
rect 374206 1020232 374323 1020242
rect 373978 1020208 374323 1020232
rect 373991 1020164 374191 1020208
rect 374206 1020198 374230 1020208
rect 374206 1020174 374240 1020198
rect 374251 1020174 374323 1020208
rect 374206 1020164 374323 1020174
rect 373978 1020140 374323 1020164
rect 373991 1020096 374191 1020140
rect 374206 1020130 374230 1020140
rect 374206 1020106 374240 1020130
rect 374251 1020106 374323 1020140
rect 374206 1020096 374323 1020106
rect 373978 1020072 374323 1020096
rect 373991 1020028 374191 1020072
rect 374206 1020062 374230 1020072
rect 374206 1020038 374240 1020062
rect 374251 1020038 374323 1020072
rect 374206 1020028 374323 1020038
rect 373978 1020004 374323 1020028
rect 373991 1019960 374191 1020004
rect 374206 1019994 374230 1020004
rect 374206 1019970 374240 1019994
rect 374251 1019970 374323 1020004
rect 374206 1019960 374323 1019970
rect 373978 1019936 374323 1019960
rect 373991 1019892 374191 1019936
rect 374206 1019926 374230 1019936
rect 374206 1019902 374240 1019926
rect 374251 1019902 374323 1019936
rect 374206 1019892 374323 1019902
rect 373978 1019868 374323 1019892
rect 373991 1019824 374191 1019868
rect 374206 1019858 374230 1019868
rect 374206 1019834 374240 1019858
rect 374251 1019834 374323 1019868
rect 374206 1019824 374323 1019834
rect 373978 1019800 374323 1019824
rect 373991 1019756 374191 1019800
rect 374206 1019790 374230 1019800
rect 374206 1019766 374240 1019790
rect 374251 1019766 374323 1019800
rect 374206 1019756 374323 1019766
rect 373978 1019732 374323 1019756
rect 373991 1019688 374191 1019732
rect 374206 1019722 374230 1019732
rect 374206 1019698 374240 1019722
rect 374251 1019698 374323 1019732
rect 374206 1019688 374323 1019698
rect 373978 1019664 374323 1019688
rect 373991 1019620 374191 1019664
rect 374206 1019654 374230 1019664
rect 374206 1019630 374240 1019654
rect 374251 1019630 374323 1019664
rect 374206 1019620 374323 1019630
rect 373978 1019596 374323 1019620
rect 373991 1019552 374191 1019596
rect 374206 1019586 374230 1019596
rect 374206 1019562 374240 1019586
rect 374251 1019562 374323 1019596
rect 374206 1019552 374323 1019562
rect 373978 1019528 374323 1019552
rect 373991 1019484 374191 1019528
rect 374206 1019518 374230 1019528
rect 374206 1019494 374240 1019518
rect 374251 1019494 374323 1019528
rect 374206 1019484 374323 1019494
rect 373978 1019460 374323 1019484
rect 373991 1019416 374191 1019460
rect 374206 1019450 374230 1019460
rect 374206 1019426 374240 1019450
rect 374251 1019426 374323 1019460
rect 374206 1019416 374323 1019426
rect 373978 1019392 374323 1019416
rect 373991 1019322 374191 1019392
rect 374206 1019368 374230 1019392
rect 374251 1019322 374323 1019392
rect 374553 1019322 374609 1020322
rect 374625 1019322 374681 1020322
rect 374983 1020300 375183 1020322
rect 375198 1020310 375232 1020334
rect 375986 1020322 376020 1020334
rect 375243 1020310 375315 1020322
rect 375198 1020300 375315 1020310
rect 374970 1020276 375315 1020300
rect 374983 1020232 375183 1020276
rect 375198 1020266 375222 1020276
rect 375198 1020242 375232 1020266
rect 375243 1020242 375315 1020276
rect 375198 1020232 375315 1020242
rect 374970 1020208 375315 1020232
rect 374983 1020164 375183 1020208
rect 375198 1020198 375222 1020208
rect 375198 1020174 375232 1020198
rect 375243 1020174 375315 1020208
rect 375198 1020164 375315 1020174
rect 374970 1020140 375315 1020164
rect 374983 1020096 375183 1020140
rect 375198 1020130 375222 1020140
rect 375198 1020106 375232 1020130
rect 375243 1020106 375315 1020140
rect 375198 1020096 375315 1020106
rect 374970 1020072 375315 1020096
rect 374983 1020028 375183 1020072
rect 375198 1020062 375222 1020072
rect 375198 1020038 375232 1020062
rect 375243 1020038 375315 1020072
rect 375198 1020028 375315 1020038
rect 374970 1020004 375315 1020028
rect 374983 1019960 375183 1020004
rect 375198 1019994 375222 1020004
rect 375198 1019970 375232 1019994
rect 375243 1019970 375315 1020004
rect 375198 1019960 375315 1019970
rect 374970 1019936 375315 1019960
rect 374983 1019892 375183 1019936
rect 375198 1019926 375222 1019936
rect 375198 1019902 375232 1019926
rect 375243 1019902 375315 1019936
rect 375198 1019892 375315 1019902
rect 374970 1019868 375315 1019892
rect 374983 1019824 375183 1019868
rect 375198 1019858 375222 1019868
rect 375198 1019834 375232 1019858
rect 375243 1019834 375315 1019868
rect 375198 1019824 375315 1019834
rect 374970 1019800 375315 1019824
rect 374983 1019756 375183 1019800
rect 375198 1019790 375222 1019800
rect 375198 1019766 375232 1019790
rect 375243 1019766 375315 1019800
rect 375198 1019756 375315 1019766
rect 374970 1019732 375315 1019756
rect 374983 1019688 375183 1019732
rect 375198 1019722 375222 1019732
rect 375198 1019698 375232 1019722
rect 375243 1019698 375315 1019732
rect 375198 1019688 375315 1019698
rect 374970 1019664 375315 1019688
rect 374983 1019620 375183 1019664
rect 375198 1019654 375222 1019664
rect 375198 1019630 375232 1019654
rect 375243 1019630 375315 1019664
rect 375198 1019620 375315 1019630
rect 374970 1019596 375315 1019620
rect 374983 1019552 375183 1019596
rect 375198 1019586 375222 1019596
rect 375198 1019562 375232 1019586
rect 375243 1019562 375315 1019596
rect 375198 1019552 375315 1019562
rect 374970 1019528 375315 1019552
rect 374983 1019484 375183 1019528
rect 375198 1019518 375222 1019528
rect 375198 1019494 375232 1019518
rect 375243 1019494 375315 1019528
rect 375198 1019484 375315 1019494
rect 374970 1019460 375315 1019484
rect 374983 1019416 375183 1019460
rect 375198 1019450 375222 1019460
rect 375198 1019426 375232 1019450
rect 375243 1019426 375315 1019460
rect 375198 1019416 375315 1019426
rect 374970 1019392 375315 1019416
rect 374983 1019322 375183 1019392
rect 375198 1019368 375222 1019392
rect 375243 1019322 375315 1019392
rect 375545 1019322 375601 1020322
rect 375617 1019322 375673 1020322
rect 375975 1020300 376175 1020322
rect 376190 1020310 376224 1020334
rect 376978 1020322 377012 1020334
rect 376235 1020310 376307 1020322
rect 376190 1020300 376307 1020310
rect 375962 1020276 376307 1020300
rect 375975 1020232 376175 1020276
rect 376190 1020266 376214 1020276
rect 376190 1020242 376224 1020266
rect 376235 1020242 376307 1020276
rect 376190 1020232 376307 1020242
rect 375962 1020208 376307 1020232
rect 375975 1020164 376175 1020208
rect 376190 1020198 376214 1020208
rect 376190 1020174 376224 1020198
rect 376235 1020174 376307 1020208
rect 376190 1020164 376307 1020174
rect 375962 1020140 376307 1020164
rect 375975 1020096 376175 1020140
rect 376190 1020130 376214 1020140
rect 376190 1020106 376224 1020130
rect 376235 1020106 376307 1020140
rect 376190 1020096 376307 1020106
rect 375962 1020072 376307 1020096
rect 375975 1020028 376175 1020072
rect 376190 1020062 376214 1020072
rect 376190 1020038 376224 1020062
rect 376235 1020038 376307 1020072
rect 376190 1020028 376307 1020038
rect 375962 1020004 376307 1020028
rect 375975 1019960 376175 1020004
rect 376190 1019994 376214 1020004
rect 376190 1019970 376224 1019994
rect 376235 1019970 376307 1020004
rect 376190 1019960 376307 1019970
rect 375962 1019936 376307 1019960
rect 375975 1019892 376175 1019936
rect 376190 1019926 376214 1019936
rect 376190 1019902 376224 1019926
rect 376235 1019902 376307 1019936
rect 376190 1019892 376307 1019902
rect 375962 1019868 376307 1019892
rect 375975 1019824 376175 1019868
rect 376190 1019858 376214 1019868
rect 376190 1019834 376224 1019858
rect 376235 1019834 376307 1019868
rect 376190 1019824 376307 1019834
rect 375962 1019800 376307 1019824
rect 375975 1019756 376175 1019800
rect 376190 1019790 376214 1019800
rect 376190 1019766 376224 1019790
rect 376235 1019766 376307 1019800
rect 376190 1019756 376307 1019766
rect 375962 1019732 376307 1019756
rect 375975 1019688 376175 1019732
rect 376190 1019722 376214 1019732
rect 376190 1019698 376224 1019722
rect 376235 1019698 376307 1019732
rect 376190 1019688 376307 1019698
rect 375962 1019664 376307 1019688
rect 375975 1019620 376175 1019664
rect 376190 1019654 376214 1019664
rect 376190 1019630 376224 1019654
rect 376235 1019630 376307 1019664
rect 376190 1019620 376307 1019630
rect 375962 1019596 376307 1019620
rect 375975 1019552 376175 1019596
rect 376190 1019586 376214 1019596
rect 376190 1019562 376224 1019586
rect 376235 1019562 376307 1019596
rect 376190 1019552 376307 1019562
rect 375962 1019528 376307 1019552
rect 375975 1019484 376175 1019528
rect 376190 1019518 376214 1019528
rect 376190 1019494 376224 1019518
rect 376235 1019494 376307 1019528
rect 376190 1019484 376307 1019494
rect 375962 1019460 376307 1019484
rect 375975 1019416 376175 1019460
rect 376190 1019450 376214 1019460
rect 376190 1019426 376224 1019450
rect 376235 1019426 376307 1019460
rect 376190 1019416 376307 1019426
rect 375962 1019392 376307 1019416
rect 375975 1019322 376175 1019392
rect 376190 1019368 376214 1019392
rect 376235 1019322 376307 1019392
rect 376537 1019322 376593 1020322
rect 376609 1019322 376665 1020322
rect 376967 1020300 377167 1020322
rect 377182 1020310 377216 1020334
rect 377970 1020322 378004 1020334
rect 377227 1020310 377299 1020322
rect 377182 1020300 377299 1020310
rect 376954 1020276 377299 1020300
rect 376967 1020232 377167 1020276
rect 377182 1020266 377206 1020276
rect 377182 1020242 377216 1020266
rect 377227 1020242 377299 1020276
rect 377182 1020232 377299 1020242
rect 376954 1020208 377299 1020232
rect 376967 1020164 377167 1020208
rect 377182 1020198 377206 1020208
rect 377182 1020174 377216 1020198
rect 377227 1020174 377299 1020208
rect 377182 1020164 377299 1020174
rect 376954 1020140 377299 1020164
rect 376967 1020096 377167 1020140
rect 377182 1020130 377206 1020140
rect 377182 1020106 377216 1020130
rect 377227 1020106 377299 1020140
rect 377182 1020096 377299 1020106
rect 376954 1020072 377299 1020096
rect 376967 1020028 377167 1020072
rect 377182 1020062 377206 1020072
rect 377182 1020038 377216 1020062
rect 377227 1020038 377299 1020072
rect 377182 1020028 377299 1020038
rect 376954 1020004 377299 1020028
rect 376967 1019960 377167 1020004
rect 377182 1019994 377206 1020004
rect 377182 1019970 377216 1019994
rect 377227 1019970 377299 1020004
rect 377182 1019960 377299 1019970
rect 376954 1019936 377299 1019960
rect 376967 1019892 377167 1019936
rect 377182 1019926 377206 1019936
rect 377182 1019902 377216 1019926
rect 377227 1019902 377299 1019936
rect 377182 1019892 377299 1019902
rect 376954 1019868 377299 1019892
rect 376967 1019824 377167 1019868
rect 377182 1019858 377206 1019868
rect 377182 1019834 377216 1019858
rect 377227 1019834 377299 1019868
rect 377182 1019824 377299 1019834
rect 376954 1019800 377299 1019824
rect 376967 1019756 377167 1019800
rect 377182 1019790 377206 1019800
rect 377182 1019766 377216 1019790
rect 377227 1019766 377299 1019800
rect 377182 1019756 377299 1019766
rect 376954 1019732 377299 1019756
rect 376967 1019688 377167 1019732
rect 377182 1019722 377206 1019732
rect 377182 1019698 377216 1019722
rect 377227 1019698 377299 1019732
rect 377182 1019688 377299 1019698
rect 376954 1019664 377299 1019688
rect 376967 1019620 377167 1019664
rect 377182 1019654 377206 1019664
rect 377182 1019630 377216 1019654
rect 377227 1019630 377299 1019664
rect 377182 1019620 377299 1019630
rect 376954 1019596 377299 1019620
rect 376967 1019552 377167 1019596
rect 377182 1019586 377206 1019596
rect 377182 1019562 377216 1019586
rect 377227 1019562 377299 1019596
rect 377182 1019552 377299 1019562
rect 376954 1019528 377299 1019552
rect 376967 1019484 377167 1019528
rect 377182 1019518 377206 1019528
rect 377182 1019494 377216 1019518
rect 377227 1019494 377299 1019528
rect 377182 1019484 377299 1019494
rect 376954 1019460 377299 1019484
rect 376967 1019416 377167 1019460
rect 377182 1019450 377206 1019460
rect 377182 1019426 377216 1019450
rect 377227 1019426 377299 1019460
rect 377182 1019416 377299 1019426
rect 376954 1019392 377299 1019416
rect 376967 1019322 377167 1019392
rect 377182 1019368 377206 1019392
rect 377227 1019322 377299 1019392
rect 377529 1019322 377585 1020322
rect 377601 1019322 377657 1020322
rect 377959 1020300 378159 1020322
rect 378174 1020310 378208 1020334
rect 378962 1020322 378996 1020334
rect 378219 1020310 378291 1020322
rect 378174 1020300 378291 1020310
rect 377946 1020276 378291 1020300
rect 377959 1020232 378159 1020276
rect 378174 1020266 378198 1020276
rect 378174 1020242 378208 1020266
rect 378219 1020242 378291 1020276
rect 378174 1020232 378291 1020242
rect 377946 1020208 378291 1020232
rect 377959 1020164 378159 1020208
rect 378174 1020198 378198 1020208
rect 378174 1020174 378208 1020198
rect 378219 1020174 378291 1020208
rect 378174 1020164 378291 1020174
rect 377946 1020140 378291 1020164
rect 377959 1020096 378159 1020140
rect 378174 1020130 378198 1020140
rect 378174 1020106 378208 1020130
rect 378219 1020106 378291 1020140
rect 378174 1020096 378291 1020106
rect 377946 1020072 378291 1020096
rect 377959 1020028 378159 1020072
rect 378174 1020062 378198 1020072
rect 378174 1020038 378208 1020062
rect 378219 1020038 378291 1020072
rect 378174 1020028 378291 1020038
rect 377946 1020004 378291 1020028
rect 377959 1019960 378159 1020004
rect 378174 1019994 378198 1020004
rect 378174 1019970 378208 1019994
rect 378219 1019970 378291 1020004
rect 378174 1019960 378291 1019970
rect 377946 1019936 378291 1019960
rect 377959 1019892 378159 1019936
rect 378174 1019926 378198 1019936
rect 378174 1019902 378208 1019926
rect 378219 1019902 378291 1019936
rect 378174 1019892 378291 1019902
rect 377946 1019868 378291 1019892
rect 377959 1019824 378159 1019868
rect 378174 1019858 378198 1019868
rect 378174 1019834 378208 1019858
rect 378219 1019834 378291 1019868
rect 378174 1019824 378291 1019834
rect 377946 1019800 378291 1019824
rect 377959 1019756 378159 1019800
rect 378174 1019790 378198 1019800
rect 378174 1019766 378208 1019790
rect 378219 1019766 378291 1019800
rect 378174 1019756 378291 1019766
rect 377946 1019732 378291 1019756
rect 377959 1019688 378159 1019732
rect 378174 1019722 378198 1019732
rect 378174 1019698 378208 1019722
rect 378219 1019698 378291 1019732
rect 378174 1019688 378291 1019698
rect 377946 1019664 378291 1019688
rect 377959 1019620 378159 1019664
rect 378174 1019654 378198 1019664
rect 378174 1019630 378208 1019654
rect 378219 1019630 378291 1019664
rect 378174 1019620 378291 1019630
rect 377946 1019596 378291 1019620
rect 377959 1019552 378159 1019596
rect 378174 1019586 378198 1019596
rect 378174 1019562 378208 1019586
rect 378219 1019562 378291 1019596
rect 378174 1019552 378291 1019562
rect 377946 1019528 378291 1019552
rect 377959 1019484 378159 1019528
rect 378174 1019518 378198 1019528
rect 378174 1019494 378208 1019518
rect 378219 1019494 378291 1019528
rect 378174 1019484 378291 1019494
rect 377946 1019460 378291 1019484
rect 377959 1019416 378159 1019460
rect 378174 1019450 378198 1019460
rect 378174 1019426 378208 1019450
rect 378219 1019426 378291 1019460
rect 378174 1019416 378291 1019426
rect 377946 1019392 378291 1019416
rect 377959 1019322 378159 1019392
rect 378174 1019368 378198 1019392
rect 378219 1019322 378291 1019392
rect 378521 1019322 378577 1020322
rect 378593 1019322 378649 1020322
rect 378951 1020300 379151 1020322
rect 379166 1020310 379200 1020334
rect 379211 1020310 379283 1020322
rect 379166 1020300 379283 1020310
rect 378938 1020276 379283 1020300
rect 378951 1020232 379151 1020276
rect 379166 1020266 379190 1020276
rect 379166 1020242 379200 1020266
rect 379211 1020242 379283 1020276
rect 379166 1020232 379283 1020242
rect 378938 1020208 379283 1020232
rect 378951 1020164 379151 1020208
rect 379166 1020198 379190 1020208
rect 379166 1020174 379200 1020198
rect 379211 1020174 379283 1020208
rect 379166 1020164 379283 1020174
rect 378938 1020140 379283 1020164
rect 378951 1020096 379151 1020140
rect 379166 1020130 379190 1020140
rect 379166 1020106 379200 1020130
rect 379211 1020106 379283 1020140
rect 379166 1020096 379283 1020106
rect 378938 1020072 379283 1020096
rect 378951 1020028 379151 1020072
rect 379166 1020062 379190 1020072
rect 379166 1020038 379200 1020062
rect 379211 1020038 379283 1020072
rect 379166 1020028 379283 1020038
rect 378938 1020004 379283 1020028
rect 378951 1019960 379151 1020004
rect 379166 1019994 379190 1020004
rect 379166 1019970 379200 1019994
rect 379211 1019970 379283 1020004
rect 379166 1019960 379283 1019970
rect 378938 1019936 379283 1019960
rect 378951 1019892 379151 1019936
rect 379166 1019926 379190 1019936
rect 379166 1019902 379200 1019926
rect 379211 1019902 379283 1019936
rect 379166 1019892 379283 1019902
rect 378938 1019868 379283 1019892
rect 378951 1019824 379151 1019868
rect 379166 1019858 379190 1019868
rect 379166 1019834 379200 1019858
rect 379211 1019834 379283 1019868
rect 379166 1019824 379283 1019834
rect 378938 1019800 379283 1019824
rect 378951 1019756 379151 1019800
rect 379166 1019790 379190 1019800
rect 379166 1019766 379200 1019790
rect 379211 1019766 379283 1019800
rect 379166 1019756 379283 1019766
rect 378938 1019732 379283 1019756
rect 378951 1019688 379151 1019732
rect 379166 1019722 379190 1019732
rect 379166 1019698 379200 1019722
rect 379211 1019698 379283 1019732
rect 379166 1019688 379283 1019698
rect 378938 1019664 379283 1019688
rect 378951 1019620 379151 1019664
rect 379166 1019654 379190 1019664
rect 379166 1019630 379200 1019654
rect 379211 1019630 379283 1019664
rect 379166 1019620 379283 1019630
rect 378938 1019596 379283 1019620
rect 378951 1019552 379151 1019596
rect 379166 1019586 379190 1019596
rect 379166 1019562 379200 1019586
rect 379211 1019562 379283 1019596
rect 379166 1019552 379283 1019562
rect 378938 1019528 379283 1019552
rect 378951 1019484 379151 1019528
rect 379166 1019518 379190 1019528
rect 379166 1019494 379200 1019518
rect 379211 1019494 379283 1019528
rect 379166 1019484 379283 1019494
rect 378938 1019460 379283 1019484
rect 378951 1019416 379151 1019460
rect 379166 1019450 379190 1019460
rect 379166 1019426 379200 1019450
rect 379211 1019426 379283 1019460
rect 379166 1019416 379283 1019426
rect 378938 1019392 379283 1019416
rect 378951 1019322 379151 1019392
rect 379166 1019368 379190 1019392
rect 379211 1019322 379283 1019392
rect 379472 1019322 379544 1020322
rect 379610 1019322 379627 1020322
rect 379797 1019322 379830 1020322
rect 413561 1018210 413668 1022756
rect 414356 1020922 414406 1021922
rect 414617 1020922 414673 1021922
rect 414689 1020922 414745 1021922
rect 415107 1020922 415247 1021922
rect 426521 1020922 426577 1021922
rect 426593 1020922 426649 1021922
rect 427011 1020922 427151 1021922
rect 427473 1020922 427544 1021922
rect 427610 1020922 427627 1021922
rect 427797 1020922 427830 1021922
rect 427953 1021730 428025 1021760
rect 427953 1021692 427987 1021722
rect 414356 1019322 414406 1020322
rect 414617 1019322 414673 1020322
rect 414689 1019322 414745 1020322
rect 415107 1019322 415247 1020322
rect 426521 1019322 426577 1020322
rect 426593 1019322 426649 1020322
rect 427011 1019322 427151 1020322
rect 427473 1019322 427544 1020322
rect 427610 1019322 427627 1020322
rect 427797 1019322 427830 1020322
rect 465561 1018210 465668 1022756
rect 466356 1020922 466406 1021922
rect 466617 1020922 466673 1021922
rect 466689 1020922 466745 1021922
rect 467047 1021842 467247 1021922
rect 467262 1021852 467296 1021876
rect 467307 1021852 467379 1021922
rect 467262 1021842 467379 1021852
rect 467034 1021818 467379 1021842
rect 467047 1021774 467247 1021818
rect 467262 1021808 467286 1021818
rect 467262 1021784 467296 1021808
rect 467307 1021784 467379 1021818
rect 467262 1021774 467379 1021784
rect 467034 1021750 467379 1021774
rect 467047 1021706 467247 1021750
rect 467262 1021740 467286 1021750
rect 467262 1021716 467296 1021740
rect 467307 1021716 467379 1021750
rect 467262 1021706 467379 1021716
rect 467034 1021682 467379 1021706
rect 467047 1021638 467247 1021682
rect 467262 1021672 467286 1021682
rect 467262 1021648 467296 1021672
rect 467307 1021648 467379 1021682
rect 467262 1021638 467379 1021648
rect 467034 1021614 467379 1021638
rect 467047 1021570 467247 1021614
rect 467262 1021604 467286 1021614
rect 467262 1021580 467296 1021604
rect 467307 1021580 467379 1021614
rect 467262 1021570 467379 1021580
rect 467034 1021546 467379 1021570
rect 467047 1021502 467247 1021546
rect 467262 1021536 467286 1021546
rect 467262 1021512 467296 1021536
rect 467307 1021512 467379 1021546
rect 467262 1021502 467379 1021512
rect 467034 1021478 467379 1021502
rect 467047 1021434 467247 1021478
rect 467262 1021468 467286 1021478
rect 467262 1021444 467296 1021468
rect 467307 1021444 467379 1021478
rect 467262 1021434 467379 1021444
rect 467034 1021410 467379 1021434
rect 467047 1021366 467247 1021410
rect 467262 1021400 467286 1021410
rect 467262 1021376 467296 1021400
rect 467307 1021376 467379 1021410
rect 467262 1021366 467379 1021376
rect 467034 1021342 467379 1021366
rect 467047 1021298 467247 1021342
rect 467262 1021332 467286 1021342
rect 467262 1021308 467296 1021332
rect 467307 1021308 467379 1021342
rect 467262 1021298 467379 1021308
rect 467034 1021274 467379 1021298
rect 467047 1021230 467247 1021274
rect 467262 1021264 467286 1021274
rect 467262 1021240 467296 1021264
rect 467307 1021240 467379 1021274
rect 467262 1021230 467379 1021240
rect 467034 1021206 467379 1021230
rect 467047 1021162 467247 1021206
rect 467262 1021196 467286 1021206
rect 467262 1021172 467296 1021196
rect 467307 1021172 467379 1021206
rect 467262 1021162 467379 1021172
rect 467034 1021138 467379 1021162
rect 467047 1021094 467247 1021138
rect 467262 1021128 467286 1021138
rect 467262 1021104 467296 1021128
rect 467307 1021104 467379 1021138
rect 467262 1021094 467379 1021104
rect 467034 1021070 467379 1021094
rect 467047 1021026 467247 1021070
rect 467262 1021060 467286 1021070
rect 467262 1021036 467296 1021060
rect 467307 1021036 467379 1021070
rect 467262 1021026 467379 1021036
rect 467034 1021002 467379 1021026
rect 467047 1020958 467247 1021002
rect 467262 1020992 467286 1021002
rect 467262 1020968 467296 1020992
rect 467307 1020968 467379 1021002
rect 467262 1020958 467379 1020968
rect 467034 1020934 467379 1020958
rect 467047 1020922 467247 1020934
rect 467058 1020910 467082 1020922
rect 467262 1020910 467286 1020934
rect 467307 1020922 467379 1020934
rect 467609 1020922 467665 1021922
rect 467681 1020922 467737 1021922
rect 468039 1021842 468239 1021922
rect 468254 1021852 468288 1021876
rect 468299 1021852 468371 1021922
rect 468254 1021842 468371 1021852
rect 468026 1021818 468371 1021842
rect 468039 1021774 468239 1021818
rect 468254 1021808 468278 1021818
rect 468254 1021784 468288 1021808
rect 468299 1021784 468371 1021818
rect 468254 1021774 468371 1021784
rect 468026 1021750 468371 1021774
rect 468039 1021706 468239 1021750
rect 468254 1021740 468278 1021750
rect 468254 1021716 468288 1021740
rect 468299 1021716 468371 1021750
rect 468254 1021706 468371 1021716
rect 468026 1021682 468371 1021706
rect 468039 1021638 468239 1021682
rect 468254 1021672 468278 1021682
rect 468254 1021648 468288 1021672
rect 468299 1021648 468371 1021682
rect 468254 1021638 468371 1021648
rect 468026 1021614 468371 1021638
rect 468039 1021570 468239 1021614
rect 468254 1021604 468278 1021614
rect 468254 1021580 468288 1021604
rect 468299 1021580 468371 1021614
rect 468254 1021570 468371 1021580
rect 468026 1021546 468371 1021570
rect 468039 1021502 468239 1021546
rect 468254 1021536 468278 1021546
rect 468254 1021512 468288 1021536
rect 468299 1021512 468371 1021546
rect 468254 1021502 468371 1021512
rect 468026 1021478 468371 1021502
rect 468039 1021434 468239 1021478
rect 468254 1021468 468278 1021478
rect 468254 1021444 468288 1021468
rect 468299 1021444 468371 1021478
rect 468254 1021434 468371 1021444
rect 468026 1021410 468371 1021434
rect 468039 1021366 468239 1021410
rect 468254 1021400 468278 1021410
rect 468254 1021376 468288 1021400
rect 468299 1021376 468371 1021410
rect 468254 1021366 468371 1021376
rect 468026 1021342 468371 1021366
rect 468039 1021298 468239 1021342
rect 468254 1021332 468278 1021342
rect 468254 1021308 468288 1021332
rect 468299 1021308 468371 1021342
rect 468254 1021298 468371 1021308
rect 468026 1021274 468371 1021298
rect 468039 1021230 468239 1021274
rect 468254 1021264 468278 1021274
rect 468254 1021240 468288 1021264
rect 468299 1021240 468371 1021274
rect 468254 1021230 468371 1021240
rect 468026 1021206 468371 1021230
rect 468039 1021162 468239 1021206
rect 468254 1021196 468278 1021206
rect 468254 1021172 468288 1021196
rect 468299 1021172 468371 1021206
rect 468254 1021162 468371 1021172
rect 468026 1021138 468371 1021162
rect 468039 1021094 468239 1021138
rect 468254 1021128 468278 1021138
rect 468254 1021104 468288 1021128
rect 468299 1021104 468371 1021138
rect 468254 1021094 468371 1021104
rect 468026 1021070 468371 1021094
rect 468039 1021026 468239 1021070
rect 468254 1021060 468278 1021070
rect 468254 1021036 468288 1021060
rect 468299 1021036 468371 1021070
rect 468254 1021026 468371 1021036
rect 468026 1021002 468371 1021026
rect 468039 1020958 468239 1021002
rect 468254 1020992 468278 1021002
rect 468254 1020968 468288 1020992
rect 468299 1020968 468371 1021002
rect 468254 1020958 468371 1020968
rect 468026 1020934 468371 1020958
rect 468039 1020922 468239 1020934
rect 468050 1020910 468074 1020922
rect 468254 1020910 468278 1020934
rect 468299 1020922 468371 1020934
rect 468601 1020922 468657 1021922
rect 468673 1020922 468729 1021922
rect 469031 1021842 469231 1021922
rect 469246 1021852 469280 1021876
rect 469291 1021852 469363 1021922
rect 469246 1021842 469363 1021852
rect 469018 1021818 469363 1021842
rect 469031 1021774 469231 1021818
rect 469246 1021808 469270 1021818
rect 469246 1021784 469280 1021808
rect 469291 1021784 469363 1021818
rect 469246 1021774 469363 1021784
rect 469018 1021750 469363 1021774
rect 469031 1021706 469231 1021750
rect 469246 1021740 469270 1021750
rect 469246 1021716 469280 1021740
rect 469291 1021716 469363 1021750
rect 469246 1021706 469363 1021716
rect 469018 1021682 469363 1021706
rect 469031 1021638 469231 1021682
rect 469246 1021672 469270 1021682
rect 469246 1021648 469280 1021672
rect 469291 1021648 469363 1021682
rect 469246 1021638 469363 1021648
rect 469018 1021614 469363 1021638
rect 469031 1021570 469231 1021614
rect 469246 1021604 469270 1021614
rect 469246 1021580 469280 1021604
rect 469291 1021580 469363 1021614
rect 469246 1021570 469363 1021580
rect 469018 1021546 469363 1021570
rect 469031 1021502 469231 1021546
rect 469246 1021536 469270 1021546
rect 469246 1021512 469280 1021536
rect 469291 1021512 469363 1021546
rect 469246 1021502 469363 1021512
rect 469018 1021478 469363 1021502
rect 469031 1021434 469231 1021478
rect 469246 1021468 469270 1021478
rect 469246 1021444 469280 1021468
rect 469291 1021444 469363 1021478
rect 469246 1021434 469363 1021444
rect 469018 1021410 469363 1021434
rect 469031 1021366 469231 1021410
rect 469246 1021400 469270 1021410
rect 469246 1021376 469280 1021400
rect 469291 1021376 469363 1021410
rect 469246 1021366 469363 1021376
rect 469018 1021342 469363 1021366
rect 469031 1021298 469231 1021342
rect 469246 1021332 469270 1021342
rect 469246 1021308 469280 1021332
rect 469291 1021308 469363 1021342
rect 469246 1021298 469363 1021308
rect 469018 1021274 469363 1021298
rect 469031 1021230 469231 1021274
rect 469246 1021264 469270 1021274
rect 469246 1021240 469280 1021264
rect 469291 1021240 469363 1021274
rect 469246 1021230 469363 1021240
rect 469018 1021206 469363 1021230
rect 469031 1021162 469231 1021206
rect 469246 1021196 469270 1021206
rect 469246 1021172 469280 1021196
rect 469291 1021172 469363 1021206
rect 469246 1021162 469363 1021172
rect 469018 1021138 469363 1021162
rect 469031 1021094 469231 1021138
rect 469246 1021128 469270 1021138
rect 469246 1021104 469280 1021128
rect 469291 1021104 469363 1021138
rect 469246 1021094 469363 1021104
rect 469018 1021070 469363 1021094
rect 469031 1021026 469231 1021070
rect 469246 1021060 469270 1021070
rect 469246 1021036 469280 1021060
rect 469291 1021036 469363 1021070
rect 469246 1021026 469363 1021036
rect 469018 1021002 469363 1021026
rect 469031 1020958 469231 1021002
rect 469246 1020992 469270 1021002
rect 469246 1020968 469280 1020992
rect 469291 1020968 469363 1021002
rect 469246 1020958 469363 1020968
rect 469018 1020934 469363 1020958
rect 469031 1020922 469231 1020934
rect 469042 1020910 469066 1020922
rect 469246 1020910 469270 1020934
rect 469291 1020922 469363 1020934
rect 469593 1020922 469649 1021922
rect 469665 1020922 469721 1021922
rect 470023 1021842 470223 1021922
rect 470238 1021852 470272 1021876
rect 470283 1021852 470355 1021922
rect 470238 1021842 470355 1021852
rect 470010 1021818 470355 1021842
rect 470023 1021774 470223 1021818
rect 470238 1021808 470262 1021818
rect 470238 1021784 470272 1021808
rect 470283 1021784 470355 1021818
rect 470238 1021774 470355 1021784
rect 470010 1021750 470355 1021774
rect 470023 1021706 470223 1021750
rect 470238 1021740 470262 1021750
rect 470238 1021716 470272 1021740
rect 470283 1021716 470355 1021750
rect 470238 1021706 470355 1021716
rect 470010 1021682 470355 1021706
rect 470023 1021638 470223 1021682
rect 470238 1021672 470262 1021682
rect 470238 1021648 470272 1021672
rect 470283 1021648 470355 1021682
rect 470238 1021638 470355 1021648
rect 470010 1021614 470355 1021638
rect 470023 1021570 470223 1021614
rect 470238 1021604 470262 1021614
rect 470238 1021580 470272 1021604
rect 470283 1021580 470355 1021614
rect 470238 1021570 470355 1021580
rect 470010 1021546 470355 1021570
rect 470023 1021502 470223 1021546
rect 470238 1021536 470262 1021546
rect 470238 1021512 470272 1021536
rect 470283 1021512 470355 1021546
rect 470238 1021502 470355 1021512
rect 470010 1021478 470355 1021502
rect 470023 1021434 470223 1021478
rect 470238 1021468 470262 1021478
rect 470238 1021444 470272 1021468
rect 470283 1021444 470355 1021478
rect 470238 1021434 470355 1021444
rect 470010 1021410 470355 1021434
rect 470023 1021366 470223 1021410
rect 470238 1021400 470262 1021410
rect 470238 1021376 470272 1021400
rect 470283 1021376 470355 1021410
rect 470238 1021366 470355 1021376
rect 470010 1021342 470355 1021366
rect 470023 1021298 470223 1021342
rect 470238 1021332 470262 1021342
rect 470238 1021308 470272 1021332
rect 470283 1021308 470355 1021342
rect 470238 1021298 470355 1021308
rect 470010 1021274 470355 1021298
rect 470023 1021230 470223 1021274
rect 470238 1021264 470262 1021274
rect 470238 1021240 470272 1021264
rect 470283 1021240 470355 1021274
rect 470238 1021230 470355 1021240
rect 470010 1021206 470355 1021230
rect 470023 1021162 470223 1021206
rect 470238 1021196 470262 1021206
rect 470238 1021172 470272 1021196
rect 470283 1021172 470355 1021206
rect 470238 1021162 470355 1021172
rect 470010 1021138 470355 1021162
rect 470023 1021094 470223 1021138
rect 470238 1021128 470262 1021138
rect 470238 1021104 470272 1021128
rect 470283 1021104 470355 1021138
rect 470238 1021094 470355 1021104
rect 470010 1021070 470355 1021094
rect 470023 1021026 470223 1021070
rect 470238 1021060 470262 1021070
rect 470238 1021036 470272 1021060
rect 470283 1021036 470355 1021070
rect 470238 1021026 470355 1021036
rect 470010 1021002 470355 1021026
rect 470023 1020958 470223 1021002
rect 470238 1020992 470262 1021002
rect 470238 1020968 470272 1020992
rect 470283 1020968 470355 1021002
rect 470238 1020958 470355 1020968
rect 470010 1020934 470355 1020958
rect 470023 1020922 470223 1020934
rect 470034 1020910 470058 1020922
rect 470238 1020910 470262 1020934
rect 470283 1020922 470355 1020934
rect 470585 1020922 470641 1021922
rect 470657 1020922 470713 1021922
rect 471015 1021842 471215 1021922
rect 471230 1021852 471264 1021876
rect 471275 1021852 471347 1021922
rect 471230 1021842 471347 1021852
rect 471002 1021818 471347 1021842
rect 471015 1021774 471215 1021818
rect 471230 1021808 471254 1021818
rect 471230 1021784 471264 1021808
rect 471275 1021784 471347 1021818
rect 471230 1021774 471347 1021784
rect 471002 1021750 471347 1021774
rect 471015 1021706 471215 1021750
rect 471230 1021740 471254 1021750
rect 471230 1021716 471264 1021740
rect 471275 1021716 471347 1021750
rect 471230 1021706 471347 1021716
rect 471002 1021682 471347 1021706
rect 471015 1021638 471215 1021682
rect 471230 1021672 471254 1021682
rect 471230 1021648 471264 1021672
rect 471275 1021648 471347 1021682
rect 471230 1021638 471347 1021648
rect 471002 1021614 471347 1021638
rect 471015 1021570 471215 1021614
rect 471230 1021604 471254 1021614
rect 471230 1021580 471264 1021604
rect 471275 1021580 471347 1021614
rect 471230 1021570 471347 1021580
rect 471002 1021546 471347 1021570
rect 471015 1021502 471215 1021546
rect 471230 1021536 471254 1021546
rect 471230 1021512 471264 1021536
rect 471275 1021512 471347 1021546
rect 471230 1021502 471347 1021512
rect 471002 1021478 471347 1021502
rect 471015 1021434 471215 1021478
rect 471230 1021468 471254 1021478
rect 471230 1021444 471264 1021468
rect 471275 1021444 471347 1021478
rect 471230 1021434 471347 1021444
rect 471002 1021410 471347 1021434
rect 471015 1021366 471215 1021410
rect 471230 1021400 471254 1021410
rect 471230 1021376 471264 1021400
rect 471275 1021376 471347 1021410
rect 471230 1021366 471347 1021376
rect 471002 1021342 471347 1021366
rect 471015 1021298 471215 1021342
rect 471230 1021332 471254 1021342
rect 471230 1021308 471264 1021332
rect 471275 1021308 471347 1021342
rect 471230 1021298 471347 1021308
rect 471002 1021274 471347 1021298
rect 471015 1021230 471215 1021274
rect 471230 1021264 471254 1021274
rect 471230 1021240 471264 1021264
rect 471275 1021240 471347 1021274
rect 471230 1021230 471347 1021240
rect 471002 1021206 471347 1021230
rect 471015 1021162 471215 1021206
rect 471230 1021196 471254 1021206
rect 471230 1021172 471264 1021196
rect 471275 1021172 471347 1021206
rect 471230 1021162 471347 1021172
rect 471002 1021138 471347 1021162
rect 471015 1021094 471215 1021138
rect 471230 1021128 471254 1021138
rect 471230 1021104 471264 1021128
rect 471275 1021104 471347 1021138
rect 471230 1021094 471347 1021104
rect 471002 1021070 471347 1021094
rect 471015 1021026 471215 1021070
rect 471230 1021060 471254 1021070
rect 471230 1021036 471264 1021060
rect 471275 1021036 471347 1021070
rect 471230 1021026 471347 1021036
rect 471002 1021002 471347 1021026
rect 471015 1020958 471215 1021002
rect 471230 1020992 471254 1021002
rect 471230 1020968 471264 1020992
rect 471275 1020968 471347 1021002
rect 471230 1020958 471347 1020968
rect 471002 1020934 471347 1020958
rect 471015 1020922 471215 1020934
rect 471026 1020910 471050 1020922
rect 471230 1020910 471254 1020934
rect 471275 1020922 471347 1020934
rect 471577 1020922 471633 1021922
rect 471649 1020922 471705 1021922
rect 472007 1021842 472207 1021922
rect 472222 1021852 472256 1021876
rect 472267 1021852 472339 1021922
rect 472222 1021842 472339 1021852
rect 471994 1021818 472339 1021842
rect 472007 1021774 472207 1021818
rect 472222 1021808 472246 1021818
rect 472222 1021784 472256 1021808
rect 472267 1021784 472339 1021818
rect 472222 1021774 472339 1021784
rect 471994 1021750 472339 1021774
rect 472007 1021706 472207 1021750
rect 472222 1021740 472246 1021750
rect 472222 1021716 472256 1021740
rect 472267 1021716 472339 1021750
rect 472222 1021706 472339 1021716
rect 471994 1021682 472339 1021706
rect 472007 1021638 472207 1021682
rect 472222 1021672 472246 1021682
rect 472222 1021648 472256 1021672
rect 472267 1021648 472339 1021682
rect 472222 1021638 472339 1021648
rect 471994 1021614 472339 1021638
rect 472007 1021570 472207 1021614
rect 472222 1021604 472246 1021614
rect 472222 1021580 472256 1021604
rect 472267 1021580 472339 1021614
rect 472222 1021570 472339 1021580
rect 471994 1021546 472339 1021570
rect 472007 1021502 472207 1021546
rect 472222 1021536 472246 1021546
rect 472222 1021512 472256 1021536
rect 472267 1021512 472339 1021546
rect 472222 1021502 472339 1021512
rect 471994 1021478 472339 1021502
rect 472007 1021434 472207 1021478
rect 472222 1021468 472246 1021478
rect 472222 1021444 472256 1021468
rect 472267 1021444 472339 1021478
rect 472222 1021434 472339 1021444
rect 471994 1021410 472339 1021434
rect 472007 1021366 472207 1021410
rect 472222 1021400 472246 1021410
rect 472222 1021376 472256 1021400
rect 472267 1021376 472339 1021410
rect 472222 1021366 472339 1021376
rect 471994 1021342 472339 1021366
rect 472007 1021298 472207 1021342
rect 472222 1021332 472246 1021342
rect 472222 1021308 472256 1021332
rect 472267 1021308 472339 1021342
rect 472222 1021298 472339 1021308
rect 471994 1021274 472339 1021298
rect 472007 1021230 472207 1021274
rect 472222 1021264 472246 1021274
rect 472222 1021240 472256 1021264
rect 472267 1021240 472339 1021274
rect 472222 1021230 472339 1021240
rect 471994 1021206 472339 1021230
rect 472007 1021162 472207 1021206
rect 472222 1021196 472246 1021206
rect 472222 1021172 472256 1021196
rect 472267 1021172 472339 1021206
rect 472222 1021162 472339 1021172
rect 471994 1021138 472339 1021162
rect 472007 1021094 472207 1021138
rect 472222 1021128 472246 1021138
rect 472222 1021104 472256 1021128
rect 472267 1021104 472339 1021138
rect 472222 1021094 472339 1021104
rect 471994 1021070 472339 1021094
rect 472007 1021026 472207 1021070
rect 472222 1021060 472246 1021070
rect 472222 1021036 472256 1021060
rect 472267 1021036 472339 1021070
rect 472222 1021026 472339 1021036
rect 471994 1021002 472339 1021026
rect 472007 1020958 472207 1021002
rect 472222 1020992 472246 1021002
rect 472222 1020968 472256 1020992
rect 472267 1020968 472339 1021002
rect 472222 1020958 472339 1020968
rect 471994 1020934 472339 1020958
rect 472007 1020922 472207 1020934
rect 472018 1020910 472042 1020922
rect 472222 1020910 472246 1020934
rect 472267 1020922 472339 1020934
rect 472569 1020922 472625 1021922
rect 472641 1020922 472697 1021922
rect 472999 1021842 473199 1021922
rect 473214 1021852 473248 1021876
rect 473259 1021852 473331 1021922
rect 473214 1021842 473331 1021852
rect 472986 1021818 473331 1021842
rect 472999 1021774 473199 1021818
rect 473214 1021808 473238 1021818
rect 473214 1021784 473248 1021808
rect 473259 1021784 473331 1021818
rect 473214 1021774 473331 1021784
rect 472986 1021750 473331 1021774
rect 472999 1021706 473199 1021750
rect 473214 1021740 473238 1021750
rect 473214 1021716 473248 1021740
rect 473259 1021716 473331 1021750
rect 473214 1021706 473331 1021716
rect 472986 1021682 473331 1021706
rect 472999 1021638 473199 1021682
rect 473214 1021672 473238 1021682
rect 473214 1021648 473248 1021672
rect 473259 1021648 473331 1021682
rect 473214 1021638 473331 1021648
rect 472986 1021614 473331 1021638
rect 472999 1021570 473199 1021614
rect 473214 1021604 473238 1021614
rect 473214 1021580 473248 1021604
rect 473259 1021580 473331 1021614
rect 473214 1021570 473331 1021580
rect 472986 1021546 473331 1021570
rect 472999 1021502 473199 1021546
rect 473214 1021536 473238 1021546
rect 473214 1021512 473248 1021536
rect 473259 1021512 473331 1021546
rect 473214 1021502 473331 1021512
rect 472986 1021478 473331 1021502
rect 472999 1021434 473199 1021478
rect 473214 1021468 473238 1021478
rect 473214 1021444 473248 1021468
rect 473259 1021444 473331 1021478
rect 473214 1021434 473331 1021444
rect 472986 1021410 473331 1021434
rect 472999 1021366 473199 1021410
rect 473214 1021400 473238 1021410
rect 473214 1021376 473248 1021400
rect 473259 1021376 473331 1021410
rect 473214 1021366 473331 1021376
rect 472986 1021342 473331 1021366
rect 472999 1021298 473199 1021342
rect 473214 1021332 473238 1021342
rect 473214 1021308 473248 1021332
rect 473259 1021308 473331 1021342
rect 473214 1021298 473331 1021308
rect 472986 1021274 473331 1021298
rect 472999 1021230 473199 1021274
rect 473214 1021264 473238 1021274
rect 473214 1021240 473248 1021264
rect 473259 1021240 473331 1021274
rect 473214 1021230 473331 1021240
rect 472986 1021206 473331 1021230
rect 472999 1021162 473199 1021206
rect 473214 1021196 473238 1021206
rect 473214 1021172 473248 1021196
rect 473259 1021172 473331 1021206
rect 473214 1021162 473331 1021172
rect 472986 1021138 473331 1021162
rect 472999 1021094 473199 1021138
rect 473214 1021128 473238 1021138
rect 473214 1021104 473248 1021128
rect 473259 1021104 473331 1021138
rect 473214 1021094 473331 1021104
rect 472986 1021070 473331 1021094
rect 472999 1021026 473199 1021070
rect 473214 1021060 473238 1021070
rect 473214 1021036 473248 1021060
rect 473259 1021036 473331 1021070
rect 473214 1021026 473331 1021036
rect 472986 1021002 473331 1021026
rect 472999 1020958 473199 1021002
rect 473214 1020992 473238 1021002
rect 473214 1020968 473248 1020992
rect 473259 1020968 473331 1021002
rect 473214 1020958 473331 1020968
rect 472986 1020934 473331 1020958
rect 472999 1020922 473199 1020934
rect 473010 1020910 473034 1020922
rect 473214 1020910 473238 1020934
rect 473259 1020922 473331 1020934
rect 473561 1020922 473617 1021922
rect 473633 1020922 473689 1021922
rect 473991 1021842 474191 1021922
rect 474206 1021852 474240 1021876
rect 474251 1021852 474323 1021922
rect 474206 1021842 474323 1021852
rect 473978 1021818 474323 1021842
rect 473991 1021774 474191 1021818
rect 474206 1021808 474230 1021818
rect 474206 1021784 474240 1021808
rect 474251 1021784 474323 1021818
rect 474206 1021774 474323 1021784
rect 473978 1021750 474323 1021774
rect 473991 1021706 474191 1021750
rect 474206 1021740 474230 1021750
rect 474206 1021716 474240 1021740
rect 474251 1021716 474323 1021750
rect 474206 1021706 474323 1021716
rect 473978 1021682 474323 1021706
rect 473991 1021638 474191 1021682
rect 474206 1021672 474230 1021682
rect 474206 1021648 474240 1021672
rect 474251 1021648 474323 1021682
rect 474206 1021638 474323 1021648
rect 473978 1021614 474323 1021638
rect 473991 1021570 474191 1021614
rect 474206 1021604 474230 1021614
rect 474206 1021580 474240 1021604
rect 474251 1021580 474323 1021614
rect 474206 1021570 474323 1021580
rect 473978 1021546 474323 1021570
rect 473991 1021502 474191 1021546
rect 474206 1021536 474230 1021546
rect 474206 1021512 474240 1021536
rect 474251 1021512 474323 1021546
rect 474206 1021502 474323 1021512
rect 473978 1021478 474323 1021502
rect 473991 1021434 474191 1021478
rect 474206 1021468 474230 1021478
rect 474206 1021444 474240 1021468
rect 474251 1021444 474323 1021478
rect 474206 1021434 474323 1021444
rect 473978 1021410 474323 1021434
rect 473991 1021366 474191 1021410
rect 474206 1021400 474230 1021410
rect 474206 1021376 474240 1021400
rect 474251 1021376 474323 1021410
rect 474206 1021366 474323 1021376
rect 473978 1021342 474323 1021366
rect 473991 1021298 474191 1021342
rect 474206 1021332 474230 1021342
rect 474206 1021308 474240 1021332
rect 474251 1021308 474323 1021342
rect 474206 1021298 474323 1021308
rect 473978 1021274 474323 1021298
rect 473991 1021230 474191 1021274
rect 474206 1021264 474230 1021274
rect 474206 1021240 474240 1021264
rect 474251 1021240 474323 1021274
rect 474206 1021230 474323 1021240
rect 473978 1021206 474323 1021230
rect 473991 1021162 474191 1021206
rect 474206 1021196 474230 1021206
rect 474206 1021172 474240 1021196
rect 474251 1021172 474323 1021206
rect 474206 1021162 474323 1021172
rect 473978 1021138 474323 1021162
rect 473991 1021094 474191 1021138
rect 474206 1021128 474230 1021138
rect 474206 1021104 474240 1021128
rect 474251 1021104 474323 1021138
rect 474206 1021094 474323 1021104
rect 473978 1021070 474323 1021094
rect 473991 1021026 474191 1021070
rect 474206 1021060 474230 1021070
rect 474206 1021036 474240 1021060
rect 474251 1021036 474323 1021070
rect 474206 1021026 474323 1021036
rect 473978 1021002 474323 1021026
rect 473991 1020958 474191 1021002
rect 474206 1020992 474230 1021002
rect 474206 1020968 474240 1020992
rect 474251 1020968 474323 1021002
rect 474206 1020958 474323 1020968
rect 473978 1020934 474323 1020958
rect 473991 1020922 474191 1020934
rect 474002 1020910 474026 1020922
rect 474206 1020910 474230 1020934
rect 474251 1020922 474323 1020934
rect 474553 1020922 474609 1021922
rect 474625 1020922 474681 1021922
rect 474983 1021842 475183 1021922
rect 475198 1021852 475232 1021876
rect 475243 1021852 475315 1021922
rect 475198 1021842 475315 1021852
rect 474970 1021818 475315 1021842
rect 474983 1021774 475183 1021818
rect 475198 1021808 475222 1021818
rect 475198 1021784 475232 1021808
rect 475243 1021784 475315 1021818
rect 475198 1021774 475315 1021784
rect 474970 1021750 475315 1021774
rect 474983 1021706 475183 1021750
rect 475198 1021740 475222 1021750
rect 475198 1021716 475232 1021740
rect 475243 1021716 475315 1021750
rect 475198 1021706 475315 1021716
rect 474970 1021682 475315 1021706
rect 474983 1021638 475183 1021682
rect 475198 1021672 475222 1021682
rect 475198 1021648 475232 1021672
rect 475243 1021648 475315 1021682
rect 475198 1021638 475315 1021648
rect 474970 1021614 475315 1021638
rect 474983 1021570 475183 1021614
rect 475198 1021604 475222 1021614
rect 475198 1021580 475232 1021604
rect 475243 1021580 475315 1021614
rect 475198 1021570 475315 1021580
rect 474970 1021546 475315 1021570
rect 474983 1021502 475183 1021546
rect 475198 1021536 475222 1021546
rect 475198 1021512 475232 1021536
rect 475243 1021512 475315 1021546
rect 475198 1021502 475315 1021512
rect 474970 1021478 475315 1021502
rect 474983 1021434 475183 1021478
rect 475198 1021468 475222 1021478
rect 475198 1021444 475232 1021468
rect 475243 1021444 475315 1021478
rect 475198 1021434 475315 1021444
rect 474970 1021410 475315 1021434
rect 474983 1021366 475183 1021410
rect 475198 1021400 475222 1021410
rect 475198 1021376 475232 1021400
rect 475243 1021376 475315 1021410
rect 475198 1021366 475315 1021376
rect 474970 1021342 475315 1021366
rect 474983 1021298 475183 1021342
rect 475198 1021332 475222 1021342
rect 475198 1021308 475232 1021332
rect 475243 1021308 475315 1021342
rect 475198 1021298 475315 1021308
rect 474970 1021274 475315 1021298
rect 474983 1021230 475183 1021274
rect 475198 1021264 475222 1021274
rect 475198 1021240 475232 1021264
rect 475243 1021240 475315 1021274
rect 475198 1021230 475315 1021240
rect 474970 1021206 475315 1021230
rect 474983 1021162 475183 1021206
rect 475198 1021196 475222 1021206
rect 475198 1021172 475232 1021196
rect 475243 1021172 475315 1021206
rect 475198 1021162 475315 1021172
rect 474970 1021138 475315 1021162
rect 474983 1021094 475183 1021138
rect 475198 1021128 475222 1021138
rect 475198 1021104 475232 1021128
rect 475243 1021104 475315 1021138
rect 475198 1021094 475315 1021104
rect 474970 1021070 475315 1021094
rect 474983 1021026 475183 1021070
rect 475198 1021060 475222 1021070
rect 475198 1021036 475232 1021060
rect 475243 1021036 475315 1021070
rect 475198 1021026 475315 1021036
rect 474970 1021002 475315 1021026
rect 474983 1020958 475183 1021002
rect 475198 1020992 475222 1021002
rect 475198 1020968 475232 1020992
rect 475243 1020968 475315 1021002
rect 475198 1020958 475315 1020968
rect 474970 1020934 475315 1020958
rect 474983 1020922 475183 1020934
rect 474994 1020910 475018 1020922
rect 475198 1020910 475222 1020934
rect 475243 1020922 475315 1020934
rect 475545 1020922 475601 1021922
rect 475617 1020922 475673 1021922
rect 475975 1021842 476175 1021922
rect 476190 1021852 476224 1021876
rect 476235 1021852 476307 1021922
rect 476190 1021842 476307 1021852
rect 475962 1021818 476307 1021842
rect 475975 1021774 476175 1021818
rect 476190 1021808 476214 1021818
rect 476190 1021784 476224 1021808
rect 476235 1021784 476307 1021818
rect 476190 1021774 476307 1021784
rect 475962 1021750 476307 1021774
rect 475975 1021706 476175 1021750
rect 476190 1021740 476214 1021750
rect 476190 1021716 476224 1021740
rect 476235 1021716 476307 1021750
rect 476190 1021706 476307 1021716
rect 475962 1021682 476307 1021706
rect 475975 1021638 476175 1021682
rect 476190 1021672 476214 1021682
rect 476190 1021648 476224 1021672
rect 476235 1021648 476307 1021682
rect 476190 1021638 476307 1021648
rect 475962 1021614 476307 1021638
rect 475975 1021570 476175 1021614
rect 476190 1021604 476214 1021614
rect 476190 1021580 476224 1021604
rect 476235 1021580 476307 1021614
rect 476190 1021570 476307 1021580
rect 475962 1021546 476307 1021570
rect 475975 1021502 476175 1021546
rect 476190 1021536 476214 1021546
rect 476190 1021512 476224 1021536
rect 476235 1021512 476307 1021546
rect 476190 1021502 476307 1021512
rect 475962 1021478 476307 1021502
rect 475975 1021434 476175 1021478
rect 476190 1021468 476214 1021478
rect 476190 1021444 476224 1021468
rect 476235 1021444 476307 1021478
rect 476190 1021434 476307 1021444
rect 475962 1021410 476307 1021434
rect 475975 1021366 476175 1021410
rect 476190 1021400 476214 1021410
rect 476190 1021376 476224 1021400
rect 476235 1021376 476307 1021410
rect 476190 1021366 476307 1021376
rect 475962 1021342 476307 1021366
rect 475975 1021298 476175 1021342
rect 476190 1021332 476214 1021342
rect 476190 1021308 476224 1021332
rect 476235 1021308 476307 1021342
rect 476190 1021298 476307 1021308
rect 475962 1021274 476307 1021298
rect 475975 1021230 476175 1021274
rect 476190 1021264 476214 1021274
rect 476190 1021240 476224 1021264
rect 476235 1021240 476307 1021274
rect 476190 1021230 476307 1021240
rect 475962 1021206 476307 1021230
rect 475975 1021162 476175 1021206
rect 476190 1021196 476214 1021206
rect 476190 1021172 476224 1021196
rect 476235 1021172 476307 1021206
rect 476190 1021162 476307 1021172
rect 475962 1021138 476307 1021162
rect 475975 1021094 476175 1021138
rect 476190 1021128 476214 1021138
rect 476190 1021104 476224 1021128
rect 476235 1021104 476307 1021138
rect 476190 1021094 476307 1021104
rect 475962 1021070 476307 1021094
rect 475975 1021026 476175 1021070
rect 476190 1021060 476214 1021070
rect 476190 1021036 476224 1021060
rect 476235 1021036 476307 1021070
rect 476190 1021026 476307 1021036
rect 475962 1021002 476307 1021026
rect 475975 1020958 476175 1021002
rect 476190 1020992 476214 1021002
rect 476190 1020968 476224 1020992
rect 476235 1020968 476307 1021002
rect 476190 1020958 476307 1020968
rect 475962 1020934 476307 1020958
rect 475975 1020922 476175 1020934
rect 475986 1020910 476010 1020922
rect 476190 1020910 476214 1020934
rect 476235 1020922 476307 1020934
rect 476537 1020922 476593 1021922
rect 476609 1020922 476665 1021922
rect 476967 1021842 477167 1021922
rect 477182 1021852 477216 1021876
rect 477227 1021852 477299 1021922
rect 477182 1021842 477299 1021852
rect 476954 1021818 477299 1021842
rect 476967 1021774 477167 1021818
rect 477182 1021808 477206 1021818
rect 477182 1021784 477216 1021808
rect 477227 1021784 477299 1021818
rect 477182 1021774 477299 1021784
rect 476954 1021750 477299 1021774
rect 476967 1021706 477167 1021750
rect 477182 1021740 477206 1021750
rect 477182 1021716 477216 1021740
rect 477227 1021716 477299 1021750
rect 477182 1021706 477299 1021716
rect 476954 1021682 477299 1021706
rect 476967 1021638 477167 1021682
rect 477182 1021672 477206 1021682
rect 477182 1021648 477216 1021672
rect 477227 1021648 477299 1021682
rect 477182 1021638 477299 1021648
rect 476954 1021614 477299 1021638
rect 476967 1021570 477167 1021614
rect 477182 1021604 477206 1021614
rect 477182 1021580 477216 1021604
rect 477227 1021580 477299 1021614
rect 477182 1021570 477299 1021580
rect 476954 1021546 477299 1021570
rect 476967 1021502 477167 1021546
rect 477182 1021536 477206 1021546
rect 477182 1021512 477216 1021536
rect 477227 1021512 477299 1021546
rect 477182 1021502 477299 1021512
rect 476954 1021478 477299 1021502
rect 476967 1021434 477167 1021478
rect 477182 1021468 477206 1021478
rect 477182 1021444 477216 1021468
rect 477227 1021444 477299 1021478
rect 477182 1021434 477299 1021444
rect 476954 1021410 477299 1021434
rect 476967 1021366 477167 1021410
rect 477182 1021400 477206 1021410
rect 477182 1021376 477216 1021400
rect 477227 1021376 477299 1021410
rect 477182 1021366 477299 1021376
rect 476954 1021342 477299 1021366
rect 476967 1021298 477167 1021342
rect 477182 1021332 477206 1021342
rect 477182 1021308 477216 1021332
rect 477227 1021308 477299 1021342
rect 477182 1021298 477299 1021308
rect 476954 1021274 477299 1021298
rect 476967 1021230 477167 1021274
rect 477182 1021264 477206 1021274
rect 477182 1021240 477216 1021264
rect 477227 1021240 477299 1021274
rect 477182 1021230 477299 1021240
rect 476954 1021206 477299 1021230
rect 476967 1021162 477167 1021206
rect 477182 1021196 477206 1021206
rect 477182 1021172 477216 1021196
rect 477227 1021172 477299 1021206
rect 477182 1021162 477299 1021172
rect 476954 1021138 477299 1021162
rect 476967 1021094 477167 1021138
rect 477182 1021128 477206 1021138
rect 477182 1021104 477216 1021128
rect 477227 1021104 477299 1021138
rect 477182 1021094 477299 1021104
rect 476954 1021070 477299 1021094
rect 476967 1021026 477167 1021070
rect 477182 1021060 477206 1021070
rect 477182 1021036 477216 1021060
rect 477227 1021036 477299 1021070
rect 477182 1021026 477299 1021036
rect 476954 1021002 477299 1021026
rect 476967 1020958 477167 1021002
rect 477182 1020992 477206 1021002
rect 477182 1020968 477216 1020992
rect 477227 1020968 477299 1021002
rect 477182 1020958 477299 1020968
rect 476954 1020934 477299 1020958
rect 476967 1020922 477167 1020934
rect 476978 1020910 477002 1020922
rect 477182 1020910 477206 1020934
rect 477227 1020922 477299 1020934
rect 477529 1020922 477585 1021922
rect 477601 1020922 477657 1021922
rect 477959 1021842 478159 1021922
rect 478174 1021852 478208 1021876
rect 478219 1021852 478291 1021922
rect 478174 1021842 478291 1021852
rect 477946 1021818 478291 1021842
rect 477959 1021774 478159 1021818
rect 478174 1021808 478198 1021818
rect 478174 1021784 478208 1021808
rect 478219 1021784 478291 1021818
rect 478174 1021774 478291 1021784
rect 477946 1021750 478291 1021774
rect 477959 1021706 478159 1021750
rect 478174 1021740 478198 1021750
rect 478174 1021716 478208 1021740
rect 478219 1021716 478291 1021750
rect 478174 1021706 478291 1021716
rect 477946 1021682 478291 1021706
rect 477959 1021638 478159 1021682
rect 478174 1021672 478198 1021682
rect 478174 1021648 478208 1021672
rect 478219 1021648 478291 1021682
rect 478174 1021638 478291 1021648
rect 477946 1021614 478291 1021638
rect 477959 1021570 478159 1021614
rect 478174 1021604 478198 1021614
rect 478174 1021580 478208 1021604
rect 478219 1021580 478291 1021614
rect 478174 1021570 478291 1021580
rect 477946 1021546 478291 1021570
rect 477959 1021502 478159 1021546
rect 478174 1021536 478198 1021546
rect 478174 1021512 478208 1021536
rect 478219 1021512 478291 1021546
rect 478174 1021502 478291 1021512
rect 477946 1021478 478291 1021502
rect 477959 1021434 478159 1021478
rect 478174 1021468 478198 1021478
rect 478174 1021444 478208 1021468
rect 478219 1021444 478291 1021478
rect 478174 1021434 478291 1021444
rect 477946 1021410 478291 1021434
rect 477959 1021366 478159 1021410
rect 478174 1021400 478198 1021410
rect 478174 1021376 478208 1021400
rect 478219 1021376 478291 1021410
rect 478174 1021366 478291 1021376
rect 477946 1021342 478291 1021366
rect 477959 1021298 478159 1021342
rect 478174 1021332 478198 1021342
rect 478174 1021308 478208 1021332
rect 478219 1021308 478291 1021342
rect 478174 1021298 478291 1021308
rect 477946 1021274 478291 1021298
rect 477959 1021230 478159 1021274
rect 478174 1021264 478198 1021274
rect 478174 1021240 478208 1021264
rect 478219 1021240 478291 1021274
rect 478174 1021230 478291 1021240
rect 477946 1021206 478291 1021230
rect 477959 1021162 478159 1021206
rect 478174 1021196 478198 1021206
rect 478174 1021172 478208 1021196
rect 478219 1021172 478291 1021206
rect 478174 1021162 478291 1021172
rect 477946 1021138 478291 1021162
rect 477959 1021094 478159 1021138
rect 478174 1021128 478198 1021138
rect 478174 1021104 478208 1021128
rect 478219 1021104 478291 1021138
rect 478174 1021094 478291 1021104
rect 477946 1021070 478291 1021094
rect 477959 1021026 478159 1021070
rect 478174 1021060 478198 1021070
rect 478174 1021036 478208 1021060
rect 478219 1021036 478291 1021070
rect 478174 1021026 478291 1021036
rect 477946 1021002 478291 1021026
rect 477959 1020958 478159 1021002
rect 478174 1020992 478198 1021002
rect 478174 1020968 478208 1020992
rect 478219 1020968 478291 1021002
rect 478174 1020958 478291 1020968
rect 477946 1020934 478291 1020958
rect 477959 1020922 478159 1020934
rect 477970 1020910 477994 1020922
rect 478174 1020910 478198 1020934
rect 478219 1020922 478291 1020934
rect 478521 1020922 478577 1021922
rect 478593 1020922 478649 1021922
rect 478951 1021842 479151 1021922
rect 479166 1021852 479200 1021876
rect 479211 1021852 479283 1021922
rect 479166 1021842 479283 1021852
rect 478938 1021818 479283 1021842
rect 478951 1021774 479151 1021818
rect 479166 1021808 479190 1021818
rect 479166 1021784 479200 1021808
rect 479211 1021784 479283 1021818
rect 479166 1021774 479283 1021784
rect 478938 1021750 479283 1021774
rect 478951 1021706 479151 1021750
rect 479166 1021740 479190 1021750
rect 479166 1021716 479200 1021740
rect 479211 1021716 479283 1021750
rect 479166 1021706 479283 1021716
rect 478938 1021682 479283 1021706
rect 478951 1021638 479151 1021682
rect 479166 1021672 479190 1021682
rect 479166 1021648 479200 1021672
rect 479211 1021648 479283 1021682
rect 479166 1021638 479283 1021648
rect 478938 1021614 479283 1021638
rect 478951 1021570 479151 1021614
rect 479166 1021604 479190 1021614
rect 479166 1021580 479200 1021604
rect 479211 1021580 479283 1021614
rect 479166 1021570 479283 1021580
rect 478938 1021546 479283 1021570
rect 478951 1021502 479151 1021546
rect 479166 1021536 479190 1021546
rect 479166 1021512 479200 1021536
rect 479211 1021512 479283 1021546
rect 479166 1021502 479283 1021512
rect 478938 1021478 479283 1021502
rect 478951 1021434 479151 1021478
rect 479166 1021468 479190 1021478
rect 479166 1021444 479200 1021468
rect 479211 1021444 479283 1021478
rect 479166 1021434 479283 1021444
rect 478938 1021410 479283 1021434
rect 478951 1021366 479151 1021410
rect 479166 1021400 479190 1021410
rect 479166 1021376 479200 1021400
rect 479211 1021376 479283 1021410
rect 479166 1021366 479283 1021376
rect 478938 1021342 479283 1021366
rect 478951 1021298 479151 1021342
rect 479166 1021332 479190 1021342
rect 479166 1021308 479200 1021332
rect 479211 1021308 479283 1021342
rect 479166 1021298 479283 1021308
rect 478938 1021274 479283 1021298
rect 478951 1021230 479151 1021274
rect 479166 1021264 479190 1021274
rect 479166 1021240 479200 1021264
rect 479211 1021240 479283 1021274
rect 479166 1021230 479283 1021240
rect 478938 1021206 479283 1021230
rect 478951 1021162 479151 1021206
rect 479166 1021196 479190 1021206
rect 479166 1021172 479200 1021196
rect 479211 1021172 479283 1021206
rect 479166 1021162 479283 1021172
rect 478938 1021138 479283 1021162
rect 478951 1021094 479151 1021138
rect 479166 1021128 479190 1021138
rect 479166 1021104 479200 1021128
rect 479211 1021104 479283 1021138
rect 479166 1021094 479283 1021104
rect 478938 1021070 479283 1021094
rect 478951 1021026 479151 1021070
rect 479166 1021060 479190 1021070
rect 479166 1021036 479200 1021060
rect 479211 1021036 479283 1021070
rect 479166 1021026 479283 1021036
rect 478938 1021002 479283 1021026
rect 478951 1020958 479151 1021002
rect 479166 1020992 479190 1021002
rect 479166 1020968 479200 1020992
rect 479211 1020968 479283 1021002
rect 479166 1020958 479283 1020968
rect 478938 1020934 479283 1020958
rect 478951 1020922 479151 1020934
rect 478962 1020910 478986 1020922
rect 479166 1020910 479190 1020934
rect 479211 1020922 479283 1020934
rect 479472 1020922 479544 1021922
rect 479610 1020922 479627 1021922
rect 479797 1020922 479830 1021922
rect 479953 1021730 480025 1021760
rect 479953 1021692 479987 1021722
rect 467058 1020322 467092 1020334
rect 466356 1019322 466406 1020322
rect 466617 1019322 466673 1020322
rect 466689 1019322 466745 1020322
rect 467047 1020300 467247 1020322
rect 467262 1020310 467296 1020334
rect 468050 1020322 468084 1020334
rect 467307 1020310 467379 1020322
rect 467262 1020300 467379 1020310
rect 467034 1020276 467379 1020300
rect 467047 1020232 467247 1020276
rect 467262 1020266 467286 1020276
rect 467262 1020242 467296 1020266
rect 467307 1020242 467379 1020276
rect 467262 1020232 467379 1020242
rect 467034 1020208 467379 1020232
rect 467047 1020164 467247 1020208
rect 467262 1020198 467286 1020208
rect 467262 1020174 467296 1020198
rect 467307 1020174 467379 1020208
rect 467262 1020164 467379 1020174
rect 467034 1020140 467379 1020164
rect 467047 1020096 467247 1020140
rect 467262 1020130 467286 1020140
rect 467262 1020106 467296 1020130
rect 467307 1020106 467379 1020140
rect 467262 1020096 467379 1020106
rect 467034 1020072 467379 1020096
rect 467047 1020028 467247 1020072
rect 467262 1020062 467286 1020072
rect 467262 1020038 467296 1020062
rect 467307 1020038 467379 1020072
rect 467262 1020028 467379 1020038
rect 467034 1020004 467379 1020028
rect 467047 1019960 467247 1020004
rect 467262 1019994 467286 1020004
rect 467262 1019970 467296 1019994
rect 467307 1019970 467379 1020004
rect 467262 1019960 467379 1019970
rect 467034 1019936 467379 1019960
rect 467047 1019892 467247 1019936
rect 467262 1019926 467286 1019936
rect 467262 1019902 467296 1019926
rect 467307 1019902 467379 1019936
rect 467262 1019892 467379 1019902
rect 467034 1019868 467379 1019892
rect 467047 1019824 467247 1019868
rect 467262 1019858 467286 1019868
rect 467262 1019834 467296 1019858
rect 467307 1019834 467379 1019868
rect 467262 1019824 467379 1019834
rect 467034 1019800 467379 1019824
rect 467047 1019756 467247 1019800
rect 467262 1019790 467286 1019800
rect 467262 1019766 467296 1019790
rect 467307 1019766 467379 1019800
rect 467262 1019756 467379 1019766
rect 467034 1019732 467379 1019756
rect 467047 1019688 467247 1019732
rect 467262 1019722 467286 1019732
rect 467262 1019698 467296 1019722
rect 467307 1019698 467379 1019732
rect 467262 1019688 467379 1019698
rect 467034 1019664 467379 1019688
rect 467047 1019620 467247 1019664
rect 467262 1019654 467286 1019664
rect 467262 1019630 467296 1019654
rect 467307 1019630 467379 1019664
rect 467262 1019620 467379 1019630
rect 467034 1019596 467379 1019620
rect 467047 1019552 467247 1019596
rect 467262 1019586 467286 1019596
rect 467262 1019562 467296 1019586
rect 467307 1019562 467379 1019596
rect 467262 1019552 467379 1019562
rect 467034 1019528 467379 1019552
rect 467047 1019484 467247 1019528
rect 467262 1019518 467286 1019528
rect 467262 1019494 467296 1019518
rect 467307 1019494 467379 1019528
rect 467262 1019484 467379 1019494
rect 467034 1019460 467379 1019484
rect 467047 1019416 467247 1019460
rect 467262 1019450 467286 1019460
rect 467262 1019426 467296 1019450
rect 467307 1019426 467379 1019460
rect 467262 1019416 467379 1019426
rect 467034 1019392 467379 1019416
rect 467047 1019322 467247 1019392
rect 467262 1019368 467286 1019392
rect 467307 1019322 467379 1019392
rect 467609 1019322 467665 1020322
rect 467681 1019322 467737 1020322
rect 468039 1020300 468239 1020322
rect 468254 1020310 468288 1020334
rect 469042 1020322 469076 1020334
rect 468299 1020310 468371 1020322
rect 468254 1020300 468371 1020310
rect 468026 1020276 468371 1020300
rect 468039 1020232 468239 1020276
rect 468254 1020266 468278 1020276
rect 468254 1020242 468288 1020266
rect 468299 1020242 468371 1020276
rect 468254 1020232 468371 1020242
rect 468026 1020208 468371 1020232
rect 468039 1020164 468239 1020208
rect 468254 1020198 468278 1020208
rect 468254 1020174 468288 1020198
rect 468299 1020174 468371 1020208
rect 468254 1020164 468371 1020174
rect 468026 1020140 468371 1020164
rect 468039 1020096 468239 1020140
rect 468254 1020130 468278 1020140
rect 468254 1020106 468288 1020130
rect 468299 1020106 468371 1020140
rect 468254 1020096 468371 1020106
rect 468026 1020072 468371 1020096
rect 468039 1020028 468239 1020072
rect 468254 1020062 468278 1020072
rect 468254 1020038 468288 1020062
rect 468299 1020038 468371 1020072
rect 468254 1020028 468371 1020038
rect 468026 1020004 468371 1020028
rect 468039 1019960 468239 1020004
rect 468254 1019994 468278 1020004
rect 468254 1019970 468288 1019994
rect 468299 1019970 468371 1020004
rect 468254 1019960 468371 1019970
rect 468026 1019936 468371 1019960
rect 468039 1019892 468239 1019936
rect 468254 1019926 468278 1019936
rect 468254 1019902 468288 1019926
rect 468299 1019902 468371 1019936
rect 468254 1019892 468371 1019902
rect 468026 1019868 468371 1019892
rect 468039 1019824 468239 1019868
rect 468254 1019858 468278 1019868
rect 468254 1019834 468288 1019858
rect 468299 1019834 468371 1019868
rect 468254 1019824 468371 1019834
rect 468026 1019800 468371 1019824
rect 468039 1019756 468239 1019800
rect 468254 1019790 468278 1019800
rect 468254 1019766 468288 1019790
rect 468299 1019766 468371 1019800
rect 468254 1019756 468371 1019766
rect 468026 1019732 468371 1019756
rect 468039 1019688 468239 1019732
rect 468254 1019722 468278 1019732
rect 468254 1019698 468288 1019722
rect 468299 1019698 468371 1019732
rect 468254 1019688 468371 1019698
rect 468026 1019664 468371 1019688
rect 468039 1019620 468239 1019664
rect 468254 1019654 468278 1019664
rect 468254 1019630 468288 1019654
rect 468299 1019630 468371 1019664
rect 468254 1019620 468371 1019630
rect 468026 1019596 468371 1019620
rect 468039 1019552 468239 1019596
rect 468254 1019586 468278 1019596
rect 468254 1019562 468288 1019586
rect 468299 1019562 468371 1019596
rect 468254 1019552 468371 1019562
rect 468026 1019528 468371 1019552
rect 468039 1019484 468239 1019528
rect 468254 1019518 468278 1019528
rect 468254 1019494 468288 1019518
rect 468299 1019494 468371 1019528
rect 468254 1019484 468371 1019494
rect 468026 1019460 468371 1019484
rect 468039 1019416 468239 1019460
rect 468254 1019450 468278 1019460
rect 468254 1019426 468288 1019450
rect 468299 1019426 468371 1019460
rect 468254 1019416 468371 1019426
rect 468026 1019392 468371 1019416
rect 468039 1019322 468239 1019392
rect 468254 1019368 468278 1019392
rect 468299 1019322 468371 1019392
rect 468601 1019322 468657 1020322
rect 468673 1019322 468729 1020322
rect 469031 1020300 469231 1020322
rect 469246 1020310 469280 1020334
rect 470034 1020322 470068 1020334
rect 469291 1020310 469363 1020322
rect 469246 1020300 469363 1020310
rect 469018 1020276 469363 1020300
rect 469031 1020232 469231 1020276
rect 469246 1020266 469270 1020276
rect 469246 1020242 469280 1020266
rect 469291 1020242 469363 1020276
rect 469246 1020232 469363 1020242
rect 469018 1020208 469363 1020232
rect 469031 1020164 469231 1020208
rect 469246 1020198 469270 1020208
rect 469246 1020174 469280 1020198
rect 469291 1020174 469363 1020208
rect 469246 1020164 469363 1020174
rect 469018 1020140 469363 1020164
rect 469031 1020096 469231 1020140
rect 469246 1020130 469270 1020140
rect 469246 1020106 469280 1020130
rect 469291 1020106 469363 1020140
rect 469246 1020096 469363 1020106
rect 469018 1020072 469363 1020096
rect 469031 1020028 469231 1020072
rect 469246 1020062 469270 1020072
rect 469246 1020038 469280 1020062
rect 469291 1020038 469363 1020072
rect 469246 1020028 469363 1020038
rect 469018 1020004 469363 1020028
rect 469031 1019960 469231 1020004
rect 469246 1019994 469270 1020004
rect 469246 1019970 469280 1019994
rect 469291 1019970 469363 1020004
rect 469246 1019960 469363 1019970
rect 469018 1019936 469363 1019960
rect 469031 1019892 469231 1019936
rect 469246 1019926 469270 1019936
rect 469246 1019902 469280 1019926
rect 469291 1019902 469363 1019936
rect 469246 1019892 469363 1019902
rect 469018 1019868 469363 1019892
rect 469031 1019824 469231 1019868
rect 469246 1019858 469270 1019868
rect 469246 1019834 469280 1019858
rect 469291 1019834 469363 1019868
rect 469246 1019824 469363 1019834
rect 469018 1019800 469363 1019824
rect 469031 1019756 469231 1019800
rect 469246 1019790 469270 1019800
rect 469246 1019766 469280 1019790
rect 469291 1019766 469363 1019800
rect 469246 1019756 469363 1019766
rect 469018 1019732 469363 1019756
rect 469031 1019688 469231 1019732
rect 469246 1019722 469270 1019732
rect 469246 1019698 469280 1019722
rect 469291 1019698 469363 1019732
rect 469246 1019688 469363 1019698
rect 469018 1019664 469363 1019688
rect 469031 1019620 469231 1019664
rect 469246 1019654 469270 1019664
rect 469246 1019630 469280 1019654
rect 469291 1019630 469363 1019664
rect 469246 1019620 469363 1019630
rect 469018 1019596 469363 1019620
rect 469031 1019552 469231 1019596
rect 469246 1019586 469270 1019596
rect 469246 1019562 469280 1019586
rect 469291 1019562 469363 1019596
rect 469246 1019552 469363 1019562
rect 469018 1019528 469363 1019552
rect 469031 1019484 469231 1019528
rect 469246 1019518 469270 1019528
rect 469246 1019494 469280 1019518
rect 469291 1019494 469363 1019528
rect 469246 1019484 469363 1019494
rect 469018 1019460 469363 1019484
rect 469031 1019416 469231 1019460
rect 469246 1019450 469270 1019460
rect 469246 1019426 469280 1019450
rect 469291 1019426 469363 1019460
rect 469246 1019416 469363 1019426
rect 469018 1019392 469363 1019416
rect 469031 1019322 469231 1019392
rect 469246 1019368 469270 1019392
rect 469291 1019322 469363 1019392
rect 469593 1019322 469649 1020322
rect 469665 1019322 469721 1020322
rect 470023 1020300 470223 1020322
rect 470238 1020310 470272 1020334
rect 471026 1020322 471060 1020334
rect 470283 1020310 470355 1020322
rect 470238 1020300 470355 1020310
rect 470010 1020276 470355 1020300
rect 470023 1020232 470223 1020276
rect 470238 1020266 470262 1020276
rect 470238 1020242 470272 1020266
rect 470283 1020242 470355 1020276
rect 470238 1020232 470355 1020242
rect 470010 1020208 470355 1020232
rect 470023 1020164 470223 1020208
rect 470238 1020198 470262 1020208
rect 470238 1020174 470272 1020198
rect 470283 1020174 470355 1020208
rect 470238 1020164 470355 1020174
rect 470010 1020140 470355 1020164
rect 470023 1020096 470223 1020140
rect 470238 1020130 470262 1020140
rect 470238 1020106 470272 1020130
rect 470283 1020106 470355 1020140
rect 470238 1020096 470355 1020106
rect 470010 1020072 470355 1020096
rect 470023 1020028 470223 1020072
rect 470238 1020062 470262 1020072
rect 470238 1020038 470272 1020062
rect 470283 1020038 470355 1020072
rect 470238 1020028 470355 1020038
rect 470010 1020004 470355 1020028
rect 470023 1019960 470223 1020004
rect 470238 1019994 470262 1020004
rect 470238 1019970 470272 1019994
rect 470283 1019970 470355 1020004
rect 470238 1019960 470355 1019970
rect 470010 1019936 470355 1019960
rect 470023 1019892 470223 1019936
rect 470238 1019926 470262 1019936
rect 470238 1019902 470272 1019926
rect 470283 1019902 470355 1019936
rect 470238 1019892 470355 1019902
rect 470010 1019868 470355 1019892
rect 470023 1019824 470223 1019868
rect 470238 1019858 470262 1019868
rect 470238 1019834 470272 1019858
rect 470283 1019834 470355 1019868
rect 470238 1019824 470355 1019834
rect 470010 1019800 470355 1019824
rect 470023 1019756 470223 1019800
rect 470238 1019790 470262 1019800
rect 470238 1019766 470272 1019790
rect 470283 1019766 470355 1019800
rect 470238 1019756 470355 1019766
rect 470010 1019732 470355 1019756
rect 470023 1019688 470223 1019732
rect 470238 1019722 470262 1019732
rect 470238 1019698 470272 1019722
rect 470283 1019698 470355 1019732
rect 470238 1019688 470355 1019698
rect 470010 1019664 470355 1019688
rect 470023 1019620 470223 1019664
rect 470238 1019654 470262 1019664
rect 470238 1019630 470272 1019654
rect 470283 1019630 470355 1019664
rect 470238 1019620 470355 1019630
rect 470010 1019596 470355 1019620
rect 470023 1019552 470223 1019596
rect 470238 1019586 470262 1019596
rect 470238 1019562 470272 1019586
rect 470283 1019562 470355 1019596
rect 470238 1019552 470355 1019562
rect 470010 1019528 470355 1019552
rect 470023 1019484 470223 1019528
rect 470238 1019518 470262 1019528
rect 470238 1019494 470272 1019518
rect 470283 1019494 470355 1019528
rect 470238 1019484 470355 1019494
rect 470010 1019460 470355 1019484
rect 470023 1019416 470223 1019460
rect 470238 1019450 470262 1019460
rect 470238 1019426 470272 1019450
rect 470283 1019426 470355 1019460
rect 470238 1019416 470355 1019426
rect 470010 1019392 470355 1019416
rect 470023 1019322 470223 1019392
rect 470238 1019368 470262 1019392
rect 470283 1019322 470355 1019392
rect 470585 1019322 470641 1020322
rect 470657 1019322 470713 1020322
rect 471015 1020300 471215 1020322
rect 471230 1020310 471264 1020334
rect 472018 1020322 472052 1020334
rect 471275 1020310 471347 1020322
rect 471230 1020300 471347 1020310
rect 471002 1020276 471347 1020300
rect 471015 1020232 471215 1020276
rect 471230 1020266 471254 1020276
rect 471230 1020242 471264 1020266
rect 471275 1020242 471347 1020276
rect 471230 1020232 471347 1020242
rect 471002 1020208 471347 1020232
rect 471015 1020164 471215 1020208
rect 471230 1020198 471254 1020208
rect 471230 1020174 471264 1020198
rect 471275 1020174 471347 1020208
rect 471230 1020164 471347 1020174
rect 471002 1020140 471347 1020164
rect 471015 1020096 471215 1020140
rect 471230 1020130 471254 1020140
rect 471230 1020106 471264 1020130
rect 471275 1020106 471347 1020140
rect 471230 1020096 471347 1020106
rect 471002 1020072 471347 1020096
rect 471015 1020028 471215 1020072
rect 471230 1020062 471254 1020072
rect 471230 1020038 471264 1020062
rect 471275 1020038 471347 1020072
rect 471230 1020028 471347 1020038
rect 471002 1020004 471347 1020028
rect 471015 1019960 471215 1020004
rect 471230 1019994 471254 1020004
rect 471230 1019970 471264 1019994
rect 471275 1019970 471347 1020004
rect 471230 1019960 471347 1019970
rect 471002 1019936 471347 1019960
rect 471015 1019892 471215 1019936
rect 471230 1019926 471254 1019936
rect 471230 1019902 471264 1019926
rect 471275 1019902 471347 1019936
rect 471230 1019892 471347 1019902
rect 471002 1019868 471347 1019892
rect 471015 1019824 471215 1019868
rect 471230 1019858 471254 1019868
rect 471230 1019834 471264 1019858
rect 471275 1019834 471347 1019868
rect 471230 1019824 471347 1019834
rect 471002 1019800 471347 1019824
rect 471015 1019756 471215 1019800
rect 471230 1019790 471254 1019800
rect 471230 1019766 471264 1019790
rect 471275 1019766 471347 1019800
rect 471230 1019756 471347 1019766
rect 471002 1019732 471347 1019756
rect 471015 1019688 471215 1019732
rect 471230 1019722 471254 1019732
rect 471230 1019698 471264 1019722
rect 471275 1019698 471347 1019732
rect 471230 1019688 471347 1019698
rect 471002 1019664 471347 1019688
rect 471015 1019620 471215 1019664
rect 471230 1019654 471254 1019664
rect 471230 1019630 471264 1019654
rect 471275 1019630 471347 1019664
rect 471230 1019620 471347 1019630
rect 471002 1019596 471347 1019620
rect 471015 1019552 471215 1019596
rect 471230 1019586 471254 1019596
rect 471230 1019562 471264 1019586
rect 471275 1019562 471347 1019596
rect 471230 1019552 471347 1019562
rect 471002 1019528 471347 1019552
rect 471015 1019484 471215 1019528
rect 471230 1019518 471254 1019528
rect 471230 1019494 471264 1019518
rect 471275 1019494 471347 1019528
rect 471230 1019484 471347 1019494
rect 471002 1019460 471347 1019484
rect 471015 1019416 471215 1019460
rect 471230 1019450 471254 1019460
rect 471230 1019426 471264 1019450
rect 471275 1019426 471347 1019460
rect 471230 1019416 471347 1019426
rect 471002 1019392 471347 1019416
rect 471015 1019322 471215 1019392
rect 471230 1019368 471254 1019392
rect 471275 1019322 471347 1019392
rect 471577 1019322 471633 1020322
rect 471649 1019322 471705 1020322
rect 472007 1020300 472207 1020322
rect 472222 1020310 472256 1020334
rect 473010 1020322 473044 1020334
rect 472267 1020310 472339 1020322
rect 472222 1020300 472339 1020310
rect 471994 1020276 472339 1020300
rect 472007 1020232 472207 1020276
rect 472222 1020266 472246 1020276
rect 472222 1020242 472256 1020266
rect 472267 1020242 472339 1020276
rect 472222 1020232 472339 1020242
rect 471994 1020208 472339 1020232
rect 472007 1020164 472207 1020208
rect 472222 1020198 472246 1020208
rect 472222 1020174 472256 1020198
rect 472267 1020174 472339 1020208
rect 472222 1020164 472339 1020174
rect 471994 1020140 472339 1020164
rect 472007 1020096 472207 1020140
rect 472222 1020130 472246 1020140
rect 472222 1020106 472256 1020130
rect 472267 1020106 472339 1020140
rect 472222 1020096 472339 1020106
rect 471994 1020072 472339 1020096
rect 472007 1020028 472207 1020072
rect 472222 1020062 472246 1020072
rect 472222 1020038 472256 1020062
rect 472267 1020038 472339 1020072
rect 472222 1020028 472339 1020038
rect 471994 1020004 472339 1020028
rect 472007 1019960 472207 1020004
rect 472222 1019994 472246 1020004
rect 472222 1019970 472256 1019994
rect 472267 1019970 472339 1020004
rect 472222 1019960 472339 1019970
rect 471994 1019936 472339 1019960
rect 472007 1019892 472207 1019936
rect 472222 1019926 472246 1019936
rect 472222 1019902 472256 1019926
rect 472267 1019902 472339 1019936
rect 472222 1019892 472339 1019902
rect 471994 1019868 472339 1019892
rect 472007 1019824 472207 1019868
rect 472222 1019858 472246 1019868
rect 472222 1019834 472256 1019858
rect 472267 1019834 472339 1019868
rect 472222 1019824 472339 1019834
rect 471994 1019800 472339 1019824
rect 472007 1019756 472207 1019800
rect 472222 1019790 472246 1019800
rect 472222 1019766 472256 1019790
rect 472267 1019766 472339 1019800
rect 472222 1019756 472339 1019766
rect 471994 1019732 472339 1019756
rect 472007 1019688 472207 1019732
rect 472222 1019722 472246 1019732
rect 472222 1019698 472256 1019722
rect 472267 1019698 472339 1019732
rect 472222 1019688 472339 1019698
rect 471994 1019664 472339 1019688
rect 472007 1019620 472207 1019664
rect 472222 1019654 472246 1019664
rect 472222 1019630 472256 1019654
rect 472267 1019630 472339 1019664
rect 472222 1019620 472339 1019630
rect 471994 1019596 472339 1019620
rect 472007 1019552 472207 1019596
rect 472222 1019586 472246 1019596
rect 472222 1019562 472256 1019586
rect 472267 1019562 472339 1019596
rect 472222 1019552 472339 1019562
rect 471994 1019528 472339 1019552
rect 472007 1019484 472207 1019528
rect 472222 1019518 472246 1019528
rect 472222 1019494 472256 1019518
rect 472267 1019494 472339 1019528
rect 472222 1019484 472339 1019494
rect 471994 1019460 472339 1019484
rect 472007 1019416 472207 1019460
rect 472222 1019450 472246 1019460
rect 472222 1019426 472256 1019450
rect 472267 1019426 472339 1019460
rect 472222 1019416 472339 1019426
rect 471994 1019392 472339 1019416
rect 472007 1019322 472207 1019392
rect 472222 1019368 472246 1019392
rect 472267 1019322 472339 1019392
rect 472569 1019322 472625 1020322
rect 472641 1019322 472697 1020322
rect 472999 1020300 473199 1020322
rect 473214 1020310 473248 1020334
rect 474002 1020322 474036 1020334
rect 473259 1020310 473331 1020322
rect 473214 1020300 473331 1020310
rect 472986 1020276 473331 1020300
rect 472999 1020232 473199 1020276
rect 473214 1020266 473238 1020276
rect 473214 1020242 473248 1020266
rect 473259 1020242 473331 1020276
rect 473214 1020232 473331 1020242
rect 472986 1020208 473331 1020232
rect 472999 1020164 473199 1020208
rect 473214 1020198 473238 1020208
rect 473214 1020174 473248 1020198
rect 473259 1020174 473331 1020208
rect 473214 1020164 473331 1020174
rect 472986 1020140 473331 1020164
rect 472999 1020096 473199 1020140
rect 473214 1020130 473238 1020140
rect 473214 1020106 473248 1020130
rect 473259 1020106 473331 1020140
rect 473214 1020096 473331 1020106
rect 472986 1020072 473331 1020096
rect 472999 1020028 473199 1020072
rect 473214 1020062 473238 1020072
rect 473214 1020038 473248 1020062
rect 473259 1020038 473331 1020072
rect 473214 1020028 473331 1020038
rect 472986 1020004 473331 1020028
rect 472999 1019960 473199 1020004
rect 473214 1019994 473238 1020004
rect 473214 1019970 473248 1019994
rect 473259 1019970 473331 1020004
rect 473214 1019960 473331 1019970
rect 472986 1019936 473331 1019960
rect 472999 1019892 473199 1019936
rect 473214 1019926 473238 1019936
rect 473214 1019902 473248 1019926
rect 473259 1019902 473331 1019936
rect 473214 1019892 473331 1019902
rect 472986 1019868 473331 1019892
rect 472999 1019824 473199 1019868
rect 473214 1019858 473238 1019868
rect 473214 1019834 473248 1019858
rect 473259 1019834 473331 1019868
rect 473214 1019824 473331 1019834
rect 472986 1019800 473331 1019824
rect 472999 1019756 473199 1019800
rect 473214 1019790 473238 1019800
rect 473214 1019766 473248 1019790
rect 473259 1019766 473331 1019800
rect 473214 1019756 473331 1019766
rect 472986 1019732 473331 1019756
rect 472999 1019688 473199 1019732
rect 473214 1019722 473238 1019732
rect 473214 1019698 473248 1019722
rect 473259 1019698 473331 1019732
rect 473214 1019688 473331 1019698
rect 472986 1019664 473331 1019688
rect 472999 1019620 473199 1019664
rect 473214 1019654 473238 1019664
rect 473214 1019630 473248 1019654
rect 473259 1019630 473331 1019664
rect 473214 1019620 473331 1019630
rect 472986 1019596 473331 1019620
rect 472999 1019552 473199 1019596
rect 473214 1019586 473238 1019596
rect 473214 1019562 473248 1019586
rect 473259 1019562 473331 1019596
rect 473214 1019552 473331 1019562
rect 472986 1019528 473331 1019552
rect 472999 1019484 473199 1019528
rect 473214 1019518 473238 1019528
rect 473214 1019494 473248 1019518
rect 473259 1019494 473331 1019528
rect 473214 1019484 473331 1019494
rect 472986 1019460 473331 1019484
rect 472999 1019416 473199 1019460
rect 473214 1019450 473238 1019460
rect 473214 1019426 473248 1019450
rect 473259 1019426 473331 1019460
rect 473214 1019416 473331 1019426
rect 472986 1019392 473331 1019416
rect 472999 1019322 473199 1019392
rect 473214 1019368 473238 1019392
rect 473259 1019322 473331 1019392
rect 473561 1019322 473617 1020322
rect 473633 1019322 473689 1020322
rect 473991 1020300 474191 1020322
rect 474206 1020310 474240 1020334
rect 474994 1020322 475028 1020334
rect 474251 1020310 474323 1020322
rect 474206 1020300 474323 1020310
rect 473978 1020276 474323 1020300
rect 473991 1020232 474191 1020276
rect 474206 1020266 474230 1020276
rect 474206 1020242 474240 1020266
rect 474251 1020242 474323 1020276
rect 474206 1020232 474323 1020242
rect 473978 1020208 474323 1020232
rect 473991 1020164 474191 1020208
rect 474206 1020198 474230 1020208
rect 474206 1020174 474240 1020198
rect 474251 1020174 474323 1020208
rect 474206 1020164 474323 1020174
rect 473978 1020140 474323 1020164
rect 473991 1020096 474191 1020140
rect 474206 1020130 474230 1020140
rect 474206 1020106 474240 1020130
rect 474251 1020106 474323 1020140
rect 474206 1020096 474323 1020106
rect 473978 1020072 474323 1020096
rect 473991 1020028 474191 1020072
rect 474206 1020062 474230 1020072
rect 474206 1020038 474240 1020062
rect 474251 1020038 474323 1020072
rect 474206 1020028 474323 1020038
rect 473978 1020004 474323 1020028
rect 473991 1019960 474191 1020004
rect 474206 1019994 474230 1020004
rect 474206 1019970 474240 1019994
rect 474251 1019970 474323 1020004
rect 474206 1019960 474323 1019970
rect 473978 1019936 474323 1019960
rect 473991 1019892 474191 1019936
rect 474206 1019926 474230 1019936
rect 474206 1019902 474240 1019926
rect 474251 1019902 474323 1019936
rect 474206 1019892 474323 1019902
rect 473978 1019868 474323 1019892
rect 473991 1019824 474191 1019868
rect 474206 1019858 474230 1019868
rect 474206 1019834 474240 1019858
rect 474251 1019834 474323 1019868
rect 474206 1019824 474323 1019834
rect 473978 1019800 474323 1019824
rect 473991 1019756 474191 1019800
rect 474206 1019790 474230 1019800
rect 474206 1019766 474240 1019790
rect 474251 1019766 474323 1019800
rect 474206 1019756 474323 1019766
rect 473978 1019732 474323 1019756
rect 473991 1019688 474191 1019732
rect 474206 1019722 474230 1019732
rect 474206 1019698 474240 1019722
rect 474251 1019698 474323 1019732
rect 474206 1019688 474323 1019698
rect 473978 1019664 474323 1019688
rect 473991 1019620 474191 1019664
rect 474206 1019654 474230 1019664
rect 474206 1019630 474240 1019654
rect 474251 1019630 474323 1019664
rect 474206 1019620 474323 1019630
rect 473978 1019596 474323 1019620
rect 473991 1019552 474191 1019596
rect 474206 1019586 474230 1019596
rect 474206 1019562 474240 1019586
rect 474251 1019562 474323 1019596
rect 474206 1019552 474323 1019562
rect 473978 1019528 474323 1019552
rect 473991 1019484 474191 1019528
rect 474206 1019518 474230 1019528
rect 474206 1019494 474240 1019518
rect 474251 1019494 474323 1019528
rect 474206 1019484 474323 1019494
rect 473978 1019460 474323 1019484
rect 473991 1019416 474191 1019460
rect 474206 1019450 474230 1019460
rect 474206 1019426 474240 1019450
rect 474251 1019426 474323 1019460
rect 474206 1019416 474323 1019426
rect 473978 1019392 474323 1019416
rect 473991 1019322 474191 1019392
rect 474206 1019368 474230 1019392
rect 474251 1019322 474323 1019392
rect 474553 1019322 474609 1020322
rect 474625 1019322 474681 1020322
rect 474983 1020300 475183 1020322
rect 475198 1020310 475232 1020334
rect 475986 1020322 476020 1020334
rect 475243 1020310 475315 1020322
rect 475198 1020300 475315 1020310
rect 474970 1020276 475315 1020300
rect 474983 1020232 475183 1020276
rect 475198 1020266 475222 1020276
rect 475198 1020242 475232 1020266
rect 475243 1020242 475315 1020276
rect 475198 1020232 475315 1020242
rect 474970 1020208 475315 1020232
rect 474983 1020164 475183 1020208
rect 475198 1020198 475222 1020208
rect 475198 1020174 475232 1020198
rect 475243 1020174 475315 1020208
rect 475198 1020164 475315 1020174
rect 474970 1020140 475315 1020164
rect 474983 1020096 475183 1020140
rect 475198 1020130 475222 1020140
rect 475198 1020106 475232 1020130
rect 475243 1020106 475315 1020140
rect 475198 1020096 475315 1020106
rect 474970 1020072 475315 1020096
rect 474983 1020028 475183 1020072
rect 475198 1020062 475222 1020072
rect 475198 1020038 475232 1020062
rect 475243 1020038 475315 1020072
rect 475198 1020028 475315 1020038
rect 474970 1020004 475315 1020028
rect 474983 1019960 475183 1020004
rect 475198 1019994 475222 1020004
rect 475198 1019970 475232 1019994
rect 475243 1019970 475315 1020004
rect 475198 1019960 475315 1019970
rect 474970 1019936 475315 1019960
rect 474983 1019892 475183 1019936
rect 475198 1019926 475222 1019936
rect 475198 1019902 475232 1019926
rect 475243 1019902 475315 1019936
rect 475198 1019892 475315 1019902
rect 474970 1019868 475315 1019892
rect 474983 1019824 475183 1019868
rect 475198 1019858 475222 1019868
rect 475198 1019834 475232 1019858
rect 475243 1019834 475315 1019868
rect 475198 1019824 475315 1019834
rect 474970 1019800 475315 1019824
rect 474983 1019756 475183 1019800
rect 475198 1019790 475222 1019800
rect 475198 1019766 475232 1019790
rect 475243 1019766 475315 1019800
rect 475198 1019756 475315 1019766
rect 474970 1019732 475315 1019756
rect 474983 1019688 475183 1019732
rect 475198 1019722 475222 1019732
rect 475198 1019698 475232 1019722
rect 475243 1019698 475315 1019732
rect 475198 1019688 475315 1019698
rect 474970 1019664 475315 1019688
rect 474983 1019620 475183 1019664
rect 475198 1019654 475222 1019664
rect 475198 1019630 475232 1019654
rect 475243 1019630 475315 1019664
rect 475198 1019620 475315 1019630
rect 474970 1019596 475315 1019620
rect 474983 1019552 475183 1019596
rect 475198 1019586 475222 1019596
rect 475198 1019562 475232 1019586
rect 475243 1019562 475315 1019596
rect 475198 1019552 475315 1019562
rect 474970 1019528 475315 1019552
rect 474983 1019484 475183 1019528
rect 475198 1019518 475222 1019528
rect 475198 1019494 475232 1019518
rect 475243 1019494 475315 1019528
rect 475198 1019484 475315 1019494
rect 474970 1019460 475315 1019484
rect 474983 1019416 475183 1019460
rect 475198 1019450 475222 1019460
rect 475198 1019426 475232 1019450
rect 475243 1019426 475315 1019460
rect 475198 1019416 475315 1019426
rect 474970 1019392 475315 1019416
rect 474983 1019322 475183 1019392
rect 475198 1019368 475222 1019392
rect 475243 1019322 475315 1019392
rect 475545 1019322 475601 1020322
rect 475617 1019322 475673 1020322
rect 475975 1020300 476175 1020322
rect 476190 1020310 476224 1020334
rect 476978 1020322 477012 1020334
rect 476235 1020310 476307 1020322
rect 476190 1020300 476307 1020310
rect 475962 1020276 476307 1020300
rect 475975 1020232 476175 1020276
rect 476190 1020266 476214 1020276
rect 476190 1020242 476224 1020266
rect 476235 1020242 476307 1020276
rect 476190 1020232 476307 1020242
rect 475962 1020208 476307 1020232
rect 475975 1020164 476175 1020208
rect 476190 1020198 476214 1020208
rect 476190 1020174 476224 1020198
rect 476235 1020174 476307 1020208
rect 476190 1020164 476307 1020174
rect 475962 1020140 476307 1020164
rect 475975 1020096 476175 1020140
rect 476190 1020130 476214 1020140
rect 476190 1020106 476224 1020130
rect 476235 1020106 476307 1020140
rect 476190 1020096 476307 1020106
rect 475962 1020072 476307 1020096
rect 475975 1020028 476175 1020072
rect 476190 1020062 476214 1020072
rect 476190 1020038 476224 1020062
rect 476235 1020038 476307 1020072
rect 476190 1020028 476307 1020038
rect 475962 1020004 476307 1020028
rect 475975 1019960 476175 1020004
rect 476190 1019994 476214 1020004
rect 476190 1019970 476224 1019994
rect 476235 1019970 476307 1020004
rect 476190 1019960 476307 1019970
rect 475962 1019936 476307 1019960
rect 475975 1019892 476175 1019936
rect 476190 1019926 476214 1019936
rect 476190 1019902 476224 1019926
rect 476235 1019902 476307 1019936
rect 476190 1019892 476307 1019902
rect 475962 1019868 476307 1019892
rect 475975 1019824 476175 1019868
rect 476190 1019858 476214 1019868
rect 476190 1019834 476224 1019858
rect 476235 1019834 476307 1019868
rect 476190 1019824 476307 1019834
rect 475962 1019800 476307 1019824
rect 475975 1019756 476175 1019800
rect 476190 1019790 476214 1019800
rect 476190 1019766 476224 1019790
rect 476235 1019766 476307 1019800
rect 476190 1019756 476307 1019766
rect 475962 1019732 476307 1019756
rect 475975 1019688 476175 1019732
rect 476190 1019722 476214 1019732
rect 476190 1019698 476224 1019722
rect 476235 1019698 476307 1019732
rect 476190 1019688 476307 1019698
rect 475962 1019664 476307 1019688
rect 475975 1019620 476175 1019664
rect 476190 1019654 476214 1019664
rect 476190 1019630 476224 1019654
rect 476235 1019630 476307 1019664
rect 476190 1019620 476307 1019630
rect 475962 1019596 476307 1019620
rect 475975 1019552 476175 1019596
rect 476190 1019586 476214 1019596
rect 476190 1019562 476224 1019586
rect 476235 1019562 476307 1019596
rect 476190 1019552 476307 1019562
rect 475962 1019528 476307 1019552
rect 475975 1019484 476175 1019528
rect 476190 1019518 476214 1019528
rect 476190 1019494 476224 1019518
rect 476235 1019494 476307 1019528
rect 476190 1019484 476307 1019494
rect 475962 1019460 476307 1019484
rect 475975 1019416 476175 1019460
rect 476190 1019450 476214 1019460
rect 476190 1019426 476224 1019450
rect 476235 1019426 476307 1019460
rect 476190 1019416 476307 1019426
rect 475962 1019392 476307 1019416
rect 475975 1019322 476175 1019392
rect 476190 1019368 476214 1019392
rect 476235 1019322 476307 1019392
rect 476537 1019322 476593 1020322
rect 476609 1019322 476665 1020322
rect 476967 1020300 477167 1020322
rect 477182 1020310 477216 1020334
rect 477970 1020322 478004 1020334
rect 477227 1020310 477299 1020322
rect 477182 1020300 477299 1020310
rect 476954 1020276 477299 1020300
rect 476967 1020232 477167 1020276
rect 477182 1020266 477206 1020276
rect 477182 1020242 477216 1020266
rect 477227 1020242 477299 1020276
rect 477182 1020232 477299 1020242
rect 476954 1020208 477299 1020232
rect 476967 1020164 477167 1020208
rect 477182 1020198 477206 1020208
rect 477182 1020174 477216 1020198
rect 477227 1020174 477299 1020208
rect 477182 1020164 477299 1020174
rect 476954 1020140 477299 1020164
rect 476967 1020096 477167 1020140
rect 477182 1020130 477206 1020140
rect 477182 1020106 477216 1020130
rect 477227 1020106 477299 1020140
rect 477182 1020096 477299 1020106
rect 476954 1020072 477299 1020096
rect 476967 1020028 477167 1020072
rect 477182 1020062 477206 1020072
rect 477182 1020038 477216 1020062
rect 477227 1020038 477299 1020072
rect 477182 1020028 477299 1020038
rect 476954 1020004 477299 1020028
rect 476967 1019960 477167 1020004
rect 477182 1019994 477206 1020004
rect 477182 1019970 477216 1019994
rect 477227 1019970 477299 1020004
rect 477182 1019960 477299 1019970
rect 476954 1019936 477299 1019960
rect 476967 1019892 477167 1019936
rect 477182 1019926 477206 1019936
rect 477182 1019902 477216 1019926
rect 477227 1019902 477299 1019936
rect 477182 1019892 477299 1019902
rect 476954 1019868 477299 1019892
rect 476967 1019824 477167 1019868
rect 477182 1019858 477206 1019868
rect 477182 1019834 477216 1019858
rect 477227 1019834 477299 1019868
rect 477182 1019824 477299 1019834
rect 476954 1019800 477299 1019824
rect 476967 1019756 477167 1019800
rect 477182 1019790 477206 1019800
rect 477182 1019766 477216 1019790
rect 477227 1019766 477299 1019800
rect 477182 1019756 477299 1019766
rect 476954 1019732 477299 1019756
rect 476967 1019688 477167 1019732
rect 477182 1019722 477206 1019732
rect 477182 1019698 477216 1019722
rect 477227 1019698 477299 1019732
rect 477182 1019688 477299 1019698
rect 476954 1019664 477299 1019688
rect 476967 1019620 477167 1019664
rect 477182 1019654 477206 1019664
rect 477182 1019630 477216 1019654
rect 477227 1019630 477299 1019664
rect 477182 1019620 477299 1019630
rect 476954 1019596 477299 1019620
rect 476967 1019552 477167 1019596
rect 477182 1019586 477206 1019596
rect 477182 1019562 477216 1019586
rect 477227 1019562 477299 1019596
rect 477182 1019552 477299 1019562
rect 476954 1019528 477299 1019552
rect 476967 1019484 477167 1019528
rect 477182 1019518 477206 1019528
rect 477182 1019494 477216 1019518
rect 477227 1019494 477299 1019528
rect 477182 1019484 477299 1019494
rect 476954 1019460 477299 1019484
rect 476967 1019416 477167 1019460
rect 477182 1019450 477206 1019460
rect 477182 1019426 477216 1019450
rect 477227 1019426 477299 1019460
rect 477182 1019416 477299 1019426
rect 476954 1019392 477299 1019416
rect 476967 1019322 477167 1019392
rect 477182 1019368 477206 1019392
rect 477227 1019322 477299 1019392
rect 477529 1019322 477585 1020322
rect 477601 1019322 477657 1020322
rect 477959 1020300 478159 1020322
rect 478174 1020310 478208 1020334
rect 478962 1020322 478996 1020334
rect 478219 1020310 478291 1020322
rect 478174 1020300 478291 1020310
rect 477946 1020276 478291 1020300
rect 477959 1020232 478159 1020276
rect 478174 1020266 478198 1020276
rect 478174 1020242 478208 1020266
rect 478219 1020242 478291 1020276
rect 478174 1020232 478291 1020242
rect 477946 1020208 478291 1020232
rect 477959 1020164 478159 1020208
rect 478174 1020198 478198 1020208
rect 478174 1020174 478208 1020198
rect 478219 1020174 478291 1020208
rect 478174 1020164 478291 1020174
rect 477946 1020140 478291 1020164
rect 477959 1020096 478159 1020140
rect 478174 1020130 478198 1020140
rect 478174 1020106 478208 1020130
rect 478219 1020106 478291 1020140
rect 478174 1020096 478291 1020106
rect 477946 1020072 478291 1020096
rect 477959 1020028 478159 1020072
rect 478174 1020062 478198 1020072
rect 478174 1020038 478208 1020062
rect 478219 1020038 478291 1020072
rect 478174 1020028 478291 1020038
rect 477946 1020004 478291 1020028
rect 477959 1019960 478159 1020004
rect 478174 1019994 478198 1020004
rect 478174 1019970 478208 1019994
rect 478219 1019970 478291 1020004
rect 478174 1019960 478291 1019970
rect 477946 1019936 478291 1019960
rect 477959 1019892 478159 1019936
rect 478174 1019926 478198 1019936
rect 478174 1019902 478208 1019926
rect 478219 1019902 478291 1019936
rect 478174 1019892 478291 1019902
rect 477946 1019868 478291 1019892
rect 477959 1019824 478159 1019868
rect 478174 1019858 478198 1019868
rect 478174 1019834 478208 1019858
rect 478219 1019834 478291 1019868
rect 478174 1019824 478291 1019834
rect 477946 1019800 478291 1019824
rect 477959 1019756 478159 1019800
rect 478174 1019790 478198 1019800
rect 478174 1019766 478208 1019790
rect 478219 1019766 478291 1019800
rect 478174 1019756 478291 1019766
rect 477946 1019732 478291 1019756
rect 477959 1019688 478159 1019732
rect 478174 1019722 478198 1019732
rect 478174 1019698 478208 1019722
rect 478219 1019698 478291 1019732
rect 478174 1019688 478291 1019698
rect 477946 1019664 478291 1019688
rect 477959 1019620 478159 1019664
rect 478174 1019654 478198 1019664
rect 478174 1019630 478208 1019654
rect 478219 1019630 478291 1019664
rect 478174 1019620 478291 1019630
rect 477946 1019596 478291 1019620
rect 477959 1019552 478159 1019596
rect 478174 1019586 478198 1019596
rect 478174 1019562 478208 1019586
rect 478219 1019562 478291 1019596
rect 478174 1019552 478291 1019562
rect 477946 1019528 478291 1019552
rect 477959 1019484 478159 1019528
rect 478174 1019518 478198 1019528
rect 478174 1019494 478208 1019518
rect 478219 1019494 478291 1019528
rect 478174 1019484 478291 1019494
rect 477946 1019460 478291 1019484
rect 477959 1019416 478159 1019460
rect 478174 1019450 478198 1019460
rect 478174 1019426 478208 1019450
rect 478219 1019426 478291 1019460
rect 478174 1019416 478291 1019426
rect 477946 1019392 478291 1019416
rect 477959 1019322 478159 1019392
rect 478174 1019368 478198 1019392
rect 478219 1019322 478291 1019392
rect 478521 1019322 478577 1020322
rect 478593 1019322 478649 1020322
rect 478951 1020300 479151 1020322
rect 479166 1020310 479200 1020334
rect 479211 1020310 479283 1020322
rect 479166 1020300 479283 1020310
rect 478938 1020276 479283 1020300
rect 478951 1020232 479151 1020276
rect 479166 1020266 479190 1020276
rect 479166 1020242 479200 1020266
rect 479211 1020242 479283 1020276
rect 479166 1020232 479283 1020242
rect 478938 1020208 479283 1020232
rect 478951 1020164 479151 1020208
rect 479166 1020198 479190 1020208
rect 479166 1020174 479200 1020198
rect 479211 1020174 479283 1020208
rect 479166 1020164 479283 1020174
rect 478938 1020140 479283 1020164
rect 478951 1020096 479151 1020140
rect 479166 1020130 479190 1020140
rect 479166 1020106 479200 1020130
rect 479211 1020106 479283 1020140
rect 479166 1020096 479283 1020106
rect 478938 1020072 479283 1020096
rect 478951 1020028 479151 1020072
rect 479166 1020062 479190 1020072
rect 479166 1020038 479200 1020062
rect 479211 1020038 479283 1020072
rect 479166 1020028 479283 1020038
rect 478938 1020004 479283 1020028
rect 478951 1019960 479151 1020004
rect 479166 1019994 479190 1020004
rect 479166 1019970 479200 1019994
rect 479211 1019970 479283 1020004
rect 479166 1019960 479283 1019970
rect 478938 1019936 479283 1019960
rect 478951 1019892 479151 1019936
rect 479166 1019926 479190 1019936
rect 479166 1019902 479200 1019926
rect 479211 1019902 479283 1019936
rect 479166 1019892 479283 1019902
rect 478938 1019868 479283 1019892
rect 478951 1019824 479151 1019868
rect 479166 1019858 479190 1019868
rect 479166 1019834 479200 1019858
rect 479211 1019834 479283 1019868
rect 479166 1019824 479283 1019834
rect 478938 1019800 479283 1019824
rect 478951 1019756 479151 1019800
rect 479166 1019790 479190 1019800
rect 479166 1019766 479200 1019790
rect 479211 1019766 479283 1019800
rect 479166 1019756 479283 1019766
rect 478938 1019732 479283 1019756
rect 478951 1019688 479151 1019732
rect 479166 1019722 479190 1019732
rect 479166 1019698 479200 1019722
rect 479211 1019698 479283 1019732
rect 479166 1019688 479283 1019698
rect 478938 1019664 479283 1019688
rect 478951 1019620 479151 1019664
rect 479166 1019654 479190 1019664
rect 479166 1019630 479200 1019654
rect 479211 1019630 479283 1019664
rect 479166 1019620 479283 1019630
rect 478938 1019596 479283 1019620
rect 478951 1019552 479151 1019596
rect 479166 1019586 479190 1019596
rect 479166 1019562 479200 1019586
rect 479211 1019562 479283 1019596
rect 479166 1019552 479283 1019562
rect 478938 1019528 479283 1019552
rect 478951 1019484 479151 1019528
rect 479166 1019518 479190 1019528
rect 479166 1019494 479200 1019518
rect 479211 1019494 479283 1019528
rect 479166 1019484 479283 1019494
rect 478938 1019460 479283 1019484
rect 478951 1019416 479151 1019460
rect 479166 1019450 479190 1019460
rect 479166 1019426 479200 1019450
rect 479211 1019426 479283 1019460
rect 479166 1019416 479283 1019426
rect 478938 1019392 479283 1019416
rect 478951 1019322 479151 1019392
rect 479166 1019368 479190 1019392
rect 479211 1019322 479283 1019392
rect 479472 1019322 479544 1020322
rect 479610 1019322 479627 1020322
rect 479797 1019322 479830 1020322
rect 517561 1018210 517668 1022756
rect 518356 1020922 518406 1021922
rect 518617 1020922 518673 1021922
rect 518689 1020922 518745 1021922
rect 519107 1020922 519247 1021922
rect 530521 1020922 530577 1021922
rect 530593 1020922 530649 1021922
rect 531011 1020922 531151 1021922
rect 531473 1020922 531544 1021922
rect 531610 1020922 531627 1021922
rect 531797 1020922 531830 1021922
rect 531953 1021730 532025 1021760
rect 531953 1021692 531987 1021722
rect 518356 1019322 518406 1020322
rect 518617 1019322 518673 1020322
rect 518689 1019322 518745 1020322
rect 519107 1019322 519247 1020322
rect 530521 1019322 530577 1020322
rect 530593 1019322 530649 1020322
rect 531011 1019322 531151 1020322
rect 531473 1019322 531544 1020322
rect 531610 1019322 531627 1020322
rect 531797 1019322 531830 1020322
rect 569561 1018210 569668 1022756
rect 570356 1020922 570406 1021922
rect 570617 1020922 570673 1021922
rect 570689 1020922 570745 1021922
rect 571047 1021842 571247 1021922
rect 571262 1021852 571296 1021876
rect 571307 1021852 571379 1021922
rect 571262 1021842 571379 1021852
rect 571034 1021818 571379 1021842
rect 571047 1021774 571247 1021818
rect 571262 1021808 571286 1021818
rect 571262 1021784 571296 1021808
rect 571307 1021784 571379 1021818
rect 571262 1021774 571379 1021784
rect 571034 1021750 571379 1021774
rect 571047 1021706 571247 1021750
rect 571262 1021740 571286 1021750
rect 571262 1021716 571296 1021740
rect 571307 1021716 571379 1021750
rect 571262 1021706 571379 1021716
rect 571034 1021682 571379 1021706
rect 571047 1021638 571247 1021682
rect 571262 1021672 571286 1021682
rect 571262 1021648 571296 1021672
rect 571307 1021648 571379 1021682
rect 571262 1021638 571379 1021648
rect 571034 1021614 571379 1021638
rect 571047 1021570 571247 1021614
rect 571262 1021604 571286 1021614
rect 571262 1021580 571296 1021604
rect 571307 1021580 571379 1021614
rect 571262 1021570 571379 1021580
rect 571034 1021546 571379 1021570
rect 571047 1021502 571247 1021546
rect 571262 1021536 571286 1021546
rect 571262 1021512 571296 1021536
rect 571307 1021512 571379 1021546
rect 571262 1021502 571379 1021512
rect 571034 1021478 571379 1021502
rect 571047 1021434 571247 1021478
rect 571262 1021468 571286 1021478
rect 571262 1021444 571296 1021468
rect 571307 1021444 571379 1021478
rect 571262 1021434 571379 1021444
rect 571034 1021410 571379 1021434
rect 571047 1021366 571247 1021410
rect 571262 1021400 571286 1021410
rect 571262 1021376 571296 1021400
rect 571307 1021376 571379 1021410
rect 571262 1021366 571379 1021376
rect 571034 1021342 571379 1021366
rect 571047 1021298 571247 1021342
rect 571262 1021332 571286 1021342
rect 571262 1021308 571296 1021332
rect 571307 1021308 571379 1021342
rect 571262 1021298 571379 1021308
rect 571034 1021274 571379 1021298
rect 571047 1021230 571247 1021274
rect 571262 1021264 571286 1021274
rect 571262 1021240 571296 1021264
rect 571307 1021240 571379 1021274
rect 571262 1021230 571379 1021240
rect 571034 1021206 571379 1021230
rect 571047 1021162 571247 1021206
rect 571262 1021196 571286 1021206
rect 571262 1021172 571296 1021196
rect 571307 1021172 571379 1021206
rect 571262 1021162 571379 1021172
rect 571034 1021138 571379 1021162
rect 571047 1021094 571247 1021138
rect 571262 1021128 571286 1021138
rect 571262 1021104 571296 1021128
rect 571307 1021104 571379 1021138
rect 571262 1021094 571379 1021104
rect 571034 1021070 571379 1021094
rect 571047 1021026 571247 1021070
rect 571262 1021060 571286 1021070
rect 571262 1021036 571296 1021060
rect 571307 1021036 571379 1021070
rect 571262 1021026 571379 1021036
rect 571034 1021002 571379 1021026
rect 571047 1020958 571247 1021002
rect 571262 1020992 571286 1021002
rect 571262 1020968 571296 1020992
rect 571307 1020968 571379 1021002
rect 571262 1020958 571379 1020968
rect 571034 1020934 571379 1020958
rect 571047 1020922 571247 1020934
rect 571058 1020910 571082 1020922
rect 571262 1020910 571286 1020934
rect 571307 1020922 571379 1020934
rect 571609 1020922 571665 1021922
rect 571681 1020922 571737 1021922
rect 572039 1021842 572239 1021922
rect 572254 1021852 572288 1021876
rect 572299 1021852 572371 1021922
rect 572254 1021842 572371 1021852
rect 572026 1021818 572371 1021842
rect 572039 1021774 572239 1021818
rect 572254 1021808 572278 1021818
rect 572254 1021784 572288 1021808
rect 572299 1021784 572371 1021818
rect 572254 1021774 572371 1021784
rect 572026 1021750 572371 1021774
rect 572039 1021706 572239 1021750
rect 572254 1021740 572278 1021750
rect 572254 1021716 572288 1021740
rect 572299 1021716 572371 1021750
rect 572254 1021706 572371 1021716
rect 572026 1021682 572371 1021706
rect 572039 1021638 572239 1021682
rect 572254 1021672 572278 1021682
rect 572254 1021648 572288 1021672
rect 572299 1021648 572371 1021682
rect 572254 1021638 572371 1021648
rect 572026 1021614 572371 1021638
rect 572039 1021570 572239 1021614
rect 572254 1021604 572278 1021614
rect 572254 1021580 572288 1021604
rect 572299 1021580 572371 1021614
rect 572254 1021570 572371 1021580
rect 572026 1021546 572371 1021570
rect 572039 1021502 572239 1021546
rect 572254 1021536 572278 1021546
rect 572254 1021512 572288 1021536
rect 572299 1021512 572371 1021546
rect 572254 1021502 572371 1021512
rect 572026 1021478 572371 1021502
rect 572039 1021434 572239 1021478
rect 572254 1021468 572278 1021478
rect 572254 1021444 572288 1021468
rect 572299 1021444 572371 1021478
rect 572254 1021434 572371 1021444
rect 572026 1021410 572371 1021434
rect 572039 1021366 572239 1021410
rect 572254 1021400 572278 1021410
rect 572254 1021376 572288 1021400
rect 572299 1021376 572371 1021410
rect 572254 1021366 572371 1021376
rect 572026 1021342 572371 1021366
rect 572039 1021298 572239 1021342
rect 572254 1021332 572278 1021342
rect 572254 1021308 572288 1021332
rect 572299 1021308 572371 1021342
rect 572254 1021298 572371 1021308
rect 572026 1021274 572371 1021298
rect 572039 1021230 572239 1021274
rect 572254 1021264 572278 1021274
rect 572254 1021240 572288 1021264
rect 572299 1021240 572371 1021274
rect 572254 1021230 572371 1021240
rect 572026 1021206 572371 1021230
rect 572039 1021162 572239 1021206
rect 572254 1021196 572278 1021206
rect 572254 1021172 572288 1021196
rect 572299 1021172 572371 1021206
rect 572254 1021162 572371 1021172
rect 572026 1021138 572371 1021162
rect 572039 1021094 572239 1021138
rect 572254 1021128 572278 1021138
rect 572254 1021104 572288 1021128
rect 572299 1021104 572371 1021138
rect 572254 1021094 572371 1021104
rect 572026 1021070 572371 1021094
rect 572039 1021026 572239 1021070
rect 572254 1021060 572278 1021070
rect 572254 1021036 572288 1021060
rect 572299 1021036 572371 1021070
rect 572254 1021026 572371 1021036
rect 572026 1021002 572371 1021026
rect 572039 1020958 572239 1021002
rect 572254 1020992 572278 1021002
rect 572254 1020968 572288 1020992
rect 572299 1020968 572371 1021002
rect 572254 1020958 572371 1020968
rect 572026 1020934 572371 1020958
rect 572039 1020922 572239 1020934
rect 572050 1020910 572074 1020922
rect 572254 1020910 572278 1020934
rect 572299 1020922 572371 1020934
rect 572601 1020922 572657 1021922
rect 572673 1020922 572729 1021922
rect 573031 1021842 573231 1021922
rect 573246 1021852 573280 1021876
rect 573291 1021852 573363 1021922
rect 573246 1021842 573363 1021852
rect 573018 1021818 573363 1021842
rect 573031 1021774 573231 1021818
rect 573246 1021808 573270 1021818
rect 573246 1021784 573280 1021808
rect 573291 1021784 573363 1021818
rect 573246 1021774 573363 1021784
rect 573018 1021750 573363 1021774
rect 573031 1021706 573231 1021750
rect 573246 1021740 573270 1021750
rect 573246 1021716 573280 1021740
rect 573291 1021716 573363 1021750
rect 573246 1021706 573363 1021716
rect 573018 1021682 573363 1021706
rect 573031 1021638 573231 1021682
rect 573246 1021672 573270 1021682
rect 573246 1021648 573280 1021672
rect 573291 1021648 573363 1021682
rect 573246 1021638 573363 1021648
rect 573018 1021614 573363 1021638
rect 573031 1021570 573231 1021614
rect 573246 1021604 573270 1021614
rect 573246 1021580 573280 1021604
rect 573291 1021580 573363 1021614
rect 573246 1021570 573363 1021580
rect 573018 1021546 573363 1021570
rect 573031 1021502 573231 1021546
rect 573246 1021536 573270 1021546
rect 573246 1021512 573280 1021536
rect 573291 1021512 573363 1021546
rect 573246 1021502 573363 1021512
rect 573018 1021478 573363 1021502
rect 573031 1021434 573231 1021478
rect 573246 1021468 573270 1021478
rect 573246 1021444 573280 1021468
rect 573291 1021444 573363 1021478
rect 573246 1021434 573363 1021444
rect 573018 1021410 573363 1021434
rect 573031 1021366 573231 1021410
rect 573246 1021400 573270 1021410
rect 573246 1021376 573280 1021400
rect 573291 1021376 573363 1021410
rect 573246 1021366 573363 1021376
rect 573018 1021342 573363 1021366
rect 573031 1021298 573231 1021342
rect 573246 1021332 573270 1021342
rect 573246 1021308 573280 1021332
rect 573291 1021308 573363 1021342
rect 573246 1021298 573363 1021308
rect 573018 1021274 573363 1021298
rect 573031 1021230 573231 1021274
rect 573246 1021264 573270 1021274
rect 573246 1021240 573280 1021264
rect 573291 1021240 573363 1021274
rect 573246 1021230 573363 1021240
rect 573018 1021206 573363 1021230
rect 573031 1021162 573231 1021206
rect 573246 1021196 573270 1021206
rect 573246 1021172 573280 1021196
rect 573291 1021172 573363 1021206
rect 573246 1021162 573363 1021172
rect 573018 1021138 573363 1021162
rect 573031 1021094 573231 1021138
rect 573246 1021128 573270 1021138
rect 573246 1021104 573280 1021128
rect 573291 1021104 573363 1021138
rect 573246 1021094 573363 1021104
rect 573018 1021070 573363 1021094
rect 573031 1021026 573231 1021070
rect 573246 1021060 573270 1021070
rect 573246 1021036 573280 1021060
rect 573291 1021036 573363 1021070
rect 573246 1021026 573363 1021036
rect 573018 1021002 573363 1021026
rect 573031 1020958 573231 1021002
rect 573246 1020992 573270 1021002
rect 573246 1020968 573280 1020992
rect 573291 1020968 573363 1021002
rect 573246 1020958 573363 1020968
rect 573018 1020934 573363 1020958
rect 573031 1020922 573231 1020934
rect 573042 1020910 573066 1020922
rect 573246 1020910 573270 1020934
rect 573291 1020922 573363 1020934
rect 573593 1020922 573649 1021922
rect 573665 1020922 573721 1021922
rect 574023 1021842 574223 1021922
rect 574238 1021852 574272 1021876
rect 574283 1021852 574355 1021922
rect 574238 1021842 574355 1021852
rect 574010 1021818 574355 1021842
rect 574023 1021774 574223 1021818
rect 574238 1021808 574262 1021818
rect 574238 1021784 574272 1021808
rect 574283 1021784 574355 1021818
rect 574238 1021774 574355 1021784
rect 574010 1021750 574355 1021774
rect 574023 1021706 574223 1021750
rect 574238 1021740 574262 1021750
rect 574238 1021716 574272 1021740
rect 574283 1021716 574355 1021750
rect 574238 1021706 574355 1021716
rect 574010 1021682 574355 1021706
rect 574023 1021638 574223 1021682
rect 574238 1021672 574262 1021682
rect 574238 1021648 574272 1021672
rect 574283 1021648 574355 1021682
rect 574238 1021638 574355 1021648
rect 574010 1021614 574355 1021638
rect 574023 1021570 574223 1021614
rect 574238 1021604 574262 1021614
rect 574238 1021580 574272 1021604
rect 574283 1021580 574355 1021614
rect 574238 1021570 574355 1021580
rect 574010 1021546 574355 1021570
rect 574023 1021502 574223 1021546
rect 574238 1021536 574262 1021546
rect 574238 1021512 574272 1021536
rect 574283 1021512 574355 1021546
rect 574238 1021502 574355 1021512
rect 574010 1021478 574355 1021502
rect 574023 1021434 574223 1021478
rect 574238 1021468 574262 1021478
rect 574238 1021444 574272 1021468
rect 574283 1021444 574355 1021478
rect 574238 1021434 574355 1021444
rect 574010 1021410 574355 1021434
rect 574023 1021366 574223 1021410
rect 574238 1021400 574262 1021410
rect 574238 1021376 574272 1021400
rect 574283 1021376 574355 1021410
rect 574238 1021366 574355 1021376
rect 574010 1021342 574355 1021366
rect 574023 1021298 574223 1021342
rect 574238 1021332 574262 1021342
rect 574238 1021308 574272 1021332
rect 574283 1021308 574355 1021342
rect 574238 1021298 574355 1021308
rect 574010 1021274 574355 1021298
rect 574023 1021230 574223 1021274
rect 574238 1021264 574262 1021274
rect 574238 1021240 574272 1021264
rect 574283 1021240 574355 1021274
rect 574238 1021230 574355 1021240
rect 574010 1021206 574355 1021230
rect 574023 1021162 574223 1021206
rect 574238 1021196 574262 1021206
rect 574238 1021172 574272 1021196
rect 574283 1021172 574355 1021206
rect 574238 1021162 574355 1021172
rect 574010 1021138 574355 1021162
rect 574023 1021094 574223 1021138
rect 574238 1021128 574262 1021138
rect 574238 1021104 574272 1021128
rect 574283 1021104 574355 1021138
rect 574238 1021094 574355 1021104
rect 574010 1021070 574355 1021094
rect 574023 1021026 574223 1021070
rect 574238 1021060 574262 1021070
rect 574238 1021036 574272 1021060
rect 574283 1021036 574355 1021070
rect 574238 1021026 574355 1021036
rect 574010 1021002 574355 1021026
rect 574023 1020958 574223 1021002
rect 574238 1020992 574262 1021002
rect 574238 1020968 574272 1020992
rect 574283 1020968 574355 1021002
rect 574238 1020958 574355 1020968
rect 574010 1020934 574355 1020958
rect 574023 1020922 574223 1020934
rect 574034 1020910 574058 1020922
rect 574238 1020910 574262 1020934
rect 574283 1020922 574355 1020934
rect 574585 1020922 574641 1021922
rect 574657 1020922 574713 1021922
rect 575015 1021842 575215 1021922
rect 575230 1021852 575264 1021876
rect 575275 1021852 575347 1021922
rect 575230 1021842 575347 1021852
rect 575002 1021818 575347 1021842
rect 575015 1021774 575215 1021818
rect 575230 1021808 575254 1021818
rect 575230 1021784 575264 1021808
rect 575275 1021784 575347 1021818
rect 575230 1021774 575347 1021784
rect 575002 1021750 575347 1021774
rect 575015 1021706 575215 1021750
rect 575230 1021740 575254 1021750
rect 575230 1021716 575264 1021740
rect 575275 1021716 575347 1021750
rect 575230 1021706 575347 1021716
rect 575002 1021682 575347 1021706
rect 575015 1021638 575215 1021682
rect 575230 1021672 575254 1021682
rect 575230 1021648 575264 1021672
rect 575275 1021648 575347 1021682
rect 575230 1021638 575347 1021648
rect 575002 1021614 575347 1021638
rect 575015 1021570 575215 1021614
rect 575230 1021604 575254 1021614
rect 575230 1021580 575264 1021604
rect 575275 1021580 575347 1021614
rect 575230 1021570 575347 1021580
rect 575002 1021546 575347 1021570
rect 575015 1021502 575215 1021546
rect 575230 1021536 575254 1021546
rect 575230 1021512 575264 1021536
rect 575275 1021512 575347 1021546
rect 575230 1021502 575347 1021512
rect 575002 1021478 575347 1021502
rect 575015 1021434 575215 1021478
rect 575230 1021468 575254 1021478
rect 575230 1021444 575264 1021468
rect 575275 1021444 575347 1021478
rect 575230 1021434 575347 1021444
rect 575002 1021410 575347 1021434
rect 575015 1021366 575215 1021410
rect 575230 1021400 575254 1021410
rect 575230 1021376 575264 1021400
rect 575275 1021376 575347 1021410
rect 575230 1021366 575347 1021376
rect 575002 1021342 575347 1021366
rect 575015 1021298 575215 1021342
rect 575230 1021332 575254 1021342
rect 575230 1021308 575264 1021332
rect 575275 1021308 575347 1021342
rect 575230 1021298 575347 1021308
rect 575002 1021274 575347 1021298
rect 575015 1021230 575215 1021274
rect 575230 1021264 575254 1021274
rect 575230 1021240 575264 1021264
rect 575275 1021240 575347 1021274
rect 575230 1021230 575347 1021240
rect 575002 1021206 575347 1021230
rect 575015 1021162 575215 1021206
rect 575230 1021196 575254 1021206
rect 575230 1021172 575264 1021196
rect 575275 1021172 575347 1021206
rect 575230 1021162 575347 1021172
rect 575002 1021138 575347 1021162
rect 575015 1021094 575215 1021138
rect 575230 1021128 575254 1021138
rect 575230 1021104 575264 1021128
rect 575275 1021104 575347 1021138
rect 575230 1021094 575347 1021104
rect 575002 1021070 575347 1021094
rect 575015 1021026 575215 1021070
rect 575230 1021060 575254 1021070
rect 575230 1021036 575264 1021060
rect 575275 1021036 575347 1021070
rect 575230 1021026 575347 1021036
rect 575002 1021002 575347 1021026
rect 575015 1020958 575215 1021002
rect 575230 1020992 575254 1021002
rect 575230 1020968 575264 1020992
rect 575275 1020968 575347 1021002
rect 575230 1020958 575347 1020968
rect 575002 1020934 575347 1020958
rect 575015 1020922 575215 1020934
rect 575026 1020910 575050 1020922
rect 575230 1020910 575254 1020934
rect 575275 1020922 575347 1020934
rect 575577 1020922 575633 1021922
rect 575649 1020922 575705 1021922
rect 576007 1021842 576207 1021922
rect 576222 1021852 576256 1021876
rect 576267 1021852 576339 1021922
rect 576222 1021842 576339 1021852
rect 575994 1021818 576339 1021842
rect 576007 1021774 576207 1021818
rect 576222 1021808 576246 1021818
rect 576222 1021784 576256 1021808
rect 576267 1021784 576339 1021818
rect 576222 1021774 576339 1021784
rect 575994 1021750 576339 1021774
rect 576007 1021706 576207 1021750
rect 576222 1021740 576246 1021750
rect 576222 1021716 576256 1021740
rect 576267 1021716 576339 1021750
rect 576222 1021706 576339 1021716
rect 575994 1021682 576339 1021706
rect 576007 1021638 576207 1021682
rect 576222 1021672 576246 1021682
rect 576222 1021648 576256 1021672
rect 576267 1021648 576339 1021682
rect 576222 1021638 576339 1021648
rect 575994 1021614 576339 1021638
rect 576007 1021570 576207 1021614
rect 576222 1021604 576246 1021614
rect 576222 1021580 576256 1021604
rect 576267 1021580 576339 1021614
rect 576222 1021570 576339 1021580
rect 575994 1021546 576339 1021570
rect 576007 1021502 576207 1021546
rect 576222 1021536 576246 1021546
rect 576222 1021512 576256 1021536
rect 576267 1021512 576339 1021546
rect 576222 1021502 576339 1021512
rect 575994 1021478 576339 1021502
rect 576007 1021434 576207 1021478
rect 576222 1021468 576246 1021478
rect 576222 1021444 576256 1021468
rect 576267 1021444 576339 1021478
rect 576222 1021434 576339 1021444
rect 575994 1021410 576339 1021434
rect 576007 1021366 576207 1021410
rect 576222 1021400 576246 1021410
rect 576222 1021376 576256 1021400
rect 576267 1021376 576339 1021410
rect 576222 1021366 576339 1021376
rect 575994 1021342 576339 1021366
rect 576007 1021298 576207 1021342
rect 576222 1021332 576246 1021342
rect 576222 1021308 576256 1021332
rect 576267 1021308 576339 1021342
rect 576222 1021298 576339 1021308
rect 575994 1021274 576339 1021298
rect 576007 1021230 576207 1021274
rect 576222 1021264 576246 1021274
rect 576222 1021240 576256 1021264
rect 576267 1021240 576339 1021274
rect 576222 1021230 576339 1021240
rect 575994 1021206 576339 1021230
rect 576007 1021162 576207 1021206
rect 576222 1021196 576246 1021206
rect 576222 1021172 576256 1021196
rect 576267 1021172 576339 1021206
rect 576222 1021162 576339 1021172
rect 575994 1021138 576339 1021162
rect 576007 1021094 576207 1021138
rect 576222 1021128 576246 1021138
rect 576222 1021104 576256 1021128
rect 576267 1021104 576339 1021138
rect 576222 1021094 576339 1021104
rect 575994 1021070 576339 1021094
rect 576007 1021026 576207 1021070
rect 576222 1021060 576246 1021070
rect 576222 1021036 576256 1021060
rect 576267 1021036 576339 1021070
rect 576222 1021026 576339 1021036
rect 575994 1021002 576339 1021026
rect 576007 1020958 576207 1021002
rect 576222 1020992 576246 1021002
rect 576222 1020968 576256 1020992
rect 576267 1020968 576339 1021002
rect 576222 1020958 576339 1020968
rect 575994 1020934 576339 1020958
rect 576007 1020922 576207 1020934
rect 576018 1020910 576042 1020922
rect 576222 1020910 576246 1020934
rect 576267 1020922 576339 1020934
rect 576569 1020922 576625 1021922
rect 576641 1020922 576697 1021922
rect 576999 1021842 577199 1021922
rect 577214 1021852 577248 1021876
rect 577259 1021852 577331 1021922
rect 577214 1021842 577331 1021852
rect 576986 1021818 577331 1021842
rect 576999 1021774 577199 1021818
rect 577214 1021808 577238 1021818
rect 577214 1021784 577248 1021808
rect 577259 1021784 577331 1021818
rect 577214 1021774 577331 1021784
rect 576986 1021750 577331 1021774
rect 576999 1021706 577199 1021750
rect 577214 1021740 577238 1021750
rect 577214 1021716 577248 1021740
rect 577259 1021716 577331 1021750
rect 577214 1021706 577331 1021716
rect 576986 1021682 577331 1021706
rect 576999 1021638 577199 1021682
rect 577214 1021672 577238 1021682
rect 577214 1021648 577248 1021672
rect 577259 1021648 577331 1021682
rect 577214 1021638 577331 1021648
rect 576986 1021614 577331 1021638
rect 576999 1021570 577199 1021614
rect 577214 1021604 577238 1021614
rect 577214 1021580 577248 1021604
rect 577259 1021580 577331 1021614
rect 577214 1021570 577331 1021580
rect 576986 1021546 577331 1021570
rect 576999 1021502 577199 1021546
rect 577214 1021536 577238 1021546
rect 577214 1021512 577248 1021536
rect 577259 1021512 577331 1021546
rect 577214 1021502 577331 1021512
rect 576986 1021478 577331 1021502
rect 576999 1021434 577199 1021478
rect 577214 1021468 577238 1021478
rect 577214 1021444 577248 1021468
rect 577259 1021444 577331 1021478
rect 577214 1021434 577331 1021444
rect 576986 1021410 577331 1021434
rect 576999 1021366 577199 1021410
rect 577214 1021400 577238 1021410
rect 577214 1021376 577248 1021400
rect 577259 1021376 577331 1021410
rect 577214 1021366 577331 1021376
rect 576986 1021342 577331 1021366
rect 576999 1021298 577199 1021342
rect 577214 1021332 577238 1021342
rect 577214 1021308 577248 1021332
rect 577259 1021308 577331 1021342
rect 577214 1021298 577331 1021308
rect 576986 1021274 577331 1021298
rect 576999 1021230 577199 1021274
rect 577214 1021264 577238 1021274
rect 577214 1021240 577248 1021264
rect 577259 1021240 577331 1021274
rect 577214 1021230 577331 1021240
rect 576986 1021206 577331 1021230
rect 576999 1021162 577199 1021206
rect 577214 1021196 577238 1021206
rect 577214 1021172 577248 1021196
rect 577259 1021172 577331 1021206
rect 577214 1021162 577331 1021172
rect 576986 1021138 577331 1021162
rect 576999 1021094 577199 1021138
rect 577214 1021128 577238 1021138
rect 577214 1021104 577248 1021128
rect 577259 1021104 577331 1021138
rect 577214 1021094 577331 1021104
rect 576986 1021070 577331 1021094
rect 576999 1021026 577199 1021070
rect 577214 1021060 577238 1021070
rect 577214 1021036 577248 1021060
rect 577259 1021036 577331 1021070
rect 577214 1021026 577331 1021036
rect 576986 1021002 577331 1021026
rect 576999 1020958 577199 1021002
rect 577214 1020992 577238 1021002
rect 577214 1020968 577248 1020992
rect 577259 1020968 577331 1021002
rect 577214 1020958 577331 1020968
rect 576986 1020934 577331 1020958
rect 576999 1020922 577199 1020934
rect 577010 1020910 577034 1020922
rect 577214 1020910 577238 1020934
rect 577259 1020922 577331 1020934
rect 577561 1020922 577617 1021922
rect 577633 1020922 577689 1021922
rect 577991 1021842 578191 1021922
rect 578206 1021852 578240 1021876
rect 578251 1021852 578323 1021922
rect 578206 1021842 578323 1021852
rect 577978 1021818 578323 1021842
rect 577991 1021774 578191 1021818
rect 578206 1021808 578230 1021818
rect 578206 1021784 578240 1021808
rect 578251 1021784 578323 1021818
rect 578206 1021774 578323 1021784
rect 577978 1021750 578323 1021774
rect 577991 1021706 578191 1021750
rect 578206 1021740 578230 1021750
rect 578206 1021716 578240 1021740
rect 578251 1021716 578323 1021750
rect 578206 1021706 578323 1021716
rect 577978 1021682 578323 1021706
rect 577991 1021638 578191 1021682
rect 578206 1021672 578230 1021682
rect 578206 1021648 578240 1021672
rect 578251 1021648 578323 1021682
rect 578206 1021638 578323 1021648
rect 577978 1021614 578323 1021638
rect 577991 1021570 578191 1021614
rect 578206 1021604 578230 1021614
rect 578206 1021580 578240 1021604
rect 578251 1021580 578323 1021614
rect 578206 1021570 578323 1021580
rect 577978 1021546 578323 1021570
rect 577991 1021502 578191 1021546
rect 578206 1021536 578230 1021546
rect 578206 1021512 578240 1021536
rect 578251 1021512 578323 1021546
rect 578206 1021502 578323 1021512
rect 577978 1021478 578323 1021502
rect 577991 1021434 578191 1021478
rect 578206 1021468 578230 1021478
rect 578206 1021444 578240 1021468
rect 578251 1021444 578323 1021478
rect 578206 1021434 578323 1021444
rect 577978 1021410 578323 1021434
rect 577991 1021366 578191 1021410
rect 578206 1021400 578230 1021410
rect 578206 1021376 578240 1021400
rect 578251 1021376 578323 1021410
rect 578206 1021366 578323 1021376
rect 577978 1021342 578323 1021366
rect 577991 1021298 578191 1021342
rect 578206 1021332 578230 1021342
rect 578206 1021308 578240 1021332
rect 578251 1021308 578323 1021342
rect 578206 1021298 578323 1021308
rect 577978 1021274 578323 1021298
rect 577991 1021230 578191 1021274
rect 578206 1021264 578230 1021274
rect 578206 1021240 578240 1021264
rect 578251 1021240 578323 1021274
rect 578206 1021230 578323 1021240
rect 577978 1021206 578323 1021230
rect 577991 1021162 578191 1021206
rect 578206 1021196 578230 1021206
rect 578206 1021172 578240 1021196
rect 578251 1021172 578323 1021206
rect 578206 1021162 578323 1021172
rect 577978 1021138 578323 1021162
rect 577991 1021094 578191 1021138
rect 578206 1021128 578230 1021138
rect 578206 1021104 578240 1021128
rect 578251 1021104 578323 1021138
rect 578206 1021094 578323 1021104
rect 577978 1021070 578323 1021094
rect 577991 1021026 578191 1021070
rect 578206 1021060 578230 1021070
rect 578206 1021036 578240 1021060
rect 578251 1021036 578323 1021070
rect 578206 1021026 578323 1021036
rect 577978 1021002 578323 1021026
rect 577991 1020958 578191 1021002
rect 578206 1020992 578230 1021002
rect 578206 1020968 578240 1020992
rect 578251 1020968 578323 1021002
rect 578206 1020958 578323 1020968
rect 577978 1020934 578323 1020958
rect 577991 1020922 578191 1020934
rect 578002 1020910 578026 1020922
rect 578206 1020910 578230 1020934
rect 578251 1020922 578323 1020934
rect 578553 1020922 578609 1021922
rect 578625 1020922 578681 1021922
rect 578983 1021842 579183 1021922
rect 579198 1021852 579232 1021876
rect 579243 1021852 579315 1021922
rect 579198 1021842 579315 1021852
rect 578970 1021818 579315 1021842
rect 578983 1021774 579183 1021818
rect 579198 1021808 579222 1021818
rect 579198 1021784 579232 1021808
rect 579243 1021784 579315 1021818
rect 579198 1021774 579315 1021784
rect 578970 1021750 579315 1021774
rect 578983 1021706 579183 1021750
rect 579198 1021740 579222 1021750
rect 579198 1021716 579232 1021740
rect 579243 1021716 579315 1021750
rect 579198 1021706 579315 1021716
rect 578970 1021682 579315 1021706
rect 578983 1021638 579183 1021682
rect 579198 1021672 579222 1021682
rect 579198 1021648 579232 1021672
rect 579243 1021648 579315 1021682
rect 579198 1021638 579315 1021648
rect 578970 1021614 579315 1021638
rect 578983 1021570 579183 1021614
rect 579198 1021604 579222 1021614
rect 579198 1021580 579232 1021604
rect 579243 1021580 579315 1021614
rect 579198 1021570 579315 1021580
rect 578970 1021546 579315 1021570
rect 578983 1021502 579183 1021546
rect 579198 1021536 579222 1021546
rect 579198 1021512 579232 1021536
rect 579243 1021512 579315 1021546
rect 579198 1021502 579315 1021512
rect 578970 1021478 579315 1021502
rect 578983 1021434 579183 1021478
rect 579198 1021468 579222 1021478
rect 579198 1021444 579232 1021468
rect 579243 1021444 579315 1021478
rect 579198 1021434 579315 1021444
rect 578970 1021410 579315 1021434
rect 578983 1021366 579183 1021410
rect 579198 1021400 579222 1021410
rect 579198 1021376 579232 1021400
rect 579243 1021376 579315 1021410
rect 579198 1021366 579315 1021376
rect 578970 1021342 579315 1021366
rect 578983 1021298 579183 1021342
rect 579198 1021332 579222 1021342
rect 579198 1021308 579232 1021332
rect 579243 1021308 579315 1021342
rect 579198 1021298 579315 1021308
rect 578970 1021274 579315 1021298
rect 578983 1021230 579183 1021274
rect 579198 1021264 579222 1021274
rect 579198 1021240 579232 1021264
rect 579243 1021240 579315 1021274
rect 579198 1021230 579315 1021240
rect 578970 1021206 579315 1021230
rect 578983 1021162 579183 1021206
rect 579198 1021196 579222 1021206
rect 579198 1021172 579232 1021196
rect 579243 1021172 579315 1021206
rect 579198 1021162 579315 1021172
rect 578970 1021138 579315 1021162
rect 578983 1021094 579183 1021138
rect 579198 1021128 579222 1021138
rect 579198 1021104 579232 1021128
rect 579243 1021104 579315 1021138
rect 579198 1021094 579315 1021104
rect 578970 1021070 579315 1021094
rect 578983 1021026 579183 1021070
rect 579198 1021060 579222 1021070
rect 579198 1021036 579232 1021060
rect 579243 1021036 579315 1021070
rect 579198 1021026 579315 1021036
rect 578970 1021002 579315 1021026
rect 578983 1020958 579183 1021002
rect 579198 1020992 579222 1021002
rect 579198 1020968 579232 1020992
rect 579243 1020968 579315 1021002
rect 579198 1020958 579315 1020968
rect 578970 1020934 579315 1020958
rect 578983 1020922 579183 1020934
rect 578994 1020910 579018 1020922
rect 579198 1020910 579222 1020934
rect 579243 1020922 579315 1020934
rect 579545 1020922 579601 1021922
rect 579617 1020922 579673 1021922
rect 579975 1021842 580175 1021922
rect 580190 1021852 580224 1021876
rect 580235 1021852 580307 1021922
rect 580190 1021842 580307 1021852
rect 579962 1021818 580307 1021842
rect 579975 1021774 580175 1021818
rect 580190 1021808 580214 1021818
rect 580190 1021784 580224 1021808
rect 580235 1021784 580307 1021818
rect 580190 1021774 580307 1021784
rect 579962 1021750 580307 1021774
rect 579975 1021706 580175 1021750
rect 580190 1021740 580214 1021750
rect 580190 1021716 580224 1021740
rect 580235 1021716 580307 1021750
rect 580190 1021706 580307 1021716
rect 579962 1021682 580307 1021706
rect 579975 1021638 580175 1021682
rect 580190 1021672 580214 1021682
rect 580190 1021648 580224 1021672
rect 580235 1021648 580307 1021682
rect 580190 1021638 580307 1021648
rect 579962 1021614 580307 1021638
rect 579975 1021570 580175 1021614
rect 580190 1021604 580214 1021614
rect 580190 1021580 580224 1021604
rect 580235 1021580 580307 1021614
rect 580190 1021570 580307 1021580
rect 579962 1021546 580307 1021570
rect 579975 1021502 580175 1021546
rect 580190 1021536 580214 1021546
rect 580190 1021512 580224 1021536
rect 580235 1021512 580307 1021546
rect 580190 1021502 580307 1021512
rect 579962 1021478 580307 1021502
rect 579975 1021434 580175 1021478
rect 580190 1021468 580214 1021478
rect 580190 1021444 580224 1021468
rect 580235 1021444 580307 1021478
rect 580190 1021434 580307 1021444
rect 579962 1021410 580307 1021434
rect 579975 1021366 580175 1021410
rect 580190 1021400 580214 1021410
rect 580190 1021376 580224 1021400
rect 580235 1021376 580307 1021410
rect 580190 1021366 580307 1021376
rect 579962 1021342 580307 1021366
rect 579975 1021298 580175 1021342
rect 580190 1021332 580214 1021342
rect 580190 1021308 580224 1021332
rect 580235 1021308 580307 1021342
rect 580190 1021298 580307 1021308
rect 579962 1021274 580307 1021298
rect 579975 1021230 580175 1021274
rect 580190 1021264 580214 1021274
rect 580190 1021240 580224 1021264
rect 580235 1021240 580307 1021274
rect 580190 1021230 580307 1021240
rect 579962 1021206 580307 1021230
rect 579975 1021162 580175 1021206
rect 580190 1021196 580214 1021206
rect 580190 1021172 580224 1021196
rect 580235 1021172 580307 1021206
rect 580190 1021162 580307 1021172
rect 579962 1021138 580307 1021162
rect 579975 1021094 580175 1021138
rect 580190 1021128 580214 1021138
rect 580190 1021104 580224 1021128
rect 580235 1021104 580307 1021138
rect 580190 1021094 580307 1021104
rect 579962 1021070 580307 1021094
rect 579975 1021026 580175 1021070
rect 580190 1021060 580214 1021070
rect 580190 1021036 580224 1021060
rect 580235 1021036 580307 1021070
rect 580190 1021026 580307 1021036
rect 579962 1021002 580307 1021026
rect 579975 1020958 580175 1021002
rect 580190 1020992 580214 1021002
rect 580190 1020968 580224 1020992
rect 580235 1020968 580307 1021002
rect 580190 1020958 580307 1020968
rect 579962 1020934 580307 1020958
rect 579975 1020922 580175 1020934
rect 579986 1020910 580010 1020922
rect 580190 1020910 580214 1020934
rect 580235 1020922 580307 1020934
rect 580537 1020922 580593 1021922
rect 580609 1020922 580665 1021922
rect 580967 1021842 581167 1021922
rect 581182 1021852 581216 1021876
rect 581227 1021852 581299 1021922
rect 581182 1021842 581299 1021852
rect 580954 1021818 581299 1021842
rect 580967 1021774 581167 1021818
rect 581182 1021808 581206 1021818
rect 581182 1021784 581216 1021808
rect 581227 1021784 581299 1021818
rect 581182 1021774 581299 1021784
rect 580954 1021750 581299 1021774
rect 580967 1021706 581167 1021750
rect 581182 1021740 581206 1021750
rect 581182 1021716 581216 1021740
rect 581227 1021716 581299 1021750
rect 581182 1021706 581299 1021716
rect 580954 1021682 581299 1021706
rect 580967 1021638 581167 1021682
rect 581182 1021672 581206 1021682
rect 581182 1021648 581216 1021672
rect 581227 1021648 581299 1021682
rect 581182 1021638 581299 1021648
rect 580954 1021614 581299 1021638
rect 580967 1021570 581167 1021614
rect 581182 1021604 581206 1021614
rect 581182 1021580 581216 1021604
rect 581227 1021580 581299 1021614
rect 581182 1021570 581299 1021580
rect 580954 1021546 581299 1021570
rect 580967 1021502 581167 1021546
rect 581182 1021536 581206 1021546
rect 581182 1021512 581216 1021536
rect 581227 1021512 581299 1021546
rect 581182 1021502 581299 1021512
rect 580954 1021478 581299 1021502
rect 580967 1021434 581167 1021478
rect 581182 1021468 581206 1021478
rect 581182 1021444 581216 1021468
rect 581227 1021444 581299 1021478
rect 581182 1021434 581299 1021444
rect 580954 1021410 581299 1021434
rect 580967 1021366 581167 1021410
rect 581182 1021400 581206 1021410
rect 581182 1021376 581216 1021400
rect 581227 1021376 581299 1021410
rect 581182 1021366 581299 1021376
rect 580954 1021342 581299 1021366
rect 580967 1021298 581167 1021342
rect 581182 1021332 581206 1021342
rect 581182 1021308 581216 1021332
rect 581227 1021308 581299 1021342
rect 581182 1021298 581299 1021308
rect 580954 1021274 581299 1021298
rect 580967 1021230 581167 1021274
rect 581182 1021264 581206 1021274
rect 581182 1021240 581216 1021264
rect 581227 1021240 581299 1021274
rect 581182 1021230 581299 1021240
rect 580954 1021206 581299 1021230
rect 580967 1021162 581167 1021206
rect 581182 1021196 581206 1021206
rect 581182 1021172 581216 1021196
rect 581227 1021172 581299 1021206
rect 581182 1021162 581299 1021172
rect 580954 1021138 581299 1021162
rect 580967 1021094 581167 1021138
rect 581182 1021128 581206 1021138
rect 581182 1021104 581216 1021128
rect 581227 1021104 581299 1021138
rect 581182 1021094 581299 1021104
rect 580954 1021070 581299 1021094
rect 580967 1021026 581167 1021070
rect 581182 1021060 581206 1021070
rect 581182 1021036 581216 1021060
rect 581227 1021036 581299 1021070
rect 581182 1021026 581299 1021036
rect 580954 1021002 581299 1021026
rect 580967 1020958 581167 1021002
rect 581182 1020992 581206 1021002
rect 581182 1020968 581216 1020992
rect 581227 1020968 581299 1021002
rect 581182 1020958 581299 1020968
rect 580954 1020934 581299 1020958
rect 580967 1020922 581167 1020934
rect 580978 1020910 581002 1020922
rect 581182 1020910 581206 1020934
rect 581227 1020922 581299 1020934
rect 581529 1020922 581585 1021922
rect 581601 1020922 581657 1021922
rect 581959 1021842 582159 1021922
rect 582174 1021852 582208 1021876
rect 582219 1021852 582291 1021922
rect 582174 1021842 582291 1021852
rect 581946 1021818 582291 1021842
rect 581959 1021774 582159 1021818
rect 582174 1021808 582198 1021818
rect 582174 1021784 582208 1021808
rect 582219 1021784 582291 1021818
rect 582174 1021774 582291 1021784
rect 581946 1021750 582291 1021774
rect 581959 1021706 582159 1021750
rect 582174 1021740 582198 1021750
rect 582174 1021716 582208 1021740
rect 582219 1021716 582291 1021750
rect 582174 1021706 582291 1021716
rect 581946 1021682 582291 1021706
rect 581959 1021638 582159 1021682
rect 582174 1021672 582198 1021682
rect 582174 1021648 582208 1021672
rect 582219 1021648 582291 1021682
rect 582174 1021638 582291 1021648
rect 581946 1021614 582291 1021638
rect 581959 1021570 582159 1021614
rect 582174 1021604 582198 1021614
rect 582174 1021580 582208 1021604
rect 582219 1021580 582291 1021614
rect 582174 1021570 582291 1021580
rect 581946 1021546 582291 1021570
rect 581959 1021502 582159 1021546
rect 582174 1021536 582198 1021546
rect 582174 1021512 582208 1021536
rect 582219 1021512 582291 1021546
rect 582174 1021502 582291 1021512
rect 581946 1021478 582291 1021502
rect 581959 1021434 582159 1021478
rect 582174 1021468 582198 1021478
rect 582174 1021444 582208 1021468
rect 582219 1021444 582291 1021478
rect 582174 1021434 582291 1021444
rect 581946 1021410 582291 1021434
rect 581959 1021366 582159 1021410
rect 582174 1021400 582198 1021410
rect 582174 1021376 582208 1021400
rect 582219 1021376 582291 1021410
rect 582174 1021366 582291 1021376
rect 581946 1021342 582291 1021366
rect 581959 1021298 582159 1021342
rect 582174 1021332 582198 1021342
rect 582174 1021308 582208 1021332
rect 582219 1021308 582291 1021342
rect 582174 1021298 582291 1021308
rect 581946 1021274 582291 1021298
rect 581959 1021230 582159 1021274
rect 582174 1021264 582198 1021274
rect 582174 1021240 582208 1021264
rect 582219 1021240 582291 1021274
rect 582174 1021230 582291 1021240
rect 581946 1021206 582291 1021230
rect 581959 1021162 582159 1021206
rect 582174 1021196 582198 1021206
rect 582174 1021172 582208 1021196
rect 582219 1021172 582291 1021206
rect 582174 1021162 582291 1021172
rect 581946 1021138 582291 1021162
rect 581959 1021094 582159 1021138
rect 582174 1021128 582198 1021138
rect 582174 1021104 582208 1021128
rect 582219 1021104 582291 1021138
rect 582174 1021094 582291 1021104
rect 581946 1021070 582291 1021094
rect 581959 1021026 582159 1021070
rect 582174 1021060 582198 1021070
rect 582174 1021036 582208 1021060
rect 582219 1021036 582291 1021070
rect 582174 1021026 582291 1021036
rect 581946 1021002 582291 1021026
rect 581959 1020958 582159 1021002
rect 582174 1020992 582198 1021002
rect 582174 1020968 582208 1020992
rect 582219 1020968 582291 1021002
rect 582174 1020958 582291 1020968
rect 581946 1020934 582291 1020958
rect 581959 1020922 582159 1020934
rect 581970 1020910 581994 1020922
rect 582174 1020910 582198 1020934
rect 582219 1020922 582291 1020934
rect 582521 1020922 582577 1021922
rect 582593 1020922 582649 1021922
rect 582951 1021842 583151 1021922
rect 583166 1021852 583200 1021876
rect 583211 1021852 583283 1021922
rect 583166 1021842 583283 1021852
rect 582938 1021818 583283 1021842
rect 582951 1021774 583151 1021818
rect 583166 1021808 583190 1021818
rect 583166 1021784 583200 1021808
rect 583211 1021784 583283 1021818
rect 583166 1021774 583283 1021784
rect 582938 1021750 583283 1021774
rect 582951 1021706 583151 1021750
rect 583166 1021740 583190 1021750
rect 583166 1021716 583200 1021740
rect 583211 1021716 583283 1021750
rect 583166 1021706 583283 1021716
rect 582938 1021682 583283 1021706
rect 582951 1021638 583151 1021682
rect 583166 1021672 583190 1021682
rect 583166 1021648 583200 1021672
rect 583211 1021648 583283 1021682
rect 583166 1021638 583283 1021648
rect 582938 1021614 583283 1021638
rect 582951 1021570 583151 1021614
rect 583166 1021604 583190 1021614
rect 583166 1021580 583200 1021604
rect 583211 1021580 583283 1021614
rect 583166 1021570 583283 1021580
rect 582938 1021546 583283 1021570
rect 582951 1021502 583151 1021546
rect 583166 1021536 583190 1021546
rect 583166 1021512 583200 1021536
rect 583211 1021512 583283 1021546
rect 583166 1021502 583283 1021512
rect 582938 1021478 583283 1021502
rect 582951 1021434 583151 1021478
rect 583166 1021468 583190 1021478
rect 583166 1021444 583200 1021468
rect 583211 1021444 583283 1021478
rect 583166 1021434 583283 1021444
rect 582938 1021410 583283 1021434
rect 582951 1021366 583151 1021410
rect 583166 1021400 583190 1021410
rect 583166 1021376 583200 1021400
rect 583211 1021376 583283 1021410
rect 583166 1021366 583283 1021376
rect 582938 1021342 583283 1021366
rect 582951 1021298 583151 1021342
rect 583166 1021332 583190 1021342
rect 583166 1021308 583200 1021332
rect 583211 1021308 583283 1021342
rect 583166 1021298 583283 1021308
rect 582938 1021274 583283 1021298
rect 582951 1021230 583151 1021274
rect 583166 1021264 583190 1021274
rect 583166 1021240 583200 1021264
rect 583211 1021240 583283 1021274
rect 583166 1021230 583283 1021240
rect 582938 1021206 583283 1021230
rect 582951 1021162 583151 1021206
rect 583166 1021196 583190 1021206
rect 583166 1021172 583200 1021196
rect 583211 1021172 583283 1021206
rect 583166 1021162 583283 1021172
rect 582938 1021138 583283 1021162
rect 582951 1021094 583151 1021138
rect 583166 1021128 583190 1021138
rect 583166 1021104 583200 1021128
rect 583211 1021104 583283 1021138
rect 583166 1021094 583283 1021104
rect 582938 1021070 583283 1021094
rect 582951 1021026 583151 1021070
rect 583166 1021060 583190 1021070
rect 583166 1021036 583200 1021060
rect 583211 1021036 583283 1021070
rect 583166 1021026 583283 1021036
rect 582938 1021002 583283 1021026
rect 582951 1020958 583151 1021002
rect 583166 1020992 583190 1021002
rect 583166 1020968 583200 1020992
rect 583211 1020968 583283 1021002
rect 583166 1020958 583283 1020968
rect 582938 1020934 583283 1020958
rect 582951 1020922 583151 1020934
rect 582962 1020910 582986 1020922
rect 583166 1020910 583190 1020934
rect 583211 1020922 583283 1020934
rect 583472 1020922 583544 1021922
rect 583610 1020922 583627 1021922
rect 583797 1020922 583830 1021922
rect 583953 1021730 584025 1021760
rect 583953 1021692 583987 1021722
rect 571058 1020322 571092 1020334
rect 570356 1019322 570406 1020322
rect 570617 1019322 570673 1020322
rect 570689 1019322 570745 1020322
rect 571047 1020300 571247 1020322
rect 571262 1020310 571296 1020334
rect 572050 1020322 572084 1020334
rect 571307 1020310 571379 1020322
rect 571262 1020300 571379 1020310
rect 571034 1020276 571379 1020300
rect 571047 1020232 571247 1020276
rect 571262 1020266 571286 1020276
rect 571262 1020242 571296 1020266
rect 571307 1020242 571379 1020276
rect 571262 1020232 571379 1020242
rect 571034 1020208 571379 1020232
rect 571047 1020164 571247 1020208
rect 571262 1020198 571286 1020208
rect 571262 1020174 571296 1020198
rect 571307 1020174 571379 1020208
rect 571262 1020164 571379 1020174
rect 571034 1020140 571379 1020164
rect 571047 1020096 571247 1020140
rect 571262 1020130 571286 1020140
rect 571262 1020106 571296 1020130
rect 571307 1020106 571379 1020140
rect 571262 1020096 571379 1020106
rect 571034 1020072 571379 1020096
rect 571047 1020028 571247 1020072
rect 571262 1020062 571286 1020072
rect 571262 1020038 571296 1020062
rect 571307 1020038 571379 1020072
rect 571262 1020028 571379 1020038
rect 571034 1020004 571379 1020028
rect 571047 1019960 571247 1020004
rect 571262 1019994 571286 1020004
rect 571262 1019970 571296 1019994
rect 571307 1019970 571379 1020004
rect 571262 1019960 571379 1019970
rect 571034 1019936 571379 1019960
rect 571047 1019892 571247 1019936
rect 571262 1019926 571286 1019936
rect 571262 1019902 571296 1019926
rect 571307 1019902 571379 1019936
rect 571262 1019892 571379 1019902
rect 571034 1019868 571379 1019892
rect 571047 1019824 571247 1019868
rect 571262 1019858 571286 1019868
rect 571262 1019834 571296 1019858
rect 571307 1019834 571379 1019868
rect 571262 1019824 571379 1019834
rect 571034 1019800 571379 1019824
rect 571047 1019756 571247 1019800
rect 571262 1019790 571286 1019800
rect 571262 1019766 571296 1019790
rect 571307 1019766 571379 1019800
rect 571262 1019756 571379 1019766
rect 571034 1019732 571379 1019756
rect 571047 1019688 571247 1019732
rect 571262 1019722 571286 1019732
rect 571262 1019698 571296 1019722
rect 571307 1019698 571379 1019732
rect 571262 1019688 571379 1019698
rect 571034 1019664 571379 1019688
rect 571047 1019620 571247 1019664
rect 571262 1019654 571286 1019664
rect 571262 1019630 571296 1019654
rect 571307 1019630 571379 1019664
rect 571262 1019620 571379 1019630
rect 571034 1019596 571379 1019620
rect 571047 1019552 571247 1019596
rect 571262 1019586 571286 1019596
rect 571262 1019562 571296 1019586
rect 571307 1019562 571379 1019596
rect 571262 1019552 571379 1019562
rect 571034 1019528 571379 1019552
rect 571047 1019484 571247 1019528
rect 571262 1019518 571286 1019528
rect 571262 1019494 571296 1019518
rect 571307 1019494 571379 1019528
rect 571262 1019484 571379 1019494
rect 571034 1019460 571379 1019484
rect 571047 1019416 571247 1019460
rect 571262 1019450 571286 1019460
rect 571262 1019426 571296 1019450
rect 571307 1019426 571379 1019460
rect 571262 1019416 571379 1019426
rect 571034 1019392 571379 1019416
rect 571047 1019322 571247 1019392
rect 571262 1019368 571286 1019392
rect 571307 1019322 571379 1019392
rect 571609 1019322 571665 1020322
rect 571681 1019322 571737 1020322
rect 572039 1020300 572239 1020322
rect 572254 1020310 572288 1020334
rect 573042 1020322 573076 1020334
rect 572299 1020310 572371 1020322
rect 572254 1020300 572371 1020310
rect 572026 1020276 572371 1020300
rect 572039 1020232 572239 1020276
rect 572254 1020266 572278 1020276
rect 572254 1020242 572288 1020266
rect 572299 1020242 572371 1020276
rect 572254 1020232 572371 1020242
rect 572026 1020208 572371 1020232
rect 572039 1020164 572239 1020208
rect 572254 1020198 572278 1020208
rect 572254 1020174 572288 1020198
rect 572299 1020174 572371 1020208
rect 572254 1020164 572371 1020174
rect 572026 1020140 572371 1020164
rect 572039 1020096 572239 1020140
rect 572254 1020130 572278 1020140
rect 572254 1020106 572288 1020130
rect 572299 1020106 572371 1020140
rect 572254 1020096 572371 1020106
rect 572026 1020072 572371 1020096
rect 572039 1020028 572239 1020072
rect 572254 1020062 572278 1020072
rect 572254 1020038 572288 1020062
rect 572299 1020038 572371 1020072
rect 572254 1020028 572371 1020038
rect 572026 1020004 572371 1020028
rect 572039 1019960 572239 1020004
rect 572254 1019994 572278 1020004
rect 572254 1019970 572288 1019994
rect 572299 1019970 572371 1020004
rect 572254 1019960 572371 1019970
rect 572026 1019936 572371 1019960
rect 572039 1019892 572239 1019936
rect 572254 1019926 572278 1019936
rect 572254 1019902 572288 1019926
rect 572299 1019902 572371 1019936
rect 572254 1019892 572371 1019902
rect 572026 1019868 572371 1019892
rect 572039 1019824 572239 1019868
rect 572254 1019858 572278 1019868
rect 572254 1019834 572288 1019858
rect 572299 1019834 572371 1019868
rect 572254 1019824 572371 1019834
rect 572026 1019800 572371 1019824
rect 572039 1019756 572239 1019800
rect 572254 1019790 572278 1019800
rect 572254 1019766 572288 1019790
rect 572299 1019766 572371 1019800
rect 572254 1019756 572371 1019766
rect 572026 1019732 572371 1019756
rect 572039 1019688 572239 1019732
rect 572254 1019722 572278 1019732
rect 572254 1019698 572288 1019722
rect 572299 1019698 572371 1019732
rect 572254 1019688 572371 1019698
rect 572026 1019664 572371 1019688
rect 572039 1019620 572239 1019664
rect 572254 1019654 572278 1019664
rect 572254 1019630 572288 1019654
rect 572299 1019630 572371 1019664
rect 572254 1019620 572371 1019630
rect 572026 1019596 572371 1019620
rect 572039 1019552 572239 1019596
rect 572254 1019586 572278 1019596
rect 572254 1019562 572288 1019586
rect 572299 1019562 572371 1019596
rect 572254 1019552 572371 1019562
rect 572026 1019528 572371 1019552
rect 572039 1019484 572239 1019528
rect 572254 1019518 572278 1019528
rect 572254 1019494 572288 1019518
rect 572299 1019494 572371 1019528
rect 572254 1019484 572371 1019494
rect 572026 1019460 572371 1019484
rect 572039 1019416 572239 1019460
rect 572254 1019450 572278 1019460
rect 572254 1019426 572288 1019450
rect 572299 1019426 572371 1019460
rect 572254 1019416 572371 1019426
rect 572026 1019392 572371 1019416
rect 572039 1019322 572239 1019392
rect 572254 1019368 572278 1019392
rect 572299 1019322 572371 1019392
rect 572601 1019322 572657 1020322
rect 572673 1019322 572729 1020322
rect 573031 1020300 573231 1020322
rect 573246 1020310 573280 1020334
rect 574034 1020322 574068 1020334
rect 573291 1020310 573363 1020322
rect 573246 1020300 573363 1020310
rect 573018 1020276 573363 1020300
rect 573031 1020232 573231 1020276
rect 573246 1020266 573270 1020276
rect 573246 1020242 573280 1020266
rect 573291 1020242 573363 1020276
rect 573246 1020232 573363 1020242
rect 573018 1020208 573363 1020232
rect 573031 1020164 573231 1020208
rect 573246 1020198 573270 1020208
rect 573246 1020174 573280 1020198
rect 573291 1020174 573363 1020208
rect 573246 1020164 573363 1020174
rect 573018 1020140 573363 1020164
rect 573031 1020096 573231 1020140
rect 573246 1020130 573270 1020140
rect 573246 1020106 573280 1020130
rect 573291 1020106 573363 1020140
rect 573246 1020096 573363 1020106
rect 573018 1020072 573363 1020096
rect 573031 1020028 573231 1020072
rect 573246 1020062 573270 1020072
rect 573246 1020038 573280 1020062
rect 573291 1020038 573363 1020072
rect 573246 1020028 573363 1020038
rect 573018 1020004 573363 1020028
rect 573031 1019960 573231 1020004
rect 573246 1019994 573270 1020004
rect 573246 1019970 573280 1019994
rect 573291 1019970 573363 1020004
rect 573246 1019960 573363 1019970
rect 573018 1019936 573363 1019960
rect 573031 1019892 573231 1019936
rect 573246 1019926 573270 1019936
rect 573246 1019902 573280 1019926
rect 573291 1019902 573363 1019936
rect 573246 1019892 573363 1019902
rect 573018 1019868 573363 1019892
rect 573031 1019824 573231 1019868
rect 573246 1019858 573270 1019868
rect 573246 1019834 573280 1019858
rect 573291 1019834 573363 1019868
rect 573246 1019824 573363 1019834
rect 573018 1019800 573363 1019824
rect 573031 1019756 573231 1019800
rect 573246 1019790 573270 1019800
rect 573246 1019766 573280 1019790
rect 573291 1019766 573363 1019800
rect 573246 1019756 573363 1019766
rect 573018 1019732 573363 1019756
rect 573031 1019688 573231 1019732
rect 573246 1019722 573270 1019732
rect 573246 1019698 573280 1019722
rect 573291 1019698 573363 1019732
rect 573246 1019688 573363 1019698
rect 573018 1019664 573363 1019688
rect 573031 1019620 573231 1019664
rect 573246 1019654 573270 1019664
rect 573246 1019630 573280 1019654
rect 573291 1019630 573363 1019664
rect 573246 1019620 573363 1019630
rect 573018 1019596 573363 1019620
rect 573031 1019552 573231 1019596
rect 573246 1019586 573270 1019596
rect 573246 1019562 573280 1019586
rect 573291 1019562 573363 1019596
rect 573246 1019552 573363 1019562
rect 573018 1019528 573363 1019552
rect 573031 1019484 573231 1019528
rect 573246 1019518 573270 1019528
rect 573246 1019494 573280 1019518
rect 573291 1019494 573363 1019528
rect 573246 1019484 573363 1019494
rect 573018 1019460 573363 1019484
rect 573031 1019416 573231 1019460
rect 573246 1019450 573270 1019460
rect 573246 1019426 573280 1019450
rect 573291 1019426 573363 1019460
rect 573246 1019416 573363 1019426
rect 573018 1019392 573363 1019416
rect 573031 1019322 573231 1019392
rect 573246 1019368 573270 1019392
rect 573291 1019322 573363 1019392
rect 573593 1019322 573649 1020322
rect 573665 1019322 573721 1020322
rect 574023 1020300 574223 1020322
rect 574238 1020310 574272 1020334
rect 575026 1020322 575060 1020334
rect 574283 1020310 574355 1020322
rect 574238 1020300 574355 1020310
rect 574010 1020276 574355 1020300
rect 574023 1020232 574223 1020276
rect 574238 1020266 574262 1020276
rect 574238 1020242 574272 1020266
rect 574283 1020242 574355 1020276
rect 574238 1020232 574355 1020242
rect 574010 1020208 574355 1020232
rect 574023 1020164 574223 1020208
rect 574238 1020198 574262 1020208
rect 574238 1020174 574272 1020198
rect 574283 1020174 574355 1020208
rect 574238 1020164 574355 1020174
rect 574010 1020140 574355 1020164
rect 574023 1020096 574223 1020140
rect 574238 1020130 574262 1020140
rect 574238 1020106 574272 1020130
rect 574283 1020106 574355 1020140
rect 574238 1020096 574355 1020106
rect 574010 1020072 574355 1020096
rect 574023 1020028 574223 1020072
rect 574238 1020062 574262 1020072
rect 574238 1020038 574272 1020062
rect 574283 1020038 574355 1020072
rect 574238 1020028 574355 1020038
rect 574010 1020004 574355 1020028
rect 574023 1019960 574223 1020004
rect 574238 1019994 574262 1020004
rect 574238 1019970 574272 1019994
rect 574283 1019970 574355 1020004
rect 574238 1019960 574355 1019970
rect 574010 1019936 574355 1019960
rect 574023 1019892 574223 1019936
rect 574238 1019926 574262 1019936
rect 574238 1019902 574272 1019926
rect 574283 1019902 574355 1019936
rect 574238 1019892 574355 1019902
rect 574010 1019868 574355 1019892
rect 574023 1019824 574223 1019868
rect 574238 1019858 574262 1019868
rect 574238 1019834 574272 1019858
rect 574283 1019834 574355 1019868
rect 574238 1019824 574355 1019834
rect 574010 1019800 574355 1019824
rect 574023 1019756 574223 1019800
rect 574238 1019790 574262 1019800
rect 574238 1019766 574272 1019790
rect 574283 1019766 574355 1019800
rect 574238 1019756 574355 1019766
rect 574010 1019732 574355 1019756
rect 574023 1019688 574223 1019732
rect 574238 1019722 574262 1019732
rect 574238 1019698 574272 1019722
rect 574283 1019698 574355 1019732
rect 574238 1019688 574355 1019698
rect 574010 1019664 574355 1019688
rect 574023 1019620 574223 1019664
rect 574238 1019654 574262 1019664
rect 574238 1019630 574272 1019654
rect 574283 1019630 574355 1019664
rect 574238 1019620 574355 1019630
rect 574010 1019596 574355 1019620
rect 574023 1019552 574223 1019596
rect 574238 1019586 574262 1019596
rect 574238 1019562 574272 1019586
rect 574283 1019562 574355 1019596
rect 574238 1019552 574355 1019562
rect 574010 1019528 574355 1019552
rect 574023 1019484 574223 1019528
rect 574238 1019518 574262 1019528
rect 574238 1019494 574272 1019518
rect 574283 1019494 574355 1019528
rect 574238 1019484 574355 1019494
rect 574010 1019460 574355 1019484
rect 574023 1019416 574223 1019460
rect 574238 1019450 574262 1019460
rect 574238 1019426 574272 1019450
rect 574283 1019426 574355 1019460
rect 574238 1019416 574355 1019426
rect 574010 1019392 574355 1019416
rect 574023 1019322 574223 1019392
rect 574238 1019368 574262 1019392
rect 574283 1019322 574355 1019392
rect 574585 1019322 574641 1020322
rect 574657 1019322 574713 1020322
rect 575015 1020300 575215 1020322
rect 575230 1020310 575264 1020334
rect 576018 1020322 576052 1020334
rect 575275 1020310 575347 1020322
rect 575230 1020300 575347 1020310
rect 575002 1020276 575347 1020300
rect 575015 1020232 575215 1020276
rect 575230 1020266 575254 1020276
rect 575230 1020242 575264 1020266
rect 575275 1020242 575347 1020276
rect 575230 1020232 575347 1020242
rect 575002 1020208 575347 1020232
rect 575015 1020164 575215 1020208
rect 575230 1020198 575254 1020208
rect 575230 1020174 575264 1020198
rect 575275 1020174 575347 1020208
rect 575230 1020164 575347 1020174
rect 575002 1020140 575347 1020164
rect 575015 1020096 575215 1020140
rect 575230 1020130 575254 1020140
rect 575230 1020106 575264 1020130
rect 575275 1020106 575347 1020140
rect 575230 1020096 575347 1020106
rect 575002 1020072 575347 1020096
rect 575015 1020028 575215 1020072
rect 575230 1020062 575254 1020072
rect 575230 1020038 575264 1020062
rect 575275 1020038 575347 1020072
rect 575230 1020028 575347 1020038
rect 575002 1020004 575347 1020028
rect 575015 1019960 575215 1020004
rect 575230 1019994 575254 1020004
rect 575230 1019970 575264 1019994
rect 575275 1019970 575347 1020004
rect 575230 1019960 575347 1019970
rect 575002 1019936 575347 1019960
rect 575015 1019892 575215 1019936
rect 575230 1019926 575254 1019936
rect 575230 1019902 575264 1019926
rect 575275 1019902 575347 1019936
rect 575230 1019892 575347 1019902
rect 575002 1019868 575347 1019892
rect 575015 1019824 575215 1019868
rect 575230 1019858 575254 1019868
rect 575230 1019834 575264 1019858
rect 575275 1019834 575347 1019868
rect 575230 1019824 575347 1019834
rect 575002 1019800 575347 1019824
rect 575015 1019756 575215 1019800
rect 575230 1019790 575254 1019800
rect 575230 1019766 575264 1019790
rect 575275 1019766 575347 1019800
rect 575230 1019756 575347 1019766
rect 575002 1019732 575347 1019756
rect 575015 1019688 575215 1019732
rect 575230 1019722 575254 1019732
rect 575230 1019698 575264 1019722
rect 575275 1019698 575347 1019732
rect 575230 1019688 575347 1019698
rect 575002 1019664 575347 1019688
rect 575015 1019620 575215 1019664
rect 575230 1019654 575254 1019664
rect 575230 1019630 575264 1019654
rect 575275 1019630 575347 1019664
rect 575230 1019620 575347 1019630
rect 575002 1019596 575347 1019620
rect 575015 1019552 575215 1019596
rect 575230 1019586 575254 1019596
rect 575230 1019562 575264 1019586
rect 575275 1019562 575347 1019596
rect 575230 1019552 575347 1019562
rect 575002 1019528 575347 1019552
rect 575015 1019484 575215 1019528
rect 575230 1019518 575254 1019528
rect 575230 1019494 575264 1019518
rect 575275 1019494 575347 1019528
rect 575230 1019484 575347 1019494
rect 575002 1019460 575347 1019484
rect 575015 1019416 575215 1019460
rect 575230 1019450 575254 1019460
rect 575230 1019426 575264 1019450
rect 575275 1019426 575347 1019460
rect 575230 1019416 575347 1019426
rect 575002 1019392 575347 1019416
rect 575015 1019322 575215 1019392
rect 575230 1019368 575254 1019392
rect 575275 1019322 575347 1019392
rect 575577 1019322 575633 1020322
rect 575649 1019322 575705 1020322
rect 576007 1020300 576207 1020322
rect 576222 1020310 576256 1020334
rect 577010 1020322 577044 1020334
rect 576267 1020310 576339 1020322
rect 576222 1020300 576339 1020310
rect 575994 1020276 576339 1020300
rect 576007 1020232 576207 1020276
rect 576222 1020266 576246 1020276
rect 576222 1020242 576256 1020266
rect 576267 1020242 576339 1020276
rect 576222 1020232 576339 1020242
rect 575994 1020208 576339 1020232
rect 576007 1020164 576207 1020208
rect 576222 1020198 576246 1020208
rect 576222 1020174 576256 1020198
rect 576267 1020174 576339 1020208
rect 576222 1020164 576339 1020174
rect 575994 1020140 576339 1020164
rect 576007 1020096 576207 1020140
rect 576222 1020130 576246 1020140
rect 576222 1020106 576256 1020130
rect 576267 1020106 576339 1020140
rect 576222 1020096 576339 1020106
rect 575994 1020072 576339 1020096
rect 576007 1020028 576207 1020072
rect 576222 1020062 576246 1020072
rect 576222 1020038 576256 1020062
rect 576267 1020038 576339 1020072
rect 576222 1020028 576339 1020038
rect 575994 1020004 576339 1020028
rect 576007 1019960 576207 1020004
rect 576222 1019994 576246 1020004
rect 576222 1019970 576256 1019994
rect 576267 1019970 576339 1020004
rect 576222 1019960 576339 1019970
rect 575994 1019936 576339 1019960
rect 576007 1019892 576207 1019936
rect 576222 1019926 576246 1019936
rect 576222 1019902 576256 1019926
rect 576267 1019902 576339 1019936
rect 576222 1019892 576339 1019902
rect 575994 1019868 576339 1019892
rect 576007 1019824 576207 1019868
rect 576222 1019858 576246 1019868
rect 576222 1019834 576256 1019858
rect 576267 1019834 576339 1019868
rect 576222 1019824 576339 1019834
rect 575994 1019800 576339 1019824
rect 576007 1019756 576207 1019800
rect 576222 1019790 576246 1019800
rect 576222 1019766 576256 1019790
rect 576267 1019766 576339 1019800
rect 576222 1019756 576339 1019766
rect 575994 1019732 576339 1019756
rect 576007 1019688 576207 1019732
rect 576222 1019722 576246 1019732
rect 576222 1019698 576256 1019722
rect 576267 1019698 576339 1019732
rect 576222 1019688 576339 1019698
rect 575994 1019664 576339 1019688
rect 576007 1019620 576207 1019664
rect 576222 1019654 576246 1019664
rect 576222 1019630 576256 1019654
rect 576267 1019630 576339 1019664
rect 576222 1019620 576339 1019630
rect 575994 1019596 576339 1019620
rect 576007 1019552 576207 1019596
rect 576222 1019586 576246 1019596
rect 576222 1019562 576256 1019586
rect 576267 1019562 576339 1019596
rect 576222 1019552 576339 1019562
rect 575994 1019528 576339 1019552
rect 576007 1019484 576207 1019528
rect 576222 1019518 576246 1019528
rect 576222 1019494 576256 1019518
rect 576267 1019494 576339 1019528
rect 576222 1019484 576339 1019494
rect 575994 1019460 576339 1019484
rect 576007 1019416 576207 1019460
rect 576222 1019450 576246 1019460
rect 576222 1019426 576256 1019450
rect 576267 1019426 576339 1019460
rect 576222 1019416 576339 1019426
rect 575994 1019392 576339 1019416
rect 576007 1019322 576207 1019392
rect 576222 1019368 576246 1019392
rect 576267 1019322 576339 1019392
rect 576569 1019322 576625 1020322
rect 576641 1019322 576697 1020322
rect 576999 1020300 577199 1020322
rect 577214 1020310 577248 1020334
rect 578002 1020322 578036 1020334
rect 577259 1020310 577331 1020322
rect 577214 1020300 577331 1020310
rect 576986 1020276 577331 1020300
rect 576999 1020232 577199 1020276
rect 577214 1020266 577238 1020276
rect 577214 1020242 577248 1020266
rect 577259 1020242 577331 1020276
rect 577214 1020232 577331 1020242
rect 576986 1020208 577331 1020232
rect 576999 1020164 577199 1020208
rect 577214 1020198 577238 1020208
rect 577214 1020174 577248 1020198
rect 577259 1020174 577331 1020208
rect 577214 1020164 577331 1020174
rect 576986 1020140 577331 1020164
rect 576999 1020096 577199 1020140
rect 577214 1020130 577238 1020140
rect 577214 1020106 577248 1020130
rect 577259 1020106 577331 1020140
rect 577214 1020096 577331 1020106
rect 576986 1020072 577331 1020096
rect 576999 1020028 577199 1020072
rect 577214 1020062 577238 1020072
rect 577214 1020038 577248 1020062
rect 577259 1020038 577331 1020072
rect 577214 1020028 577331 1020038
rect 576986 1020004 577331 1020028
rect 576999 1019960 577199 1020004
rect 577214 1019994 577238 1020004
rect 577214 1019970 577248 1019994
rect 577259 1019970 577331 1020004
rect 577214 1019960 577331 1019970
rect 576986 1019936 577331 1019960
rect 576999 1019892 577199 1019936
rect 577214 1019926 577238 1019936
rect 577214 1019902 577248 1019926
rect 577259 1019902 577331 1019936
rect 577214 1019892 577331 1019902
rect 576986 1019868 577331 1019892
rect 576999 1019824 577199 1019868
rect 577214 1019858 577238 1019868
rect 577214 1019834 577248 1019858
rect 577259 1019834 577331 1019868
rect 577214 1019824 577331 1019834
rect 576986 1019800 577331 1019824
rect 576999 1019756 577199 1019800
rect 577214 1019790 577238 1019800
rect 577214 1019766 577248 1019790
rect 577259 1019766 577331 1019800
rect 577214 1019756 577331 1019766
rect 576986 1019732 577331 1019756
rect 576999 1019688 577199 1019732
rect 577214 1019722 577238 1019732
rect 577214 1019698 577248 1019722
rect 577259 1019698 577331 1019732
rect 577214 1019688 577331 1019698
rect 576986 1019664 577331 1019688
rect 576999 1019620 577199 1019664
rect 577214 1019654 577238 1019664
rect 577214 1019630 577248 1019654
rect 577259 1019630 577331 1019664
rect 577214 1019620 577331 1019630
rect 576986 1019596 577331 1019620
rect 576999 1019552 577199 1019596
rect 577214 1019586 577238 1019596
rect 577214 1019562 577248 1019586
rect 577259 1019562 577331 1019596
rect 577214 1019552 577331 1019562
rect 576986 1019528 577331 1019552
rect 576999 1019484 577199 1019528
rect 577214 1019518 577238 1019528
rect 577214 1019494 577248 1019518
rect 577259 1019494 577331 1019528
rect 577214 1019484 577331 1019494
rect 576986 1019460 577331 1019484
rect 576999 1019416 577199 1019460
rect 577214 1019450 577238 1019460
rect 577214 1019426 577248 1019450
rect 577259 1019426 577331 1019460
rect 577214 1019416 577331 1019426
rect 576986 1019392 577331 1019416
rect 576999 1019322 577199 1019392
rect 577214 1019368 577238 1019392
rect 577259 1019322 577331 1019392
rect 577561 1019322 577617 1020322
rect 577633 1019322 577689 1020322
rect 577991 1020300 578191 1020322
rect 578206 1020310 578240 1020334
rect 578994 1020322 579028 1020334
rect 578251 1020310 578323 1020322
rect 578206 1020300 578323 1020310
rect 577978 1020276 578323 1020300
rect 577991 1020232 578191 1020276
rect 578206 1020266 578230 1020276
rect 578206 1020242 578240 1020266
rect 578251 1020242 578323 1020276
rect 578206 1020232 578323 1020242
rect 577978 1020208 578323 1020232
rect 577991 1020164 578191 1020208
rect 578206 1020198 578230 1020208
rect 578206 1020174 578240 1020198
rect 578251 1020174 578323 1020208
rect 578206 1020164 578323 1020174
rect 577978 1020140 578323 1020164
rect 577991 1020096 578191 1020140
rect 578206 1020130 578230 1020140
rect 578206 1020106 578240 1020130
rect 578251 1020106 578323 1020140
rect 578206 1020096 578323 1020106
rect 577978 1020072 578323 1020096
rect 577991 1020028 578191 1020072
rect 578206 1020062 578230 1020072
rect 578206 1020038 578240 1020062
rect 578251 1020038 578323 1020072
rect 578206 1020028 578323 1020038
rect 577978 1020004 578323 1020028
rect 577991 1019960 578191 1020004
rect 578206 1019994 578230 1020004
rect 578206 1019970 578240 1019994
rect 578251 1019970 578323 1020004
rect 578206 1019960 578323 1019970
rect 577978 1019936 578323 1019960
rect 577991 1019892 578191 1019936
rect 578206 1019926 578230 1019936
rect 578206 1019902 578240 1019926
rect 578251 1019902 578323 1019936
rect 578206 1019892 578323 1019902
rect 577978 1019868 578323 1019892
rect 577991 1019824 578191 1019868
rect 578206 1019858 578230 1019868
rect 578206 1019834 578240 1019858
rect 578251 1019834 578323 1019868
rect 578206 1019824 578323 1019834
rect 577978 1019800 578323 1019824
rect 577991 1019756 578191 1019800
rect 578206 1019790 578230 1019800
rect 578206 1019766 578240 1019790
rect 578251 1019766 578323 1019800
rect 578206 1019756 578323 1019766
rect 577978 1019732 578323 1019756
rect 577991 1019688 578191 1019732
rect 578206 1019722 578230 1019732
rect 578206 1019698 578240 1019722
rect 578251 1019698 578323 1019732
rect 578206 1019688 578323 1019698
rect 577978 1019664 578323 1019688
rect 577991 1019620 578191 1019664
rect 578206 1019654 578230 1019664
rect 578206 1019630 578240 1019654
rect 578251 1019630 578323 1019664
rect 578206 1019620 578323 1019630
rect 577978 1019596 578323 1019620
rect 577991 1019552 578191 1019596
rect 578206 1019586 578230 1019596
rect 578206 1019562 578240 1019586
rect 578251 1019562 578323 1019596
rect 578206 1019552 578323 1019562
rect 577978 1019528 578323 1019552
rect 577991 1019484 578191 1019528
rect 578206 1019518 578230 1019528
rect 578206 1019494 578240 1019518
rect 578251 1019494 578323 1019528
rect 578206 1019484 578323 1019494
rect 577978 1019460 578323 1019484
rect 577991 1019416 578191 1019460
rect 578206 1019450 578230 1019460
rect 578206 1019426 578240 1019450
rect 578251 1019426 578323 1019460
rect 578206 1019416 578323 1019426
rect 577978 1019392 578323 1019416
rect 577991 1019322 578191 1019392
rect 578206 1019368 578230 1019392
rect 578251 1019322 578323 1019392
rect 578553 1019322 578609 1020322
rect 578625 1019322 578681 1020322
rect 578983 1020300 579183 1020322
rect 579198 1020310 579232 1020334
rect 579986 1020322 580020 1020334
rect 579243 1020310 579315 1020322
rect 579198 1020300 579315 1020310
rect 578970 1020276 579315 1020300
rect 578983 1020232 579183 1020276
rect 579198 1020266 579222 1020276
rect 579198 1020242 579232 1020266
rect 579243 1020242 579315 1020276
rect 579198 1020232 579315 1020242
rect 578970 1020208 579315 1020232
rect 578983 1020164 579183 1020208
rect 579198 1020198 579222 1020208
rect 579198 1020174 579232 1020198
rect 579243 1020174 579315 1020208
rect 579198 1020164 579315 1020174
rect 578970 1020140 579315 1020164
rect 578983 1020096 579183 1020140
rect 579198 1020130 579222 1020140
rect 579198 1020106 579232 1020130
rect 579243 1020106 579315 1020140
rect 579198 1020096 579315 1020106
rect 578970 1020072 579315 1020096
rect 578983 1020028 579183 1020072
rect 579198 1020062 579222 1020072
rect 579198 1020038 579232 1020062
rect 579243 1020038 579315 1020072
rect 579198 1020028 579315 1020038
rect 578970 1020004 579315 1020028
rect 578983 1019960 579183 1020004
rect 579198 1019994 579222 1020004
rect 579198 1019970 579232 1019994
rect 579243 1019970 579315 1020004
rect 579198 1019960 579315 1019970
rect 578970 1019936 579315 1019960
rect 578983 1019892 579183 1019936
rect 579198 1019926 579222 1019936
rect 579198 1019902 579232 1019926
rect 579243 1019902 579315 1019936
rect 579198 1019892 579315 1019902
rect 578970 1019868 579315 1019892
rect 578983 1019824 579183 1019868
rect 579198 1019858 579222 1019868
rect 579198 1019834 579232 1019858
rect 579243 1019834 579315 1019868
rect 579198 1019824 579315 1019834
rect 578970 1019800 579315 1019824
rect 578983 1019756 579183 1019800
rect 579198 1019790 579222 1019800
rect 579198 1019766 579232 1019790
rect 579243 1019766 579315 1019800
rect 579198 1019756 579315 1019766
rect 578970 1019732 579315 1019756
rect 578983 1019688 579183 1019732
rect 579198 1019722 579222 1019732
rect 579198 1019698 579232 1019722
rect 579243 1019698 579315 1019732
rect 579198 1019688 579315 1019698
rect 578970 1019664 579315 1019688
rect 578983 1019620 579183 1019664
rect 579198 1019654 579222 1019664
rect 579198 1019630 579232 1019654
rect 579243 1019630 579315 1019664
rect 579198 1019620 579315 1019630
rect 578970 1019596 579315 1019620
rect 578983 1019552 579183 1019596
rect 579198 1019586 579222 1019596
rect 579198 1019562 579232 1019586
rect 579243 1019562 579315 1019596
rect 579198 1019552 579315 1019562
rect 578970 1019528 579315 1019552
rect 578983 1019484 579183 1019528
rect 579198 1019518 579222 1019528
rect 579198 1019494 579232 1019518
rect 579243 1019494 579315 1019528
rect 579198 1019484 579315 1019494
rect 578970 1019460 579315 1019484
rect 578983 1019416 579183 1019460
rect 579198 1019450 579222 1019460
rect 579198 1019426 579232 1019450
rect 579243 1019426 579315 1019460
rect 579198 1019416 579315 1019426
rect 578970 1019392 579315 1019416
rect 578983 1019322 579183 1019392
rect 579198 1019368 579222 1019392
rect 579243 1019322 579315 1019392
rect 579545 1019322 579601 1020322
rect 579617 1019322 579673 1020322
rect 579975 1020300 580175 1020322
rect 580190 1020310 580224 1020334
rect 580978 1020322 581012 1020334
rect 580235 1020310 580307 1020322
rect 580190 1020300 580307 1020310
rect 579962 1020276 580307 1020300
rect 579975 1020232 580175 1020276
rect 580190 1020266 580214 1020276
rect 580190 1020242 580224 1020266
rect 580235 1020242 580307 1020276
rect 580190 1020232 580307 1020242
rect 579962 1020208 580307 1020232
rect 579975 1020164 580175 1020208
rect 580190 1020198 580214 1020208
rect 580190 1020174 580224 1020198
rect 580235 1020174 580307 1020208
rect 580190 1020164 580307 1020174
rect 579962 1020140 580307 1020164
rect 579975 1020096 580175 1020140
rect 580190 1020130 580214 1020140
rect 580190 1020106 580224 1020130
rect 580235 1020106 580307 1020140
rect 580190 1020096 580307 1020106
rect 579962 1020072 580307 1020096
rect 579975 1020028 580175 1020072
rect 580190 1020062 580214 1020072
rect 580190 1020038 580224 1020062
rect 580235 1020038 580307 1020072
rect 580190 1020028 580307 1020038
rect 579962 1020004 580307 1020028
rect 579975 1019960 580175 1020004
rect 580190 1019994 580214 1020004
rect 580190 1019970 580224 1019994
rect 580235 1019970 580307 1020004
rect 580190 1019960 580307 1019970
rect 579962 1019936 580307 1019960
rect 579975 1019892 580175 1019936
rect 580190 1019926 580214 1019936
rect 580190 1019902 580224 1019926
rect 580235 1019902 580307 1019936
rect 580190 1019892 580307 1019902
rect 579962 1019868 580307 1019892
rect 579975 1019824 580175 1019868
rect 580190 1019858 580214 1019868
rect 580190 1019834 580224 1019858
rect 580235 1019834 580307 1019868
rect 580190 1019824 580307 1019834
rect 579962 1019800 580307 1019824
rect 579975 1019756 580175 1019800
rect 580190 1019790 580214 1019800
rect 580190 1019766 580224 1019790
rect 580235 1019766 580307 1019800
rect 580190 1019756 580307 1019766
rect 579962 1019732 580307 1019756
rect 579975 1019688 580175 1019732
rect 580190 1019722 580214 1019732
rect 580190 1019698 580224 1019722
rect 580235 1019698 580307 1019732
rect 580190 1019688 580307 1019698
rect 579962 1019664 580307 1019688
rect 579975 1019620 580175 1019664
rect 580190 1019654 580214 1019664
rect 580190 1019630 580224 1019654
rect 580235 1019630 580307 1019664
rect 580190 1019620 580307 1019630
rect 579962 1019596 580307 1019620
rect 579975 1019552 580175 1019596
rect 580190 1019586 580214 1019596
rect 580190 1019562 580224 1019586
rect 580235 1019562 580307 1019596
rect 580190 1019552 580307 1019562
rect 579962 1019528 580307 1019552
rect 579975 1019484 580175 1019528
rect 580190 1019518 580214 1019528
rect 580190 1019494 580224 1019518
rect 580235 1019494 580307 1019528
rect 580190 1019484 580307 1019494
rect 579962 1019460 580307 1019484
rect 579975 1019416 580175 1019460
rect 580190 1019450 580214 1019460
rect 580190 1019426 580224 1019450
rect 580235 1019426 580307 1019460
rect 580190 1019416 580307 1019426
rect 579962 1019392 580307 1019416
rect 579975 1019322 580175 1019392
rect 580190 1019368 580214 1019392
rect 580235 1019322 580307 1019392
rect 580537 1019322 580593 1020322
rect 580609 1019322 580665 1020322
rect 580967 1020300 581167 1020322
rect 581182 1020310 581216 1020334
rect 581970 1020322 582004 1020334
rect 581227 1020310 581299 1020322
rect 581182 1020300 581299 1020310
rect 580954 1020276 581299 1020300
rect 580967 1020232 581167 1020276
rect 581182 1020266 581206 1020276
rect 581182 1020242 581216 1020266
rect 581227 1020242 581299 1020276
rect 581182 1020232 581299 1020242
rect 580954 1020208 581299 1020232
rect 580967 1020164 581167 1020208
rect 581182 1020198 581206 1020208
rect 581182 1020174 581216 1020198
rect 581227 1020174 581299 1020208
rect 581182 1020164 581299 1020174
rect 580954 1020140 581299 1020164
rect 580967 1020096 581167 1020140
rect 581182 1020130 581206 1020140
rect 581182 1020106 581216 1020130
rect 581227 1020106 581299 1020140
rect 581182 1020096 581299 1020106
rect 580954 1020072 581299 1020096
rect 580967 1020028 581167 1020072
rect 581182 1020062 581206 1020072
rect 581182 1020038 581216 1020062
rect 581227 1020038 581299 1020072
rect 581182 1020028 581299 1020038
rect 580954 1020004 581299 1020028
rect 580967 1019960 581167 1020004
rect 581182 1019994 581206 1020004
rect 581182 1019970 581216 1019994
rect 581227 1019970 581299 1020004
rect 581182 1019960 581299 1019970
rect 580954 1019936 581299 1019960
rect 580967 1019892 581167 1019936
rect 581182 1019926 581206 1019936
rect 581182 1019902 581216 1019926
rect 581227 1019902 581299 1019936
rect 581182 1019892 581299 1019902
rect 580954 1019868 581299 1019892
rect 580967 1019824 581167 1019868
rect 581182 1019858 581206 1019868
rect 581182 1019834 581216 1019858
rect 581227 1019834 581299 1019868
rect 581182 1019824 581299 1019834
rect 580954 1019800 581299 1019824
rect 580967 1019756 581167 1019800
rect 581182 1019790 581206 1019800
rect 581182 1019766 581216 1019790
rect 581227 1019766 581299 1019800
rect 581182 1019756 581299 1019766
rect 580954 1019732 581299 1019756
rect 580967 1019688 581167 1019732
rect 581182 1019722 581206 1019732
rect 581182 1019698 581216 1019722
rect 581227 1019698 581299 1019732
rect 581182 1019688 581299 1019698
rect 580954 1019664 581299 1019688
rect 580967 1019620 581167 1019664
rect 581182 1019654 581206 1019664
rect 581182 1019630 581216 1019654
rect 581227 1019630 581299 1019664
rect 581182 1019620 581299 1019630
rect 580954 1019596 581299 1019620
rect 580967 1019552 581167 1019596
rect 581182 1019586 581206 1019596
rect 581182 1019562 581216 1019586
rect 581227 1019562 581299 1019596
rect 581182 1019552 581299 1019562
rect 580954 1019528 581299 1019552
rect 580967 1019484 581167 1019528
rect 581182 1019518 581206 1019528
rect 581182 1019494 581216 1019518
rect 581227 1019494 581299 1019528
rect 581182 1019484 581299 1019494
rect 580954 1019460 581299 1019484
rect 580967 1019416 581167 1019460
rect 581182 1019450 581206 1019460
rect 581182 1019426 581216 1019450
rect 581227 1019426 581299 1019460
rect 581182 1019416 581299 1019426
rect 580954 1019392 581299 1019416
rect 580967 1019322 581167 1019392
rect 581182 1019368 581206 1019392
rect 581227 1019322 581299 1019392
rect 581529 1019322 581585 1020322
rect 581601 1019322 581657 1020322
rect 581959 1020300 582159 1020322
rect 582174 1020310 582208 1020334
rect 582962 1020322 582996 1020334
rect 582219 1020310 582291 1020322
rect 582174 1020300 582291 1020310
rect 581946 1020276 582291 1020300
rect 581959 1020232 582159 1020276
rect 582174 1020266 582198 1020276
rect 582174 1020242 582208 1020266
rect 582219 1020242 582291 1020276
rect 582174 1020232 582291 1020242
rect 581946 1020208 582291 1020232
rect 581959 1020164 582159 1020208
rect 582174 1020198 582198 1020208
rect 582174 1020174 582208 1020198
rect 582219 1020174 582291 1020208
rect 582174 1020164 582291 1020174
rect 581946 1020140 582291 1020164
rect 581959 1020096 582159 1020140
rect 582174 1020130 582198 1020140
rect 582174 1020106 582208 1020130
rect 582219 1020106 582291 1020140
rect 582174 1020096 582291 1020106
rect 581946 1020072 582291 1020096
rect 581959 1020028 582159 1020072
rect 582174 1020062 582198 1020072
rect 582174 1020038 582208 1020062
rect 582219 1020038 582291 1020072
rect 582174 1020028 582291 1020038
rect 581946 1020004 582291 1020028
rect 581959 1019960 582159 1020004
rect 582174 1019994 582198 1020004
rect 582174 1019970 582208 1019994
rect 582219 1019970 582291 1020004
rect 582174 1019960 582291 1019970
rect 581946 1019936 582291 1019960
rect 581959 1019892 582159 1019936
rect 582174 1019926 582198 1019936
rect 582174 1019902 582208 1019926
rect 582219 1019902 582291 1019936
rect 582174 1019892 582291 1019902
rect 581946 1019868 582291 1019892
rect 581959 1019824 582159 1019868
rect 582174 1019858 582198 1019868
rect 582174 1019834 582208 1019858
rect 582219 1019834 582291 1019868
rect 582174 1019824 582291 1019834
rect 581946 1019800 582291 1019824
rect 581959 1019756 582159 1019800
rect 582174 1019790 582198 1019800
rect 582174 1019766 582208 1019790
rect 582219 1019766 582291 1019800
rect 582174 1019756 582291 1019766
rect 581946 1019732 582291 1019756
rect 581959 1019688 582159 1019732
rect 582174 1019722 582198 1019732
rect 582174 1019698 582208 1019722
rect 582219 1019698 582291 1019732
rect 582174 1019688 582291 1019698
rect 581946 1019664 582291 1019688
rect 581959 1019620 582159 1019664
rect 582174 1019654 582198 1019664
rect 582174 1019630 582208 1019654
rect 582219 1019630 582291 1019664
rect 582174 1019620 582291 1019630
rect 581946 1019596 582291 1019620
rect 581959 1019552 582159 1019596
rect 582174 1019586 582198 1019596
rect 582174 1019562 582208 1019586
rect 582219 1019562 582291 1019596
rect 582174 1019552 582291 1019562
rect 581946 1019528 582291 1019552
rect 581959 1019484 582159 1019528
rect 582174 1019518 582198 1019528
rect 582174 1019494 582208 1019518
rect 582219 1019494 582291 1019528
rect 582174 1019484 582291 1019494
rect 581946 1019460 582291 1019484
rect 581959 1019416 582159 1019460
rect 582174 1019450 582198 1019460
rect 582174 1019426 582208 1019450
rect 582219 1019426 582291 1019460
rect 582174 1019416 582291 1019426
rect 581946 1019392 582291 1019416
rect 581959 1019322 582159 1019392
rect 582174 1019368 582198 1019392
rect 582219 1019322 582291 1019392
rect 582521 1019322 582577 1020322
rect 582593 1019322 582649 1020322
rect 582951 1020300 583151 1020322
rect 583166 1020310 583200 1020334
rect 583211 1020310 583283 1020322
rect 583166 1020300 583283 1020310
rect 582938 1020276 583283 1020300
rect 582951 1020232 583151 1020276
rect 583166 1020266 583190 1020276
rect 583166 1020242 583200 1020266
rect 583211 1020242 583283 1020276
rect 583166 1020232 583283 1020242
rect 582938 1020208 583283 1020232
rect 582951 1020164 583151 1020208
rect 583166 1020198 583190 1020208
rect 583166 1020174 583200 1020198
rect 583211 1020174 583283 1020208
rect 583166 1020164 583283 1020174
rect 582938 1020140 583283 1020164
rect 582951 1020096 583151 1020140
rect 583166 1020130 583190 1020140
rect 583166 1020106 583200 1020130
rect 583211 1020106 583283 1020140
rect 583166 1020096 583283 1020106
rect 582938 1020072 583283 1020096
rect 582951 1020028 583151 1020072
rect 583166 1020062 583190 1020072
rect 583166 1020038 583200 1020062
rect 583211 1020038 583283 1020072
rect 583166 1020028 583283 1020038
rect 582938 1020004 583283 1020028
rect 582951 1019960 583151 1020004
rect 583166 1019994 583190 1020004
rect 583166 1019970 583200 1019994
rect 583211 1019970 583283 1020004
rect 583166 1019960 583283 1019970
rect 582938 1019936 583283 1019960
rect 582951 1019892 583151 1019936
rect 583166 1019926 583190 1019936
rect 583166 1019902 583200 1019926
rect 583211 1019902 583283 1019936
rect 583166 1019892 583283 1019902
rect 582938 1019868 583283 1019892
rect 582951 1019824 583151 1019868
rect 583166 1019858 583190 1019868
rect 583166 1019834 583200 1019858
rect 583211 1019834 583283 1019868
rect 583166 1019824 583283 1019834
rect 582938 1019800 583283 1019824
rect 582951 1019756 583151 1019800
rect 583166 1019790 583190 1019800
rect 583166 1019766 583200 1019790
rect 583211 1019766 583283 1019800
rect 583166 1019756 583283 1019766
rect 582938 1019732 583283 1019756
rect 582951 1019688 583151 1019732
rect 583166 1019722 583190 1019732
rect 583166 1019698 583200 1019722
rect 583211 1019698 583283 1019732
rect 583166 1019688 583283 1019698
rect 582938 1019664 583283 1019688
rect 582951 1019620 583151 1019664
rect 583166 1019654 583190 1019664
rect 583166 1019630 583200 1019654
rect 583211 1019630 583283 1019664
rect 583166 1019620 583283 1019630
rect 582938 1019596 583283 1019620
rect 582951 1019552 583151 1019596
rect 583166 1019586 583190 1019596
rect 583166 1019562 583200 1019586
rect 583211 1019562 583283 1019596
rect 583166 1019552 583283 1019562
rect 582938 1019528 583283 1019552
rect 582951 1019484 583151 1019528
rect 583166 1019518 583190 1019528
rect 583166 1019494 583200 1019518
rect 583211 1019494 583283 1019528
rect 583166 1019484 583283 1019494
rect 582938 1019460 583283 1019484
rect 582951 1019416 583151 1019460
rect 583166 1019450 583190 1019460
rect 583166 1019426 583200 1019450
rect 583211 1019426 583283 1019460
rect 583166 1019416 583283 1019426
rect 582938 1019392 583283 1019416
rect 582951 1019322 583151 1019392
rect 583166 1019368 583190 1019392
rect 583211 1019322 583283 1019392
rect 583472 1019322 583544 1020322
rect 583610 1019322 583627 1020322
rect 583797 1019322 583830 1020322
rect 61561 1018120 61716 1018210
rect 109561 1018120 109716 1018210
rect 161561 1018120 161716 1018210
rect 213561 1018120 213716 1018210
rect 261561 1018120 261716 1018210
rect 313561 1018120 313716 1018210
rect 365561 1018120 365716 1018210
rect 413561 1018120 413716 1018210
rect 465561 1018120 465716 1018210
rect 517561 1018120 517716 1018210
rect 569561 1018120 569716 1018210
rect 61561 1018084 68702 1018120
rect 109561 1018084 109993 1018120
rect 161561 1018084 168702 1018120
rect 213561 1018084 213993 1018120
rect 261561 1018084 261993 1018120
rect 313561 1018084 313993 1018120
rect 365561 1018084 372702 1018120
rect 413561 1018084 413993 1018120
rect 465561 1018084 472702 1018120
rect 517561 1018084 517993 1018120
rect 569561 1018084 576702 1018120
rect 61680 1018053 61716 1018084
rect 61795 1018053 61829 1018077
rect 61863 1018053 61897 1018077
rect 61931 1018053 61965 1018077
rect 61999 1018053 62033 1018077
rect 62067 1018053 62101 1018077
rect 62135 1018053 62169 1018077
rect 62203 1018053 62237 1018077
rect 62271 1018053 62305 1018077
rect 62339 1018053 62373 1018077
rect 62407 1018053 62441 1018077
rect 62475 1018053 62509 1018077
rect 62543 1018053 62577 1018077
rect 62611 1018053 62645 1018077
rect 62679 1018053 62713 1018077
rect 62747 1018053 62781 1018077
rect 62815 1018053 62849 1018077
rect 62883 1018053 62917 1018077
rect 62951 1018053 62985 1018077
rect 63019 1018053 63053 1018077
rect 63087 1018053 63121 1018077
rect 63155 1018053 63189 1018077
rect 63223 1018053 63257 1018077
rect 63291 1018053 63325 1018077
rect 63359 1018053 63393 1018077
rect 63427 1018053 63461 1018077
rect 63495 1018053 63529 1018077
rect 63563 1018053 63597 1018077
rect 63631 1018053 63665 1018077
rect 63699 1018053 63733 1018077
rect 63767 1018053 63801 1018077
rect 63835 1018053 63869 1018077
rect 63903 1018053 63937 1018077
rect 63971 1018053 64005 1018077
rect 64039 1018053 64073 1018077
rect 64107 1018053 64141 1018077
rect 64175 1018053 64209 1018077
rect 64243 1018053 64277 1018077
rect 64311 1018053 64345 1018077
rect 64379 1018053 64413 1018077
rect 64447 1018053 64481 1018077
rect 64515 1018053 64549 1018077
rect 64583 1018053 64617 1018077
rect 64651 1018053 64685 1018077
rect 64719 1018053 64753 1018077
rect 64787 1018053 64821 1018077
rect 64855 1018053 64889 1018077
rect 64923 1018053 64957 1018077
rect 64991 1018053 65025 1018077
rect 65059 1018053 65093 1018077
rect 65127 1018053 65161 1018077
rect 65225 1018053 65259 1018077
rect 65293 1018053 65327 1018077
rect 65361 1018053 65395 1018077
rect 65429 1018053 65463 1018077
rect 65497 1018053 65531 1018077
rect 65565 1018053 65599 1018077
rect 65633 1018053 65667 1018077
rect 65701 1018053 65735 1018077
rect 65769 1018053 65803 1018077
rect 65837 1018053 65871 1018077
rect 65905 1018053 65939 1018077
rect 65973 1018053 66007 1018077
rect 66041 1018053 66075 1018077
rect 66109 1018053 66143 1018077
rect 66177 1018053 66211 1018077
rect 66245 1018053 66279 1018077
rect 66313 1018053 66347 1018077
rect 66381 1018053 66415 1018077
rect 66449 1018053 66483 1018077
rect 66517 1018053 66551 1018077
rect 66585 1018053 66619 1018077
rect 66653 1018053 66687 1018077
rect 66721 1018053 66755 1018077
rect 66789 1018053 66823 1018077
rect 66857 1018053 66891 1018077
rect 66925 1018053 66959 1018077
rect 66993 1018053 67027 1018077
rect 67061 1018053 67095 1018077
rect 67129 1018053 67163 1018077
rect 67197 1018053 67231 1018077
rect 67265 1018053 67299 1018077
rect 67333 1018053 67367 1018077
rect 67401 1018053 67435 1018077
rect 67469 1018053 67503 1018077
rect 67537 1018053 67571 1018077
rect 67605 1018053 67639 1018077
rect 67673 1018053 67707 1018077
rect 67741 1018053 67775 1018077
rect 67809 1018053 67843 1018077
rect 67877 1018053 67911 1018077
rect 67945 1018053 67979 1018077
rect 68013 1018053 68047 1018077
rect 68081 1018053 68115 1018077
rect 68149 1018053 68183 1018077
rect 68217 1018053 68251 1018077
rect 68285 1018053 68319 1018077
rect 68353 1018053 68387 1018077
rect 68421 1018053 68455 1018077
rect 68489 1018053 68523 1018077
rect 68557 1018053 68591 1018077
rect 68666 1018053 68702 1018084
rect 61680 1018030 68702 1018053
rect 61680 1018017 61795 1018030
rect 61829 1018017 61863 1018030
rect 61897 1018017 61931 1018030
rect 61965 1018017 61999 1018030
rect 62033 1018017 62067 1018030
rect 62101 1018017 62135 1018030
rect 62169 1018017 62203 1018030
rect 62237 1018017 62271 1018030
rect 62305 1018017 62339 1018030
rect 62373 1018017 62407 1018030
rect 62441 1018017 62475 1018030
rect 62509 1018017 62543 1018030
rect 62577 1018017 62611 1018030
rect 62645 1018017 62679 1018030
rect 62713 1018017 62747 1018030
rect 62781 1018017 62815 1018030
rect 62849 1018017 62883 1018030
rect 62917 1018017 62951 1018030
rect 62985 1018017 63019 1018030
rect 63053 1018017 63087 1018030
rect 63121 1018017 63155 1018030
rect 63189 1018017 63223 1018030
rect 63257 1018017 63291 1018030
rect 63325 1018017 63359 1018030
rect 63393 1018017 63427 1018030
rect 63461 1018017 63495 1018030
rect 63529 1018017 63563 1018030
rect 63597 1018017 63631 1018030
rect 63665 1018017 63699 1018030
rect 63733 1018017 63767 1018030
rect 63801 1018017 63835 1018030
rect 63869 1018017 63903 1018030
rect 63937 1018017 63971 1018030
rect 64005 1018017 64039 1018030
rect 64073 1018017 64107 1018030
rect 64141 1018017 64175 1018030
rect 64209 1018017 64243 1018030
rect 64277 1018017 64311 1018030
rect 64345 1018017 64379 1018030
rect 64413 1018017 64447 1018030
rect 64481 1018017 64515 1018030
rect 64549 1018017 64583 1018030
rect 64617 1018017 64651 1018030
rect 64685 1018017 64719 1018030
rect 64753 1018017 64787 1018030
rect 64821 1018017 64855 1018030
rect 64889 1018017 64923 1018030
rect 64957 1018017 64991 1018030
rect 65025 1018017 65059 1018030
rect 65093 1018017 65127 1018030
rect 65161 1018017 65225 1018030
rect 65259 1018017 65293 1018030
rect 65327 1018017 65361 1018030
rect 65395 1018017 65429 1018030
rect 65463 1018017 65497 1018030
rect 65531 1018017 65565 1018030
rect 65599 1018017 65633 1018030
rect 65667 1018017 65701 1018030
rect 65735 1018017 65769 1018030
rect 65803 1018017 65837 1018030
rect 65871 1018017 65905 1018030
rect 65939 1018017 65973 1018030
rect 66007 1018017 66041 1018030
rect 66075 1018017 66109 1018030
rect 66143 1018017 66177 1018030
rect 66211 1018017 66245 1018030
rect 66279 1018017 66313 1018030
rect 66347 1018017 66381 1018030
rect 66415 1018017 66449 1018030
rect 66483 1018017 66517 1018030
rect 66551 1018017 66585 1018030
rect 66619 1018017 66653 1018030
rect 66687 1018017 66721 1018030
rect 66755 1018017 66789 1018030
rect 66823 1018017 66857 1018030
rect 66891 1018017 66925 1018030
rect 66959 1018017 66993 1018030
rect 67027 1018017 67061 1018030
rect 67095 1018017 67129 1018030
rect 67163 1018017 67197 1018030
rect 67231 1018017 67265 1018030
rect 67299 1018017 67333 1018030
rect 67367 1018017 67401 1018030
rect 67435 1018017 67469 1018030
rect 67503 1018017 67537 1018030
rect 67571 1018017 67605 1018030
rect 67639 1018017 67673 1018030
rect 67707 1018017 67741 1018030
rect 67775 1018017 67809 1018030
rect 67843 1018017 67877 1018030
rect 67911 1018017 67945 1018030
rect 67979 1018017 68013 1018030
rect 68047 1018017 68081 1018030
rect 68115 1018017 68149 1018030
rect 68183 1018017 68217 1018030
rect 68251 1018017 68285 1018030
rect 68319 1018017 68353 1018030
rect 68387 1018017 68421 1018030
rect 68455 1018017 68489 1018030
rect 68523 1018017 68557 1018030
rect 68591 1018017 68702 1018030
rect 109680 1018053 109716 1018084
rect 109795 1018053 109829 1018077
rect 109863 1018053 109897 1018077
rect 109931 1018053 109965 1018077
rect 161680 1018053 161716 1018084
rect 161795 1018053 161829 1018077
rect 161863 1018053 161897 1018077
rect 161931 1018053 161965 1018077
rect 161999 1018053 162033 1018077
rect 162067 1018053 162101 1018077
rect 162135 1018053 162169 1018077
rect 162203 1018053 162237 1018077
rect 162271 1018053 162305 1018077
rect 162339 1018053 162373 1018077
rect 162407 1018053 162441 1018077
rect 162475 1018053 162509 1018077
rect 162543 1018053 162577 1018077
rect 162611 1018053 162645 1018077
rect 162679 1018053 162713 1018077
rect 162747 1018053 162781 1018077
rect 162815 1018053 162849 1018077
rect 162883 1018053 162917 1018077
rect 162951 1018053 162985 1018077
rect 163019 1018053 163053 1018077
rect 163087 1018053 163121 1018077
rect 163155 1018053 163189 1018077
rect 163223 1018053 163257 1018077
rect 163291 1018053 163325 1018077
rect 163359 1018053 163393 1018077
rect 163427 1018053 163461 1018077
rect 163495 1018053 163529 1018077
rect 163563 1018053 163597 1018077
rect 163631 1018053 163665 1018077
rect 163699 1018053 163733 1018077
rect 163767 1018053 163801 1018077
rect 163835 1018053 163869 1018077
rect 163903 1018053 163937 1018077
rect 163971 1018053 164005 1018077
rect 164039 1018053 164073 1018077
rect 164107 1018053 164141 1018077
rect 164175 1018053 164209 1018077
rect 164243 1018053 164277 1018077
rect 164311 1018053 164345 1018077
rect 164379 1018053 164413 1018077
rect 164447 1018053 164481 1018077
rect 164515 1018053 164549 1018077
rect 164583 1018053 164617 1018077
rect 164651 1018053 164685 1018077
rect 164719 1018053 164753 1018077
rect 164787 1018053 164821 1018077
rect 164855 1018053 164889 1018077
rect 164923 1018053 164957 1018077
rect 164991 1018053 165025 1018077
rect 165059 1018053 165093 1018077
rect 165127 1018053 165161 1018077
rect 165225 1018053 165259 1018077
rect 165293 1018053 165327 1018077
rect 165361 1018053 165395 1018077
rect 165429 1018053 165463 1018077
rect 165497 1018053 165531 1018077
rect 165565 1018053 165599 1018077
rect 165633 1018053 165667 1018077
rect 165701 1018053 165735 1018077
rect 165769 1018053 165803 1018077
rect 165837 1018053 165871 1018077
rect 165905 1018053 165939 1018077
rect 165973 1018053 166007 1018077
rect 166041 1018053 166075 1018077
rect 166109 1018053 166143 1018077
rect 166177 1018053 166211 1018077
rect 166245 1018053 166279 1018077
rect 166313 1018053 166347 1018077
rect 166381 1018053 166415 1018077
rect 166449 1018053 166483 1018077
rect 166517 1018053 166551 1018077
rect 166585 1018053 166619 1018077
rect 166653 1018053 166687 1018077
rect 166721 1018053 166755 1018077
rect 166789 1018053 166823 1018077
rect 166857 1018053 166891 1018077
rect 166925 1018053 166959 1018077
rect 166993 1018053 167027 1018077
rect 167061 1018053 167095 1018077
rect 167129 1018053 167163 1018077
rect 167197 1018053 167231 1018077
rect 167265 1018053 167299 1018077
rect 167333 1018053 167367 1018077
rect 167401 1018053 167435 1018077
rect 167469 1018053 167503 1018077
rect 167537 1018053 167571 1018077
rect 167605 1018053 167639 1018077
rect 167673 1018053 167707 1018077
rect 167741 1018053 167775 1018077
rect 167809 1018053 167843 1018077
rect 167877 1018053 167911 1018077
rect 167945 1018053 167979 1018077
rect 168013 1018053 168047 1018077
rect 168081 1018053 168115 1018077
rect 168149 1018053 168183 1018077
rect 168217 1018053 168251 1018077
rect 168285 1018053 168319 1018077
rect 168353 1018053 168387 1018077
rect 168421 1018053 168455 1018077
rect 168489 1018053 168523 1018077
rect 168557 1018053 168591 1018077
rect 168666 1018053 168702 1018084
rect 109680 1018030 109993 1018053
rect 109680 1018017 109795 1018030
rect 109829 1018017 109863 1018030
rect 109897 1018017 109931 1018030
rect 109965 1018017 109993 1018030
rect 161680 1018030 168702 1018053
rect 161680 1018017 161795 1018030
rect 161829 1018017 161863 1018030
rect 161897 1018017 161931 1018030
rect 161965 1018017 161999 1018030
rect 162033 1018017 162067 1018030
rect 162101 1018017 162135 1018030
rect 162169 1018017 162203 1018030
rect 162237 1018017 162271 1018030
rect 162305 1018017 162339 1018030
rect 162373 1018017 162407 1018030
rect 162441 1018017 162475 1018030
rect 162509 1018017 162543 1018030
rect 162577 1018017 162611 1018030
rect 162645 1018017 162679 1018030
rect 162713 1018017 162747 1018030
rect 162781 1018017 162815 1018030
rect 162849 1018017 162883 1018030
rect 162917 1018017 162951 1018030
rect 162985 1018017 163019 1018030
rect 163053 1018017 163087 1018030
rect 163121 1018017 163155 1018030
rect 163189 1018017 163223 1018030
rect 163257 1018017 163291 1018030
rect 163325 1018017 163359 1018030
rect 163393 1018017 163427 1018030
rect 163461 1018017 163495 1018030
rect 163529 1018017 163563 1018030
rect 163597 1018017 163631 1018030
rect 163665 1018017 163699 1018030
rect 163733 1018017 163767 1018030
rect 163801 1018017 163835 1018030
rect 163869 1018017 163903 1018030
rect 163937 1018017 163971 1018030
rect 164005 1018017 164039 1018030
rect 164073 1018017 164107 1018030
rect 164141 1018017 164175 1018030
rect 164209 1018017 164243 1018030
rect 164277 1018017 164311 1018030
rect 164345 1018017 164379 1018030
rect 164413 1018017 164447 1018030
rect 164481 1018017 164515 1018030
rect 164549 1018017 164583 1018030
rect 164617 1018017 164651 1018030
rect 164685 1018017 164719 1018030
rect 164753 1018017 164787 1018030
rect 164821 1018017 164855 1018030
rect 164889 1018017 164923 1018030
rect 164957 1018017 164991 1018030
rect 165025 1018017 165059 1018030
rect 165093 1018017 165127 1018030
rect 165161 1018017 165225 1018030
rect 165259 1018017 165293 1018030
rect 165327 1018017 165361 1018030
rect 165395 1018017 165429 1018030
rect 165463 1018017 165497 1018030
rect 165531 1018017 165565 1018030
rect 165599 1018017 165633 1018030
rect 165667 1018017 165701 1018030
rect 165735 1018017 165769 1018030
rect 165803 1018017 165837 1018030
rect 165871 1018017 165905 1018030
rect 165939 1018017 165973 1018030
rect 166007 1018017 166041 1018030
rect 166075 1018017 166109 1018030
rect 166143 1018017 166177 1018030
rect 166211 1018017 166245 1018030
rect 166279 1018017 166313 1018030
rect 166347 1018017 166381 1018030
rect 166415 1018017 166449 1018030
rect 166483 1018017 166517 1018030
rect 166551 1018017 166585 1018030
rect 166619 1018017 166653 1018030
rect 166687 1018017 166721 1018030
rect 166755 1018017 166789 1018030
rect 166823 1018017 166857 1018030
rect 166891 1018017 166925 1018030
rect 166959 1018017 166993 1018030
rect 167027 1018017 167061 1018030
rect 167095 1018017 167129 1018030
rect 167163 1018017 167197 1018030
rect 167231 1018017 167265 1018030
rect 167299 1018017 167333 1018030
rect 167367 1018017 167401 1018030
rect 167435 1018017 167469 1018030
rect 167503 1018017 167537 1018030
rect 167571 1018017 167605 1018030
rect 167639 1018017 167673 1018030
rect 167707 1018017 167741 1018030
rect 167775 1018017 167809 1018030
rect 167843 1018017 167877 1018030
rect 167911 1018017 167945 1018030
rect 167979 1018017 168013 1018030
rect 168047 1018017 168081 1018030
rect 168115 1018017 168149 1018030
rect 168183 1018017 168217 1018030
rect 168251 1018017 168285 1018030
rect 168319 1018017 168353 1018030
rect 168387 1018017 168421 1018030
rect 168455 1018017 168489 1018030
rect 168523 1018017 168557 1018030
rect 168591 1018017 168702 1018030
rect 213680 1018053 213716 1018084
rect 213795 1018053 213829 1018077
rect 213863 1018053 213897 1018077
rect 213931 1018053 213965 1018077
rect 261680 1018053 261716 1018084
rect 261795 1018053 261829 1018077
rect 261863 1018053 261897 1018077
rect 261931 1018053 261965 1018077
rect 313680 1018053 313716 1018084
rect 313795 1018053 313829 1018077
rect 313863 1018053 313897 1018077
rect 313931 1018053 313965 1018077
rect 365680 1018053 365716 1018084
rect 365795 1018053 365829 1018077
rect 365863 1018053 365897 1018077
rect 365931 1018053 365965 1018077
rect 365999 1018053 366033 1018077
rect 366067 1018053 366101 1018077
rect 366135 1018053 366169 1018077
rect 366203 1018053 366237 1018077
rect 366271 1018053 366305 1018077
rect 366339 1018053 366373 1018077
rect 366407 1018053 366441 1018077
rect 366475 1018053 366509 1018077
rect 366543 1018053 366577 1018077
rect 366611 1018053 366645 1018077
rect 366679 1018053 366713 1018077
rect 366747 1018053 366781 1018077
rect 366815 1018053 366849 1018077
rect 366883 1018053 366917 1018077
rect 366951 1018053 366985 1018077
rect 367019 1018053 367053 1018077
rect 367087 1018053 367121 1018077
rect 367155 1018053 367189 1018077
rect 367223 1018053 367257 1018077
rect 367291 1018053 367325 1018077
rect 367359 1018053 367393 1018077
rect 367427 1018053 367461 1018077
rect 367495 1018053 367529 1018077
rect 367563 1018053 367597 1018077
rect 367631 1018053 367665 1018077
rect 367699 1018053 367733 1018077
rect 367767 1018053 367801 1018077
rect 367835 1018053 367869 1018077
rect 367903 1018053 367937 1018077
rect 367971 1018053 368005 1018077
rect 368039 1018053 368073 1018077
rect 368107 1018053 368141 1018077
rect 368175 1018053 368209 1018077
rect 368243 1018053 368277 1018077
rect 368311 1018053 368345 1018077
rect 368379 1018053 368413 1018077
rect 368447 1018053 368481 1018077
rect 368515 1018053 368549 1018077
rect 368583 1018053 368617 1018077
rect 368651 1018053 368685 1018077
rect 368719 1018053 368753 1018077
rect 368787 1018053 368821 1018077
rect 368855 1018053 368889 1018077
rect 368923 1018053 368957 1018077
rect 368991 1018053 369025 1018077
rect 369059 1018053 369093 1018077
rect 369127 1018053 369161 1018077
rect 369225 1018053 369259 1018077
rect 369293 1018053 369327 1018077
rect 369361 1018053 369395 1018077
rect 369429 1018053 369463 1018077
rect 369497 1018053 369531 1018077
rect 369565 1018053 369599 1018077
rect 369633 1018053 369667 1018077
rect 369701 1018053 369735 1018077
rect 369769 1018053 369803 1018077
rect 369837 1018053 369871 1018077
rect 369905 1018053 369939 1018077
rect 369973 1018053 370007 1018077
rect 370041 1018053 370075 1018077
rect 370109 1018053 370143 1018077
rect 370177 1018053 370211 1018077
rect 370245 1018053 370279 1018077
rect 370313 1018053 370347 1018077
rect 370381 1018053 370415 1018077
rect 370449 1018053 370483 1018077
rect 370517 1018053 370551 1018077
rect 370585 1018053 370619 1018077
rect 370653 1018053 370687 1018077
rect 370721 1018053 370755 1018077
rect 370789 1018053 370823 1018077
rect 370857 1018053 370891 1018077
rect 370925 1018053 370959 1018077
rect 370993 1018053 371027 1018077
rect 371061 1018053 371095 1018077
rect 371129 1018053 371163 1018077
rect 371197 1018053 371231 1018077
rect 371265 1018053 371299 1018077
rect 371333 1018053 371367 1018077
rect 371401 1018053 371435 1018077
rect 371469 1018053 371503 1018077
rect 371537 1018053 371571 1018077
rect 371605 1018053 371639 1018077
rect 371673 1018053 371707 1018077
rect 371741 1018053 371775 1018077
rect 371809 1018053 371843 1018077
rect 371877 1018053 371911 1018077
rect 371945 1018053 371979 1018077
rect 372013 1018053 372047 1018077
rect 372081 1018053 372115 1018077
rect 372149 1018053 372183 1018077
rect 372217 1018053 372251 1018077
rect 372285 1018053 372319 1018077
rect 372353 1018053 372387 1018077
rect 372421 1018053 372455 1018077
rect 372489 1018053 372523 1018077
rect 372557 1018053 372591 1018077
rect 372666 1018053 372702 1018084
rect 213680 1018030 213993 1018053
rect 213680 1018017 213795 1018030
rect 213829 1018017 213863 1018030
rect 213897 1018017 213931 1018030
rect 213965 1018017 213993 1018030
rect 261680 1018030 261993 1018053
rect 261680 1018017 261795 1018030
rect 261829 1018017 261863 1018030
rect 261897 1018017 261931 1018030
rect 261965 1018017 261993 1018030
rect 313680 1018030 313993 1018053
rect 313680 1018017 313795 1018030
rect 313829 1018017 313863 1018030
rect 313897 1018017 313931 1018030
rect 313965 1018017 313993 1018030
rect 365680 1018030 372702 1018053
rect 365680 1018017 365795 1018030
rect 365829 1018017 365863 1018030
rect 365897 1018017 365931 1018030
rect 365965 1018017 365999 1018030
rect 366033 1018017 366067 1018030
rect 366101 1018017 366135 1018030
rect 366169 1018017 366203 1018030
rect 366237 1018017 366271 1018030
rect 366305 1018017 366339 1018030
rect 366373 1018017 366407 1018030
rect 366441 1018017 366475 1018030
rect 366509 1018017 366543 1018030
rect 366577 1018017 366611 1018030
rect 366645 1018017 366679 1018030
rect 366713 1018017 366747 1018030
rect 366781 1018017 366815 1018030
rect 366849 1018017 366883 1018030
rect 366917 1018017 366951 1018030
rect 366985 1018017 367019 1018030
rect 367053 1018017 367087 1018030
rect 367121 1018017 367155 1018030
rect 367189 1018017 367223 1018030
rect 367257 1018017 367291 1018030
rect 367325 1018017 367359 1018030
rect 367393 1018017 367427 1018030
rect 367461 1018017 367495 1018030
rect 367529 1018017 367563 1018030
rect 367597 1018017 367631 1018030
rect 367665 1018017 367699 1018030
rect 367733 1018017 367767 1018030
rect 367801 1018017 367835 1018030
rect 367869 1018017 367903 1018030
rect 367937 1018017 367971 1018030
rect 368005 1018017 368039 1018030
rect 368073 1018017 368107 1018030
rect 368141 1018017 368175 1018030
rect 368209 1018017 368243 1018030
rect 368277 1018017 368311 1018030
rect 368345 1018017 368379 1018030
rect 368413 1018017 368447 1018030
rect 368481 1018017 368515 1018030
rect 368549 1018017 368583 1018030
rect 368617 1018017 368651 1018030
rect 368685 1018017 368719 1018030
rect 368753 1018017 368787 1018030
rect 368821 1018017 368855 1018030
rect 368889 1018017 368923 1018030
rect 368957 1018017 368991 1018030
rect 369025 1018017 369059 1018030
rect 369093 1018017 369127 1018030
rect 369161 1018017 369225 1018030
rect 369259 1018017 369293 1018030
rect 369327 1018017 369361 1018030
rect 369395 1018017 369429 1018030
rect 369463 1018017 369497 1018030
rect 369531 1018017 369565 1018030
rect 369599 1018017 369633 1018030
rect 369667 1018017 369701 1018030
rect 369735 1018017 369769 1018030
rect 369803 1018017 369837 1018030
rect 369871 1018017 369905 1018030
rect 369939 1018017 369973 1018030
rect 370007 1018017 370041 1018030
rect 370075 1018017 370109 1018030
rect 370143 1018017 370177 1018030
rect 370211 1018017 370245 1018030
rect 370279 1018017 370313 1018030
rect 370347 1018017 370381 1018030
rect 370415 1018017 370449 1018030
rect 370483 1018017 370517 1018030
rect 370551 1018017 370585 1018030
rect 370619 1018017 370653 1018030
rect 370687 1018017 370721 1018030
rect 370755 1018017 370789 1018030
rect 370823 1018017 370857 1018030
rect 370891 1018017 370925 1018030
rect 370959 1018017 370993 1018030
rect 371027 1018017 371061 1018030
rect 371095 1018017 371129 1018030
rect 371163 1018017 371197 1018030
rect 371231 1018017 371265 1018030
rect 371299 1018017 371333 1018030
rect 371367 1018017 371401 1018030
rect 371435 1018017 371469 1018030
rect 371503 1018017 371537 1018030
rect 371571 1018017 371605 1018030
rect 371639 1018017 371673 1018030
rect 371707 1018017 371741 1018030
rect 371775 1018017 371809 1018030
rect 371843 1018017 371877 1018030
rect 371911 1018017 371945 1018030
rect 371979 1018017 372013 1018030
rect 372047 1018017 372081 1018030
rect 372115 1018017 372149 1018030
rect 372183 1018017 372217 1018030
rect 372251 1018017 372285 1018030
rect 372319 1018017 372353 1018030
rect 372387 1018017 372421 1018030
rect 372455 1018017 372489 1018030
rect 372523 1018017 372557 1018030
rect 372591 1018017 372702 1018030
rect 413680 1018053 413716 1018084
rect 413795 1018053 413829 1018077
rect 413863 1018053 413897 1018077
rect 413931 1018053 413965 1018077
rect 465680 1018053 465716 1018084
rect 465795 1018053 465829 1018077
rect 465863 1018053 465897 1018077
rect 465931 1018053 465965 1018077
rect 465999 1018053 466033 1018077
rect 466067 1018053 466101 1018077
rect 466135 1018053 466169 1018077
rect 466203 1018053 466237 1018077
rect 466271 1018053 466305 1018077
rect 466339 1018053 466373 1018077
rect 466407 1018053 466441 1018077
rect 466475 1018053 466509 1018077
rect 466543 1018053 466577 1018077
rect 466611 1018053 466645 1018077
rect 466679 1018053 466713 1018077
rect 466747 1018053 466781 1018077
rect 466815 1018053 466849 1018077
rect 466883 1018053 466917 1018077
rect 466951 1018053 466985 1018077
rect 467019 1018053 467053 1018077
rect 467087 1018053 467121 1018077
rect 467155 1018053 467189 1018077
rect 467223 1018053 467257 1018077
rect 467291 1018053 467325 1018077
rect 467359 1018053 467393 1018077
rect 467427 1018053 467461 1018077
rect 467495 1018053 467529 1018077
rect 467563 1018053 467597 1018077
rect 467631 1018053 467665 1018077
rect 467699 1018053 467733 1018077
rect 467767 1018053 467801 1018077
rect 467835 1018053 467869 1018077
rect 467903 1018053 467937 1018077
rect 467971 1018053 468005 1018077
rect 468039 1018053 468073 1018077
rect 468107 1018053 468141 1018077
rect 468175 1018053 468209 1018077
rect 468243 1018053 468277 1018077
rect 468311 1018053 468345 1018077
rect 468379 1018053 468413 1018077
rect 468447 1018053 468481 1018077
rect 468515 1018053 468549 1018077
rect 468583 1018053 468617 1018077
rect 468651 1018053 468685 1018077
rect 468719 1018053 468753 1018077
rect 468787 1018053 468821 1018077
rect 468855 1018053 468889 1018077
rect 468923 1018053 468957 1018077
rect 468991 1018053 469025 1018077
rect 469059 1018053 469093 1018077
rect 469127 1018053 469161 1018077
rect 469225 1018053 469259 1018077
rect 469293 1018053 469327 1018077
rect 469361 1018053 469395 1018077
rect 469429 1018053 469463 1018077
rect 469497 1018053 469531 1018077
rect 469565 1018053 469599 1018077
rect 469633 1018053 469667 1018077
rect 469701 1018053 469735 1018077
rect 469769 1018053 469803 1018077
rect 469837 1018053 469871 1018077
rect 469905 1018053 469939 1018077
rect 469973 1018053 470007 1018077
rect 470041 1018053 470075 1018077
rect 470109 1018053 470143 1018077
rect 470177 1018053 470211 1018077
rect 470245 1018053 470279 1018077
rect 470313 1018053 470347 1018077
rect 470381 1018053 470415 1018077
rect 470449 1018053 470483 1018077
rect 470517 1018053 470551 1018077
rect 470585 1018053 470619 1018077
rect 470653 1018053 470687 1018077
rect 470721 1018053 470755 1018077
rect 470789 1018053 470823 1018077
rect 470857 1018053 470891 1018077
rect 470925 1018053 470959 1018077
rect 470993 1018053 471027 1018077
rect 471061 1018053 471095 1018077
rect 471129 1018053 471163 1018077
rect 471197 1018053 471231 1018077
rect 471265 1018053 471299 1018077
rect 471333 1018053 471367 1018077
rect 471401 1018053 471435 1018077
rect 471469 1018053 471503 1018077
rect 471537 1018053 471571 1018077
rect 471605 1018053 471639 1018077
rect 471673 1018053 471707 1018077
rect 471741 1018053 471775 1018077
rect 471809 1018053 471843 1018077
rect 471877 1018053 471911 1018077
rect 471945 1018053 471979 1018077
rect 472013 1018053 472047 1018077
rect 472081 1018053 472115 1018077
rect 472149 1018053 472183 1018077
rect 472217 1018053 472251 1018077
rect 472285 1018053 472319 1018077
rect 472353 1018053 472387 1018077
rect 472421 1018053 472455 1018077
rect 472489 1018053 472523 1018077
rect 472557 1018053 472591 1018077
rect 472666 1018053 472702 1018084
rect 413680 1018030 413993 1018053
rect 413680 1018017 413795 1018030
rect 413829 1018017 413863 1018030
rect 413897 1018017 413931 1018030
rect 413965 1018017 413993 1018030
rect 465680 1018030 472702 1018053
rect 465680 1018017 465795 1018030
rect 465829 1018017 465863 1018030
rect 465897 1018017 465931 1018030
rect 465965 1018017 465999 1018030
rect 466033 1018017 466067 1018030
rect 466101 1018017 466135 1018030
rect 466169 1018017 466203 1018030
rect 466237 1018017 466271 1018030
rect 466305 1018017 466339 1018030
rect 466373 1018017 466407 1018030
rect 466441 1018017 466475 1018030
rect 466509 1018017 466543 1018030
rect 466577 1018017 466611 1018030
rect 466645 1018017 466679 1018030
rect 466713 1018017 466747 1018030
rect 466781 1018017 466815 1018030
rect 466849 1018017 466883 1018030
rect 466917 1018017 466951 1018030
rect 466985 1018017 467019 1018030
rect 467053 1018017 467087 1018030
rect 467121 1018017 467155 1018030
rect 467189 1018017 467223 1018030
rect 467257 1018017 467291 1018030
rect 467325 1018017 467359 1018030
rect 467393 1018017 467427 1018030
rect 467461 1018017 467495 1018030
rect 467529 1018017 467563 1018030
rect 467597 1018017 467631 1018030
rect 467665 1018017 467699 1018030
rect 467733 1018017 467767 1018030
rect 467801 1018017 467835 1018030
rect 467869 1018017 467903 1018030
rect 467937 1018017 467971 1018030
rect 468005 1018017 468039 1018030
rect 468073 1018017 468107 1018030
rect 468141 1018017 468175 1018030
rect 468209 1018017 468243 1018030
rect 468277 1018017 468311 1018030
rect 468345 1018017 468379 1018030
rect 468413 1018017 468447 1018030
rect 468481 1018017 468515 1018030
rect 468549 1018017 468583 1018030
rect 468617 1018017 468651 1018030
rect 468685 1018017 468719 1018030
rect 468753 1018017 468787 1018030
rect 468821 1018017 468855 1018030
rect 468889 1018017 468923 1018030
rect 468957 1018017 468991 1018030
rect 469025 1018017 469059 1018030
rect 469093 1018017 469127 1018030
rect 469161 1018017 469225 1018030
rect 469259 1018017 469293 1018030
rect 469327 1018017 469361 1018030
rect 469395 1018017 469429 1018030
rect 469463 1018017 469497 1018030
rect 469531 1018017 469565 1018030
rect 469599 1018017 469633 1018030
rect 469667 1018017 469701 1018030
rect 469735 1018017 469769 1018030
rect 469803 1018017 469837 1018030
rect 469871 1018017 469905 1018030
rect 469939 1018017 469973 1018030
rect 470007 1018017 470041 1018030
rect 470075 1018017 470109 1018030
rect 470143 1018017 470177 1018030
rect 470211 1018017 470245 1018030
rect 470279 1018017 470313 1018030
rect 470347 1018017 470381 1018030
rect 470415 1018017 470449 1018030
rect 470483 1018017 470517 1018030
rect 470551 1018017 470585 1018030
rect 470619 1018017 470653 1018030
rect 470687 1018017 470721 1018030
rect 470755 1018017 470789 1018030
rect 470823 1018017 470857 1018030
rect 470891 1018017 470925 1018030
rect 470959 1018017 470993 1018030
rect 471027 1018017 471061 1018030
rect 471095 1018017 471129 1018030
rect 471163 1018017 471197 1018030
rect 471231 1018017 471265 1018030
rect 471299 1018017 471333 1018030
rect 471367 1018017 471401 1018030
rect 471435 1018017 471469 1018030
rect 471503 1018017 471537 1018030
rect 471571 1018017 471605 1018030
rect 471639 1018017 471673 1018030
rect 471707 1018017 471741 1018030
rect 471775 1018017 471809 1018030
rect 471843 1018017 471877 1018030
rect 471911 1018017 471945 1018030
rect 471979 1018017 472013 1018030
rect 472047 1018017 472081 1018030
rect 472115 1018017 472149 1018030
rect 472183 1018017 472217 1018030
rect 472251 1018017 472285 1018030
rect 472319 1018017 472353 1018030
rect 472387 1018017 472421 1018030
rect 472455 1018017 472489 1018030
rect 472523 1018017 472557 1018030
rect 472591 1018017 472702 1018030
rect 517680 1018053 517716 1018084
rect 517795 1018053 517829 1018077
rect 517863 1018053 517897 1018077
rect 517931 1018053 517965 1018077
rect 569680 1018053 569716 1018084
rect 569795 1018053 569829 1018077
rect 569863 1018053 569897 1018077
rect 569931 1018053 569965 1018077
rect 569999 1018053 570033 1018077
rect 570067 1018053 570101 1018077
rect 570135 1018053 570169 1018077
rect 570203 1018053 570237 1018077
rect 570271 1018053 570305 1018077
rect 570339 1018053 570373 1018077
rect 570407 1018053 570441 1018077
rect 570475 1018053 570509 1018077
rect 570543 1018053 570577 1018077
rect 570611 1018053 570645 1018077
rect 570679 1018053 570713 1018077
rect 570747 1018053 570781 1018077
rect 570815 1018053 570849 1018077
rect 570883 1018053 570917 1018077
rect 570951 1018053 570985 1018077
rect 571019 1018053 571053 1018077
rect 571087 1018053 571121 1018077
rect 571155 1018053 571189 1018077
rect 571223 1018053 571257 1018077
rect 571291 1018053 571325 1018077
rect 571359 1018053 571393 1018077
rect 571427 1018053 571461 1018077
rect 571495 1018053 571529 1018077
rect 571563 1018053 571597 1018077
rect 571631 1018053 571665 1018077
rect 571699 1018053 571733 1018077
rect 571767 1018053 571801 1018077
rect 571835 1018053 571869 1018077
rect 571903 1018053 571937 1018077
rect 571971 1018053 572005 1018077
rect 572039 1018053 572073 1018077
rect 572107 1018053 572141 1018077
rect 572175 1018053 572209 1018077
rect 572243 1018053 572277 1018077
rect 572311 1018053 572345 1018077
rect 572379 1018053 572413 1018077
rect 572447 1018053 572481 1018077
rect 572515 1018053 572549 1018077
rect 572583 1018053 572617 1018077
rect 572651 1018053 572685 1018077
rect 572719 1018053 572753 1018077
rect 572787 1018053 572821 1018077
rect 572855 1018053 572889 1018077
rect 572923 1018053 572957 1018077
rect 572991 1018053 573025 1018077
rect 573059 1018053 573093 1018077
rect 573127 1018053 573161 1018077
rect 573225 1018053 573259 1018077
rect 573293 1018053 573327 1018077
rect 573361 1018053 573395 1018077
rect 573429 1018053 573463 1018077
rect 573497 1018053 573531 1018077
rect 573565 1018053 573599 1018077
rect 573633 1018053 573667 1018077
rect 573701 1018053 573735 1018077
rect 573769 1018053 573803 1018077
rect 573837 1018053 573871 1018077
rect 573905 1018053 573939 1018077
rect 573973 1018053 574007 1018077
rect 574041 1018053 574075 1018077
rect 574109 1018053 574143 1018077
rect 574177 1018053 574211 1018077
rect 574245 1018053 574279 1018077
rect 574313 1018053 574347 1018077
rect 574381 1018053 574415 1018077
rect 574449 1018053 574483 1018077
rect 574517 1018053 574551 1018077
rect 574585 1018053 574619 1018077
rect 574653 1018053 574687 1018077
rect 574721 1018053 574755 1018077
rect 574789 1018053 574823 1018077
rect 574857 1018053 574891 1018077
rect 574925 1018053 574959 1018077
rect 574993 1018053 575027 1018077
rect 575061 1018053 575095 1018077
rect 575129 1018053 575163 1018077
rect 575197 1018053 575231 1018077
rect 575265 1018053 575299 1018077
rect 575333 1018053 575367 1018077
rect 575401 1018053 575435 1018077
rect 575469 1018053 575503 1018077
rect 575537 1018053 575571 1018077
rect 575605 1018053 575639 1018077
rect 575673 1018053 575707 1018077
rect 575741 1018053 575775 1018077
rect 575809 1018053 575843 1018077
rect 575877 1018053 575911 1018077
rect 575945 1018053 575979 1018077
rect 576013 1018053 576047 1018077
rect 576081 1018053 576115 1018077
rect 576149 1018053 576183 1018077
rect 576217 1018053 576251 1018077
rect 576285 1018053 576319 1018077
rect 576353 1018053 576387 1018077
rect 576421 1018053 576455 1018077
rect 576489 1018053 576523 1018077
rect 576557 1018053 576591 1018077
rect 576666 1018053 576702 1018084
rect 517680 1018030 517993 1018053
rect 517680 1018017 517795 1018030
rect 517829 1018017 517863 1018030
rect 517897 1018017 517931 1018030
rect 517965 1018017 517993 1018030
rect 569680 1018030 576702 1018053
rect 569680 1018017 569795 1018030
rect 569829 1018017 569863 1018030
rect 569897 1018017 569931 1018030
rect 569965 1018017 569999 1018030
rect 570033 1018017 570067 1018030
rect 570101 1018017 570135 1018030
rect 570169 1018017 570203 1018030
rect 570237 1018017 570271 1018030
rect 570305 1018017 570339 1018030
rect 570373 1018017 570407 1018030
rect 570441 1018017 570475 1018030
rect 570509 1018017 570543 1018030
rect 570577 1018017 570611 1018030
rect 570645 1018017 570679 1018030
rect 570713 1018017 570747 1018030
rect 570781 1018017 570815 1018030
rect 570849 1018017 570883 1018030
rect 570917 1018017 570951 1018030
rect 570985 1018017 571019 1018030
rect 571053 1018017 571087 1018030
rect 571121 1018017 571155 1018030
rect 571189 1018017 571223 1018030
rect 571257 1018017 571291 1018030
rect 571325 1018017 571359 1018030
rect 571393 1018017 571427 1018030
rect 571461 1018017 571495 1018030
rect 571529 1018017 571563 1018030
rect 571597 1018017 571631 1018030
rect 571665 1018017 571699 1018030
rect 571733 1018017 571767 1018030
rect 571801 1018017 571835 1018030
rect 571869 1018017 571903 1018030
rect 571937 1018017 571971 1018030
rect 572005 1018017 572039 1018030
rect 572073 1018017 572107 1018030
rect 572141 1018017 572175 1018030
rect 572209 1018017 572243 1018030
rect 572277 1018017 572311 1018030
rect 572345 1018017 572379 1018030
rect 572413 1018017 572447 1018030
rect 572481 1018017 572515 1018030
rect 572549 1018017 572583 1018030
rect 572617 1018017 572651 1018030
rect 572685 1018017 572719 1018030
rect 572753 1018017 572787 1018030
rect 572821 1018017 572855 1018030
rect 572889 1018017 572923 1018030
rect 572957 1018017 572991 1018030
rect 573025 1018017 573059 1018030
rect 573093 1018017 573127 1018030
rect 573161 1018017 573225 1018030
rect 573259 1018017 573293 1018030
rect 573327 1018017 573361 1018030
rect 573395 1018017 573429 1018030
rect 573463 1018017 573497 1018030
rect 573531 1018017 573565 1018030
rect 573599 1018017 573633 1018030
rect 573667 1018017 573701 1018030
rect 573735 1018017 573769 1018030
rect 573803 1018017 573837 1018030
rect 573871 1018017 573905 1018030
rect 573939 1018017 573973 1018030
rect 574007 1018017 574041 1018030
rect 574075 1018017 574109 1018030
rect 574143 1018017 574177 1018030
rect 574211 1018017 574245 1018030
rect 574279 1018017 574313 1018030
rect 574347 1018017 574381 1018030
rect 574415 1018017 574449 1018030
rect 574483 1018017 574517 1018030
rect 574551 1018017 574585 1018030
rect 574619 1018017 574653 1018030
rect 574687 1018017 574721 1018030
rect 574755 1018017 574789 1018030
rect 574823 1018017 574857 1018030
rect 574891 1018017 574925 1018030
rect 574959 1018017 574993 1018030
rect 575027 1018017 575061 1018030
rect 575095 1018017 575129 1018030
rect 575163 1018017 575197 1018030
rect 575231 1018017 575265 1018030
rect 575299 1018017 575333 1018030
rect 575367 1018017 575401 1018030
rect 575435 1018017 575469 1018030
rect 575503 1018017 575537 1018030
rect 575571 1018017 575605 1018030
rect 575639 1018017 575673 1018030
rect 575707 1018017 575741 1018030
rect 575775 1018017 575809 1018030
rect 575843 1018017 575877 1018030
rect 575911 1018017 575945 1018030
rect 575979 1018017 576013 1018030
rect 576047 1018017 576081 1018030
rect 576115 1018017 576149 1018030
rect 576183 1018017 576217 1018030
rect 576251 1018017 576285 1018030
rect 576319 1018017 576353 1018030
rect 576387 1018017 576421 1018030
rect 576455 1018017 576489 1018030
rect 576523 1018017 576557 1018030
rect 576591 1018017 576702 1018030
rect 62482 1017706 63482 1017756
rect 63612 1017706 65012 1017756
rect 65374 1017706 66774 1017756
rect 66904 1017706 68304 1017756
rect 110482 1017706 111253 1017756
rect 162482 1017706 163482 1017756
rect 163612 1017706 165012 1017756
rect 165374 1017706 166774 1017756
rect 166904 1017706 168304 1017756
rect 214482 1017706 215253 1017756
rect 314482 1017706 315253 1017756
rect 366482 1017706 367482 1017756
rect 367612 1017706 369012 1017756
rect 369374 1017706 370774 1017756
rect 370904 1017706 372304 1017756
rect 414482 1017706 415253 1017756
rect 466482 1017706 467482 1017756
rect 467612 1017706 469012 1017756
rect 469374 1017706 470774 1017756
rect 470904 1017706 472304 1017756
rect 518482 1017706 519253 1017756
rect 570482 1017706 571482 1017756
rect 571612 1017706 573012 1017756
rect 573374 1017706 574774 1017756
rect 574904 1017706 576304 1017756
rect 62482 1017550 63482 1017678
rect 63612 1017550 65012 1017678
rect 65374 1017550 66774 1017678
rect 66904 1017550 68304 1017678
rect 62482 1017394 63482 1017522
rect 63612 1017394 65012 1017522
rect 65374 1017394 66774 1017522
rect 66904 1017394 68304 1017522
rect 62482 1017238 63482 1017366
rect 63612 1017238 65012 1017366
rect 65374 1017238 66774 1017366
rect 66904 1017238 68304 1017366
rect 70315 1017314 70485 1017620
rect 162482 1017550 163482 1017678
rect 163612 1017550 165012 1017678
rect 165374 1017550 166774 1017678
rect 166904 1017550 168304 1017678
rect 162482 1017394 163482 1017522
rect 163612 1017394 165012 1017522
rect 165374 1017394 166774 1017522
rect 166904 1017394 168304 1017522
rect 73603 1017284 73619 1017350
rect 75627 1017284 75643 1017350
rect 123627 1017284 123643 1017350
rect 162482 1017238 163482 1017366
rect 163612 1017238 165012 1017366
rect 165374 1017238 166774 1017366
rect 166904 1017238 168304 1017366
rect 170315 1017314 170485 1017620
rect 366482 1017550 367482 1017678
rect 367612 1017550 369012 1017678
rect 369374 1017550 370774 1017678
rect 370904 1017550 372304 1017678
rect 366482 1017394 367482 1017522
rect 367612 1017394 369012 1017522
rect 369374 1017394 370774 1017522
rect 370904 1017394 372304 1017522
rect 173603 1017284 173619 1017350
rect 175627 1017284 175643 1017350
rect 227627 1017284 227643 1017350
rect 275627 1017284 275643 1017350
rect 327627 1017284 327643 1017350
rect 366482 1017238 367482 1017366
rect 367612 1017238 369012 1017366
rect 369374 1017238 370774 1017366
rect 370904 1017238 372304 1017366
rect 374315 1017314 374485 1017620
rect 466482 1017550 467482 1017678
rect 467612 1017550 469012 1017678
rect 469374 1017550 470774 1017678
rect 470904 1017550 472304 1017678
rect 466482 1017394 467482 1017522
rect 467612 1017394 469012 1017522
rect 469374 1017394 470774 1017522
rect 470904 1017394 472304 1017522
rect 377603 1017284 377619 1017350
rect 379627 1017284 379643 1017350
rect 427627 1017284 427643 1017350
rect 466482 1017238 467482 1017366
rect 467612 1017238 469012 1017366
rect 469374 1017238 470774 1017366
rect 470904 1017238 472304 1017366
rect 474315 1017314 474485 1017620
rect 570482 1017550 571482 1017678
rect 571612 1017550 573012 1017678
rect 573374 1017550 574774 1017678
rect 574904 1017550 576304 1017678
rect 570482 1017394 571482 1017522
rect 571612 1017394 573012 1017522
rect 573374 1017394 574774 1017522
rect 574904 1017394 576304 1017522
rect 477603 1017284 477619 1017350
rect 479627 1017284 479643 1017350
rect 531627 1017284 531643 1017350
rect 570482 1017238 571482 1017366
rect 571612 1017238 573012 1017366
rect 573374 1017238 574774 1017366
rect 574904 1017238 576304 1017366
rect 578315 1017314 578485 1017620
rect 581603 1017284 581619 1017350
rect 583627 1017284 583643 1017350
rect 62482 1017088 63482 1017138
rect 63612 1017088 65012 1017138
rect 65374 1017088 66774 1017138
rect 66904 1017088 68304 1017138
rect 110482 1017088 111253 1017138
rect 162482 1017088 163482 1017138
rect 163612 1017088 165012 1017138
rect 165374 1017088 166774 1017138
rect 166904 1017088 168304 1017138
rect 214482 1017088 215253 1017138
rect 314482 1017088 315253 1017138
rect 366482 1017088 367482 1017138
rect 367612 1017088 369012 1017138
rect 369374 1017088 370774 1017138
rect 370904 1017088 372304 1017138
rect 414482 1017088 415253 1017138
rect 466482 1017088 467482 1017138
rect 467612 1017088 469012 1017138
rect 469374 1017088 470774 1017138
rect 470904 1017088 472304 1017138
rect 518482 1017088 519253 1017138
rect 570482 1017088 571482 1017138
rect 571612 1017088 573012 1017138
rect 573374 1017088 574774 1017138
rect 574904 1017088 576304 1017138
rect 62640 1016651 62674 1016675
rect 62708 1016651 62742 1016675
rect 62776 1016651 62810 1016675
rect 62844 1016651 62878 1016675
rect 62912 1016651 62946 1016675
rect 62980 1016651 63014 1016675
rect 63048 1016651 63082 1016675
rect 63116 1016651 63150 1016675
rect 63184 1016651 63218 1016675
rect 63252 1016651 63286 1016675
rect 63320 1016651 63354 1016675
rect 63388 1016651 63422 1016675
rect 63456 1016651 63490 1016675
rect 63524 1016651 63558 1016675
rect 63592 1016651 63626 1016675
rect 63660 1016651 63694 1016675
rect 63728 1016651 63762 1016675
rect 63796 1016651 63830 1016675
rect 63864 1016651 63898 1016675
rect 63932 1016651 63966 1016675
rect 64000 1016651 64034 1016675
rect 64068 1016651 64102 1016675
rect 64136 1016651 64170 1016675
rect 64204 1016651 64238 1016675
rect 64272 1016651 64306 1016675
rect 64340 1016651 64374 1016675
rect 64408 1016651 64442 1016675
rect 64476 1016651 64510 1016675
rect 64544 1016651 64578 1016675
rect 64612 1016651 64646 1016675
rect 64680 1016651 64714 1016675
rect 64748 1016651 64782 1016675
rect 64816 1016651 64850 1016675
rect 64884 1016651 64918 1016675
rect 64952 1016651 64986 1016675
rect 65020 1016651 65054 1016675
rect 65088 1016651 65122 1016675
rect 65156 1016651 65190 1016675
rect 65224 1016651 65258 1016675
rect 65292 1016651 65326 1016675
rect 65360 1016651 65394 1016675
rect 65428 1016651 65462 1016675
rect 65496 1016651 65530 1016675
rect 65564 1016651 65598 1016675
rect 65632 1016651 65666 1016675
rect 65700 1016651 65734 1016675
rect 65768 1016651 65802 1016675
rect 65836 1016651 65870 1016675
rect 65904 1016651 65938 1016675
rect 65972 1016651 66006 1016675
rect 66040 1016651 66074 1016675
rect 66108 1016651 66142 1016675
rect 66176 1016651 66210 1016675
rect 66244 1016651 66278 1016675
rect 66312 1016651 66346 1016675
rect 66380 1016651 66414 1016675
rect 66448 1016660 66482 1016675
rect 66430 1016651 66482 1016660
rect 66430 1016626 66448 1016651
rect 66464 1016626 66482 1016651
rect 66505 1016626 66506 1016651
rect 66464 1016617 66506 1016626
rect 40933 1016597 41053 1016600
rect 60733 1016597 60853 1016600
rect 63015 1016287 66015 1016337
rect 63015 1016131 66015 1016259
rect 66464 1016215 66566 1016239
rect 66464 1016191 66488 1016215
rect 66542 1016191 66566 1016215
rect 67947 1016191 67981 1016249
rect 68136 1016215 68170 1016249
rect 68208 1016215 68242 1016249
rect 68280 1016215 68314 1016249
rect 68352 1016215 68386 1016249
rect 68136 1016191 68160 1016215
rect 68362 1016191 68386 1016215
rect 68540 1016215 68642 1016239
rect 69770 1016228 69794 1016252
rect 69668 1016215 69692 1016218
rect 68540 1016191 68564 1016215
rect 68618 1016191 68642 1016215
rect 69746 1016204 69770 1016218
rect 69923 1016215 70025 1016239
rect 63015 1015975 66015 1016103
rect 63015 1015819 66015 1015947
rect 63015 1015663 66015 1015791
rect 63015 1015507 66015 1015635
rect 63015 1015351 66015 1015479
rect 63015 1015201 66015 1015251
rect 66852 1014787 66895 1016187
rect 67002 1014787 67130 1016187
rect 67165 1014787 67293 1016187
rect 67328 1014787 67456 1016187
rect 67491 1014787 67619 1016187
rect 67654 1014787 67782 1016187
rect 67817 1014787 67860 1016187
rect 68729 1014787 68779 1016187
rect 68886 1014787 69014 1016187
rect 69049 1014787 69177 1016187
rect 69212 1014787 69340 1016187
rect 69375 1014787 69503 1016187
rect 69538 1014787 69581 1016187
rect 69644 1016170 69668 1016194
rect 69770 1016170 69794 1016194
rect 69923 1016191 69947 1016215
rect 70001 1016191 70025 1016215
rect 63508 1014388 63678 1014694
rect 64308 1014388 64478 1014694
rect 65108 1014388 65278 1014694
rect 63508 1013888 63678 1014194
rect 64308 1013888 64478 1014194
rect 65108 1013888 65278 1014194
rect 60965 1012428 61015 1013028
rect 61115 1012428 61243 1013028
rect 61271 1012428 61399 1013028
rect 61427 1012428 61483 1013028
rect 61583 1012428 61711 1013028
rect 61739 1012428 61867 1013028
rect 61895 1012428 61945 1013028
rect 62025 1012428 62075 1013028
rect 62175 1012428 62225 1013028
rect 62663 1012427 62713 1013027
rect 62813 1012427 62941 1013027
rect 62969 1012427 63097 1013027
rect 63125 1012427 63181 1013027
rect 63281 1012427 63409 1013027
rect 63437 1012427 63565 1013027
rect 63593 1012427 63643 1013027
rect 63723 1012427 63773 1013027
rect 63873 1012427 63923 1013027
rect 64045 1012427 64095 1013027
rect 64195 1012427 64245 1013027
rect 64325 1012427 64375 1013027
rect 64475 1012427 64603 1013027
rect 64631 1012427 64759 1013027
rect 64787 1012427 64843 1013027
rect 64943 1012427 65071 1013027
rect 65099 1012427 65227 1013027
rect 65255 1012427 65305 1013027
rect 66852 1012515 66895 1013915
rect 67002 1012515 67130 1013915
rect 67165 1012515 67293 1013915
rect 67328 1012515 67456 1013915
rect 67491 1012515 67619 1013915
rect 67654 1012515 67782 1013915
rect 67817 1012515 67860 1013915
rect 66464 1012487 66566 1012511
rect 66542 1012463 66566 1012487
rect 67947 1012463 67981 1012521
rect 68136 1012487 68170 1012521
rect 68208 1012487 68242 1012521
rect 68280 1012487 68314 1012521
rect 68352 1012487 68386 1012521
rect 68729 1012515 68779 1013915
rect 68886 1012515 69014 1013915
rect 69049 1012515 69177 1013915
rect 69212 1012515 69340 1013915
rect 69375 1012515 69503 1013915
rect 69538 1012515 69581 1013915
rect 68136 1012463 68160 1012487
rect 68362 1012463 68386 1012487
rect 68540 1012487 68642 1012511
rect 69644 1012508 69668 1012532
rect 69770 1012508 69794 1012532
rect 68540 1012463 68564 1012487
rect 68618 1012463 68642 1012487
rect 69668 1012484 69692 1012487
rect 69746 1012484 69770 1012498
rect 69923 1012487 70025 1012511
rect 69770 1012450 69794 1012474
rect 69923 1012463 69947 1012487
rect 70001 1012463 70025 1012487
rect 70201 1012047 70737 1016655
rect 162640 1016651 162674 1016675
rect 162708 1016651 162742 1016675
rect 162776 1016651 162810 1016675
rect 162844 1016651 162878 1016675
rect 162912 1016651 162946 1016675
rect 162980 1016651 163014 1016675
rect 163048 1016651 163082 1016675
rect 163116 1016651 163150 1016675
rect 163184 1016651 163218 1016675
rect 163252 1016651 163286 1016675
rect 163320 1016651 163354 1016675
rect 163388 1016651 163422 1016675
rect 163456 1016651 163490 1016675
rect 163524 1016651 163558 1016675
rect 163592 1016651 163626 1016675
rect 163660 1016651 163694 1016675
rect 163728 1016651 163762 1016675
rect 163796 1016651 163830 1016675
rect 163864 1016651 163898 1016675
rect 163932 1016651 163966 1016675
rect 164000 1016651 164034 1016675
rect 164068 1016651 164102 1016675
rect 164136 1016651 164170 1016675
rect 164204 1016651 164238 1016675
rect 164272 1016651 164306 1016675
rect 164340 1016651 164374 1016675
rect 164408 1016651 164442 1016675
rect 164476 1016651 164510 1016675
rect 164544 1016651 164578 1016675
rect 164612 1016651 164646 1016675
rect 164680 1016651 164714 1016675
rect 164748 1016651 164782 1016675
rect 164816 1016651 164850 1016675
rect 164884 1016651 164918 1016675
rect 164952 1016651 164986 1016675
rect 165020 1016651 165054 1016675
rect 165088 1016651 165122 1016675
rect 165156 1016651 165190 1016675
rect 165224 1016651 165258 1016675
rect 165292 1016651 165326 1016675
rect 165360 1016651 165394 1016675
rect 165428 1016651 165462 1016675
rect 165496 1016651 165530 1016675
rect 165564 1016651 165598 1016675
rect 165632 1016651 165666 1016675
rect 165700 1016651 165734 1016675
rect 165768 1016651 165802 1016675
rect 165836 1016651 165870 1016675
rect 165904 1016651 165938 1016675
rect 165972 1016651 166006 1016675
rect 166040 1016651 166074 1016675
rect 166108 1016651 166142 1016675
rect 166176 1016651 166210 1016675
rect 166244 1016651 166278 1016675
rect 166312 1016651 166346 1016675
rect 166380 1016651 166414 1016675
rect 166448 1016660 166482 1016675
rect 166430 1016651 166482 1016660
rect 166430 1016626 166448 1016651
rect 166464 1016626 166482 1016651
rect 166505 1016626 166506 1016651
rect 166464 1016617 166506 1016626
rect 76933 1016597 77053 1016600
rect 108733 1016597 108853 1016600
rect 124933 1016597 125053 1016600
rect 160733 1016597 160853 1016600
rect 73496 1016414 73510 1016438
rect 73462 1016390 73486 1016414
rect 73520 1016390 73544 1016414
rect 76716 1016340 76750 1016360
rect 124716 1016340 124750 1016360
rect 111015 1016287 111253 1016337
rect 163015 1016287 166015 1016337
rect 73119 1016227 73143 1016251
rect 73177 1016227 73201 1016251
rect 73653 1016245 73687 1016249
rect 73721 1016245 73755 1016249
rect 73789 1016245 73823 1016249
rect 73857 1016245 73891 1016249
rect 73925 1016245 73959 1016249
rect 73993 1016245 74027 1016249
rect 74061 1016245 74095 1016249
rect 74129 1016245 74163 1016249
rect 74197 1016245 74231 1016249
rect 74265 1016245 74299 1016249
rect 74333 1016245 74367 1016249
rect 74401 1016245 74435 1016249
rect 74469 1016245 74503 1016249
rect 74537 1016245 74571 1016249
rect 74605 1016245 74639 1016249
rect 74673 1016245 74707 1016249
rect 74741 1016245 74775 1016249
rect 74809 1016245 74843 1016249
rect 74877 1016245 74911 1016249
rect 74945 1016245 74979 1016249
rect 75013 1016245 75047 1016249
rect 75081 1016245 75115 1016249
rect 75149 1016245 75183 1016249
rect 75217 1016245 75251 1016249
rect 75285 1016245 75319 1016249
rect 75353 1016245 75387 1016249
rect 75421 1016245 75455 1016249
rect 75489 1016245 75523 1016249
rect 75557 1016245 75591 1016249
rect 75625 1016245 75659 1016249
rect 75693 1016245 75727 1016249
rect 75761 1016245 75795 1016249
rect 75829 1016245 75863 1016249
rect 75897 1016245 75931 1016249
rect 75965 1016245 75999 1016249
rect 76033 1016245 76067 1016249
rect 76101 1016245 76135 1016249
rect 76169 1016245 76203 1016249
rect 76237 1016245 76271 1016249
rect 76305 1016245 76339 1016249
rect 76373 1016245 76407 1016249
rect 73585 1016227 76485 1016245
rect 73653 1016223 73687 1016227
rect 73721 1016223 73755 1016227
rect 73789 1016223 73823 1016227
rect 73857 1016223 73891 1016227
rect 73925 1016223 73959 1016227
rect 73993 1016223 74027 1016227
rect 74061 1016223 74095 1016227
rect 74129 1016223 74163 1016227
rect 74197 1016223 74231 1016227
rect 74265 1016223 74299 1016227
rect 74333 1016223 74367 1016227
rect 74401 1016223 74435 1016227
rect 74469 1016223 74503 1016227
rect 74537 1016223 74571 1016227
rect 74605 1016223 74639 1016227
rect 74673 1016223 74707 1016227
rect 74741 1016223 74775 1016227
rect 74809 1016223 74843 1016227
rect 74877 1016223 74911 1016227
rect 74945 1016223 74979 1016227
rect 75013 1016223 75047 1016227
rect 75081 1016223 75115 1016227
rect 75149 1016223 75183 1016227
rect 75217 1016223 75251 1016227
rect 75285 1016223 75319 1016227
rect 75353 1016223 75387 1016227
rect 75421 1016223 75455 1016227
rect 75489 1016223 75523 1016227
rect 75557 1016223 75591 1016227
rect 75625 1016223 75659 1016227
rect 75693 1016223 75727 1016227
rect 75761 1016223 75795 1016227
rect 75829 1016223 75863 1016227
rect 75897 1016223 75931 1016227
rect 75965 1016223 75999 1016227
rect 76033 1016223 76067 1016227
rect 76101 1016223 76135 1016227
rect 76169 1016223 76203 1016227
rect 76237 1016223 76271 1016227
rect 76305 1016223 76339 1016227
rect 76373 1016223 76407 1016227
rect 76624 1016224 76648 1016248
rect 123489 1016245 123523 1016249
rect 123557 1016245 123591 1016249
rect 123625 1016245 123659 1016249
rect 123693 1016245 123727 1016249
rect 123761 1016245 123795 1016249
rect 123829 1016245 123863 1016249
rect 123897 1016245 123931 1016249
rect 123965 1016245 123999 1016249
rect 124033 1016245 124067 1016249
rect 124101 1016245 124135 1016249
rect 124169 1016245 124203 1016249
rect 124237 1016245 124271 1016249
rect 124305 1016245 124339 1016249
rect 124373 1016245 124407 1016249
rect 73143 1016203 73177 1016217
rect 73589 1016215 76481 1016223
rect 73629 1016203 76431 1016215
rect 76648 1016200 76672 1016215
rect 76716 1016204 76750 1016239
rect 123473 1016227 124485 1016245
rect 123489 1016223 123523 1016227
rect 123557 1016223 123591 1016227
rect 123625 1016223 123659 1016227
rect 123693 1016223 123727 1016227
rect 123761 1016223 123795 1016227
rect 123829 1016223 123863 1016227
rect 123897 1016223 123931 1016227
rect 123965 1016223 123999 1016227
rect 124033 1016223 124067 1016227
rect 124101 1016223 124135 1016227
rect 124169 1016223 124203 1016227
rect 124237 1016223 124271 1016227
rect 124305 1016223 124339 1016227
rect 124373 1016223 124407 1016227
rect 124624 1016224 124648 1016248
rect 70771 1014787 70899 1016187
rect 70934 1014787 71062 1016187
rect 71097 1014787 71225 1016187
rect 71260 1014787 71388 1016187
rect 71423 1014787 71551 1016187
rect 71586 1014787 71714 1016187
rect 71749 1014787 71792 1016187
rect 71885 1014787 71928 1016187
rect 72035 1014787 72163 1016187
rect 72198 1014787 72326 1016187
rect 72361 1014787 72489 1016187
rect 72524 1014787 72652 1016187
rect 72687 1014787 72815 1016187
rect 72850 1014787 72978 1016187
rect 73013 1014787 73063 1016187
rect 73119 1016169 73143 1016193
rect 73177 1016169 73201 1016193
rect 76726 1016191 76750 1016204
rect 123473 1016215 124481 1016223
rect 123473 1016203 124431 1016215
rect 124648 1016200 124672 1016215
rect 124716 1016204 124750 1016239
rect 124726 1016191 124750 1016204
rect 163015 1016131 166015 1016259
rect 166464 1016215 166566 1016239
rect 166464 1016191 166488 1016215
rect 166542 1016191 166566 1016215
rect 167947 1016191 167981 1016249
rect 168136 1016215 168170 1016249
rect 168208 1016215 168242 1016249
rect 168280 1016215 168314 1016249
rect 168352 1016215 168386 1016249
rect 168136 1016191 168160 1016215
rect 168362 1016191 168386 1016215
rect 168540 1016215 168642 1016239
rect 169770 1016228 169794 1016252
rect 169668 1016215 169692 1016218
rect 168540 1016191 168564 1016215
rect 168618 1016191 168642 1016215
rect 169746 1016204 169770 1016218
rect 169923 1016215 170025 1016239
rect 73330 1014402 73432 1015966
rect 73699 1014719 73749 1016119
rect 73856 1014719 73984 1016119
rect 74019 1014719 74147 1016119
rect 74182 1014719 74310 1016119
rect 74345 1014719 74473 1016119
rect 74508 1014719 74636 1016119
rect 74671 1014719 74799 1016119
rect 74834 1014719 74877 1016119
rect 74970 1014719 75013 1016119
rect 75120 1014719 75248 1016119
rect 75283 1014719 75411 1016119
rect 75446 1014719 75574 1016119
rect 75609 1014719 75737 1016119
rect 75772 1014719 75900 1016119
rect 75935 1014719 76063 1016119
rect 76098 1014719 76226 1016119
rect 76261 1014719 76304 1016119
rect 111015 1015201 111253 1015251
rect 122834 1014719 122877 1016119
rect 122970 1014719 123013 1016119
rect 123473 1014719 123574 1016119
rect 123609 1014719 123737 1016119
rect 123772 1014719 123900 1016119
rect 123935 1014719 124063 1016119
rect 124098 1014719 124226 1016119
rect 124261 1014719 124304 1016119
rect 163015 1015975 166015 1016103
rect 163015 1015819 166015 1015947
rect 163015 1015663 166015 1015791
rect 163015 1015507 166015 1015635
rect 163015 1015351 166015 1015479
rect 163015 1015201 166015 1015251
rect 166852 1014787 166895 1016187
rect 167002 1014787 167130 1016187
rect 167165 1014787 167293 1016187
rect 167328 1014787 167456 1016187
rect 167491 1014787 167619 1016187
rect 167654 1014787 167782 1016187
rect 167817 1014787 167860 1016187
rect 168729 1014787 168779 1016187
rect 168886 1014787 169014 1016187
rect 169049 1014787 169177 1016187
rect 169212 1014787 169340 1016187
rect 169375 1014787 169503 1016187
rect 169538 1014787 169581 1016187
rect 169644 1016170 169668 1016194
rect 169770 1016170 169794 1016194
rect 169923 1016191 169947 1016215
rect 170001 1016191 170025 1016215
rect 73364 1014378 73398 1014402
rect 163508 1014388 163678 1014694
rect 164308 1014388 164478 1014694
rect 165108 1014388 165278 1014694
rect 73364 1014300 73398 1014324
rect 70771 1012515 70899 1013915
rect 70934 1012515 71062 1013915
rect 71097 1012515 71225 1013915
rect 71260 1012515 71388 1013915
rect 71423 1012515 71551 1013915
rect 71586 1012515 71714 1013915
rect 71749 1012515 71792 1013915
rect 71885 1012515 71928 1013915
rect 72035 1012515 72163 1013915
rect 72198 1012515 72326 1013915
rect 72361 1012515 72489 1013915
rect 72524 1012515 72652 1013915
rect 72687 1012515 72815 1013915
rect 72850 1012515 72978 1013915
rect 73013 1012515 73063 1013915
rect 73330 1012736 73432 1014300
rect 73699 1012583 73749 1013983
rect 73856 1012583 73984 1013983
rect 74019 1012583 74147 1013983
rect 74182 1012583 74310 1013983
rect 74345 1012583 74473 1013983
rect 74508 1012583 74636 1013983
rect 74671 1012583 74799 1013983
rect 74834 1012583 74877 1013983
rect 74970 1012583 75013 1013983
rect 75120 1012583 75248 1013983
rect 75283 1012583 75411 1013983
rect 75446 1012583 75574 1013983
rect 75609 1012583 75737 1013983
rect 75772 1012583 75900 1013983
rect 75935 1012583 76063 1013983
rect 76098 1012583 76226 1013983
rect 76261 1012583 76304 1013983
rect 73119 1012509 73143 1012533
rect 73177 1012509 73201 1012533
rect 73653 1012517 73687 1012521
rect 73721 1012517 73755 1012521
rect 73789 1012517 73823 1012521
rect 73857 1012517 73891 1012521
rect 73925 1012517 73959 1012521
rect 73993 1012517 74027 1012521
rect 74061 1012517 74095 1012521
rect 74129 1012517 74163 1012521
rect 74197 1012517 74231 1012521
rect 74265 1012517 74299 1012521
rect 74333 1012517 74367 1012521
rect 74401 1012517 74435 1012521
rect 74469 1012517 74503 1012521
rect 74537 1012517 74571 1012521
rect 74605 1012517 74639 1012521
rect 74673 1012517 74707 1012521
rect 74741 1012517 74775 1012521
rect 74809 1012517 74843 1012521
rect 74877 1012517 74911 1012521
rect 74945 1012517 74979 1012521
rect 75013 1012517 75047 1012521
rect 75081 1012517 75115 1012521
rect 75149 1012517 75183 1012521
rect 75217 1012517 75251 1012521
rect 75285 1012517 75319 1012521
rect 75353 1012517 75387 1012521
rect 75421 1012517 75455 1012521
rect 75489 1012517 75523 1012521
rect 75557 1012517 75591 1012521
rect 75625 1012517 75659 1012521
rect 75693 1012517 75727 1012521
rect 75761 1012517 75795 1012521
rect 75829 1012517 75863 1012521
rect 75897 1012517 75931 1012521
rect 75965 1012517 75999 1012521
rect 76033 1012517 76067 1012521
rect 76101 1012517 76135 1012521
rect 76169 1012517 76203 1012521
rect 76237 1012517 76271 1012521
rect 76305 1012517 76339 1012521
rect 76373 1012517 76407 1012521
rect 73619 1012509 76451 1012517
rect 76682 1012512 76750 1012532
rect 73653 1012505 73687 1012509
rect 73721 1012505 73755 1012509
rect 73789 1012505 73823 1012509
rect 73857 1012505 73891 1012509
rect 73925 1012505 73959 1012509
rect 73993 1012505 74027 1012509
rect 74061 1012505 74095 1012509
rect 74129 1012505 74163 1012509
rect 74197 1012505 74231 1012509
rect 74265 1012505 74299 1012509
rect 74333 1012505 74367 1012509
rect 74401 1012505 74435 1012509
rect 74469 1012505 74503 1012509
rect 74537 1012505 74571 1012509
rect 74605 1012505 74639 1012509
rect 74673 1012505 74707 1012509
rect 74741 1012505 74775 1012509
rect 74809 1012505 74843 1012509
rect 74877 1012505 74911 1012509
rect 74945 1012505 74979 1012509
rect 75013 1012505 75047 1012509
rect 75081 1012505 75115 1012509
rect 75149 1012505 75183 1012509
rect 75217 1012505 75251 1012509
rect 75285 1012505 75319 1012509
rect 75353 1012505 75387 1012509
rect 75421 1012505 75455 1012509
rect 75489 1012505 75523 1012509
rect 75557 1012505 75591 1012509
rect 75625 1012505 75659 1012509
rect 75693 1012505 75727 1012509
rect 75761 1012505 75795 1012509
rect 75829 1012505 75863 1012509
rect 75897 1012505 75931 1012509
rect 75965 1012505 75999 1012509
rect 76033 1012505 76067 1012509
rect 76101 1012505 76135 1012509
rect 76169 1012505 76203 1012509
rect 76237 1012505 76271 1012509
rect 76305 1012505 76339 1012509
rect 76373 1012505 76407 1012509
rect 73143 1012485 73177 1012499
rect 73585 1012487 76485 1012505
rect 76648 1012487 76672 1012502
rect 76716 1012487 76750 1012512
rect 73629 1012485 76431 1012487
rect 73119 1012451 73143 1012475
rect 73177 1012451 73201 1012475
rect 76624 1012454 76648 1012478
rect 76726 1012463 76750 1012487
rect 108965 1012428 109015 1013028
rect 109115 1012428 109243 1013028
rect 109271 1012428 109399 1013028
rect 109427 1012428 109483 1013028
rect 109583 1012428 109711 1013028
rect 109739 1012428 109867 1013028
rect 109895 1012428 109945 1013028
rect 110025 1012428 110075 1013028
rect 110175 1012428 110225 1013028
rect 110663 1012427 110713 1013027
rect 111125 1012427 111181 1013027
rect 122834 1012583 122877 1013983
rect 122970 1012583 123013 1013983
rect 123473 1012583 123574 1013983
rect 123609 1012583 123737 1013983
rect 123772 1012583 123900 1013983
rect 123935 1012583 124063 1013983
rect 124098 1012583 124226 1013983
rect 124261 1012583 124304 1013983
rect 163508 1013888 163678 1014194
rect 164308 1013888 164478 1014194
rect 165108 1013888 165278 1014194
rect 123489 1012517 123523 1012521
rect 123557 1012517 123591 1012521
rect 123625 1012517 123659 1012521
rect 123693 1012517 123727 1012521
rect 123761 1012517 123795 1012521
rect 123829 1012517 123863 1012521
rect 123897 1012517 123931 1012521
rect 123965 1012517 123999 1012521
rect 124033 1012517 124067 1012521
rect 124101 1012517 124135 1012521
rect 124169 1012517 124203 1012521
rect 124237 1012517 124271 1012521
rect 124305 1012517 124339 1012521
rect 124373 1012517 124407 1012521
rect 123473 1012509 124451 1012517
rect 124682 1012512 124750 1012532
rect 123489 1012505 123523 1012509
rect 123557 1012505 123591 1012509
rect 123625 1012505 123659 1012509
rect 123693 1012505 123727 1012509
rect 123761 1012505 123795 1012509
rect 123829 1012505 123863 1012509
rect 123897 1012505 123931 1012509
rect 123965 1012505 123999 1012509
rect 124033 1012505 124067 1012509
rect 124101 1012505 124135 1012509
rect 124169 1012505 124203 1012509
rect 124237 1012505 124271 1012509
rect 124305 1012505 124339 1012509
rect 124373 1012505 124407 1012509
rect 123473 1012487 124485 1012505
rect 124648 1012487 124672 1012502
rect 124716 1012487 124750 1012512
rect 123473 1012485 124431 1012487
rect 124624 1012454 124648 1012478
rect 124726 1012463 124750 1012487
rect 160965 1012428 161015 1013028
rect 161115 1012428 161243 1013028
rect 161271 1012428 161399 1013028
rect 161427 1012428 161483 1013028
rect 161583 1012428 161711 1013028
rect 161739 1012428 161867 1013028
rect 161895 1012428 161945 1013028
rect 162025 1012428 162075 1013028
rect 162175 1012428 162225 1013028
rect 162663 1012427 162713 1013027
rect 162813 1012427 162941 1013027
rect 162969 1012427 163097 1013027
rect 163125 1012427 163181 1013027
rect 163281 1012427 163409 1013027
rect 163437 1012427 163565 1013027
rect 163593 1012427 163643 1013027
rect 163723 1012427 163773 1013027
rect 163873 1012427 163923 1013027
rect 164045 1012427 164095 1013027
rect 164195 1012427 164245 1013027
rect 164325 1012427 164375 1013027
rect 164475 1012427 164603 1013027
rect 164631 1012427 164759 1013027
rect 164787 1012427 164843 1013027
rect 164943 1012427 165071 1013027
rect 165099 1012427 165227 1013027
rect 165255 1012427 165305 1013027
rect 166852 1012515 166895 1013915
rect 167002 1012515 167130 1013915
rect 167165 1012515 167293 1013915
rect 167328 1012515 167456 1013915
rect 167491 1012515 167619 1013915
rect 167654 1012515 167782 1013915
rect 167817 1012515 167860 1013915
rect 166464 1012487 166566 1012511
rect 166542 1012463 166566 1012487
rect 167947 1012463 167981 1012521
rect 168136 1012487 168170 1012521
rect 168208 1012487 168242 1012521
rect 168280 1012487 168314 1012521
rect 168352 1012487 168386 1012521
rect 168729 1012515 168779 1013915
rect 168886 1012515 169014 1013915
rect 169049 1012515 169177 1013915
rect 169212 1012515 169340 1013915
rect 169375 1012515 169503 1013915
rect 169538 1012515 169581 1013915
rect 168136 1012463 168160 1012487
rect 168362 1012463 168386 1012487
rect 168540 1012487 168642 1012511
rect 169644 1012508 169668 1012532
rect 169770 1012508 169794 1012532
rect 168540 1012463 168564 1012487
rect 168618 1012463 168642 1012487
rect 169668 1012484 169692 1012487
rect 169746 1012484 169770 1012498
rect 169923 1012487 170025 1012511
rect 169770 1012450 169794 1012474
rect 169923 1012463 169947 1012487
rect 170001 1012463 170025 1012487
rect 76682 1012376 76750 1012396
rect 124682 1012376 124750 1012396
rect 73462 1012288 73486 1012312
rect 73520 1012288 73544 1012312
rect 73496 1012264 73510 1012288
rect 170201 1012047 170737 1016655
rect 366640 1016651 366674 1016675
rect 366708 1016651 366742 1016675
rect 366776 1016651 366810 1016675
rect 366844 1016651 366878 1016675
rect 366912 1016651 366946 1016675
rect 366980 1016651 367014 1016675
rect 367048 1016651 367082 1016675
rect 367116 1016651 367150 1016675
rect 367184 1016651 367218 1016675
rect 367252 1016651 367286 1016675
rect 367320 1016651 367354 1016675
rect 367388 1016651 367422 1016675
rect 367456 1016651 367490 1016675
rect 367524 1016651 367558 1016675
rect 367592 1016651 367626 1016675
rect 367660 1016651 367694 1016675
rect 367728 1016651 367762 1016675
rect 367796 1016651 367830 1016675
rect 367864 1016651 367898 1016675
rect 367932 1016651 367966 1016675
rect 368000 1016651 368034 1016675
rect 368068 1016651 368102 1016675
rect 368136 1016651 368170 1016675
rect 368204 1016651 368238 1016675
rect 368272 1016651 368306 1016675
rect 368340 1016651 368374 1016675
rect 368408 1016651 368442 1016675
rect 368476 1016651 368510 1016675
rect 368544 1016651 368578 1016675
rect 368612 1016651 368646 1016675
rect 368680 1016651 368714 1016675
rect 368748 1016651 368782 1016675
rect 368816 1016651 368850 1016675
rect 368884 1016651 368918 1016675
rect 368952 1016651 368986 1016675
rect 369020 1016651 369054 1016675
rect 369088 1016651 369122 1016675
rect 369156 1016651 369190 1016675
rect 369224 1016651 369258 1016675
rect 369292 1016651 369326 1016675
rect 369360 1016651 369394 1016675
rect 369428 1016651 369462 1016675
rect 369496 1016651 369530 1016675
rect 369564 1016651 369598 1016675
rect 369632 1016651 369666 1016675
rect 369700 1016651 369734 1016675
rect 369768 1016651 369802 1016675
rect 369836 1016651 369870 1016675
rect 369904 1016651 369938 1016675
rect 369972 1016651 370006 1016675
rect 370040 1016651 370074 1016675
rect 370108 1016651 370142 1016675
rect 370176 1016651 370210 1016675
rect 370244 1016651 370278 1016675
rect 370312 1016651 370346 1016675
rect 370380 1016651 370414 1016675
rect 370448 1016660 370482 1016675
rect 370430 1016651 370482 1016660
rect 370430 1016626 370448 1016651
rect 370464 1016626 370482 1016651
rect 370505 1016626 370506 1016651
rect 370464 1016617 370506 1016626
rect 176933 1016597 177053 1016600
rect 212733 1016597 212853 1016600
rect 228933 1016597 229053 1016600
rect 260733 1016597 260853 1016600
rect 276933 1016597 277053 1016600
rect 312733 1016597 312853 1016600
rect 328933 1016597 329053 1016600
rect 364733 1016597 364853 1016600
rect 173496 1016414 173510 1016438
rect 173462 1016390 173486 1016414
rect 173520 1016390 173544 1016414
rect 176716 1016340 176750 1016360
rect 228716 1016340 228750 1016360
rect 276716 1016340 276750 1016360
rect 328716 1016340 328750 1016360
rect 215015 1016287 215253 1016337
rect 315015 1016287 315253 1016337
rect 367015 1016287 370015 1016337
rect 173119 1016227 173143 1016251
rect 173177 1016227 173201 1016251
rect 173653 1016245 173687 1016249
rect 173721 1016245 173755 1016249
rect 173789 1016245 173823 1016249
rect 173857 1016245 173891 1016249
rect 173925 1016245 173959 1016249
rect 173993 1016245 174027 1016249
rect 174061 1016245 174095 1016249
rect 174129 1016245 174163 1016249
rect 174197 1016245 174231 1016249
rect 174265 1016245 174299 1016249
rect 174333 1016245 174367 1016249
rect 174401 1016245 174435 1016249
rect 174469 1016245 174503 1016249
rect 174537 1016245 174571 1016249
rect 174605 1016245 174639 1016249
rect 174673 1016245 174707 1016249
rect 174741 1016245 174775 1016249
rect 174809 1016245 174843 1016249
rect 174877 1016245 174911 1016249
rect 174945 1016245 174979 1016249
rect 175013 1016245 175047 1016249
rect 175081 1016245 175115 1016249
rect 175149 1016245 175183 1016249
rect 175217 1016245 175251 1016249
rect 175285 1016245 175319 1016249
rect 175353 1016245 175387 1016249
rect 175421 1016245 175455 1016249
rect 175489 1016245 175523 1016249
rect 175557 1016245 175591 1016249
rect 175625 1016245 175659 1016249
rect 175693 1016245 175727 1016249
rect 175761 1016245 175795 1016249
rect 175829 1016245 175863 1016249
rect 175897 1016245 175931 1016249
rect 175965 1016245 175999 1016249
rect 176033 1016245 176067 1016249
rect 176101 1016245 176135 1016249
rect 176169 1016245 176203 1016249
rect 176237 1016245 176271 1016249
rect 176305 1016245 176339 1016249
rect 176373 1016245 176407 1016249
rect 173585 1016227 176485 1016245
rect 173653 1016223 173687 1016227
rect 173721 1016223 173755 1016227
rect 173789 1016223 173823 1016227
rect 173857 1016223 173891 1016227
rect 173925 1016223 173959 1016227
rect 173993 1016223 174027 1016227
rect 174061 1016223 174095 1016227
rect 174129 1016223 174163 1016227
rect 174197 1016223 174231 1016227
rect 174265 1016223 174299 1016227
rect 174333 1016223 174367 1016227
rect 174401 1016223 174435 1016227
rect 174469 1016223 174503 1016227
rect 174537 1016223 174571 1016227
rect 174605 1016223 174639 1016227
rect 174673 1016223 174707 1016227
rect 174741 1016223 174775 1016227
rect 174809 1016223 174843 1016227
rect 174877 1016223 174911 1016227
rect 174945 1016223 174979 1016227
rect 175013 1016223 175047 1016227
rect 175081 1016223 175115 1016227
rect 175149 1016223 175183 1016227
rect 175217 1016223 175251 1016227
rect 175285 1016223 175319 1016227
rect 175353 1016223 175387 1016227
rect 175421 1016223 175455 1016227
rect 175489 1016223 175523 1016227
rect 175557 1016223 175591 1016227
rect 175625 1016223 175659 1016227
rect 175693 1016223 175727 1016227
rect 175761 1016223 175795 1016227
rect 175829 1016223 175863 1016227
rect 175897 1016223 175931 1016227
rect 175965 1016223 175999 1016227
rect 176033 1016223 176067 1016227
rect 176101 1016223 176135 1016227
rect 176169 1016223 176203 1016227
rect 176237 1016223 176271 1016227
rect 176305 1016223 176339 1016227
rect 176373 1016223 176407 1016227
rect 176624 1016224 176648 1016248
rect 227489 1016245 227523 1016249
rect 227557 1016245 227591 1016249
rect 227625 1016245 227659 1016249
rect 227693 1016245 227727 1016249
rect 227761 1016245 227795 1016249
rect 227829 1016245 227863 1016249
rect 227897 1016245 227931 1016249
rect 227965 1016245 227999 1016249
rect 228033 1016245 228067 1016249
rect 228101 1016245 228135 1016249
rect 228169 1016245 228203 1016249
rect 228237 1016245 228271 1016249
rect 228305 1016245 228339 1016249
rect 228373 1016245 228407 1016249
rect 173143 1016203 173177 1016217
rect 173589 1016215 176481 1016223
rect 173629 1016203 176431 1016215
rect 176648 1016200 176672 1016215
rect 176716 1016204 176750 1016239
rect 227473 1016227 228485 1016245
rect 227489 1016223 227523 1016227
rect 227557 1016223 227591 1016227
rect 227625 1016223 227659 1016227
rect 227693 1016223 227727 1016227
rect 227761 1016223 227795 1016227
rect 227829 1016223 227863 1016227
rect 227897 1016223 227931 1016227
rect 227965 1016223 227999 1016227
rect 228033 1016223 228067 1016227
rect 228101 1016223 228135 1016227
rect 228169 1016223 228203 1016227
rect 228237 1016223 228271 1016227
rect 228305 1016223 228339 1016227
rect 228373 1016223 228407 1016227
rect 228624 1016224 228648 1016248
rect 275489 1016245 275523 1016249
rect 275557 1016245 275591 1016249
rect 275625 1016245 275659 1016249
rect 275693 1016245 275727 1016249
rect 275761 1016245 275795 1016249
rect 275829 1016245 275863 1016249
rect 275897 1016245 275931 1016249
rect 275965 1016245 275999 1016249
rect 276033 1016245 276067 1016249
rect 276101 1016245 276135 1016249
rect 276169 1016245 276203 1016249
rect 276237 1016245 276271 1016249
rect 276305 1016245 276339 1016249
rect 276373 1016245 276407 1016249
rect 170771 1014787 170899 1016187
rect 170934 1014787 171062 1016187
rect 171097 1014787 171225 1016187
rect 171260 1014787 171388 1016187
rect 171423 1014787 171551 1016187
rect 171586 1014787 171714 1016187
rect 171749 1014787 171792 1016187
rect 171885 1014787 171928 1016187
rect 172035 1014787 172163 1016187
rect 172198 1014787 172326 1016187
rect 172361 1014787 172489 1016187
rect 172524 1014787 172652 1016187
rect 172687 1014787 172815 1016187
rect 172850 1014787 172978 1016187
rect 173013 1014787 173063 1016187
rect 173119 1016169 173143 1016193
rect 173177 1016169 173201 1016193
rect 176726 1016191 176750 1016204
rect 227473 1016215 228481 1016223
rect 227473 1016203 228431 1016215
rect 228648 1016200 228672 1016215
rect 228716 1016204 228750 1016239
rect 275473 1016227 276485 1016245
rect 275489 1016223 275523 1016227
rect 275557 1016223 275591 1016227
rect 275625 1016223 275659 1016227
rect 275693 1016223 275727 1016227
rect 275761 1016223 275795 1016227
rect 275829 1016223 275863 1016227
rect 275897 1016223 275931 1016227
rect 275965 1016223 275999 1016227
rect 276033 1016223 276067 1016227
rect 276101 1016223 276135 1016227
rect 276169 1016223 276203 1016227
rect 276237 1016223 276271 1016227
rect 276305 1016223 276339 1016227
rect 276373 1016223 276407 1016227
rect 276624 1016224 276648 1016248
rect 327489 1016245 327523 1016249
rect 327557 1016245 327591 1016249
rect 327625 1016245 327659 1016249
rect 327693 1016245 327727 1016249
rect 327761 1016245 327795 1016249
rect 327829 1016245 327863 1016249
rect 327897 1016245 327931 1016249
rect 327965 1016245 327999 1016249
rect 328033 1016245 328067 1016249
rect 328101 1016245 328135 1016249
rect 328169 1016245 328203 1016249
rect 328237 1016245 328271 1016249
rect 328305 1016245 328339 1016249
rect 328373 1016245 328407 1016249
rect 228726 1016191 228750 1016204
rect 275473 1016215 276481 1016223
rect 275473 1016203 276431 1016215
rect 276648 1016200 276672 1016215
rect 276716 1016204 276750 1016239
rect 327473 1016227 328485 1016245
rect 327489 1016223 327523 1016227
rect 327557 1016223 327591 1016227
rect 327625 1016223 327659 1016227
rect 327693 1016223 327727 1016227
rect 327761 1016223 327795 1016227
rect 327829 1016223 327863 1016227
rect 327897 1016223 327931 1016227
rect 327965 1016223 327999 1016227
rect 328033 1016223 328067 1016227
rect 328101 1016223 328135 1016227
rect 328169 1016223 328203 1016227
rect 328237 1016223 328271 1016227
rect 328305 1016223 328339 1016227
rect 328373 1016223 328407 1016227
rect 328624 1016224 328648 1016248
rect 276726 1016191 276750 1016204
rect 327473 1016215 328481 1016223
rect 327473 1016203 328431 1016215
rect 328648 1016200 328672 1016215
rect 328716 1016204 328750 1016239
rect 328726 1016191 328750 1016204
rect 367015 1016131 370015 1016259
rect 370464 1016215 370566 1016239
rect 370464 1016191 370488 1016215
rect 370542 1016191 370566 1016215
rect 371947 1016191 371981 1016249
rect 372136 1016215 372170 1016249
rect 372208 1016215 372242 1016249
rect 372280 1016215 372314 1016249
rect 372352 1016215 372386 1016249
rect 372136 1016191 372160 1016215
rect 372362 1016191 372386 1016215
rect 372540 1016215 372642 1016239
rect 373770 1016228 373794 1016252
rect 373668 1016215 373692 1016218
rect 372540 1016191 372564 1016215
rect 372618 1016191 372642 1016215
rect 373746 1016204 373770 1016218
rect 373923 1016215 374025 1016239
rect 173330 1014402 173432 1015966
rect 173699 1014719 173749 1016119
rect 173856 1014719 173984 1016119
rect 174019 1014719 174147 1016119
rect 174182 1014719 174310 1016119
rect 174345 1014719 174473 1016119
rect 174508 1014719 174636 1016119
rect 174671 1014719 174799 1016119
rect 174834 1014719 174877 1016119
rect 174970 1014719 175013 1016119
rect 175120 1014719 175248 1016119
rect 175283 1014719 175411 1016119
rect 175446 1014719 175574 1016119
rect 175609 1014719 175737 1016119
rect 175772 1014719 175900 1016119
rect 175935 1014719 176063 1016119
rect 176098 1014719 176226 1016119
rect 176261 1014719 176304 1016119
rect 215015 1015201 215253 1015251
rect 226834 1014719 226877 1016119
rect 226970 1014719 227013 1016119
rect 227473 1014719 227574 1016119
rect 227609 1014719 227737 1016119
rect 227772 1014719 227900 1016119
rect 227935 1014719 228063 1016119
rect 228098 1014719 228226 1016119
rect 228261 1014719 228304 1016119
rect 274834 1014719 274877 1016119
rect 274970 1014719 275013 1016119
rect 275473 1014719 275574 1016119
rect 275609 1014719 275737 1016119
rect 275772 1014719 275900 1016119
rect 275935 1014719 276063 1016119
rect 276098 1014719 276226 1016119
rect 276261 1014719 276304 1016119
rect 315015 1015201 315253 1015251
rect 326834 1014719 326877 1016119
rect 326970 1014719 327013 1016119
rect 327473 1014719 327574 1016119
rect 327609 1014719 327737 1016119
rect 327772 1014719 327900 1016119
rect 327935 1014719 328063 1016119
rect 328098 1014719 328226 1016119
rect 328261 1014719 328304 1016119
rect 367015 1015975 370015 1016103
rect 367015 1015819 370015 1015947
rect 367015 1015663 370015 1015791
rect 367015 1015507 370015 1015635
rect 367015 1015351 370015 1015479
rect 367015 1015201 370015 1015251
rect 370852 1014787 370895 1016187
rect 371002 1014787 371130 1016187
rect 371165 1014787 371293 1016187
rect 371328 1014787 371456 1016187
rect 371491 1014787 371619 1016187
rect 371654 1014787 371782 1016187
rect 371817 1014787 371860 1016187
rect 372729 1014787 372779 1016187
rect 372886 1014787 373014 1016187
rect 373049 1014787 373177 1016187
rect 373212 1014787 373340 1016187
rect 373375 1014787 373503 1016187
rect 373538 1014787 373581 1016187
rect 373644 1016170 373668 1016194
rect 373770 1016170 373794 1016194
rect 373923 1016191 373947 1016215
rect 374001 1016191 374025 1016215
rect 173364 1014378 173398 1014402
rect 367508 1014388 367678 1014694
rect 368308 1014388 368478 1014694
rect 369108 1014388 369278 1014694
rect 173364 1014300 173398 1014324
rect 170771 1012515 170899 1013915
rect 170934 1012515 171062 1013915
rect 171097 1012515 171225 1013915
rect 171260 1012515 171388 1013915
rect 171423 1012515 171551 1013915
rect 171586 1012515 171714 1013915
rect 171749 1012515 171792 1013915
rect 171885 1012515 171928 1013915
rect 172035 1012515 172163 1013915
rect 172198 1012515 172326 1013915
rect 172361 1012515 172489 1013915
rect 172524 1012515 172652 1013915
rect 172687 1012515 172815 1013915
rect 172850 1012515 172978 1013915
rect 173013 1012515 173063 1013915
rect 173330 1012736 173432 1014300
rect 173699 1012583 173749 1013983
rect 173856 1012583 173984 1013983
rect 174019 1012583 174147 1013983
rect 174182 1012583 174310 1013983
rect 174345 1012583 174473 1013983
rect 174508 1012583 174636 1013983
rect 174671 1012583 174799 1013983
rect 174834 1012583 174877 1013983
rect 174970 1012583 175013 1013983
rect 175120 1012583 175248 1013983
rect 175283 1012583 175411 1013983
rect 175446 1012583 175574 1013983
rect 175609 1012583 175737 1013983
rect 175772 1012583 175900 1013983
rect 175935 1012583 176063 1013983
rect 176098 1012583 176226 1013983
rect 176261 1012583 176304 1013983
rect 173119 1012509 173143 1012533
rect 173177 1012509 173201 1012533
rect 173653 1012517 173687 1012521
rect 173721 1012517 173755 1012521
rect 173789 1012517 173823 1012521
rect 173857 1012517 173891 1012521
rect 173925 1012517 173959 1012521
rect 173993 1012517 174027 1012521
rect 174061 1012517 174095 1012521
rect 174129 1012517 174163 1012521
rect 174197 1012517 174231 1012521
rect 174265 1012517 174299 1012521
rect 174333 1012517 174367 1012521
rect 174401 1012517 174435 1012521
rect 174469 1012517 174503 1012521
rect 174537 1012517 174571 1012521
rect 174605 1012517 174639 1012521
rect 174673 1012517 174707 1012521
rect 174741 1012517 174775 1012521
rect 174809 1012517 174843 1012521
rect 174877 1012517 174911 1012521
rect 174945 1012517 174979 1012521
rect 175013 1012517 175047 1012521
rect 175081 1012517 175115 1012521
rect 175149 1012517 175183 1012521
rect 175217 1012517 175251 1012521
rect 175285 1012517 175319 1012521
rect 175353 1012517 175387 1012521
rect 175421 1012517 175455 1012521
rect 175489 1012517 175523 1012521
rect 175557 1012517 175591 1012521
rect 175625 1012517 175659 1012521
rect 175693 1012517 175727 1012521
rect 175761 1012517 175795 1012521
rect 175829 1012517 175863 1012521
rect 175897 1012517 175931 1012521
rect 175965 1012517 175999 1012521
rect 176033 1012517 176067 1012521
rect 176101 1012517 176135 1012521
rect 176169 1012517 176203 1012521
rect 176237 1012517 176271 1012521
rect 176305 1012517 176339 1012521
rect 176373 1012517 176407 1012521
rect 173619 1012509 176451 1012517
rect 176682 1012512 176750 1012532
rect 173653 1012505 173687 1012509
rect 173721 1012505 173755 1012509
rect 173789 1012505 173823 1012509
rect 173857 1012505 173891 1012509
rect 173925 1012505 173959 1012509
rect 173993 1012505 174027 1012509
rect 174061 1012505 174095 1012509
rect 174129 1012505 174163 1012509
rect 174197 1012505 174231 1012509
rect 174265 1012505 174299 1012509
rect 174333 1012505 174367 1012509
rect 174401 1012505 174435 1012509
rect 174469 1012505 174503 1012509
rect 174537 1012505 174571 1012509
rect 174605 1012505 174639 1012509
rect 174673 1012505 174707 1012509
rect 174741 1012505 174775 1012509
rect 174809 1012505 174843 1012509
rect 174877 1012505 174911 1012509
rect 174945 1012505 174979 1012509
rect 175013 1012505 175047 1012509
rect 175081 1012505 175115 1012509
rect 175149 1012505 175183 1012509
rect 175217 1012505 175251 1012509
rect 175285 1012505 175319 1012509
rect 175353 1012505 175387 1012509
rect 175421 1012505 175455 1012509
rect 175489 1012505 175523 1012509
rect 175557 1012505 175591 1012509
rect 175625 1012505 175659 1012509
rect 175693 1012505 175727 1012509
rect 175761 1012505 175795 1012509
rect 175829 1012505 175863 1012509
rect 175897 1012505 175931 1012509
rect 175965 1012505 175999 1012509
rect 176033 1012505 176067 1012509
rect 176101 1012505 176135 1012509
rect 176169 1012505 176203 1012509
rect 176237 1012505 176271 1012509
rect 176305 1012505 176339 1012509
rect 176373 1012505 176407 1012509
rect 173143 1012485 173177 1012499
rect 173585 1012487 176485 1012505
rect 176648 1012487 176672 1012502
rect 176716 1012487 176750 1012512
rect 173629 1012485 176431 1012487
rect 173119 1012451 173143 1012475
rect 173177 1012451 173201 1012475
rect 176624 1012454 176648 1012478
rect 176726 1012463 176750 1012487
rect 212965 1012428 213015 1013028
rect 213115 1012428 213243 1013028
rect 213271 1012428 213399 1013028
rect 213427 1012428 213483 1013028
rect 213583 1012428 213711 1013028
rect 213739 1012428 213867 1013028
rect 213895 1012428 213945 1013028
rect 214025 1012428 214075 1013028
rect 214175 1012428 214225 1013028
rect 214663 1012427 214713 1013027
rect 215125 1012427 215181 1013027
rect 226834 1012583 226877 1013983
rect 226970 1012583 227013 1013983
rect 227473 1012583 227574 1013983
rect 227609 1012583 227737 1013983
rect 227772 1012583 227900 1013983
rect 227935 1012583 228063 1013983
rect 228098 1012583 228226 1013983
rect 228261 1012583 228304 1013983
rect 227489 1012517 227523 1012521
rect 227557 1012517 227591 1012521
rect 227625 1012517 227659 1012521
rect 227693 1012517 227727 1012521
rect 227761 1012517 227795 1012521
rect 227829 1012517 227863 1012521
rect 227897 1012517 227931 1012521
rect 227965 1012517 227999 1012521
rect 228033 1012517 228067 1012521
rect 228101 1012517 228135 1012521
rect 228169 1012517 228203 1012521
rect 228237 1012517 228271 1012521
rect 228305 1012517 228339 1012521
rect 228373 1012517 228407 1012521
rect 227473 1012509 228451 1012517
rect 228682 1012512 228750 1012532
rect 227489 1012505 227523 1012509
rect 227557 1012505 227591 1012509
rect 227625 1012505 227659 1012509
rect 227693 1012505 227727 1012509
rect 227761 1012505 227795 1012509
rect 227829 1012505 227863 1012509
rect 227897 1012505 227931 1012509
rect 227965 1012505 227999 1012509
rect 228033 1012505 228067 1012509
rect 228101 1012505 228135 1012509
rect 228169 1012505 228203 1012509
rect 228237 1012505 228271 1012509
rect 228305 1012505 228339 1012509
rect 228373 1012505 228407 1012509
rect 227473 1012487 228485 1012505
rect 228648 1012487 228672 1012502
rect 228716 1012487 228750 1012512
rect 227473 1012485 228431 1012487
rect 228624 1012454 228648 1012478
rect 228726 1012463 228750 1012487
rect 260965 1012428 261015 1013028
rect 261115 1012428 261243 1013028
rect 261271 1012428 261399 1013028
rect 261427 1012428 261483 1013028
rect 261583 1012428 261711 1013028
rect 261739 1012428 261867 1013028
rect 261895 1012428 261945 1013028
rect 262025 1012428 262075 1013028
rect 274834 1012583 274877 1013983
rect 274970 1012583 275013 1013983
rect 275473 1012583 275574 1013983
rect 275609 1012583 275737 1013983
rect 275772 1012583 275900 1013983
rect 275935 1012583 276063 1013983
rect 276098 1012583 276226 1013983
rect 276261 1012583 276304 1013983
rect 275489 1012517 275523 1012521
rect 275557 1012517 275591 1012521
rect 275625 1012517 275659 1012521
rect 275693 1012517 275727 1012521
rect 275761 1012517 275795 1012521
rect 275829 1012517 275863 1012521
rect 275897 1012517 275931 1012521
rect 275965 1012517 275999 1012521
rect 276033 1012517 276067 1012521
rect 276101 1012517 276135 1012521
rect 276169 1012517 276203 1012521
rect 276237 1012517 276271 1012521
rect 276305 1012517 276339 1012521
rect 276373 1012517 276407 1012521
rect 275473 1012509 276451 1012517
rect 276682 1012512 276750 1012532
rect 275489 1012505 275523 1012509
rect 275557 1012505 275591 1012509
rect 275625 1012505 275659 1012509
rect 275693 1012505 275727 1012509
rect 275761 1012505 275795 1012509
rect 275829 1012505 275863 1012509
rect 275897 1012505 275931 1012509
rect 275965 1012505 275999 1012509
rect 276033 1012505 276067 1012509
rect 276101 1012505 276135 1012509
rect 276169 1012505 276203 1012509
rect 276237 1012505 276271 1012509
rect 276305 1012505 276339 1012509
rect 276373 1012505 276407 1012509
rect 275473 1012487 276485 1012505
rect 276648 1012487 276672 1012502
rect 276716 1012487 276750 1012512
rect 275473 1012485 276431 1012487
rect 276624 1012454 276648 1012478
rect 276726 1012463 276750 1012487
rect 312965 1012428 313015 1013028
rect 313115 1012428 313243 1013028
rect 313271 1012428 313399 1013028
rect 313427 1012428 313483 1013028
rect 313583 1012428 313711 1013028
rect 313739 1012428 313867 1013028
rect 313895 1012428 313945 1013028
rect 314025 1012428 314075 1013028
rect 314175 1012428 314225 1013028
rect 314663 1012427 314713 1013027
rect 315125 1012427 315181 1013027
rect 326834 1012583 326877 1013983
rect 326970 1012583 327013 1013983
rect 327473 1012583 327574 1013983
rect 327609 1012583 327737 1013983
rect 327772 1012583 327900 1013983
rect 327935 1012583 328063 1013983
rect 328098 1012583 328226 1013983
rect 328261 1012583 328304 1013983
rect 367508 1013888 367678 1014194
rect 368308 1013888 368478 1014194
rect 369108 1013888 369278 1014194
rect 327489 1012517 327523 1012521
rect 327557 1012517 327591 1012521
rect 327625 1012517 327659 1012521
rect 327693 1012517 327727 1012521
rect 327761 1012517 327795 1012521
rect 327829 1012517 327863 1012521
rect 327897 1012517 327931 1012521
rect 327965 1012517 327999 1012521
rect 328033 1012517 328067 1012521
rect 328101 1012517 328135 1012521
rect 328169 1012517 328203 1012521
rect 328237 1012517 328271 1012521
rect 328305 1012517 328339 1012521
rect 328373 1012517 328407 1012521
rect 327473 1012509 328451 1012517
rect 328682 1012512 328750 1012532
rect 327489 1012505 327523 1012509
rect 327557 1012505 327591 1012509
rect 327625 1012505 327659 1012509
rect 327693 1012505 327727 1012509
rect 327761 1012505 327795 1012509
rect 327829 1012505 327863 1012509
rect 327897 1012505 327931 1012509
rect 327965 1012505 327999 1012509
rect 328033 1012505 328067 1012509
rect 328101 1012505 328135 1012509
rect 328169 1012505 328203 1012509
rect 328237 1012505 328271 1012509
rect 328305 1012505 328339 1012509
rect 328373 1012505 328407 1012509
rect 327473 1012487 328485 1012505
rect 328648 1012487 328672 1012502
rect 328716 1012487 328750 1012512
rect 327473 1012485 328431 1012487
rect 328624 1012454 328648 1012478
rect 328726 1012463 328750 1012487
rect 364965 1012428 365015 1013028
rect 365115 1012428 365243 1013028
rect 365271 1012428 365399 1013028
rect 365427 1012428 365483 1013028
rect 365583 1012428 365711 1013028
rect 365739 1012428 365867 1013028
rect 365895 1012428 365945 1013028
rect 366025 1012428 366075 1013028
rect 366175 1012428 366225 1013028
rect 366663 1012427 366713 1013027
rect 366813 1012427 366941 1013027
rect 366969 1012427 367097 1013027
rect 367125 1012427 367181 1013027
rect 367281 1012427 367409 1013027
rect 367437 1012427 367565 1013027
rect 367593 1012427 367643 1013027
rect 367723 1012427 367773 1013027
rect 367873 1012427 367923 1013027
rect 368045 1012427 368095 1013027
rect 368195 1012427 368245 1013027
rect 368325 1012427 368375 1013027
rect 368475 1012427 368603 1013027
rect 368631 1012427 368759 1013027
rect 368787 1012427 368843 1013027
rect 368943 1012427 369071 1013027
rect 369099 1012427 369227 1013027
rect 369255 1012427 369305 1013027
rect 370852 1012515 370895 1013915
rect 371002 1012515 371130 1013915
rect 371165 1012515 371293 1013915
rect 371328 1012515 371456 1013915
rect 371491 1012515 371619 1013915
rect 371654 1012515 371782 1013915
rect 371817 1012515 371860 1013915
rect 370464 1012487 370566 1012511
rect 370542 1012463 370566 1012487
rect 371947 1012463 371981 1012521
rect 372136 1012487 372170 1012521
rect 372208 1012487 372242 1012521
rect 372280 1012487 372314 1012521
rect 372352 1012487 372386 1012521
rect 372729 1012515 372779 1013915
rect 372886 1012515 373014 1013915
rect 373049 1012515 373177 1013915
rect 373212 1012515 373340 1013915
rect 373375 1012515 373503 1013915
rect 373538 1012515 373581 1013915
rect 372136 1012463 372160 1012487
rect 372362 1012463 372386 1012487
rect 372540 1012487 372642 1012511
rect 373644 1012508 373668 1012532
rect 373770 1012508 373794 1012532
rect 372540 1012463 372564 1012487
rect 372618 1012463 372642 1012487
rect 373668 1012484 373692 1012487
rect 373746 1012484 373770 1012498
rect 373923 1012487 374025 1012511
rect 373770 1012450 373794 1012474
rect 373923 1012463 373947 1012487
rect 374001 1012463 374025 1012487
rect 176682 1012376 176750 1012396
rect 228682 1012376 228750 1012396
rect 276682 1012376 276750 1012396
rect 328682 1012376 328750 1012396
rect 173462 1012288 173486 1012312
rect 173520 1012288 173544 1012312
rect 173496 1012264 173510 1012288
rect 374201 1012047 374737 1016655
rect 466640 1016651 466674 1016675
rect 466708 1016651 466742 1016675
rect 466776 1016651 466810 1016675
rect 466844 1016651 466878 1016675
rect 466912 1016651 466946 1016675
rect 466980 1016651 467014 1016675
rect 467048 1016651 467082 1016675
rect 467116 1016651 467150 1016675
rect 467184 1016651 467218 1016675
rect 467252 1016651 467286 1016675
rect 467320 1016651 467354 1016675
rect 467388 1016651 467422 1016675
rect 467456 1016651 467490 1016675
rect 467524 1016651 467558 1016675
rect 467592 1016651 467626 1016675
rect 467660 1016651 467694 1016675
rect 467728 1016651 467762 1016675
rect 467796 1016651 467830 1016675
rect 467864 1016651 467898 1016675
rect 467932 1016651 467966 1016675
rect 468000 1016651 468034 1016675
rect 468068 1016651 468102 1016675
rect 468136 1016651 468170 1016675
rect 468204 1016651 468238 1016675
rect 468272 1016651 468306 1016675
rect 468340 1016651 468374 1016675
rect 468408 1016651 468442 1016675
rect 468476 1016651 468510 1016675
rect 468544 1016651 468578 1016675
rect 468612 1016651 468646 1016675
rect 468680 1016651 468714 1016675
rect 468748 1016651 468782 1016675
rect 468816 1016651 468850 1016675
rect 468884 1016651 468918 1016675
rect 468952 1016651 468986 1016675
rect 469020 1016651 469054 1016675
rect 469088 1016651 469122 1016675
rect 469156 1016651 469190 1016675
rect 469224 1016651 469258 1016675
rect 469292 1016651 469326 1016675
rect 469360 1016651 469394 1016675
rect 469428 1016651 469462 1016675
rect 469496 1016651 469530 1016675
rect 469564 1016651 469598 1016675
rect 469632 1016651 469666 1016675
rect 469700 1016651 469734 1016675
rect 469768 1016651 469802 1016675
rect 469836 1016651 469870 1016675
rect 469904 1016651 469938 1016675
rect 469972 1016651 470006 1016675
rect 470040 1016651 470074 1016675
rect 470108 1016651 470142 1016675
rect 470176 1016651 470210 1016675
rect 470244 1016651 470278 1016675
rect 470312 1016651 470346 1016675
rect 470380 1016651 470414 1016675
rect 470448 1016660 470482 1016675
rect 470430 1016651 470482 1016660
rect 470430 1016626 470448 1016651
rect 470464 1016626 470482 1016651
rect 470505 1016626 470506 1016651
rect 470464 1016617 470506 1016626
rect 380933 1016597 381053 1016600
rect 412733 1016597 412853 1016600
rect 428933 1016597 429053 1016600
rect 464733 1016597 464853 1016600
rect 377496 1016414 377510 1016438
rect 377462 1016390 377486 1016414
rect 377520 1016390 377544 1016414
rect 380716 1016340 380750 1016360
rect 428716 1016340 428750 1016360
rect 415015 1016287 415253 1016337
rect 467015 1016287 470015 1016337
rect 377119 1016227 377143 1016251
rect 377177 1016227 377201 1016251
rect 377653 1016245 377687 1016249
rect 377721 1016245 377755 1016249
rect 377789 1016245 377823 1016249
rect 377857 1016245 377891 1016249
rect 377925 1016245 377959 1016249
rect 377993 1016245 378027 1016249
rect 378061 1016245 378095 1016249
rect 378129 1016245 378163 1016249
rect 378197 1016245 378231 1016249
rect 378265 1016245 378299 1016249
rect 378333 1016245 378367 1016249
rect 378401 1016245 378435 1016249
rect 378469 1016245 378503 1016249
rect 378537 1016245 378571 1016249
rect 378605 1016245 378639 1016249
rect 378673 1016245 378707 1016249
rect 378741 1016245 378775 1016249
rect 378809 1016245 378843 1016249
rect 378877 1016245 378911 1016249
rect 378945 1016245 378979 1016249
rect 379013 1016245 379047 1016249
rect 379081 1016245 379115 1016249
rect 379149 1016245 379183 1016249
rect 379217 1016245 379251 1016249
rect 379285 1016245 379319 1016249
rect 379353 1016245 379387 1016249
rect 379421 1016245 379455 1016249
rect 379489 1016245 379523 1016249
rect 379557 1016245 379591 1016249
rect 379625 1016245 379659 1016249
rect 379693 1016245 379727 1016249
rect 379761 1016245 379795 1016249
rect 379829 1016245 379863 1016249
rect 379897 1016245 379931 1016249
rect 379965 1016245 379999 1016249
rect 380033 1016245 380067 1016249
rect 380101 1016245 380135 1016249
rect 380169 1016245 380203 1016249
rect 380237 1016245 380271 1016249
rect 380305 1016245 380339 1016249
rect 380373 1016245 380407 1016249
rect 377585 1016227 380485 1016245
rect 377653 1016223 377687 1016227
rect 377721 1016223 377755 1016227
rect 377789 1016223 377823 1016227
rect 377857 1016223 377891 1016227
rect 377925 1016223 377959 1016227
rect 377993 1016223 378027 1016227
rect 378061 1016223 378095 1016227
rect 378129 1016223 378163 1016227
rect 378197 1016223 378231 1016227
rect 378265 1016223 378299 1016227
rect 378333 1016223 378367 1016227
rect 378401 1016223 378435 1016227
rect 378469 1016223 378503 1016227
rect 378537 1016223 378571 1016227
rect 378605 1016223 378639 1016227
rect 378673 1016223 378707 1016227
rect 378741 1016223 378775 1016227
rect 378809 1016223 378843 1016227
rect 378877 1016223 378911 1016227
rect 378945 1016223 378979 1016227
rect 379013 1016223 379047 1016227
rect 379081 1016223 379115 1016227
rect 379149 1016223 379183 1016227
rect 379217 1016223 379251 1016227
rect 379285 1016223 379319 1016227
rect 379353 1016223 379387 1016227
rect 379421 1016223 379455 1016227
rect 379489 1016223 379523 1016227
rect 379557 1016223 379591 1016227
rect 379625 1016223 379659 1016227
rect 379693 1016223 379727 1016227
rect 379761 1016223 379795 1016227
rect 379829 1016223 379863 1016227
rect 379897 1016223 379931 1016227
rect 379965 1016223 379999 1016227
rect 380033 1016223 380067 1016227
rect 380101 1016223 380135 1016227
rect 380169 1016223 380203 1016227
rect 380237 1016223 380271 1016227
rect 380305 1016223 380339 1016227
rect 380373 1016223 380407 1016227
rect 380624 1016224 380648 1016248
rect 427489 1016245 427523 1016249
rect 427557 1016245 427591 1016249
rect 427625 1016245 427659 1016249
rect 427693 1016245 427727 1016249
rect 427761 1016245 427795 1016249
rect 427829 1016245 427863 1016249
rect 427897 1016245 427931 1016249
rect 427965 1016245 427999 1016249
rect 428033 1016245 428067 1016249
rect 428101 1016245 428135 1016249
rect 428169 1016245 428203 1016249
rect 428237 1016245 428271 1016249
rect 428305 1016245 428339 1016249
rect 428373 1016245 428407 1016249
rect 377143 1016203 377177 1016217
rect 377589 1016215 380481 1016223
rect 377629 1016203 380431 1016215
rect 380648 1016200 380672 1016215
rect 380716 1016204 380750 1016239
rect 427473 1016227 428485 1016245
rect 427489 1016223 427523 1016227
rect 427557 1016223 427591 1016227
rect 427625 1016223 427659 1016227
rect 427693 1016223 427727 1016227
rect 427761 1016223 427795 1016227
rect 427829 1016223 427863 1016227
rect 427897 1016223 427931 1016227
rect 427965 1016223 427999 1016227
rect 428033 1016223 428067 1016227
rect 428101 1016223 428135 1016227
rect 428169 1016223 428203 1016227
rect 428237 1016223 428271 1016227
rect 428305 1016223 428339 1016227
rect 428373 1016223 428407 1016227
rect 428624 1016224 428648 1016248
rect 374771 1014787 374899 1016187
rect 374934 1014787 375062 1016187
rect 375097 1014787 375225 1016187
rect 375260 1014787 375388 1016187
rect 375423 1014787 375551 1016187
rect 375586 1014787 375714 1016187
rect 375749 1014787 375792 1016187
rect 375885 1014787 375928 1016187
rect 376035 1014787 376163 1016187
rect 376198 1014787 376326 1016187
rect 376361 1014787 376489 1016187
rect 376524 1014787 376652 1016187
rect 376687 1014787 376815 1016187
rect 376850 1014787 376978 1016187
rect 377013 1014787 377063 1016187
rect 377119 1016169 377143 1016193
rect 377177 1016169 377201 1016193
rect 380726 1016191 380750 1016204
rect 427473 1016215 428481 1016223
rect 427473 1016203 428431 1016215
rect 428648 1016200 428672 1016215
rect 428716 1016204 428750 1016239
rect 428726 1016191 428750 1016204
rect 467015 1016131 470015 1016259
rect 470464 1016215 470566 1016239
rect 470464 1016191 470488 1016215
rect 470542 1016191 470566 1016215
rect 471947 1016191 471981 1016249
rect 472136 1016215 472170 1016249
rect 472208 1016215 472242 1016249
rect 472280 1016215 472314 1016249
rect 472352 1016215 472386 1016249
rect 472136 1016191 472160 1016215
rect 472362 1016191 472386 1016215
rect 472540 1016215 472642 1016239
rect 473770 1016228 473794 1016252
rect 473668 1016215 473692 1016218
rect 472540 1016191 472564 1016215
rect 472618 1016191 472642 1016215
rect 473746 1016204 473770 1016218
rect 473923 1016215 474025 1016239
rect 377330 1014402 377432 1015966
rect 377699 1014719 377749 1016119
rect 377856 1014719 377984 1016119
rect 378019 1014719 378147 1016119
rect 378182 1014719 378310 1016119
rect 378345 1014719 378473 1016119
rect 378508 1014719 378636 1016119
rect 378671 1014719 378799 1016119
rect 378834 1014719 378877 1016119
rect 378970 1014719 379013 1016119
rect 379120 1014719 379248 1016119
rect 379283 1014719 379411 1016119
rect 379446 1014719 379574 1016119
rect 379609 1014719 379737 1016119
rect 379772 1014719 379900 1016119
rect 379935 1014719 380063 1016119
rect 380098 1014719 380226 1016119
rect 380261 1014719 380304 1016119
rect 415015 1015201 415253 1015251
rect 426834 1014719 426877 1016119
rect 426970 1014719 427013 1016119
rect 427473 1014719 427574 1016119
rect 427609 1014719 427737 1016119
rect 427772 1014719 427900 1016119
rect 427935 1014719 428063 1016119
rect 428098 1014719 428226 1016119
rect 428261 1014719 428304 1016119
rect 467015 1015975 470015 1016103
rect 467015 1015819 470015 1015947
rect 467015 1015663 470015 1015791
rect 467015 1015507 470015 1015635
rect 467015 1015351 470015 1015479
rect 467015 1015201 470015 1015251
rect 470852 1014787 470895 1016187
rect 471002 1014787 471130 1016187
rect 471165 1014787 471293 1016187
rect 471328 1014787 471456 1016187
rect 471491 1014787 471619 1016187
rect 471654 1014787 471782 1016187
rect 471817 1014787 471860 1016187
rect 472729 1014787 472779 1016187
rect 472886 1014787 473014 1016187
rect 473049 1014787 473177 1016187
rect 473212 1014787 473340 1016187
rect 473375 1014787 473503 1016187
rect 473538 1014787 473581 1016187
rect 473644 1016170 473668 1016194
rect 473770 1016170 473794 1016194
rect 473923 1016191 473947 1016215
rect 474001 1016191 474025 1016215
rect 377364 1014378 377398 1014402
rect 467508 1014388 467678 1014694
rect 468308 1014388 468478 1014694
rect 469108 1014388 469278 1014694
rect 377364 1014300 377398 1014324
rect 374771 1012515 374899 1013915
rect 374934 1012515 375062 1013915
rect 375097 1012515 375225 1013915
rect 375260 1012515 375388 1013915
rect 375423 1012515 375551 1013915
rect 375586 1012515 375714 1013915
rect 375749 1012515 375792 1013915
rect 375885 1012515 375928 1013915
rect 376035 1012515 376163 1013915
rect 376198 1012515 376326 1013915
rect 376361 1012515 376489 1013915
rect 376524 1012515 376652 1013915
rect 376687 1012515 376815 1013915
rect 376850 1012515 376978 1013915
rect 377013 1012515 377063 1013915
rect 377330 1012736 377432 1014300
rect 377699 1012583 377749 1013983
rect 377856 1012583 377984 1013983
rect 378019 1012583 378147 1013983
rect 378182 1012583 378310 1013983
rect 378345 1012583 378473 1013983
rect 378508 1012583 378636 1013983
rect 378671 1012583 378799 1013983
rect 378834 1012583 378877 1013983
rect 378970 1012583 379013 1013983
rect 379120 1012583 379248 1013983
rect 379283 1012583 379411 1013983
rect 379446 1012583 379574 1013983
rect 379609 1012583 379737 1013983
rect 379772 1012583 379900 1013983
rect 379935 1012583 380063 1013983
rect 380098 1012583 380226 1013983
rect 380261 1012583 380304 1013983
rect 377119 1012509 377143 1012533
rect 377177 1012509 377201 1012533
rect 377653 1012517 377687 1012521
rect 377721 1012517 377755 1012521
rect 377789 1012517 377823 1012521
rect 377857 1012517 377891 1012521
rect 377925 1012517 377959 1012521
rect 377993 1012517 378027 1012521
rect 378061 1012517 378095 1012521
rect 378129 1012517 378163 1012521
rect 378197 1012517 378231 1012521
rect 378265 1012517 378299 1012521
rect 378333 1012517 378367 1012521
rect 378401 1012517 378435 1012521
rect 378469 1012517 378503 1012521
rect 378537 1012517 378571 1012521
rect 378605 1012517 378639 1012521
rect 378673 1012517 378707 1012521
rect 378741 1012517 378775 1012521
rect 378809 1012517 378843 1012521
rect 378877 1012517 378911 1012521
rect 378945 1012517 378979 1012521
rect 379013 1012517 379047 1012521
rect 379081 1012517 379115 1012521
rect 379149 1012517 379183 1012521
rect 379217 1012517 379251 1012521
rect 379285 1012517 379319 1012521
rect 379353 1012517 379387 1012521
rect 379421 1012517 379455 1012521
rect 379489 1012517 379523 1012521
rect 379557 1012517 379591 1012521
rect 379625 1012517 379659 1012521
rect 379693 1012517 379727 1012521
rect 379761 1012517 379795 1012521
rect 379829 1012517 379863 1012521
rect 379897 1012517 379931 1012521
rect 379965 1012517 379999 1012521
rect 380033 1012517 380067 1012521
rect 380101 1012517 380135 1012521
rect 380169 1012517 380203 1012521
rect 380237 1012517 380271 1012521
rect 380305 1012517 380339 1012521
rect 380373 1012517 380407 1012521
rect 377619 1012509 380451 1012517
rect 380682 1012512 380750 1012532
rect 377653 1012505 377687 1012509
rect 377721 1012505 377755 1012509
rect 377789 1012505 377823 1012509
rect 377857 1012505 377891 1012509
rect 377925 1012505 377959 1012509
rect 377993 1012505 378027 1012509
rect 378061 1012505 378095 1012509
rect 378129 1012505 378163 1012509
rect 378197 1012505 378231 1012509
rect 378265 1012505 378299 1012509
rect 378333 1012505 378367 1012509
rect 378401 1012505 378435 1012509
rect 378469 1012505 378503 1012509
rect 378537 1012505 378571 1012509
rect 378605 1012505 378639 1012509
rect 378673 1012505 378707 1012509
rect 378741 1012505 378775 1012509
rect 378809 1012505 378843 1012509
rect 378877 1012505 378911 1012509
rect 378945 1012505 378979 1012509
rect 379013 1012505 379047 1012509
rect 379081 1012505 379115 1012509
rect 379149 1012505 379183 1012509
rect 379217 1012505 379251 1012509
rect 379285 1012505 379319 1012509
rect 379353 1012505 379387 1012509
rect 379421 1012505 379455 1012509
rect 379489 1012505 379523 1012509
rect 379557 1012505 379591 1012509
rect 379625 1012505 379659 1012509
rect 379693 1012505 379727 1012509
rect 379761 1012505 379795 1012509
rect 379829 1012505 379863 1012509
rect 379897 1012505 379931 1012509
rect 379965 1012505 379999 1012509
rect 380033 1012505 380067 1012509
rect 380101 1012505 380135 1012509
rect 380169 1012505 380203 1012509
rect 380237 1012505 380271 1012509
rect 380305 1012505 380339 1012509
rect 380373 1012505 380407 1012509
rect 377143 1012485 377177 1012499
rect 377585 1012487 380485 1012505
rect 380648 1012487 380672 1012502
rect 380716 1012487 380750 1012512
rect 377629 1012485 380431 1012487
rect 377119 1012451 377143 1012475
rect 377177 1012451 377201 1012475
rect 380624 1012454 380648 1012478
rect 380726 1012463 380750 1012487
rect 412965 1012428 413015 1013028
rect 413115 1012428 413243 1013028
rect 413271 1012428 413399 1013028
rect 413427 1012428 413483 1013028
rect 413583 1012428 413711 1013028
rect 413739 1012428 413867 1013028
rect 413895 1012428 413945 1013028
rect 414025 1012428 414075 1013028
rect 414175 1012428 414225 1013028
rect 414663 1012427 414713 1013027
rect 415125 1012427 415181 1013027
rect 426834 1012583 426877 1013983
rect 426970 1012583 427013 1013983
rect 427473 1012583 427574 1013983
rect 427609 1012583 427737 1013983
rect 427772 1012583 427900 1013983
rect 427935 1012583 428063 1013983
rect 428098 1012583 428226 1013983
rect 428261 1012583 428304 1013983
rect 467508 1013888 467678 1014194
rect 468308 1013888 468478 1014194
rect 469108 1013888 469278 1014194
rect 427489 1012517 427523 1012521
rect 427557 1012517 427591 1012521
rect 427625 1012517 427659 1012521
rect 427693 1012517 427727 1012521
rect 427761 1012517 427795 1012521
rect 427829 1012517 427863 1012521
rect 427897 1012517 427931 1012521
rect 427965 1012517 427999 1012521
rect 428033 1012517 428067 1012521
rect 428101 1012517 428135 1012521
rect 428169 1012517 428203 1012521
rect 428237 1012517 428271 1012521
rect 428305 1012517 428339 1012521
rect 428373 1012517 428407 1012521
rect 427473 1012509 428451 1012517
rect 428682 1012512 428750 1012532
rect 427489 1012505 427523 1012509
rect 427557 1012505 427591 1012509
rect 427625 1012505 427659 1012509
rect 427693 1012505 427727 1012509
rect 427761 1012505 427795 1012509
rect 427829 1012505 427863 1012509
rect 427897 1012505 427931 1012509
rect 427965 1012505 427999 1012509
rect 428033 1012505 428067 1012509
rect 428101 1012505 428135 1012509
rect 428169 1012505 428203 1012509
rect 428237 1012505 428271 1012509
rect 428305 1012505 428339 1012509
rect 428373 1012505 428407 1012509
rect 427473 1012487 428485 1012505
rect 428648 1012487 428672 1012502
rect 428716 1012487 428750 1012512
rect 427473 1012485 428431 1012487
rect 428624 1012454 428648 1012478
rect 428726 1012463 428750 1012487
rect 464965 1012428 465015 1013028
rect 465115 1012428 465243 1013028
rect 465271 1012428 465399 1013028
rect 465427 1012428 465483 1013028
rect 465583 1012428 465711 1013028
rect 465739 1012428 465867 1013028
rect 465895 1012428 465945 1013028
rect 466025 1012428 466075 1013028
rect 466175 1012428 466225 1013028
rect 466663 1012427 466713 1013027
rect 466813 1012427 466941 1013027
rect 466969 1012427 467097 1013027
rect 467125 1012427 467181 1013027
rect 467281 1012427 467409 1013027
rect 467437 1012427 467565 1013027
rect 467593 1012427 467643 1013027
rect 467723 1012427 467773 1013027
rect 467873 1012427 467923 1013027
rect 468045 1012427 468095 1013027
rect 468195 1012427 468245 1013027
rect 468325 1012427 468375 1013027
rect 468475 1012427 468603 1013027
rect 468631 1012427 468759 1013027
rect 468787 1012427 468843 1013027
rect 468943 1012427 469071 1013027
rect 469099 1012427 469227 1013027
rect 469255 1012427 469305 1013027
rect 470852 1012515 470895 1013915
rect 471002 1012515 471130 1013915
rect 471165 1012515 471293 1013915
rect 471328 1012515 471456 1013915
rect 471491 1012515 471619 1013915
rect 471654 1012515 471782 1013915
rect 471817 1012515 471860 1013915
rect 470464 1012487 470566 1012511
rect 470542 1012463 470566 1012487
rect 471947 1012463 471981 1012521
rect 472136 1012487 472170 1012521
rect 472208 1012487 472242 1012521
rect 472280 1012487 472314 1012521
rect 472352 1012487 472386 1012521
rect 472729 1012515 472779 1013915
rect 472886 1012515 473014 1013915
rect 473049 1012515 473177 1013915
rect 473212 1012515 473340 1013915
rect 473375 1012515 473503 1013915
rect 473538 1012515 473581 1013915
rect 472136 1012463 472160 1012487
rect 472362 1012463 472386 1012487
rect 472540 1012487 472642 1012511
rect 473644 1012508 473668 1012532
rect 473770 1012508 473794 1012532
rect 472540 1012463 472564 1012487
rect 472618 1012463 472642 1012487
rect 473668 1012484 473692 1012487
rect 473746 1012484 473770 1012498
rect 473923 1012487 474025 1012511
rect 473770 1012450 473794 1012474
rect 473923 1012463 473947 1012487
rect 474001 1012463 474025 1012487
rect 380682 1012376 380750 1012396
rect 428682 1012376 428750 1012396
rect 377462 1012288 377486 1012312
rect 377520 1012288 377544 1012312
rect 377496 1012264 377510 1012288
rect 474201 1012047 474737 1016655
rect 570640 1016651 570674 1016675
rect 570708 1016651 570742 1016675
rect 570776 1016651 570810 1016675
rect 570844 1016651 570878 1016675
rect 570912 1016651 570946 1016675
rect 570980 1016651 571014 1016675
rect 571048 1016651 571082 1016675
rect 571116 1016651 571150 1016675
rect 571184 1016651 571218 1016675
rect 571252 1016651 571286 1016675
rect 571320 1016651 571354 1016675
rect 571388 1016651 571422 1016675
rect 571456 1016651 571490 1016675
rect 571524 1016651 571558 1016675
rect 571592 1016651 571626 1016675
rect 571660 1016651 571694 1016675
rect 571728 1016651 571762 1016675
rect 571796 1016651 571830 1016675
rect 571864 1016651 571898 1016675
rect 571932 1016651 571966 1016675
rect 572000 1016651 572034 1016675
rect 572068 1016651 572102 1016675
rect 572136 1016651 572170 1016675
rect 572204 1016651 572238 1016675
rect 572272 1016651 572306 1016675
rect 572340 1016651 572374 1016675
rect 572408 1016651 572442 1016675
rect 572476 1016651 572510 1016675
rect 572544 1016651 572578 1016675
rect 572612 1016651 572646 1016675
rect 572680 1016651 572714 1016675
rect 572748 1016651 572782 1016675
rect 572816 1016651 572850 1016675
rect 572884 1016651 572918 1016675
rect 572952 1016651 572986 1016675
rect 573020 1016651 573054 1016675
rect 573088 1016651 573122 1016675
rect 573156 1016651 573190 1016675
rect 573224 1016651 573258 1016675
rect 573292 1016651 573326 1016675
rect 573360 1016651 573394 1016675
rect 573428 1016651 573462 1016675
rect 573496 1016651 573530 1016675
rect 573564 1016651 573598 1016675
rect 573632 1016651 573666 1016675
rect 573700 1016651 573734 1016675
rect 573768 1016651 573802 1016675
rect 573836 1016651 573870 1016675
rect 573904 1016651 573938 1016675
rect 573972 1016651 574006 1016675
rect 574040 1016651 574074 1016675
rect 574108 1016651 574142 1016675
rect 574176 1016651 574210 1016675
rect 574244 1016651 574278 1016675
rect 574312 1016651 574346 1016675
rect 574380 1016651 574414 1016675
rect 574448 1016660 574482 1016675
rect 574430 1016651 574482 1016660
rect 574430 1016626 574448 1016651
rect 574464 1016626 574482 1016651
rect 574505 1016626 574506 1016651
rect 574464 1016617 574506 1016626
rect 480933 1016597 481053 1016600
rect 516733 1016597 516853 1016600
rect 532933 1016597 533053 1016600
rect 568733 1016597 568853 1016600
rect 477496 1016414 477510 1016438
rect 477462 1016390 477486 1016414
rect 477520 1016390 477544 1016414
rect 480716 1016340 480750 1016360
rect 532716 1016340 532750 1016360
rect 519015 1016287 519253 1016337
rect 571015 1016287 574015 1016337
rect 477119 1016227 477143 1016251
rect 477177 1016227 477201 1016251
rect 477653 1016245 477687 1016249
rect 477721 1016245 477755 1016249
rect 477789 1016245 477823 1016249
rect 477857 1016245 477891 1016249
rect 477925 1016245 477959 1016249
rect 477993 1016245 478027 1016249
rect 478061 1016245 478095 1016249
rect 478129 1016245 478163 1016249
rect 478197 1016245 478231 1016249
rect 478265 1016245 478299 1016249
rect 478333 1016245 478367 1016249
rect 478401 1016245 478435 1016249
rect 478469 1016245 478503 1016249
rect 478537 1016245 478571 1016249
rect 478605 1016245 478639 1016249
rect 478673 1016245 478707 1016249
rect 478741 1016245 478775 1016249
rect 478809 1016245 478843 1016249
rect 478877 1016245 478911 1016249
rect 478945 1016245 478979 1016249
rect 479013 1016245 479047 1016249
rect 479081 1016245 479115 1016249
rect 479149 1016245 479183 1016249
rect 479217 1016245 479251 1016249
rect 479285 1016245 479319 1016249
rect 479353 1016245 479387 1016249
rect 479421 1016245 479455 1016249
rect 479489 1016245 479523 1016249
rect 479557 1016245 479591 1016249
rect 479625 1016245 479659 1016249
rect 479693 1016245 479727 1016249
rect 479761 1016245 479795 1016249
rect 479829 1016245 479863 1016249
rect 479897 1016245 479931 1016249
rect 479965 1016245 479999 1016249
rect 480033 1016245 480067 1016249
rect 480101 1016245 480135 1016249
rect 480169 1016245 480203 1016249
rect 480237 1016245 480271 1016249
rect 480305 1016245 480339 1016249
rect 480373 1016245 480407 1016249
rect 477585 1016227 480485 1016245
rect 477653 1016223 477687 1016227
rect 477721 1016223 477755 1016227
rect 477789 1016223 477823 1016227
rect 477857 1016223 477891 1016227
rect 477925 1016223 477959 1016227
rect 477993 1016223 478027 1016227
rect 478061 1016223 478095 1016227
rect 478129 1016223 478163 1016227
rect 478197 1016223 478231 1016227
rect 478265 1016223 478299 1016227
rect 478333 1016223 478367 1016227
rect 478401 1016223 478435 1016227
rect 478469 1016223 478503 1016227
rect 478537 1016223 478571 1016227
rect 478605 1016223 478639 1016227
rect 478673 1016223 478707 1016227
rect 478741 1016223 478775 1016227
rect 478809 1016223 478843 1016227
rect 478877 1016223 478911 1016227
rect 478945 1016223 478979 1016227
rect 479013 1016223 479047 1016227
rect 479081 1016223 479115 1016227
rect 479149 1016223 479183 1016227
rect 479217 1016223 479251 1016227
rect 479285 1016223 479319 1016227
rect 479353 1016223 479387 1016227
rect 479421 1016223 479455 1016227
rect 479489 1016223 479523 1016227
rect 479557 1016223 479591 1016227
rect 479625 1016223 479659 1016227
rect 479693 1016223 479727 1016227
rect 479761 1016223 479795 1016227
rect 479829 1016223 479863 1016227
rect 479897 1016223 479931 1016227
rect 479965 1016223 479999 1016227
rect 480033 1016223 480067 1016227
rect 480101 1016223 480135 1016227
rect 480169 1016223 480203 1016227
rect 480237 1016223 480271 1016227
rect 480305 1016223 480339 1016227
rect 480373 1016223 480407 1016227
rect 480624 1016224 480648 1016248
rect 531489 1016245 531523 1016249
rect 531557 1016245 531591 1016249
rect 531625 1016245 531659 1016249
rect 531693 1016245 531727 1016249
rect 531761 1016245 531795 1016249
rect 531829 1016245 531863 1016249
rect 531897 1016245 531931 1016249
rect 531965 1016245 531999 1016249
rect 532033 1016245 532067 1016249
rect 532101 1016245 532135 1016249
rect 532169 1016245 532203 1016249
rect 532237 1016245 532271 1016249
rect 532305 1016245 532339 1016249
rect 532373 1016245 532407 1016249
rect 477143 1016203 477177 1016217
rect 477589 1016215 480481 1016223
rect 477629 1016203 480431 1016215
rect 480648 1016200 480672 1016215
rect 480716 1016204 480750 1016239
rect 531473 1016227 532485 1016245
rect 531489 1016223 531523 1016227
rect 531557 1016223 531591 1016227
rect 531625 1016223 531659 1016227
rect 531693 1016223 531727 1016227
rect 531761 1016223 531795 1016227
rect 531829 1016223 531863 1016227
rect 531897 1016223 531931 1016227
rect 531965 1016223 531999 1016227
rect 532033 1016223 532067 1016227
rect 532101 1016223 532135 1016227
rect 532169 1016223 532203 1016227
rect 532237 1016223 532271 1016227
rect 532305 1016223 532339 1016227
rect 532373 1016223 532407 1016227
rect 532624 1016224 532648 1016248
rect 474771 1014787 474899 1016187
rect 474934 1014787 475062 1016187
rect 475097 1014787 475225 1016187
rect 475260 1014787 475388 1016187
rect 475423 1014787 475551 1016187
rect 475586 1014787 475714 1016187
rect 475749 1014787 475792 1016187
rect 475885 1014787 475928 1016187
rect 476035 1014787 476163 1016187
rect 476198 1014787 476326 1016187
rect 476361 1014787 476489 1016187
rect 476524 1014787 476652 1016187
rect 476687 1014787 476815 1016187
rect 476850 1014787 476978 1016187
rect 477013 1014787 477063 1016187
rect 477119 1016169 477143 1016193
rect 477177 1016169 477201 1016193
rect 480726 1016191 480750 1016204
rect 531473 1016215 532481 1016223
rect 531473 1016203 532431 1016215
rect 532648 1016200 532672 1016215
rect 532716 1016204 532750 1016239
rect 532726 1016191 532750 1016204
rect 571015 1016131 574015 1016259
rect 574464 1016215 574566 1016239
rect 574464 1016191 574488 1016215
rect 574542 1016191 574566 1016215
rect 575947 1016191 575981 1016249
rect 576136 1016215 576170 1016249
rect 576208 1016215 576242 1016249
rect 576280 1016215 576314 1016249
rect 576352 1016215 576386 1016249
rect 576136 1016191 576160 1016215
rect 576362 1016191 576386 1016215
rect 576540 1016215 576642 1016239
rect 577770 1016228 577794 1016252
rect 577668 1016215 577692 1016218
rect 576540 1016191 576564 1016215
rect 576618 1016191 576642 1016215
rect 577746 1016204 577770 1016218
rect 577923 1016215 578025 1016239
rect 477330 1014402 477432 1015966
rect 477699 1014719 477749 1016119
rect 477856 1014719 477984 1016119
rect 478019 1014719 478147 1016119
rect 478182 1014719 478310 1016119
rect 478345 1014719 478473 1016119
rect 478508 1014719 478636 1016119
rect 478671 1014719 478799 1016119
rect 478834 1014719 478877 1016119
rect 478970 1014719 479013 1016119
rect 479120 1014719 479248 1016119
rect 479283 1014719 479411 1016119
rect 479446 1014719 479574 1016119
rect 479609 1014719 479737 1016119
rect 479772 1014719 479900 1016119
rect 479935 1014719 480063 1016119
rect 480098 1014719 480226 1016119
rect 480261 1014719 480304 1016119
rect 519015 1015201 519253 1015251
rect 530834 1014719 530877 1016119
rect 530970 1014719 531013 1016119
rect 531473 1014719 531574 1016119
rect 531609 1014719 531737 1016119
rect 531772 1014719 531900 1016119
rect 531935 1014719 532063 1016119
rect 532098 1014719 532226 1016119
rect 532261 1014719 532304 1016119
rect 571015 1015975 574015 1016103
rect 571015 1015819 574015 1015947
rect 571015 1015663 574015 1015791
rect 571015 1015507 574015 1015635
rect 571015 1015351 574015 1015479
rect 571015 1015201 574015 1015251
rect 574852 1014787 574895 1016187
rect 575002 1014787 575130 1016187
rect 575165 1014787 575293 1016187
rect 575328 1014787 575456 1016187
rect 575491 1014787 575619 1016187
rect 575654 1014787 575782 1016187
rect 575817 1014787 575860 1016187
rect 576729 1014787 576779 1016187
rect 576886 1014787 577014 1016187
rect 577049 1014787 577177 1016187
rect 577212 1014787 577340 1016187
rect 577375 1014787 577503 1016187
rect 577538 1014787 577581 1016187
rect 577644 1016170 577668 1016194
rect 577770 1016170 577794 1016194
rect 577923 1016191 577947 1016215
rect 578001 1016191 578025 1016215
rect 477364 1014378 477398 1014402
rect 571508 1014388 571678 1014694
rect 572308 1014388 572478 1014694
rect 573108 1014388 573278 1014694
rect 477364 1014300 477398 1014324
rect 474771 1012515 474899 1013915
rect 474934 1012515 475062 1013915
rect 475097 1012515 475225 1013915
rect 475260 1012515 475388 1013915
rect 475423 1012515 475551 1013915
rect 475586 1012515 475714 1013915
rect 475749 1012515 475792 1013915
rect 475885 1012515 475928 1013915
rect 476035 1012515 476163 1013915
rect 476198 1012515 476326 1013915
rect 476361 1012515 476489 1013915
rect 476524 1012515 476652 1013915
rect 476687 1012515 476815 1013915
rect 476850 1012515 476978 1013915
rect 477013 1012515 477063 1013915
rect 477330 1012736 477432 1014300
rect 477699 1012583 477749 1013983
rect 477856 1012583 477984 1013983
rect 478019 1012583 478147 1013983
rect 478182 1012583 478310 1013983
rect 478345 1012583 478473 1013983
rect 478508 1012583 478636 1013983
rect 478671 1012583 478799 1013983
rect 478834 1012583 478877 1013983
rect 478970 1012583 479013 1013983
rect 479120 1012583 479248 1013983
rect 479283 1012583 479411 1013983
rect 479446 1012583 479574 1013983
rect 479609 1012583 479737 1013983
rect 479772 1012583 479900 1013983
rect 479935 1012583 480063 1013983
rect 480098 1012583 480226 1013983
rect 480261 1012583 480304 1013983
rect 477119 1012509 477143 1012533
rect 477177 1012509 477201 1012533
rect 477653 1012517 477687 1012521
rect 477721 1012517 477755 1012521
rect 477789 1012517 477823 1012521
rect 477857 1012517 477891 1012521
rect 477925 1012517 477959 1012521
rect 477993 1012517 478027 1012521
rect 478061 1012517 478095 1012521
rect 478129 1012517 478163 1012521
rect 478197 1012517 478231 1012521
rect 478265 1012517 478299 1012521
rect 478333 1012517 478367 1012521
rect 478401 1012517 478435 1012521
rect 478469 1012517 478503 1012521
rect 478537 1012517 478571 1012521
rect 478605 1012517 478639 1012521
rect 478673 1012517 478707 1012521
rect 478741 1012517 478775 1012521
rect 478809 1012517 478843 1012521
rect 478877 1012517 478911 1012521
rect 478945 1012517 478979 1012521
rect 479013 1012517 479047 1012521
rect 479081 1012517 479115 1012521
rect 479149 1012517 479183 1012521
rect 479217 1012517 479251 1012521
rect 479285 1012517 479319 1012521
rect 479353 1012517 479387 1012521
rect 479421 1012517 479455 1012521
rect 479489 1012517 479523 1012521
rect 479557 1012517 479591 1012521
rect 479625 1012517 479659 1012521
rect 479693 1012517 479727 1012521
rect 479761 1012517 479795 1012521
rect 479829 1012517 479863 1012521
rect 479897 1012517 479931 1012521
rect 479965 1012517 479999 1012521
rect 480033 1012517 480067 1012521
rect 480101 1012517 480135 1012521
rect 480169 1012517 480203 1012521
rect 480237 1012517 480271 1012521
rect 480305 1012517 480339 1012521
rect 480373 1012517 480407 1012521
rect 477619 1012509 480451 1012517
rect 480682 1012512 480750 1012532
rect 477653 1012505 477687 1012509
rect 477721 1012505 477755 1012509
rect 477789 1012505 477823 1012509
rect 477857 1012505 477891 1012509
rect 477925 1012505 477959 1012509
rect 477993 1012505 478027 1012509
rect 478061 1012505 478095 1012509
rect 478129 1012505 478163 1012509
rect 478197 1012505 478231 1012509
rect 478265 1012505 478299 1012509
rect 478333 1012505 478367 1012509
rect 478401 1012505 478435 1012509
rect 478469 1012505 478503 1012509
rect 478537 1012505 478571 1012509
rect 478605 1012505 478639 1012509
rect 478673 1012505 478707 1012509
rect 478741 1012505 478775 1012509
rect 478809 1012505 478843 1012509
rect 478877 1012505 478911 1012509
rect 478945 1012505 478979 1012509
rect 479013 1012505 479047 1012509
rect 479081 1012505 479115 1012509
rect 479149 1012505 479183 1012509
rect 479217 1012505 479251 1012509
rect 479285 1012505 479319 1012509
rect 479353 1012505 479387 1012509
rect 479421 1012505 479455 1012509
rect 479489 1012505 479523 1012509
rect 479557 1012505 479591 1012509
rect 479625 1012505 479659 1012509
rect 479693 1012505 479727 1012509
rect 479761 1012505 479795 1012509
rect 479829 1012505 479863 1012509
rect 479897 1012505 479931 1012509
rect 479965 1012505 479999 1012509
rect 480033 1012505 480067 1012509
rect 480101 1012505 480135 1012509
rect 480169 1012505 480203 1012509
rect 480237 1012505 480271 1012509
rect 480305 1012505 480339 1012509
rect 480373 1012505 480407 1012509
rect 477143 1012485 477177 1012499
rect 477585 1012487 480485 1012505
rect 480648 1012487 480672 1012502
rect 480716 1012487 480750 1012512
rect 477629 1012485 480431 1012487
rect 477119 1012451 477143 1012475
rect 477177 1012451 477201 1012475
rect 480624 1012454 480648 1012478
rect 480726 1012463 480750 1012487
rect 516965 1012428 517015 1013028
rect 517115 1012428 517243 1013028
rect 517271 1012428 517399 1013028
rect 517427 1012428 517483 1013028
rect 517583 1012428 517711 1013028
rect 517739 1012428 517867 1013028
rect 517895 1012428 517945 1013028
rect 518025 1012428 518075 1013028
rect 518175 1012428 518225 1013028
rect 518663 1012427 518713 1013027
rect 519125 1012427 519181 1013027
rect 530834 1012583 530877 1013983
rect 530970 1012583 531013 1013983
rect 531473 1012583 531574 1013983
rect 531609 1012583 531737 1013983
rect 531772 1012583 531900 1013983
rect 531935 1012583 532063 1013983
rect 532098 1012583 532226 1013983
rect 532261 1012583 532304 1013983
rect 571508 1013888 571678 1014194
rect 572308 1013888 572478 1014194
rect 573108 1013888 573278 1014194
rect 531489 1012517 531523 1012521
rect 531557 1012517 531591 1012521
rect 531625 1012517 531659 1012521
rect 531693 1012517 531727 1012521
rect 531761 1012517 531795 1012521
rect 531829 1012517 531863 1012521
rect 531897 1012517 531931 1012521
rect 531965 1012517 531999 1012521
rect 532033 1012517 532067 1012521
rect 532101 1012517 532135 1012521
rect 532169 1012517 532203 1012521
rect 532237 1012517 532271 1012521
rect 532305 1012517 532339 1012521
rect 532373 1012517 532407 1012521
rect 531473 1012509 532451 1012517
rect 532682 1012512 532750 1012532
rect 531489 1012505 531523 1012509
rect 531557 1012505 531591 1012509
rect 531625 1012505 531659 1012509
rect 531693 1012505 531727 1012509
rect 531761 1012505 531795 1012509
rect 531829 1012505 531863 1012509
rect 531897 1012505 531931 1012509
rect 531965 1012505 531999 1012509
rect 532033 1012505 532067 1012509
rect 532101 1012505 532135 1012509
rect 532169 1012505 532203 1012509
rect 532237 1012505 532271 1012509
rect 532305 1012505 532339 1012509
rect 532373 1012505 532407 1012509
rect 531473 1012487 532485 1012505
rect 532648 1012487 532672 1012502
rect 532716 1012487 532750 1012512
rect 531473 1012485 532431 1012487
rect 532624 1012454 532648 1012478
rect 532726 1012463 532750 1012487
rect 568965 1012428 569015 1013028
rect 569115 1012428 569243 1013028
rect 569271 1012428 569399 1013028
rect 569427 1012428 569483 1013028
rect 569583 1012428 569711 1013028
rect 569739 1012428 569867 1013028
rect 569895 1012428 569945 1013028
rect 570025 1012428 570075 1013028
rect 570175 1012428 570225 1013028
rect 570663 1012427 570713 1013027
rect 570813 1012427 570941 1013027
rect 570969 1012427 571097 1013027
rect 571125 1012427 571181 1013027
rect 571281 1012427 571409 1013027
rect 571437 1012427 571565 1013027
rect 571593 1012427 571643 1013027
rect 571723 1012427 571773 1013027
rect 571873 1012427 571923 1013027
rect 572045 1012427 572095 1013027
rect 572195 1012427 572245 1013027
rect 572325 1012427 572375 1013027
rect 572475 1012427 572603 1013027
rect 572631 1012427 572759 1013027
rect 572787 1012427 572843 1013027
rect 572943 1012427 573071 1013027
rect 573099 1012427 573227 1013027
rect 573255 1012427 573305 1013027
rect 574852 1012515 574895 1013915
rect 575002 1012515 575130 1013915
rect 575165 1012515 575293 1013915
rect 575328 1012515 575456 1013915
rect 575491 1012515 575619 1013915
rect 575654 1012515 575782 1013915
rect 575817 1012515 575860 1013915
rect 574464 1012487 574566 1012511
rect 574542 1012463 574566 1012487
rect 575947 1012463 575981 1012521
rect 576136 1012487 576170 1012521
rect 576208 1012487 576242 1012521
rect 576280 1012487 576314 1012521
rect 576352 1012487 576386 1012521
rect 576729 1012515 576779 1013915
rect 576886 1012515 577014 1013915
rect 577049 1012515 577177 1013915
rect 577212 1012515 577340 1013915
rect 577375 1012515 577503 1013915
rect 577538 1012515 577581 1013915
rect 576136 1012463 576160 1012487
rect 576362 1012463 576386 1012487
rect 576540 1012487 576642 1012511
rect 577644 1012508 577668 1012532
rect 577770 1012508 577794 1012532
rect 576540 1012463 576564 1012487
rect 576618 1012463 576642 1012487
rect 577668 1012484 577692 1012487
rect 577746 1012484 577770 1012498
rect 577923 1012487 578025 1012511
rect 577770 1012450 577794 1012474
rect 577923 1012463 577947 1012487
rect 578001 1012463 578025 1012487
rect 480682 1012376 480750 1012396
rect 532682 1012376 532750 1012396
rect 477462 1012288 477486 1012312
rect 477520 1012288 477544 1012312
rect 477496 1012264 477510 1012288
rect 578201 1012047 578737 1016655
rect 584933 1016597 585053 1016600
rect 581496 1016414 581510 1016438
rect 581462 1016390 581486 1016414
rect 581520 1016390 581544 1016414
rect 584716 1016340 584750 1016360
rect 581119 1016227 581143 1016251
rect 581177 1016227 581201 1016251
rect 581653 1016245 581687 1016249
rect 581721 1016245 581755 1016249
rect 581789 1016245 581823 1016249
rect 581857 1016245 581891 1016249
rect 581925 1016245 581959 1016249
rect 581993 1016245 582027 1016249
rect 582061 1016245 582095 1016249
rect 582129 1016245 582163 1016249
rect 582197 1016245 582231 1016249
rect 582265 1016245 582299 1016249
rect 582333 1016245 582367 1016249
rect 582401 1016245 582435 1016249
rect 582469 1016245 582503 1016249
rect 582537 1016245 582571 1016249
rect 582605 1016245 582639 1016249
rect 582673 1016245 582707 1016249
rect 582741 1016245 582775 1016249
rect 582809 1016245 582843 1016249
rect 582877 1016245 582911 1016249
rect 582945 1016245 582979 1016249
rect 583013 1016245 583047 1016249
rect 583081 1016245 583115 1016249
rect 583149 1016245 583183 1016249
rect 583217 1016245 583251 1016249
rect 583285 1016245 583319 1016249
rect 583353 1016245 583387 1016249
rect 583421 1016245 583455 1016249
rect 583489 1016245 583523 1016249
rect 583557 1016245 583591 1016249
rect 583625 1016245 583659 1016249
rect 583693 1016245 583727 1016249
rect 583761 1016245 583795 1016249
rect 583829 1016245 583863 1016249
rect 583897 1016245 583931 1016249
rect 583965 1016245 583999 1016249
rect 584033 1016245 584067 1016249
rect 584101 1016245 584135 1016249
rect 584169 1016245 584203 1016249
rect 584237 1016245 584271 1016249
rect 584305 1016245 584339 1016249
rect 584373 1016245 584407 1016249
rect 581585 1016227 584485 1016245
rect 581653 1016223 581687 1016227
rect 581721 1016223 581755 1016227
rect 581789 1016223 581823 1016227
rect 581857 1016223 581891 1016227
rect 581925 1016223 581959 1016227
rect 581993 1016223 582027 1016227
rect 582061 1016223 582095 1016227
rect 582129 1016223 582163 1016227
rect 582197 1016223 582231 1016227
rect 582265 1016223 582299 1016227
rect 582333 1016223 582367 1016227
rect 582401 1016223 582435 1016227
rect 582469 1016223 582503 1016227
rect 582537 1016223 582571 1016227
rect 582605 1016223 582639 1016227
rect 582673 1016223 582707 1016227
rect 582741 1016223 582775 1016227
rect 582809 1016223 582843 1016227
rect 582877 1016223 582911 1016227
rect 582945 1016223 582979 1016227
rect 583013 1016223 583047 1016227
rect 583081 1016223 583115 1016227
rect 583149 1016223 583183 1016227
rect 583217 1016223 583251 1016227
rect 583285 1016223 583319 1016227
rect 583353 1016223 583387 1016227
rect 583421 1016223 583455 1016227
rect 583489 1016223 583523 1016227
rect 583557 1016223 583591 1016227
rect 583625 1016223 583659 1016227
rect 583693 1016223 583727 1016227
rect 583761 1016223 583795 1016227
rect 583829 1016223 583863 1016227
rect 583897 1016223 583931 1016227
rect 583965 1016223 583999 1016227
rect 584033 1016223 584067 1016227
rect 584101 1016223 584135 1016227
rect 584169 1016223 584203 1016227
rect 584237 1016223 584271 1016227
rect 584305 1016223 584339 1016227
rect 584373 1016223 584407 1016227
rect 584624 1016224 584648 1016248
rect 581143 1016203 581177 1016217
rect 581589 1016215 584481 1016223
rect 581629 1016203 584431 1016215
rect 584648 1016200 584672 1016215
rect 584716 1016204 584750 1016239
rect 578771 1014787 578899 1016187
rect 578934 1014787 579062 1016187
rect 579097 1014787 579225 1016187
rect 579260 1014787 579388 1016187
rect 579423 1014787 579551 1016187
rect 579586 1014787 579714 1016187
rect 579749 1014787 579792 1016187
rect 579885 1014787 579928 1016187
rect 580035 1014787 580163 1016187
rect 580198 1014787 580326 1016187
rect 580361 1014787 580489 1016187
rect 580524 1014787 580652 1016187
rect 580687 1014787 580815 1016187
rect 580850 1014787 580978 1016187
rect 581013 1014787 581063 1016187
rect 581119 1016169 581143 1016193
rect 581177 1016169 581201 1016193
rect 584726 1016191 584750 1016204
rect 581330 1014402 581432 1015966
rect 581699 1014719 581749 1016119
rect 581856 1014719 581984 1016119
rect 582019 1014719 582147 1016119
rect 582182 1014719 582310 1016119
rect 582345 1014719 582473 1016119
rect 582508 1014719 582636 1016119
rect 582671 1014719 582799 1016119
rect 582834 1014719 582877 1016119
rect 582970 1014719 583013 1016119
rect 583120 1014719 583248 1016119
rect 583283 1014719 583411 1016119
rect 583446 1014719 583574 1016119
rect 583609 1014719 583737 1016119
rect 583772 1014719 583900 1016119
rect 583935 1014719 584063 1016119
rect 584098 1014719 584226 1016119
rect 584261 1014719 584304 1016119
rect 581364 1014378 581398 1014402
rect 581364 1014300 581398 1014324
rect 578771 1012515 578899 1013915
rect 578934 1012515 579062 1013915
rect 579097 1012515 579225 1013915
rect 579260 1012515 579388 1013915
rect 579423 1012515 579551 1013915
rect 579586 1012515 579714 1013915
rect 579749 1012515 579792 1013915
rect 579885 1012515 579928 1013915
rect 580035 1012515 580163 1013915
rect 580198 1012515 580326 1013915
rect 580361 1012515 580489 1013915
rect 580524 1012515 580652 1013915
rect 580687 1012515 580815 1013915
rect 580850 1012515 580978 1013915
rect 581013 1012515 581063 1013915
rect 581330 1012736 581432 1014300
rect 581699 1012583 581749 1013983
rect 581856 1012583 581984 1013983
rect 582019 1012583 582147 1013983
rect 582182 1012583 582310 1013983
rect 582345 1012583 582473 1013983
rect 582508 1012583 582636 1013983
rect 582671 1012583 582799 1013983
rect 582834 1012583 582877 1013983
rect 582970 1012583 583013 1013983
rect 583120 1012583 583248 1013983
rect 583283 1012583 583411 1013983
rect 583446 1012583 583574 1013983
rect 583609 1012583 583737 1013983
rect 583772 1012583 583900 1013983
rect 583935 1012583 584063 1013983
rect 584098 1012583 584226 1013983
rect 584261 1012583 584304 1013983
rect 581119 1012509 581143 1012533
rect 581177 1012509 581201 1012533
rect 581653 1012517 581687 1012521
rect 581721 1012517 581755 1012521
rect 581789 1012517 581823 1012521
rect 581857 1012517 581891 1012521
rect 581925 1012517 581959 1012521
rect 581993 1012517 582027 1012521
rect 582061 1012517 582095 1012521
rect 582129 1012517 582163 1012521
rect 582197 1012517 582231 1012521
rect 582265 1012517 582299 1012521
rect 582333 1012517 582367 1012521
rect 582401 1012517 582435 1012521
rect 582469 1012517 582503 1012521
rect 582537 1012517 582571 1012521
rect 582605 1012517 582639 1012521
rect 582673 1012517 582707 1012521
rect 582741 1012517 582775 1012521
rect 582809 1012517 582843 1012521
rect 582877 1012517 582911 1012521
rect 582945 1012517 582979 1012521
rect 583013 1012517 583047 1012521
rect 583081 1012517 583115 1012521
rect 583149 1012517 583183 1012521
rect 583217 1012517 583251 1012521
rect 583285 1012517 583319 1012521
rect 583353 1012517 583387 1012521
rect 583421 1012517 583455 1012521
rect 583489 1012517 583523 1012521
rect 583557 1012517 583591 1012521
rect 583625 1012517 583659 1012521
rect 583693 1012517 583727 1012521
rect 583761 1012517 583795 1012521
rect 583829 1012517 583863 1012521
rect 583897 1012517 583931 1012521
rect 583965 1012517 583999 1012521
rect 584033 1012517 584067 1012521
rect 584101 1012517 584135 1012521
rect 584169 1012517 584203 1012521
rect 584237 1012517 584271 1012521
rect 584305 1012517 584339 1012521
rect 584373 1012517 584407 1012521
rect 581619 1012509 584451 1012517
rect 584682 1012512 584750 1012532
rect 581653 1012505 581687 1012509
rect 581721 1012505 581755 1012509
rect 581789 1012505 581823 1012509
rect 581857 1012505 581891 1012509
rect 581925 1012505 581959 1012509
rect 581993 1012505 582027 1012509
rect 582061 1012505 582095 1012509
rect 582129 1012505 582163 1012509
rect 582197 1012505 582231 1012509
rect 582265 1012505 582299 1012509
rect 582333 1012505 582367 1012509
rect 582401 1012505 582435 1012509
rect 582469 1012505 582503 1012509
rect 582537 1012505 582571 1012509
rect 582605 1012505 582639 1012509
rect 582673 1012505 582707 1012509
rect 582741 1012505 582775 1012509
rect 582809 1012505 582843 1012509
rect 582877 1012505 582911 1012509
rect 582945 1012505 582979 1012509
rect 583013 1012505 583047 1012509
rect 583081 1012505 583115 1012509
rect 583149 1012505 583183 1012509
rect 583217 1012505 583251 1012509
rect 583285 1012505 583319 1012509
rect 583353 1012505 583387 1012509
rect 583421 1012505 583455 1012509
rect 583489 1012505 583523 1012509
rect 583557 1012505 583591 1012509
rect 583625 1012505 583659 1012509
rect 583693 1012505 583727 1012509
rect 583761 1012505 583795 1012509
rect 583829 1012505 583863 1012509
rect 583897 1012505 583931 1012509
rect 583965 1012505 583999 1012509
rect 584033 1012505 584067 1012509
rect 584101 1012505 584135 1012509
rect 584169 1012505 584203 1012509
rect 584237 1012505 584271 1012509
rect 584305 1012505 584339 1012509
rect 584373 1012505 584407 1012509
rect 581143 1012485 581177 1012499
rect 581585 1012487 584485 1012505
rect 584648 1012487 584672 1012502
rect 584716 1012487 584750 1012512
rect 581629 1012485 584431 1012487
rect 581119 1012451 581143 1012475
rect 581177 1012451 581201 1012475
rect 584624 1012454 584648 1012478
rect 584726 1012463 584750 1012487
rect 584682 1012376 584750 1012396
rect 581462 1012288 581486 1012312
rect 581520 1012288 581544 1012312
rect 581496 1012264 581510 1012288
rect 63361 1010910 63411 1011110
rect 63511 1010910 63567 1011110
rect 63667 1010910 63717 1011110
rect 64067 1010910 64117 1011110
rect 64217 1010910 64273 1011110
rect 64373 1010910 64423 1011110
rect 64487 1010910 64498 1011110
rect 71351 1010664 71401 1011664
rect 71501 1010664 71557 1011664
rect 71657 1010664 71713 1011664
rect 71813 1010664 71869 1011664
rect 71969 1011207 72019 1011664
rect 72433 1011207 72483 1011664
rect 71969 1011123 72022 1011207
rect 72430 1011123 72483 1011207
rect 71969 1010874 72019 1011123
rect 72433 1010874 72483 1011123
rect 71969 1010790 72022 1010874
rect 72430 1010790 72483 1010874
rect 71969 1010664 72019 1010790
rect 72433 1010664 72483 1010790
rect 72583 1010664 72639 1011664
rect 72739 1010664 72795 1011664
rect 72895 1010664 72951 1011664
rect 73051 1010664 73101 1011664
rect 75286 1011275 75336 1011875
rect 75436 1011275 75486 1011875
rect 75558 1011275 75608 1011875
rect 75708 1011275 75758 1011875
rect 75834 1011275 75884 1011875
rect 75984 1011275 76034 1011875
rect 76106 1011275 76156 1011875
rect 76256 1011275 76306 1011875
rect 123286 1011275 123336 1011875
rect 123436 1011275 123486 1011875
rect 123558 1011275 123608 1011875
rect 123708 1011275 123758 1011875
rect 123834 1011275 123884 1011875
rect 123984 1011275 124034 1011875
rect 124106 1011275 124156 1011875
rect 124256 1011275 124306 1011875
rect 74242 1010952 74548 1011122
rect 163361 1010910 163411 1011110
rect 163511 1010910 163567 1011110
rect 163667 1010910 163717 1011110
rect 164067 1010910 164117 1011110
rect 164217 1010910 164273 1011110
rect 164373 1010910 164423 1011110
rect 164487 1010910 164498 1011110
rect 171351 1010664 171401 1011664
rect 171501 1010664 171557 1011664
rect 171657 1010664 171713 1011664
rect 171813 1010664 171869 1011664
rect 171969 1011207 172019 1011664
rect 172433 1011207 172483 1011664
rect 171969 1011123 172022 1011207
rect 172430 1011123 172483 1011207
rect 171969 1010874 172019 1011123
rect 172433 1010874 172483 1011123
rect 171969 1010790 172022 1010874
rect 172430 1010790 172483 1010874
rect 171969 1010664 172019 1010790
rect 172433 1010664 172483 1010790
rect 172583 1010664 172639 1011664
rect 172739 1010664 172795 1011664
rect 172895 1010664 172951 1011664
rect 173051 1010664 173101 1011664
rect 175286 1011275 175336 1011875
rect 175436 1011275 175486 1011875
rect 175558 1011275 175608 1011875
rect 175708 1011275 175758 1011875
rect 175834 1011275 175884 1011875
rect 175984 1011275 176034 1011875
rect 176106 1011275 176156 1011875
rect 176256 1011275 176306 1011875
rect 227286 1011275 227336 1011875
rect 227436 1011275 227486 1011875
rect 227558 1011275 227608 1011875
rect 227708 1011275 227758 1011875
rect 227834 1011275 227884 1011875
rect 227984 1011275 228034 1011875
rect 228106 1011275 228156 1011875
rect 228256 1011275 228306 1011875
rect 275286 1011275 275336 1011875
rect 275436 1011275 275486 1011875
rect 275558 1011275 275608 1011875
rect 275708 1011275 275758 1011875
rect 275834 1011275 275884 1011875
rect 275984 1011275 276034 1011875
rect 276106 1011275 276156 1011875
rect 276256 1011275 276306 1011875
rect 327286 1011275 327336 1011875
rect 327436 1011275 327486 1011875
rect 327558 1011275 327608 1011875
rect 327708 1011275 327758 1011875
rect 327834 1011275 327884 1011875
rect 327984 1011275 328034 1011875
rect 328106 1011275 328156 1011875
rect 328256 1011275 328306 1011875
rect 174242 1010952 174548 1011122
rect 367361 1010910 367411 1011110
rect 367511 1010910 367567 1011110
rect 367667 1010910 367717 1011110
rect 368067 1010910 368117 1011110
rect 368217 1010910 368273 1011110
rect 368373 1010910 368423 1011110
rect 368487 1010910 368498 1011110
rect 375351 1010664 375401 1011664
rect 375501 1010664 375557 1011664
rect 375657 1010664 375713 1011664
rect 375813 1010664 375869 1011664
rect 375969 1011207 376019 1011664
rect 376433 1011207 376483 1011664
rect 375969 1011123 376022 1011207
rect 376430 1011123 376483 1011207
rect 375969 1010874 376019 1011123
rect 376433 1010874 376483 1011123
rect 375969 1010790 376022 1010874
rect 376430 1010790 376483 1010874
rect 375969 1010664 376019 1010790
rect 376433 1010664 376483 1010790
rect 376583 1010664 376639 1011664
rect 376739 1010664 376795 1011664
rect 376895 1010664 376951 1011664
rect 377051 1010664 377101 1011664
rect 379286 1011275 379336 1011875
rect 379436 1011275 379486 1011875
rect 379558 1011275 379608 1011875
rect 379708 1011275 379758 1011875
rect 379834 1011275 379884 1011875
rect 379984 1011275 380034 1011875
rect 380106 1011275 380156 1011875
rect 380256 1011275 380306 1011875
rect 427286 1011275 427336 1011875
rect 427436 1011275 427486 1011875
rect 427558 1011275 427608 1011875
rect 427708 1011275 427758 1011875
rect 427834 1011275 427884 1011875
rect 427984 1011275 428034 1011875
rect 428106 1011275 428156 1011875
rect 428256 1011275 428306 1011875
rect 378242 1010952 378548 1011122
rect 467361 1010910 467411 1011110
rect 467511 1010910 467567 1011110
rect 467667 1010910 467717 1011110
rect 468067 1010910 468117 1011110
rect 468217 1010910 468273 1011110
rect 468373 1010910 468423 1011110
rect 468487 1010910 468498 1011110
rect 475351 1010664 475401 1011664
rect 475501 1010664 475557 1011664
rect 475657 1010664 475713 1011664
rect 475813 1010664 475869 1011664
rect 475969 1011207 476019 1011664
rect 476433 1011207 476483 1011664
rect 475969 1011123 476022 1011207
rect 476430 1011123 476483 1011207
rect 475969 1010874 476019 1011123
rect 476433 1010874 476483 1011123
rect 475969 1010790 476022 1010874
rect 476430 1010790 476483 1010874
rect 475969 1010664 476019 1010790
rect 476433 1010664 476483 1010790
rect 476583 1010664 476639 1011664
rect 476739 1010664 476795 1011664
rect 476895 1010664 476951 1011664
rect 477051 1010664 477101 1011664
rect 479286 1011275 479336 1011875
rect 479436 1011275 479486 1011875
rect 479558 1011275 479608 1011875
rect 479708 1011275 479758 1011875
rect 479834 1011275 479884 1011875
rect 479984 1011275 480034 1011875
rect 480106 1011275 480156 1011875
rect 480256 1011275 480306 1011875
rect 531286 1011275 531336 1011875
rect 531436 1011275 531486 1011875
rect 531558 1011275 531608 1011875
rect 531708 1011275 531758 1011875
rect 531834 1011275 531884 1011875
rect 531984 1011275 532034 1011875
rect 532106 1011275 532156 1011875
rect 532256 1011275 532306 1011875
rect 478242 1010952 478548 1011122
rect 571361 1010910 571411 1011110
rect 571511 1010910 571567 1011110
rect 571667 1010910 571717 1011110
rect 572067 1010910 572117 1011110
rect 572217 1010910 572273 1011110
rect 572373 1010910 572423 1011110
rect 572487 1010910 572498 1011110
rect 579351 1010664 579401 1011664
rect 579501 1010664 579557 1011664
rect 579657 1010664 579713 1011664
rect 579813 1010664 579869 1011664
rect 579969 1011207 580019 1011664
rect 580433 1011207 580483 1011664
rect 579969 1011123 580022 1011207
rect 580430 1011123 580483 1011207
rect 579969 1010874 580019 1011123
rect 580433 1010874 580483 1011123
rect 579969 1010790 580022 1010874
rect 580430 1010790 580483 1010874
rect 579969 1010664 580019 1010790
rect 580433 1010664 580483 1010790
rect 580583 1010664 580639 1011664
rect 580739 1010664 580795 1011664
rect 580895 1010664 580951 1011664
rect 581051 1010664 581101 1011664
rect 583286 1011275 583336 1011875
rect 583436 1011275 583486 1011875
rect 583558 1011275 583608 1011875
rect 583708 1011275 583758 1011875
rect 583834 1011275 583884 1011875
rect 583984 1011275 584034 1011875
rect 584106 1011275 584156 1011875
rect 584256 1011275 584306 1011875
rect 582242 1010952 582548 1011122
rect 71500 1010326 71550 1010442
rect 71497 1010242 71550 1010326
rect 71670 1010242 71798 1010442
rect 71846 1010242 71902 1010442
rect 72022 1010242 72150 1010442
rect 72198 1010242 72254 1010442
rect 72374 1010242 72502 1010442
rect 72550 1010242 72606 1010442
rect 72726 1010242 72854 1010442
rect 72902 1010326 72952 1010442
rect 75363 1010388 76363 1010438
rect 123363 1010388 124363 1010438
rect 72902 1010242 72955 1010326
rect 71505 1010238 71539 1010242
rect 72913 1010238 72947 1010242
rect 75363 1010232 76363 1010360
rect 123473 1010232 124363 1010360
rect 171500 1010326 171550 1010442
rect 171497 1010242 171550 1010326
rect 171670 1010242 171798 1010442
rect 171846 1010242 171902 1010442
rect 172022 1010242 172150 1010442
rect 172198 1010242 172254 1010442
rect 172374 1010242 172502 1010442
rect 172550 1010242 172606 1010442
rect 172726 1010242 172854 1010442
rect 172902 1010326 172952 1010442
rect 175363 1010388 176363 1010438
rect 227363 1010388 228363 1010438
rect 275363 1010388 276363 1010438
rect 327363 1010388 328363 1010438
rect 172902 1010242 172955 1010326
rect 171505 1010238 171539 1010242
rect 172913 1010238 172947 1010242
rect 175363 1010232 176363 1010360
rect 227473 1010232 228363 1010360
rect 275473 1010232 276363 1010360
rect 327473 1010232 328363 1010360
rect 375500 1010326 375550 1010442
rect 375497 1010242 375550 1010326
rect 375670 1010242 375798 1010442
rect 375846 1010242 375902 1010442
rect 376022 1010242 376150 1010442
rect 376198 1010242 376254 1010442
rect 376374 1010242 376502 1010442
rect 376550 1010242 376606 1010442
rect 376726 1010242 376854 1010442
rect 376902 1010326 376952 1010442
rect 379363 1010388 380363 1010438
rect 427363 1010388 428363 1010438
rect 376902 1010242 376955 1010326
rect 375505 1010238 375539 1010242
rect 376913 1010238 376947 1010242
rect 379363 1010232 380363 1010360
rect 427473 1010232 428363 1010360
rect 475500 1010326 475550 1010442
rect 475497 1010242 475550 1010326
rect 475670 1010242 475798 1010442
rect 475846 1010242 475902 1010442
rect 476022 1010242 476150 1010442
rect 476198 1010242 476254 1010442
rect 476374 1010242 476502 1010442
rect 476550 1010242 476606 1010442
rect 476726 1010242 476854 1010442
rect 476902 1010326 476952 1010442
rect 479363 1010388 480363 1010438
rect 531363 1010388 532363 1010438
rect 476902 1010242 476955 1010326
rect 475505 1010238 475539 1010242
rect 476913 1010238 476947 1010242
rect 479363 1010232 480363 1010360
rect 531473 1010232 532363 1010360
rect 579500 1010326 579550 1010442
rect 579497 1010242 579550 1010326
rect 579670 1010242 579798 1010442
rect 579846 1010242 579902 1010442
rect 580022 1010242 580150 1010442
rect 580198 1010242 580254 1010442
rect 580374 1010242 580502 1010442
rect 580550 1010242 580606 1010442
rect 580726 1010242 580854 1010442
rect 580902 1010326 580952 1010442
rect 583363 1010388 584363 1010438
rect 580902 1010242 580955 1010326
rect 579505 1010238 579539 1010242
rect 580913 1010238 580947 1010242
rect 583363 1010232 584363 1010360
rect 75363 1010076 76363 1010204
rect 123473 1010076 124363 1010204
rect 175363 1010076 176363 1010204
rect 227473 1010076 228363 1010204
rect 275473 1010076 276363 1010204
rect 327473 1010076 328363 1010204
rect 379363 1010076 380363 1010204
rect 427473 1010076 428363 1010204
rect 479363 1010076 480363 1010204
rect 531473 1010076 532363 1010204
rect 583363 1010076 584363 1010204
rect 71438 1009928 72438 1009978
rect 73630 1009928 74630 1009978
rect 75363 1009920 76363 1010048
rect 122213 1009928 122630 1009978
rect 123473 1009920 124363 1010048
rect 171438 1009928 172438 1009978
rect 173630 1009928 174630 1009978
rect 175363 1009920 176363 1010048
rect 226213 1009928 226630 1009978
rect 227473 1009920 228363 1010048
rect 274213 1009928 274630 1009978
rect 275473 1009920 276363 1010048
rect 326213 1009928 326630 1009978
rect 327473 1009920 328363 1010048
rect 375438 1009928 376438 1009978
rect 377630 1009928 378630 1009978
rect 379363 1009920 380363 1010048
rect 426213 1009928 426630 1009978
rect 427473 1009920 428363 1010048
rect 475438 1009928 476438 1009978
rect 477630 1009928 478630 1009978
rect 479363 1009920 480363 1010048
rect 530213 1009928 530630 1009978
rect 531473 1009920 532363 1010048
rect 579438 1009928 580438 1009978
rect 581630 1009928 582630 1009978
rect 583363 1009920 584363 1010048
rect 63801 1009309 63851 1009909
rect 63951 1009309 64001 1009909
rect 64081 1009309 64131 1009909
rect 64231 1009309 64359 1009909
rect 64387 1009309 64515 1009909
rect 64543 1009309 64599 1009909
rect 64699 1009309 64827 1009909
rect 64855 1009309 64983 1009909
rect 65011 1009309 65061 1009909
rect 71438 1009772 72438 1009828
rect 73630 1009772 74630 1009828
rect 75363 1009764 76363 1009892
rect 122213 1009772 122630 1009828
rect 123473 1009764 124363 1009892
rect 72776 1009688 72860 1009691
rect 71438 1009616 72438 1009672
rect 72660 1009638 72860 1009688
rect 73208 1009688 73292 1009691
rect 73208 1009683 73408 1009688
rect 73204 1009649 73408 1009683
rect 73208 1009638 73408 1009649
rect 73630 1009616 74630 1009672
rect 75363 1009608 76363 1009736
rect 122213 1009616 122630 1009672
rect 123473 1009608 124363 1009736
rect 71438 1009460 72438 1009516
rect 72660 1009462 72860 1009590
rect 73208 1009462 73408 1009590
rect 73630 1009460 74630 1009516
rect 75363 1009452 76363 1009580
rect 122213 1009460 122630 1009516
rect 123473 1009452 124363 1009580
rect 71438 1009304 72438 1009360
rect 72660 1009286 72860 1009342
rect 73208 1009286 73408 1009342
rect 73630 1009304 74630 1009360
rect 75363 1009296 76363 1009424
rect 122213 1009304 122630 1009360
rect 123473 1009296 124363 1009424
rect 163801 1009309 163851 1009909
rect 163951 1009309 164001 1009909
rect 164081 1009309 164131 1009909
rect 164231 1009309 164359 1009909
rect 164387 1009309 164515 1009909
rect 164543 1009309 164599 1009909
rect 164699 1009309 164827 1009909
rect 164855 1009309 164983 1009909
rect 165011 1009309 165061 1009909
rect 171438 1009772 172438 1009828
rect 173630 1009772 174630 1009828
rect 175363 1009764 176363 1009892
rect 226213 1009772 226630 1009828
rect 227473 1009764 228363 1009892
rect 274213 1009772 274630 1009828
rect 275473 1009764 276363 1009892
rect 326213 1009772 326630 1009828
rect 327473 1009764 328363 1009892
rect 172776 1009688 172860 1009691
rect 171438 1009616 172438 1009672
rect 172660 1009638 172860 1009688
rect 173208 1009688 173292 1009691
rect 173208 1009683 173408 1009688
rect 173204 1009649 173408 1009683
rect 173208 1009638 173408 1009649
rect 173630 1009616 174630 1009672
rect 175363 1009608 176363 1009736
rect 226213 1009616 226630 1009672
rect 227473 1009608 228363 1009736
rect 274213 1009616 274630 1009672
rect 275473 1009608 276363 1009736
rect 326213 1009616 326630 1009672
rect 327473 1009608 328363 1009736
rect 171438 1009460 172438 1009516
rect 172660 1009462 172860 1009590
rect 173208 1009462 173408 1009590
rect 173630 1009460 174630 1009516
rect 175363 1009452 176363 1009580
rect 226213 1009460 226630 1009516
rect 227473 1009452 228363 1009580
rect 274213 1009460 274630 1009516
rect 275473 1009452 276363 1009580
rect 326213 1009460 326630 1009516
rect 327473 1009452 328363 1009580
rect 171438 1009304 172438 1009360
rect 172660 1009286 172860 1009342
rect 173208 1009286 173408 1009342
rect 173630 1009304 174630 1009360
rect 175363 1009296 176363 1009424
rect 226213 1009304 226630 1009360
rect 227473 1009296 228363 1009424
rect 274213 1009304 274630 1009360
rect 275473 1009296 276363 1009424
rect 326213 1009304 326630 1009360
rect 327473 1009296 328363 1009424
rect 367801 1009309 367851 1009909
rect 367951 1009309 368001 1009909
rect 368081 1009309 368131 1009909
rect 368231 1009309 368359 1009909
rect 368387 1009309 368515 1009909
rect 368543 1009309 368599 1009909
rect 368699 1009309 368827 1009909
rect 368855 1009309 368983 1009909
rect 369011 1009309 369061 1009909
rect 375438 1009772 376438 1009828
rect 377630 1009772 378630 1009828
rect 379363 1009764 380363 1009892
rect 426213 1009772 426630 1009828
rect 427473 1009764 428363 1009892
rect 376776 1009688 376860 1009691
rect 375438 1009616 376438 1009672
rect 376660 1009638 376860 1009688
rect 377208 1009688 377292 1009691
rect 377208 1009683 377408 1009688
rect 377204 1009649 377408 1009683
rect 377208 1009638 377408 1009649
rect 377630 1009616 378630 1009672
rect 379363 1009608 380363 1009736
rect 426213 1009616 426630 1009672
rect 427473 1009608 428363 1009736
rect 375438 1009460 376438 1009516
rect 376660 1009462 376860 1009590
rect 377208 1009462 377408 1009590
rect 377630 1009460 378630 1009516
rect 379363 1009452 380363 1009580
rect 426213 1009460 426630 1009516
rect 427473 1009452 428363 1009580
rect 375438 1009304 376438 1009360
rect 376660 1009286 376860 1009342
rect 377208 1009286 377408 1009342
rect 377630 1009304 378630 1009360
rect 379363 1009296 380363 1009424
rect 426213 1009304 426630 1009360
rect 427473 1009296 428363 1009424
rect 467801 1009309 467851 1009909
rect 467951 1009309 468001 1009909
rect 468081 1009309 468131 1009909
rect 468231 1009309 468359 1009909
rect 468387 1009309 468515 1009909
rect 468543 1009309 468599 1009909
rect 468699 1009309 468827 1009909
rect 468855 1009309 468983 1009909
rect 469011 1009309 469061 1009909
rect 475438 1009772 476438 1009828
rect 477630 1009772 478630 1009828
rect 479363 1009764 480363 1009892
rect 530213 1009772 530630 1009828
rect 531473 1009764 532363 1009892
rect 476776 1009688 476860 1009691
rect 475438 1009616 476438 1009672
rect 476660 1009638 476860 1009688
rect 477208 1009688 477292 1009691
rect 477208 1009683 477408 1009688
rect 477204 1009649 477408 1009683
rect 477208 1009638 477408 1009649
rect 477630 1009616 478630 1009672
rect 479363 1009608 480363 1009736
rect 530213 1009616 530630 1009672
rect 531473 1009608 532363 1009736
rect 475438 1009460 476438 1009516
rect 476660 1009462 476860 1009590
rect 477208 1009462 477408 1009590
rect 477630 1009460 478630 1009516
rect 479363 1009452 480363 1009580
rect 530213 1009460 530630 1009516
rect 531473 1009452 532363 1009580
rect 475438 1009304 476438 1009360
rect 476660 1009286 476860 1009342
rect 477208 1009286 477408 1009342
rect 477630 1009304 478630 1009360
rect 479363 1009296 480363 1009424
rect 530213 1009304 530630 1009360
rect 531473 1009296 532363 1009424
rect 571801 1009309 571851 1009909
rect 571951 1009309 572001 1009909
rect 572081 1009309 572131 1009909
rect 572231 1009309 572359 1009909
rect 572387 1009309 572515 1009909
rect 572543 1009309 572599 1009909
rect 572699 1009309 572827 1009909
rect 572855 1009309 572983 1009909
rect 573011 1009309 573061 1009909
rect 579438 1009772 580438 1009828
rect 581630 1009772 582630 1009828
rect 583363 1009764 584363 1009892
rect 580776 1009688 580860 1009691
rect 579438 1009616 580438 1009672
rect 580660 1009638 580860 1009688
rect 581208 1009688 581292 1009691
rect 581208 1009683 581408 1009688
rect 581204 1009649 581408 1009683
rect 581208 1009638 581408 1009649
rect 581630 1009616 582630 1009672
rect 583363 1009608 584363 1009736
rect 579438 1009460 580438 1009516
rect 580660 1009462 580860 1009590
rect 581208 1009462 581408 1009590
rect 581630 1009460 582630 1009516
rect 583363 1009452 584363 1009580
rect 579438 1009304 580438 1009360
rect 580660 1009286 580860 1009342
rect 581208 1009286 581408 1009342
rect 581630 1009304 582630 1009360
rect 583363 1009296 584363 1009424
rect 71438 1009154 72438 1009204
rect 71896 1009151 71980 1009154
rect 72228 1009151 72312 1009154
rect 72660 1009110 72860 1009238
rect 73208 1009110 73408 1009238
rect 73630 1009154 74630 1009204
rect 73756 1009151 73840 1009154
rect 74088 1009151 74172 1009154
rect 75363 1009140 76363 1009268
rect 122213 1009154 122630 1009204
rect 123473 1009140 124363 1009268
rect 171438 1009154 172438 1009204
rect 171896 1009151 171980 1009154
rect 172228 1009151 172312 1009154
rect 67102 1008917 67136 1008951
rect 67171 1008917 67205 1008951
rect 67240 1008917 67274 1008951
rect 67309 1008917 67343 1008951
rect 67378 1008917 67412 1008951
rect 67447 1008917 67481 1008951
rect 67516 1008917 67550 1008951
rect 67585 1008917 67619 1008951
rect 67654 1008917 67688 1008951
rect 67723 1008917 67757 1008951
rect 67792 1008917 67826 1008951
rect 67861 1008917 67895 1008951
rect 67930 1008917 67964 1008951
rect 67999 1008917 68033 1008951
rect 68068 1008917 68102 1008951
rect 68137 1008917 68171 1008951
rect 68206 1008917 68240 1008951
rect 68275 1008917 68309 1008951
rect 68344 1008917 68378 1008951
rect 68413 1008917 68447 1008951
rect 68482 1008917 68516 1008951
rect 68551 1008917 68585 1008951
rect 68620 1008917 68654 1008951
rect 68689 1008917 68723 1008951
rect 68758 1008917 68792 1008951
rect 68827 1008917 68861 1008951
rect 68896 1008917 68930 1008951
rect 68965 1008917 68999 1008951
rect 69034 1008917 69068 1008951
rect 69103 1008917 69137 1008951
rect 69172 1008918 69201 1008951
rect 72660 1008940 72860 1008990
rect 73208 1008940 73408 1008990
rect 75363 1008984 76363 1009112
rect 123473 1008984 124363 1009112
rect 172660 1009110 172860 1009238
rect 173208 1009110 173408 1009238
rect 173630 1009154 174630 1009204
rect 173756 1009151 173840 1009154
rect 174088 1009151 174172 1009154
rect 175363 1009140 176363 1009268
rect 226213 1009154 226630 1009204
rect 227473 1009140 228363 1009268
rect 274213 1009154 274630 1009204
rect 275473 1009140 276363 1009268
rect 326213 1009154 326630 1009204
rect 327473 1009140 328363 1009268
rect 375438 1009154 376438 1009204
rect 375896 1009151 375980 1009154
rect 376228 1009151 376312 1009154
rect 69172 1008917 69235 1008918
rect 67102 1008893 67126 1008917
rect 75363 1008828 76363 1008956
rect 123473 1008828 124363 1008956
rect 167102 1008917 167136 1008951
rect 167171 1008917 167205 1008951
rect 167240 1008917 167274 1008951
rect 167309 1008917 167343 1008951
rect 167378 1008917 167412 1008951
rect 167447 1008917 167481 1008951
rect 167516 1008917 167550 1008951
rect 167585 1008917 167619 1008951
rect 167654 1008917 167688 1008951
rect 167723 1008917 167757 1008951
rect 167792 1008917 167826 1008951
rect 167861 1008917 167895 1008951
rect 167930 1008917 167964 1008951
rect 167999 1008917 168033 1008951
rect 168068 1008917 168102 1008951
rect 168137 1008917 168171 1008951
rect 168206 1008917 168240 1008951
rect 168275 1008917 168309 1008951
rect 168344 1008917 168378 1008951
rect 168413 1008917 168447 1008951
rect 168482 1008917 168516 1008951
rect 168551 1008917 168585 1008951
rect 168620 1008917 168654 1008951
rect 168689 1008917 168723 1008951
rect 168758 1008917 168792 1008951
rect 168827 1008917 168861 1008951
rect 168896 1008917 168930 1008951
rect 168965 1008917 168999 1008951
rect 169034 1008917 169068 1008951
rect 169103 1008917 169137 1008951
rect 169172 1008918 169201 1008951
rect 172660 1008940 172860 1008990
rect 173208 1008940 173408 1008990
rect 175363 1008984 176363 1009112
rect 227473 1008984 228363 1009112
rect 275473 1008984 276363 1009112
rect 327473 1008984 328363 1009112
rect 376660 1009110 376860 1009238
rect 377208 1009110 377408 1009238
rect 377630 1009154 378630 1009204
rect 377756 1009151 377840 1009154
rect 378088 1009151 378172 1009154
rect 379363 1009140 380363 1009268
rect 426213 1009154 426630 1009204
rect 427473 1009140 428363 1009268
rect 475438 1009154 476438 1009204
rect 475896 1009151 475980 1009154
rect 476228 1009151 476312 1009154
rect 169172 1008917 169235 1008918
rect 167102 1008893 167126 1008917
rect 175363 1008828 176363 1008956
rect 227473 1008828 228363 1008956
rect 275473 1008828 276363 1008956
rect 327473 1008828 328363 1008956
rect 371102 1008917 371136 1008951
rect 371171 1008917 371205 1008951
rect 371240 1008917 371274 1008951
rect 371309 1008917 371343 1008951
rect 371378 1008917 371412 1008951
rect 371447 1008917 371481 1008951
rect 371516 1008917 371550 1008951
rect 371585 1008917 371619 1008951
rect 371654 1008917 371688 1008951
rect 371723 1008917 371757 1008951
rect 371792 1008917 371826 1008951
rect 371861 1008917 371895 1008951
rect 371930 1008917 371964 1008951
rect 371999 1008917 372033 1008951
rect 372068 1008917 372102 1008951
rect 372137 1008917 372171 1008951
rect 372206 1008917 372240 1008951
rect 372275 1008917 372309 1008951
rect 372344 1008917 372378 1008951
rect 372413 1008917 372447 1008951
rect 372482 1008917 372516 1008951
rect 372551 1008917 372585 1008951
rect 372620 1008917 372654 1008951
rect 372689 1008917 372723 1008951
rect 372758 1008917 372792 1008951
rect 372827 1008917 372861 1008951
rect 372896 1008917 372930 1008951
rect 372965 1008917 372999 1008951
rect 373034 1008917 373068 1008951
rect 373103 1008917 373137 1008951
rect 373172 1008918 373201 1008951
rect 376660 1008940 376860 1008990
rect 377208 1008940 377408 1008990
rect 379363 1008984 380363 1009112
rect 427473 1008984 428363 1009112
rect 476660 1009110 476860 1009238
rect 477208 1009110 477408 1009238
rect 477630 1009154 478630 1009204
rect 477756 1009151 477840 1009154
rect 478088 1009151 478172 1009154
rect 479363 1009140 480363 1009268
rect 530213 1009154 530630 1009204
rect 531473 1009140 532363 1009268
rect 579438 1009154 580438 1009204
rect 579896 1009151 579980 1009154
rect 580228 1009151 580312 1009154
rect 373172 1008917 373235 1008918
rect 371102 1008893 371126 1008917
rect 379363 1008828 380363 1008956
rect 427473 1008828 428363 1008956
rect 471102 1008917 471136 1008951
rect 471171 1008917 471205 1008951
rect 471240 1008917 471274 1008951
rect 471309 1008917 471343 1008951
rect 471378 1008917 471412 1008951
rect 471447 1008917 471481 1008951
rect 471516 1008917 471550 1008951
rect 471585 1008917 471619 1008951
rect 471654 1008917 471688 1008951
rect 471723 1008917 471757 1008951
rect 471792 1008917 471826 1008951
rect 471861 1008917 471895 1008951
rect 471930 1008917 471964 1008951
rect 471999 1008917 472033 1008951
rect 472068 1008917 472102 1008951
rect 472137 1008917 472171 1008951
rect 472206 1008917 472240 1008951
rect 472275 1008917 472309 1008951
rect 472344 1008917 472378 1008951
rect 472413 1008917 472447 1008951
rect 472482 1008917 472516 1008951
rect 472551 1008917 472585 1008951
rect 472620 1008917 472654 1008951
rect 472689 1008917 472723 1008951
rect 472758 1008917 472792 1008951
rect 472827 1008917 472861 1008951
rect 472896 1008917 472930 1008951
rect 472965 1008917 472999 1008951
rect 473034 1008917 473068 1008951
rect 473103 1008917 473137 1008951
rect 473172 1008918 473201 1008951
rect 476660 1008940 476860 1008990
rect 477208 1008940 477408 1008990
rect 479363 1008984 480363 1009112
rect 531473 1008984 532363 1009112
rect 580660 1009110 580860 1009238
rect 581208 1009110 581408 1009238
rect 581630 1009154 582630 1009204
rect 581756 1009151 581840 1009154
rect 582088 1009151 582172 1009154
rect 583363 1009140 584363 1009268
rect 473172 1008917 473235 1008918
rect 471102 1008893 471126 1008917
rect 479363 1008828 480363 1008956
rect 531473 1008828 532363 1008956
rect 575102 1008917 575136 1008951
rect 575171 1008917 575205 1008951
rect 575240 1008917 575274 1008951
rect 575309 1008917 575343 1008951
rect 575378 1008917 575412 1008951
rect 575447 1008917 575481 1008951
rect 575516 1008917 575550 1008951
rect 575585 1008917 575619 1008951
rect 575654 1008917 575688 1008951
rect 575723 1008917 575757 1008951
rect 575792 1008917 575826 1008951
rect 575861 1008917 575895 1008951
rect 575930 1008917 575964 1008951
rect 575999 1008917 576033 1008951
rect 576068 1008917 576102 1008951
rect 576137 1008917 576171 1008951
rect 576206 1008917 576240 1008951
rect 576275 1008917 576309 1008951
rect 576344 1008917 576378 1008951
rect 576413 1008917 576447 1008951
rect 576482 1008917 576516 1008951
rect 576551 1008917 576585 1008951
rect 576620 1008917 576654 1008951
rect 576689 1008917 576723 1008951
rect 576758 1008917 576792 1008951
rect 576827 1008917 576861 1008951
rect 576896 1008917 576930 1008951
rect 576965 1008917 576999 1008951
rect 577034 1008917 577068 1008951
rect 577103 1008917 577137 1008951
rect 577172 1008918 577201 1008951
rect 580660 1008940 580860 1008990
rect 581208 1008940 581408 1008990
rect 583363 1008984 584363 1009112
rect 577172 1008917 577235 1008918
rect 575102 1008893 575126 1008917
rect 583363 1008828 584363 1008956
rect 75363 1008672 76363 1008800
rect 123473 1008672 124363 1008800
rect 175363 1008672 176363 1008800
rect 227473 1008672 228363 1008800
rect 275473 1008672 276363 1008800
rect 327473 1008672 328363 1008800
rect 379363 1008672 380363 1008800
rect 427473 1008672 428363 1008800
rect 479363 1008672 480363 1008800
rect 531473 1008672 532363 1008800
rect 583363 1008672 584363 1008800
rect 75363 1008516 76363 1008644
rect 123473 1008516 124363 1008644
rect 175363 1008516 176363 1008644
rect 227473 1008516 228363 1008644
rect 275473 1008516 276363 1008644
rect 327473 1008516 328363 1008644
rect 379363 1008516 380363 1008644
rect 427473 1008516 428363 1008644
rect 479363 1008516 480363 1008644
rect 531473 1008516 532363 1008644
rect 583363 1008516 584363 1008644
rect 75363 1008360 76363 1008488
rect 123473 1008360 124363 1008488
rect 175363 1008360 176363 1008488
rect 227473 1008360 228363 1008488
rect 275473 1008360 276363 1008488
rect 327473 1008360 328363 1008488
rect 379363 1008360 380363 1008488
rect 427473 1008360 428363 1008488
rect 479363 1008360 480363 1008488
rect 531473 1008360 532363 1008488
rect 583363 1008360 584363 1008488
rect 75363 1008210 76363 1008260
rect 123363 1008210 124363 1008260
rect 175363 1008210 176363 1008260
rect 227363 1008210 228363 1008260
rect 275363 1008210 276363 1008260
rect 327363 1008210 328363 1008260
rect 379363 1008210 380363 1008260
rect 427363 1008210 428363 1008260
rect 479363 1008210 480363 1008260
rect 531363 1008210 532363 1008260
rect 583363 1008210 584363 1008260
rect 69814 1007798 69838 1007822
rect 69874 1007798 69898 1007822
rect 72189 1007798 72213 1007822
rect 72248 1007798 72272 1007822
rect 169814 1007798 169838 1007822
rect 169874 1007798 169898 1007822
rect 172189 1007798 172213 1007822
rect 172248 1007798 172272 1007822
rect 373814 1007798 373838 1007822
rect 373874 1007798 373898 1007822
rect 376189 1007798 376213 1007822
rect 376248 1007798 376272 1007822
rect 473814 1007798 473838 1007822
rect 473874 1007798 473898 1007822
rect 476189 1007798 476213 1007822
rect 476248 1007798 476272 1007822
rect 577814 1007798 577838 1007822
rect 577874 1007798 577898 1007822
rect 580189 1007798 580213 1007822
rect 580248 1007798 580272 1007822
rect 69850 1007774 69862 1007798
rect 72224 1007774 72237 1007798
rect 169850 1007774 169862 1007798
rect 172224 1007774 172237 1007798
rect 373850 1007774 373862 1007798
rect 376224 1007774 376237 1007798
rect 473850 1007774 473862 1007798
rect 476224 1007774 476237 1007798
rect 577850 1007774 577862 1007798
rect 580224 1007774 580237 1007798
rect 69852 1007710 69886 1007720
rect 69828 1007686 69886 1007710
rect 72234 1007686 72268 1007720
rect 72861 1007710 72895 1007720
rect 169852 1007710 169886 1007720
rect 72837 1007686 72895 1007710
rect 74571 1007685 74595 1007709
rect 169828 1007686 169886 1007710
rect 172234 1007686 172268 1007720
rect 172861 1007710 172895 1007720
rect 373852 1007710 373886 1007720
rect 172837 1007686 172895 1007710
rect 174571 1007685 174595 1007709
rect 373828 1007686 373886 1007710
rect 376234 1007686 376268 1007720
rect 376861 1007710 376895 1007720
rect 473852 1007710 473886 1007720
rect 376837 1007686 376895 1007710
rect 378571 1007685 378595 1007709
rect 473828 1007686 473886 1007710
rect 476234 1007686 476268 1007720
rect 476861 1007710 476895 1007720
rect 577852 1007710 577886 1007720
rect 476837 1007686 476895 1007710
rect 478571 1007685 478595 1007709
rect 577828 1007686 577886 1007710
rect 580234 1007686 580268 1007720
rect 580861 1007710 580895 1007720
rect 580837 1007686 580895 1007710
rect 582571 1007685 582595 1007709
rect 74500 1007669 74571 1007675
rect 174500 1007669 174571 1007675
rect 378500 1007669 378571 1007675
rect 478500 1007669 478571 1007675
rect 582500 1007669 582571 1007675
rect 74547 1007661 74571 1007669
rect 174547 1007661 174571 1007669
rect 378547 1007661 378571 1007669
rect 478547 1007661 478571 1007669
rect 582547 1007661 582571 1007669
rect 62688 1006829 62738 1007429
rect 62858 1006829 62914 1007429
rect 63034 1006829 63084 1007429
rect 61389 1006743 61413 1006767
rect 61450 1006757 61474 1006767
rect 61450 1006753 61484 1006757
rect 61521 1006753 61555 1006757
rect 61592 1006753 61626 1006757
rect 61428 1006743 61650 1006753
rect 61426 1006739 61437 1006743
rect 61450 1006739 61484 1006743
rect 61521 1006739 61555 1006743
rect 61592 1006739 61626 1006743
rect 61426 1006719 61650 1006739
rect 61450 1006699 61474 1006719
rect 63173 1006607 63223 1007607
rect 63323 1006607 63373 1007607
rect 63482 1006607 63532 1007607
rect 63632 1006607 63682 1007607
rect 63797 1007332 64007 1007347
rect 64157 1007332 64217 1007347
rect 64243 1007332 64303 1007347
rect 65817 1007332 65877 1007347
rect 65903 1007332 65963 1007347
rect 66113 1007332 66323 1007347
rect 63812 1007162 63992 1007332
rect 64172 1007162 64202 1007332
rect 64258 1007162 64288 1007332
rect 65832 1007162 65862 1007332
rect 65918 1007162 65948 1007332
rect 66128 1007162 66308 1007332
rect 63801 1007159 64003 1007162
rect 64161 1007159 64213 1007162
rect 64247 1007159 64299 1007162
rect 65821 1007159 65873 1007162
rect 65907 1007159 65959 1007162
rect 66117 1007159 66319 1007162
rect 63797 1007147 64007 1007159
rect 64157 1007147 64217 1007159
rect 64243 1007147 64303 1007159
rect 65817 1007147 65877 1007159
rect 65903 1007147 65963 1007159
rect 66113 1007147 66323 1007159
rect 63797 1007072 64007 1007087
rect 64157 1007072 64217 1007087
rect 64243 1007072 64303 1007087
rect 65817 1007072 65877 1007087
rect 65903 1007072 65963 1007087
rect 66113 1007072 66323 1007087
rect 63812 1006902 63992 1007072
rect 64172 1006902 64202 1007072
rect 64258 1006902 64288 1007072
rect 65832 1006902 65862 1007072
rect 65918 1006902 65948 1007072
rect 66128 1006902 66308 1007072
rect 63801 1006899 64003 1006902
rect 64161 1006899 64213 1006902
rect 64247 1006899 64299 1006902
rect 65821 1006899 65873 1006902
rect 65907 1006899 65959 1006902
rect 66117 1006899 66319 1006902
rect 63797 1006887 64007 1006899
rect 64157 1006887 64217 1006899
rect 64243 1006887 64303 1006899
rect 65817 1006887 65877 1006899
rect 65903 1006887 65963 1006899
rect 66113 1006887 66323 1006899
rect 63797 1006812 64007 1006827
rect 64157 1006812 64217 1006827
rect 64243 1006812 64303 1006827
rect 65817 1006812 65877 1006827
rect 65903 1006812 65963 1006827
rect 66113 1006812 66323 1006827
rect 63812 1006642 63992 1006812
rect 64172 1006807 64202 1006812
rect 64258 1006807 64288 1006812
rect 65832 1006807 65862 1006812
rect 65918 1006807 65948 1006812
rect 66128 1006642 66308 1006812
rect 63801 1006639 64003 1006642
rect 66117 1006639 66319 1006642
rect 63797 1006627 64007 1006639
rect 66113 1006627 66323 1006639
rect 66438 1006607 66488 1007607
rect 66588 1006607 66638 1007607
rect 66747 1006607 66797 1007607
rect 66897 1006607 66947 1007607
rect 68261 1007573 74010 1007585
rect 67036 1006829 67086 1007429
rect 67206 1006829 67262 1007429
rect 67382 1006829 67432 1007429
rect 68261 1006882 68287 1007573
rect 68277 1006879 68287 1006882
rect 68421 1006865 68471 1007465
rect 68591 1006865 68647 1007465
rect 68767 1006865 68817 1007465
rect 68883 1006865 68933 1007465
rect 69053 1006865 69109 1007465
rect 69229 1006865 69357 1007465
rect 69405 1006865 69533 1007465
rect 69581 1006865 69709 1007465
rect 69757 1006865 69807 1007465
rect 69873 1006865 69923 1007465
rect 70043 1006865 70171 1007465
rect 70219 1006865 70275 1007465
rect 70395 1006865 70523 1007465
rect 70571 1006865 70621 1007465
rect 70687 1006865 70737 1007465
rect 70857 1006865 70985 1007465
rect 71033 1006865 71161 1007465
rect 71209 1006865 71337 1007465
rect 71385 1006865 71513 1007465
rect 71561 1006865 71689 1007465
rect 71737 1006865 71793 1007465
rect 71913 1006865 72041 1007465
rect 72089 1006865 72217 1007465
rect 72265 1006865 72393 1007465
rect 72441 1006865 72569 1007465
rect 72617 1006865 72745 1007465
rect 72793 1006865 72849 1007465
rect 72969 1006865 73097 1007465
rect 73145 1006865 73201 1007465
rect 73321 1006865 73449 1007465
rect 73497 1006865 73553 1007465
rect 73673 1006865 73801 1007465
rect 73849 1006865 73899 1007465
rect 75309 1007343 75519 1007355
rect 75545 1007343 75755 1007355
rect 75313 1007340 75515 1007343
rect 75549 1007340 75751 1007343
rect 75324 1007170 75504 1007340
rect 75560 1007170 75740 1007340
rect 75309 1007155 75519 1007170
rect 75545 1007155 75755 1007170
rect 75309 1007042 75519 1007057
rect 75324 1007020 75504 1007042
rect 76011 1006755 76061 1007355
rect 76181 1006755 76237 1007355
rect 76357 1006755 76413 1007355
rect 76533 1006755 76583 1007355
rect 110688 1006829 110738 1007429
rect 110858 1006829 110914 1007429
rect 111034 1006829 111084 1007429
rect 109389 1006743 109413 1006767
rect 109450 1006757 109474 1006767
rect 109450 1006753 109484 1006757
rect 109521 1006753 109555 1006757
rect 109592 1006753 109626 1006757
rect 109428 1006743 109650 1006753
rect 109426 1006739 109437 1006743
rect 109450 1006739 109484 1006743
rect 109521 1006739 109555 1006743
rect 109592 1006739 109626 1006743
rect 109426 1006719 109650 1006739
rect 109450 1006699 109474 1006719
rect 111173 1006607 111223 1007607
rect 123324 1007343 123519 1007355
rect 123545 1007343 123755 1007355
rect 123324 1007340 123515 1007343
rect 123549 1007340 123751 1007343
rect 123324 1007170 123504 1007340
rect 123560 1007170 123740 1007340
rect 123324 1007155 123519 1007170
rect 123545 1007155 123755 1007170
rect 123324 1007042 123519 1007057
rect 123324 1007020 123504 1007042
rect 124011 1006755 124061 1007355
rect 124181 1006755 124237 1007355
rect 124357 1006755 124413 1007355
rect 124533 1006755 124583 1007355
rect 162688 1006829 162738 1007429
rect 162858 1006829 162914 1007429
rect 163034 1006829 163084 1007429
rect 161389 1006743 161413 1006767
rect 161450 1006757 161474 1006767
rect 161450 1006753 161484 1006757
rect 161521 1006753 161555 1006757
rect 161592 1006753 161626 1006757
rect 161428 1006743 161650 1006753
rect 161426 1006739 161437 1006743
rect 161450 1006739 161484 1006743
rect 161521 1006739 161555 1006743
rect 161592 1006739 161626 1006743
rect 161426 1006719 161650 1006739
rect 161450 1006699 161474 1006719
rect 163173 1006607 163223 1007607
rect 163323 1006607 163373 1007607
rect 163482 1006607 163532 1007607
rect 163632 1006607 163682 1007607
rect 163797 1007332 164007 1007347
rect 164157 1007332 164217 1007347
rect 164243 1007332 164303 1007347
rect 165817 1007332 165877 1007347
rect 165903 1007332 165963 1007347
rect 166113 1007332 166323 1007347
rect 163812 1007162 163992 1007332
rect 164172 1007162 164202 1007332
rect 164258 1007162 164288 1007332
rect 165832 1007162 165862 1007332
rect 165918 1007162 165948 1007332
rect 166128 1007162 166308 1007332
rect 163801 1007159 164003 1007162
rect 164161 1007159 164213 1007162
rect 164247 1007159 164299 1007162
rect 165821 1007159 165873 1007162
rect 165907 1007159 165959 1007162
rect 166117 1007159 166319 1007162
rect 163797 1007147 164007 1007159
rect 164157 1007147 164217 1007159
rect 164243 1007147 164303 1007159
rect 165817 1007147 165877 1007159
rect 165903 1007147 165963 1007159
rect 166113 1007147 166323 1007159
rect 163797 1007072 164007 1007087
rect 164157 1007072 164217 1007087
rect 164243 1007072 164303 1007087
rect 165817 1007072 165877 1007087
rect 165903 1007072 165963 1007087
rect 166113 1007072 166323 1007087
rect 163812 1006902 163992 1007072
rect 164172 1006902 164202 1007072
rect 164258 1006902 164288 1007072
rect 165832 1006902 165862 1007072
rect 165918 1006902 165948 1007072
rect 166128 1006902 166308 1007072
rect 163801 1006899 164003 1006902
rect 164161 1006899 164213 1006902
rect 164247 1006899 164299 1006902
rect 165821 1006899 165873 1006902
rect 165907 1006899 165959 1006902
rect 166117 1006899 166319 1006902
rect 163797 1006887 164007 1006899
rect 164157 1006887 164217 1006899
rect 164243 1006887 164303 1006899
rect 165817 1006887 165877 1006899
rect 165903 1006887 165963 1006899
rect 166113 1006887 166323 1006899
rect 163797 1006812 164007 1006827
rect 164157 1006812 164217 1006827
rect 164243 1006812 164303 1006827
rect 165817 1006812 165877 1006827
rect 165903 1006812 165963 1006827
rect 166113 1006812 166323 1006827
rect 163812 1006642 163992 1006812
rect 164172 1006807 164202 1006812
rect 164258 1006807 164288 1006812
rect 165832 1006807 165862 1006812
rect 165918 1006807 165948 1006812
rect 166128 1006642 166308 1006812
rect 163801 1006639 164003 1006642
rect 166117 1006639 166319 1006642
rect 163797 1006627 164007 1006639
rect 166113 1006627 166323 1006639
rect 166438 1006607 166488 1007607
rect 166588 1006607 166638 1007607
rect 166747 1006607 166797 1007607
rect 166897 1006607 166947 1007607
rect 168261 1007573 174010 1007585
rect 167036 1006829 167086 1007429
rect 167206 1006829 167262 1007429
rect 167382 1006829 167432 1007429
rect 168261 1006882 168287 1007573
rect 168277 1006879 168287 1006882
rect 168421 1006865 168471 1007465
rect 168591 1006865 168647 1007465
rect 168767 1006865 168817 1007465
rect 168883 1006865 168933 1007465
rect 169053 1006865 169109 1007465
rect 169229 1006865 169357 1007465
rect 169405 1006865 169533 1007465
rect 169581 1006865 169709 1007465
rect 169757 1006865 169807 1007465
rect 169873 1006865 169923 1007465
rect 170043 1006865 170171 1007465
rect 170219 1006865 170275 1007465
rect 170395 1006865 170523 1007465
rect 170571 1006865 170621 1007465
rect 170687 1006865 170737 1007465
rect 170857 1006865 170985 1007465
rect 171033 1006865 171161 1007465
rect 171209 1006865 171337 1007465
rect 171385 1006865 171513 1007465
rect 171561 1006865 171689 1007465
rect 171737 1006865 171793 1007465
rect 171913 1006865 172041 1007465
rect 172089 1006865 172217 1007465
rect 172265 1006865 172393 1007465
rect 172441 1006865 172569 1007465
rect 172617 1006865 172745 1007465
rect 172793 1006865 172849 1007465
rect 172969 1006865 173097 1007465
rect 173145 1006865 173201 1007465
rect 173321 1006865 173449 1007465
rect 173497 1006865 173553 1007465
rect 173673 1006865 173801 1007465
rect 173849 1006865 173899 1007465
rect 175309 1007343 175519 1007355
rect 175545 1007343 175755 1007355
rect 175313 1007340 175515 1007343
rect 175549 1007340 175751 1007343
rect 175324 1007170 175504 1007340
rect 175560 1007170 175740 1007340
rect 175309 1007155 175519 1007170
rect 175545 1007155 175755 1007170
rect 175309 1007042 175519 1007057
rect 175324 1007020 175504 1007042
rect 176011 1006755 176061 1007355
rect 176181 1006755 176237 1007355
rect 176357 1006755 176413 1007355
rect 176533 1006755 176583 1007355
rect 214688 1006829 214738 1007429
rect 214858 1006829 214914 1007429
rect 215034 1006829 215084 1007429
rect 213389 1006743 213413 1006767
rect 213450 1006757 213474 1006767
rect 213450 1006753 213484 1006757
rect 213521 1006753 213555 1006757
rect 213592 1006753 213626 1006757
rect 213428 1006743 213650 1006753
rect 213426 1006739 213437 1006743
rect 213450 1006739 213484 1006743
rect 213521 1006739 213555 1006743
rect 213592 1006739 213626 1006743
rect 213426 1006719 213650 1006739
rect 213450 1006699 213474 1006719
rect 215173 1006607 215223 1007607
rect 227324 1007343 227519 1007355
rect 227545 1007343 227755 1007355
rect 227324 1007340 227515 1007343
rect 227549 1007340 227751 1007343
rect 227324 1007170 227504 1007340
rect 227560 1007170 227740 1007340
rect 227324 1007155 227519 1007170
rect 227545 1007155 227755 1007170
rect 227324 1007042 227519 1007057
rect 227324 1007020 227504 1007042
rect 228011 1006755 228061 1007355
rect 228181 1006755 228237 1007355
rect 228357 1006755 228413 1007355
rect 228533 1006755 228583 1007355
rect 275324 1007343 275519 1007355
rect 275545 1007343 275755 1007355
rect 275324 1007340 275515 1007343
rect 275549 1007340 275751 1007343
rect 275324 1007170 275504 1007340
rect 275560 1007170 275740 1007340
rect 275324 1007155 275519 1007170
rect 275545 1007155 275755 1007170
rect 275324 1007042 275519 1007057
rect 275324 1007020 275504 1007042
rect 261389 1006743 261413 1006767
rect 261450 1006757 261474 1006767
rect 261450 1006753 261484 1006757
rect 261521 1006753 261555 1006757
rect 261592 1006753 261626 1006757
rect 276011 1006755 276061 1007355
rect 276181 1006755 276237 1007355
rect 276357 1006755 276413 1007355
rect 276533 1006755 276583 1007355
rect 314688 1006829 314738 1007429
rect 314858 1006829 314914 1007429
rect 315034 1006829 315084 1007429
rect 261428 1006743 261650 1006753
rect 313389 1006743 313413 1006767
rect 313450 1006757 313474 1006767
rect 313450 1006753 313484 1006757
rect 313521 1006753 313555 1006757
rect 313592 1006753 313626 1006757
rect 313428 1006743 313650 1006753
rect 261426 1006739 261437 1006743
rect 261450 1006739 261484 1006743
rect 261521 1006739 261555 1006743
rect 261592 1006739 261626 1006743
rect 313426 1006739 313437 1006743
rect 313450 1006739 313484 1006743
rect 313521 1006739 313555 1006743
rect 313592 1006739 313626 1006743
rect 261426 1006719 261650 1006739
rect 313426 1006719 313650 1006739
rect 261450 1006699 261474 1006719
rect 313450 1006699 313474 1006719
rect 315173 1006607 315223 1007607
rect 327324 1007343 327519 1007355
rect 327545 1007343 327755 1007355
rect 327324 1007340 327515 1007343
rect 327549 1007340 327751 1007343
rect 327324 1007170 327504 1007340
rect 327560 1007170 327740 1007340
rect 327324 1007155 327519 1007170
rect 327545 1007155 327755 1007170
rect 327324 1007042 327519 1007057
rect 327324 1007020 327504 1007042
rect 328011 1006755 328061 1007355
rect 328181 1006755 328237 1007355
rect 328357 1006755 328413 1007355
rect 328533 1006755 328583 1007355
rect 366688 1006829 366738 1007429
rect 366858 1006829 366914 1007429
rect 367034 1006829 367084 1007429
rect 365389 1006743 365413 1006767
rect 365450 1006757 365474 1006767
rect 365450 1006753 365484 1006757
rect 365521 1006753 365555 1006757
rect 365592 1006753 365626 1006757
rect 365428 1006743 365650 1006753
rect 365426 1006739 365437 1006743
rect 365450 1006739 365484 1006743
rect 365521 1006739 365555 1006743
rect 365592 1006739 365626 1006743
rect 365426 1006719 365650 1006739
rect 365450 1006699 365474 1006719
rect 367173 1006607 367223 1007607
rect 367323 1006607 367373 1007607
rect 367482 1006607 367532 1007607
rect 367632 1006607 367682 1007607
rect 367797 1007332 368007 1007347
rect 368157 1007332 368217 1007347
rect 368243 1007332 368303 1007347
rect 369817 1007332 369877 1007347
rect 369903 1007332 369963 1007347
rect 370113 1007332 370323 1007347
rect 367812 1007162 367992 1007332
rect 368172 1007162 368202 1007332
rect 368258 1007162 368288 1007332
rect 369832 1007162 369862 1007332
rect 369918 1007162 369948 1007332
rect 370128 1007162 370308 1007332
rect 367801 1007159 368003 1007162
rect 368161 1007159 368213 1007162
rect 368247 1007159 368299 1007162
rect 369821 1007159 369873 1007162
rect 369907 1007159 369959 1007162
rect 370117 1007159 370319 1007162
rect 367797 1007147 368007 1007159
rect 368157 1007147 368217 1007159
rect 368243 1007147 368303 1007159
rect 369817 1007147 369877 1007159
rect 369903 1007147 369963 1007159
rect 370113 1007147 370323 1007159
rect 367797 1007072 368007 1007087
rect 368157 1007072 368217 1007087
rect 368243 1007072 368303 1007087
rect 369817 1007072 369877 1007087
rect 369903 1007072 369963 1007087
rect 370113 1007072 370323 1007087
rect 367812 1006902 367992 1007072
rect 368172 1006902 368202 1007072
rect 368258 1006902 368288 1007072
rect 369832 1006902 369862 1007072
rect 369918 1006902 369948 1007072
rect 370128 1006902 370308 1007072
rect 367801 1006899 368003 1006902
rect 368161 1006899 368213 1006902
rect 368247 1006899 368299 1006902
rect 369821 1006899 369873 1006902
rect 369907 1006899 369959 1006902
rect 370117 1006899 370319 1006902
rect 367797 1006887 368007 1006899
rect 368157 1006887 368217 1006899
rect 368243 1006887 368303 1006899
rect 369817 1006887 369877 1006899
rect 369903 1006887 369963 1006899
rect 370113 1006887 370323 1006899
rect 367797 1006812 368007 1006827
rect 368157 1006812 368217 1006827
rect 368243 1006812 368303 1006827
rect 369817 1006812 369877 1006827
rect 369903 1006812 369963 1006827
rect 370113 1006812 370323 1006827
rect 367812 1006642 367992 1006812
rect 368172 1006807 368202 1006812
rect 368258 1006807 368288 1006812
rect 369832 1006807 369862 1006812
rect 369918 1006807 369948 1006812
rect 370128 1006642 370308 1006812
rect 367801 1006639 368003 1006642
rect 370117 1006639 370319 1006642
rect 367797 1006627 368007 1006639
rect 370113 1006627 370323 1006639
rect 370438 1006607 370488 1007607
rect 370588 1006607 370638 1007607
rect 370747 1006607 370797 1007607
rect 370897 1006607 370947 1007607
rect 372261 1007573 378010 1007585
rect 371036 1006829 371086 1007429
rect 371206 1006829 371262 1007429
rect 371382 1006829 371432 1007429
rect 372261 1006882 372287 1007573
rect 372277 1006879 372287 1006882
rect 372421 1006865 372471 1007465
rect 372591 1006865 372647 1007465
rect 372767 1006865 372817 1007465
rect 372883 1006865 372933 1007465
rect 373053 1006865 373109 1007465
rect 373229 1006865 373357 1007465
rect 373405 1006865 373533 1007465
rect 373581 1006865 373709 1007465
rect 373757 1006865 373807 1007465
rect 373873 1006865 373923 1007465
rect 374043 1006865 374171 1007465
rect 374219 1006865 374275 1007465
rect 374395 1006865 374523 1007465
rect 374571 1006865 374621 1007465
rect 374687 1006865 374737 1007465
rect 374857 1006865 374985 1007465
rect 375033 1006865 375161 1007465
rect 375209 1006865 375337 1007465
rect 375385 1006865 375513 1007465
rect 375561 1006865 375689 1007465
rect 375737 1006865 375793 1007465
rect 375913 1006865 376041 1007465
rect 376089 1006865 376217 1007465
rect 376265 1006865 376393 1007465
rect 376441 1006865 376569 1007465
rect 376617 1006865 376745 1007465
rect 376793 1006865 376849 1007465
rect 376969 1006865 377097 1007465
rect 377145 1006865 377201 1007465
rect 377321 1006865 377449 1007465
rect 377497 1006865 377553 1007465
rect 377673 1006865 377801 1007465
rect 377849 1006865 377899 1007465
rect 379309 1007343 379519 1007355
rect 379545 1007343 379755 1007355
rect 379313 1007340 379515 1007343
rect 379549 1007340 379751 1007343
rect 379324 1007170 379504 1007340
rect 379560 1007170 379740 1007340
rect 379309 1007155 379519 1007170
rect 379545 1007155 379755 1007170
rect 379309 1007042 379519 1007057
rect 379324 1007020 379504 1007042
rect 380011 1006755 380061 1007355
rect 380181 1006755 380237 1007355
rect 380357 1006755 380413 1007355
rect 380533 1006755 380583 1007355
rect 414688 1006829 414738 1007429
rect 414858 1006829 414914 1007429
rect 415034 1006829 415084 1007429
rect 413389 1006743 413413 1006767
rect 413450 1006757 413474 1006767
rect 413450 1006753 413484 1006757
rect 413521 1006753 413555 1006757
rect 413592 1006753 413626 1006757
rect 413428 1006743 413650 1006753
rect 413426 1006739 413437 1006743
rect 413450 1006739 413484 1006743
rect 413521 1006739 413555 1006743
rect 413592 1006739 413626 1006743
rect 413426 1006719 413650 1006739
rect 413450 1006699 413474 1006719
rect 415173 1006607 415223 1007607
rect 427324 1007343 427519 1007355
rect 427545 1007343 427755 1007355
rect 427324 1007340 427515 1007343
rect 427549 1007340 427751 1007343
rect 427324 1007170 427504 1007340
rect 427560 1007170 427740 1007340
rect 427324 1007155 427519 1007170
rect 427545 1007155 427755 1007170
rect 427324 1007042 427519 1007057
rect 427324 1007020 427504 1007042
rect 428011 1006755 428061 1007355
rect 428181 1006755 428237 1007355
rect 428357 1006755 428413 1007355
rect 428533 1006755 428583 1007355
rect 466688 1006829 466738 1007429
rect 466858 1006829 466914 1007429
rect 467034 1006829 467084 1007429
rect 465389 1006743 465413 1006767
rect 465450 1006757 465474 1006767
rect 465450 1006753 465484 1006757
rect 465521 1006753 465555 1006757
rect 465592 1006753 465626 1006757
rect 465428 1006743 465650 1006753
rect 465426 1006739 465437 1006743
rect 465450 1006739 465484 1006743
rect 465521 1006739 465555 1006743
rect 465592 1006739 465626 1006743
rect 465426 1006719 465650 1006739
rect 465450 1006699 465474 1006719
rect 467173 1006607 467223 1007607
rect 467323 1006607 467373 1007607
rect 467482 1006607 467532 1007607
rect 467632 1006607 467682 1007607
rect 467797 1007332 468007 1007347
rect 468157 1007332 468217 1007347
rect 468243 1007332 468303 1007347
rect 469817 1007332 469877 1007347
rect 469903 1007332 469963 1007347
rect 470113 1007332 470323 1007347
rect 467812 1007162 467992 1007332
rect 468172 1007162 468202 1007332
rect 468258 1007162 468288 1007332
rect 469832 1007162 469862 1007332
rect 469918 1007162 469948 1007332
rect 470128 1007162 470308 1007332
rect 467801 1007159 468003 1007162
rect 468161 1007159 468213 1007162
rect 468247 1007159 468299 1007162
rect 469821 1007159 469873 1007162
rect 469907 1007159 469959 1007162
rect 470117 1007159 470319 1007162
rect 467797 1007147 468007 1007159
rect 468157 1007147 468217 1007159
rect 468243 1007147 468303 1007159
rect 469817 1007147 469877 1007159
rect 469903 1007147 469963 1007159
rect 470113 1007147 470323 1007159
rect 467797 1007072 468007 1007087
rect 468157 1007072 468217 1007087
rect 468243 1007072 468303 1007087
rect 469817 1007072 469877 1007087
rect 469903 1007072 469963 1007087
rect 470113 1007072 470323 1007087
rect 467812 1006902 467992 1007072
rect 468172 1006902 468202 1007072
rect 468258 1006902 468288 1007072
rect 469832 1006902 469862 1007072
rect 469918 1006902 469948 1007072
rect 470128 1006902 470308 1007072
rect 467801 1006899 468003 1006902
rect 468161 1006899 468213 1006902
rect 468247 1006899 468299 1006902
rect 469821 1006899 469873 1006902
rect 469907 1006899 469959 1006902
rect 470117 1006899 470319 1006902
rect 467797 1006887 468007 1006899
rect 468157 1006887 468217 1006899
rect 468243 1006887 468303 1006899
rect 469817 1006887 469877 1006899
rect 469903 1006887 469963 1006899
rect 470113 1006887 470323 1006899
rect 467797 1006812 468007 1006827
rect 468157 1006812 468217 1006827
rect 468243 1006812 468303 1006827
rect 469817 1006812 469877 1006827
rect 469903 1006812 469963 1006827
rect 470113 1006812 470323 1006827
rect 467812 1006642 467992 1006812
rect 468172 1006807 468202 1006812
rect 468258 1006807 468288 1006812
rect 469832 1006807 469862 1006812
rect 469918 1006807 469948 1006812
rect 470128 1006642 470308 1006812
rect 467801 1006639 468003 1006642
rect 470117 1006639 470319 1006642
rect 467797 1006627 468007 1006639
rect 470113 1006627 470323 1006639
rect 470438 1006607 470488 1007607
rect 470588 1006607 470638 1007607
rect 470747 1006607 470797 1007607
rect 470897 1006607 470947 1007607
rect 472261 1007573 478010 1007585
rect 471036 1006829 471086 1007429
rect 471206 1006829 471262 1007429
rect 471382 1006829 471432 1007429
rect 472261 1006882 472287 1007573
rect 472277 1006879 472287 1006882
rect 472421 1006865 472471 1007465
rect 472591 1006865 472647 1007465
rect 472767 1006865 472817 1007465
rect 472883 1006865 472933 1007465
rect 473053 1006865 473109 1007465
rect 473229 1006865 473357 1007465
rect 473405 1006865 473533 1007465
rect 473581 1006865 473709 1007465
rect 473757 1006865 473807 1007465
rect 473873 1006865 473923 1007465
rect 474043 1006865 474171 1007465
rect 474219 1006865 474275 1007465
rect 474395 1006865 474523 1007465
rect 474571 1006865 474621 1007465
rect 474687 1006865 474737 1007465
rect 474857 1006865 474985 1007465
rect 475033 1006865 475161 1007465
rect 475209 1006865 475337 1007465
rect 475385 1006865 475513 1007465
rect 475561 1006865 475689 1007465
rect 475737 1006865 475793 1007465
rect 475913 1006865 476041 1007465
rect 476089 1006865 476217 1007465
rect 476265 1006865 476393 1007465
rect 476441 1006865 476569 1007465
rect 476617 1006865 476745 1007465
rect 476793 1006865 476849 1007465
rect 476969 1006865 477097 1007465
rect 477145 1006865 477201 1007465
rect 477321 1006865 477449 1007465
rect 477497 1006865 477553 1007465
rect 477673 1006865 477801 1007465
rect 477849 1006865 477899 1007465
rect 479309 1007343 479519 1007355
rect 479545 1007343 479755 1007355
rect 479313 1007340 479515 1007343
rect 479549 1007340 479751 1007343
rect 479324 1007170 479504 1007340
rect 479560 1007170 479740 1007340
rect 479309 1007155 479519 1007170
rect 479545 1007155 479755 1007170
rect 479309 1007042 479519 1007057
rect 479324 1007020 479504 1007042
rect 480011 1006755 480061 1007355
rect 480181 1006755 480237 1007355
rect 480357 1006755 480413 1007355
rect 480533 1006755 480583 1007355
rect 518688 1006829 518738 1007429
rect 518858 1006829 518914 1007429
rect 519034 1006829 519084 1007429
rect 517389 1006743 517413 1006767
rect 517450 1006757 517474 1006767
rect 517450 1006753 517484 1006757
rect 517521 1006753 517555 1006757
rect 517592 1006753 517626 1006757
rect 517428 1006743 517650 1006753
rect 517426 1006739 517437 1006743
rect 517450 1006739 517484 1006743
rect 517521 1006739 517555 1006743
rect 517592 1006739 517626 1006743
rect 517426 1006719 517650 1006739
rect 517450 1006699 517474 1006719
rect 519173 1006607 519223 1007607
rect 531324 1007343 531519 1007355
rect 531545 1007343 531755 1007355
rect 531324 1007340 531515 1007343
rect 531549 1007340 531751 1007343
rect 531324 1007170 531504 1007340
rect 531560 1007170 531740 1007340
rect 531324 1007155 531519 1007170
rect 531545 1007155 531755 1007170
rect 531324 1007042 531519 1007057
rect 531324 1007020 531504 1007042
rect 532011 1006755 532061 1007355
rect 532181 1006755 532237 1007355
rect 532357 1006755 532413 1007355
rect 532533 1006755 532583 1007355
rect 570688 1006829 570738 1007429
rect 570858 1006829 570914 1007429
rect 571034 1006829 571084 1007429
rect 569389 1006743 569413 1006767
rect 569450 1006757 569474 1006767
rect 569450 1006753 569484 1006757
rect 569521 1006753 569555 1006757
rect 569592 1006753 569626 1006757
rect 569428 1006743 569650 1006753
rect 569426 1006739 569437 1006743
rect 569450 1006739 569484 1006743
rect 569521 1006739 569555 1006743
rect 569592 1006739 569626 1006743
rect 569426 1006719 569650 1006739
rect 569450 1006699 569474 1006719
rect 571173 1006607 571223 1007607
rect 571323 1006607 571373 1007607
rect 571482 1006607 571532 1007607
rect 571632 1006607 571682 1007607
rect 571797 1007332 572007 1007347
rect 572157 1007332 572217 1007347
rect 572243 1007332 572303 1007347
rect 573817 1007332 573877 1007347
rect 573903 1007332 573963 1007347
rect 574113 1007332 574323 1007347
rect 571812 1007162 571992 1007332
rect 572172 1007162 572202 1007332
rect 572258 1007162 572288 1007332
rect 573832 1007162 573862 1007332
rect 573918 1007162 573948 1007332
rect 574128 1007162 574308 1007332
rect 571801 1007159 572003 1007162
rect 572161 1007159 572213 1007162
rect 572247 1007159 572299 1007162
rect 573821 1007159 573873 1007162
rect 573907 1007159 573959 1007162
rect 574117 1007159 574319 1007162
rect 571797 1007147 572007 1007159
rect 572157 1007147 572217 1007159
rect 572243 1007147 572303 1007159
rect 573817 1007147 573877 1007159
rect 573903 1007147 573963 1007159
rect 574113 1007147 574323 1007159
rect 571797 1007072 572007 1007087
rect 572157 1007072 572217 1007087
rect 572243 1007072 572303 1007087
rect 573817 1007072 573877 1007087
rect 573903 1007072 573963 1007087
rect 574113 1007072 574323 1007087
rect 571812 1006902 571992 1007072
rect 572172 1006902 572202 1007072
rect 572258 1006902 572288 1007072
rect 573832 1006902 573862 1007072
rect 573918 1006902 573948 1007072
rect 574128 1006902 574308 1007072
rect 571801 1006899 572003 1006902
rect 572161 1006899 572213 1006902
rect 572247 1006899 572299 1006902
rect 573821 1006899 573873 1006902
rect 573907 1006899 573959 1006902
rect 574117 1006899 574319 1006902
rect 571797 1006887 572007 1006899
rect 572157 1006887 572217 1006899
rect 572243 1006887 572303 1006899
rect 573817 1006887 573877 1006899
rect 573903 1006887 573963 1006899
rect 574113 1006887 574323 1006899
rect 571797 1006812 572007 1006827
rect 572157 1006812 572217 1006827
rect 572243 1006812 572303 1006827
rect 573817 1006812 573877 1006827
rect 573903 1006812 573963 1006827
rect 574113 1006812 574323 1006827
rect 571812 1006642 571992 1006812
rect 572172 1006807 572202 1006812
rect 572258 1006807 572288 1006812
rect 573832 1006807 573862 1006812
rect 573918 1006807 573948 1006812
rect 574128 1006642 574308 1006812
rect 571801 1006639 572003 1006642
rect 574117 1006639 574319 1006642
rect 571797 1006627 572007 1006639
rect 574113 1006627 574323 1006639
rect 574438 1006607 574488 1007607
rect 574588 1006607 574638 1007607
rect 574747 1006607 574797 1007607
rect 574897 1006607 574947 1007607
rect 576261 1007573 582010 1007585
rect 575036 1006829 575086 1007429
rect 575206 1006829 575262 1007429
rect 575382 1006829 575432 1007429
rect 576261 1006882 576287 1007573
rect 576277 1006879 576287 1006882
rect 576421 1006865 576471 1007465
rect 576591 1006865 576647 1007465
rect 576767 1006865 576817 1007465
rect 576883 1006865 576933 1007465
rect 577053 1006865 577109 1007465
rect 577229 1006865 577357 1007465
rect 577405 1006865 577533 1007465
rect 577581 1006865 577709 1007465
rect 577757 1006865 577807 1007465
rect 577873 1006865 577923 1007465
rect 578043 1006865 578171 1007465
rect 578219 1006865 578275 1007465
rect 578395 1006865 578523 1007465
rect 578571 1006865 578621 1007465
rect 578687 1006865 578737 1007465
rect 578857 1006865 578985 1007465
rect 579033 1006865 579161 1007465
rect 579209 1006865 579337 1007465
rect 579385 1006865 579513 1007465
rect 579561 1006865 579689 1007465
rect 579737 1006865 579793 1007465
rect 579913 1006865 580041 1007465
rect 580089 1006865 580217 1007465
rect 580265 1006865 580393 1007465
rect 580441 1006865 580569 1007465
rect 580617 1006865 580745 1007465
rect 580793 1006865 580849 1007465
rect 580969 1006865 581097 1007465
rect 581145 1006865 581201 1007465
rect 581321 1006865 581449 1007465
rect 581497 1006865 581553 1007465
rect 581673 1006865 581801 1007465
rect 581849 1006865 581899 1007465
rect 583309 1007343 583519 1007355
rect 583545 1007343 583755 1007355
rect 583313 1007340 583515 1007343
rect 583549 1007340 583751 1007343
rect 583324 1007170 583504 1007340
rect 583560 1007170 583740 1007340
rect 583309 1007155 583519 1007170
rect 583545 1007155 583755 1007170
rect 583309 1007042 583519 1007057
rect 583324 1007020 583504 1007042
rect 584011 1006755 584061 1007355
rect 584181 1006755 584237 1007355
rect 584357 1006755 584413 1007355
rect 584533 1006755 584583 1007355
rect 63797 1006498 64007 1006513
rect 66113 1006498 66323 1006513
rect 63812 1006328 63992 1006498
rect 66128 1006328 66308 1006498
rect 63801 1006325 64003 1006328
rect 66117 1006325 66319 1006328
rect 63797 1006313 64007 1006325
rect 66113 1006313 66323 1006325
rect 63201 1006238 63411 1006253
rect 63437 1006238 63647 1006253
rect 63797 1006238 64007 1006253
rect 64157 1006238 64217 1006253
rect 64243 1006238 64303 1006253
rect 65817 1006238 65877 1006253
rect 65903 1006238 65963 1006253
rect 66113 1006238 66323 1006253
rect 66473 1006238 66683 1006253
rect 66709 1006238 66919 1006253
rect 62176 1005537 62226 1006137
rect 62326 1005537 62382 1006137
rect 62482 1005537 62532 1006137
rect 63216 1006068 63396 1006238
rect 63452 1006068 63632 1006238
rect 63812 1006068 63992 1006238
rect 64172 1006068 64202 1006238
rect 64258 1006068 64288 1006238
rect 63205 1006065 63407 1006068
rect 63441 1006065 63643 1006068
rect 63801 1006065 64003 1006068
rect 64161 1006065 64213 1006068
rect 64247 1006065 64299 1006068
rect 63201 1006053 63411 1006065
rect 63437 1006053 63647 1006065
rect 63797 1006053 64007 1006065
rect 64157 1006053 64217 1006065
rect 64243 1006053 64303 1006065
rect 63201 1005978 63411 1005993
rect 63437 1005978 63647 1005993
rect 63797 1005978 64007 1005993
rect 64157 1005978 64217 1005993
rect 64243 1005978 64303 1005993
rect 63216 1005808 63396 1005978
rect 63452 1005808 63632 1005978
rect 63812 1005808 63992 1005978
rect 64172 1005808 64202 1005978
rect 64258 1005808 64288 1005978
rect 63205 1005805 63407 1005808
rect 63441 1005805 63643 1005808
rect 63801 1005805 64003 1005808
rect 64161 1005805 64213 1005808
rect 64247 1005805 64299 1005808
rect 63201 1005793 63411 1005805
rect 63437 1005793 63647 1005805
rect 63797 1005793 64007 1005805
rect 64157 1005793 64217 1005805
rect 64243 1005793 64303 1005805
rect 64449 1005803 64465 1006119
rect 65653 1005803 65671 1006119
rect 65832 1006068 65862 1006238
rect 65918 1006068 65948 1006238
rect 66128 1006068 66308 1006238
rect 66488 1006068 66668 1006238
rect 66724 1006068 66904 1006238
rect 65821 1006065 65873 1006068
rect 65907 1006065 65959 1006068
rect 66117 1006065 66319 1006068
rect 66477 1006065 66679 1006068
rect 66713 1006065 66915 1006068
rect 65817 1006053 65877 1006065
rect 65903 1006053 65963 1006065
rect 66113 1006053 66323 1006065
rect 66473 1006053 66683 1006065
rect 66709 1006053 66919 1006065
rect 65817 1005978 65877 1005993
rect 65903 1005978 65963 1005993
rect 66113 1005978 66323 1005993
rect 66473 1005978 66683 1005993
rect 66709 1005978 66919 1005993
rect 65832 1005808 65862 1005978
rect 65918 1005808 65948 1005978
rect 66128 1005808 66308 1005978
rect 66488 1005808 66668 1005978
rect 66724 1005808 66904 1005978
rect 65821 1005805 65873 1005808
rect 65907 1005805 65959 1005808
rect 66117 1005805 66319 1005808
rect 66477 1005805 66679 1005808
rect 66713 1005805 66915 1005808
rect 64449 1005777 64453 1005803
rect 65817 1005793 65877 1005805
rect 65903 1005793 65963 1005805
rect 66113 1005793 66323 1005805
rect 66473 1005793 66683 1005805
rect 66709 1005793 66919 1005805
rect 63797 1005718 64007 1005733
rect 64157 1005718 64217 1005733
rect 64243 1005718 64303 1005733
rect 63812 1005548 63992 1005718
rect 64172 1005679 64202 1005718
rect 64258 1005679 64288 1005718
rect 63801 1005545 64003 1005548
rect 63797 1005533 64007 1005545
rect 64415 1005539 64453 1005777
rect 65673 1005539 65705 1005777
rect 65817 1005718 65877 1005733
rect 65903 1005718 65963 1005733
rect 66113 1005718 66323 1005733
rect 65832 1005679 65862 1005718
rect 65918 1005679 65948 1005718
rect 66128 1005548 66308 1005718
rect 66117 1005545 66319 1005548
rect 64415 1005513 64449 1005539
rect 66113 1005533 66323 1005545
rect 67588 1005537 67638 1006137
rect 67738 1005537 67794 1006137
rect 67894 1005537 67944 1006137
rect 68441 1005551 68491 1006551
rect 68591 1005551 68647 1006551
rect 68747 1005551 68797 1006551
rect 68883 1005551 68933 1006551
rect 69033 1005551 69089 1006551
rect 69189 1005551 69245 1006551
rect 69345 1005551 69401 1006551
rect 69501 1005551 69551 1006551
rect 69617 1005551 69667 1006551
rect 69767 1005551 69895 1006551
rect 69923 1005551 70051 1006551
rect 70079 1005551 70207 1006551
rect 70235 1005551 70363 1006551
rect 70391 1005551 70519 1006551
rect 70547 1005551 70603 1006551
rect 70703 1005551 70831 1006551
rect 70859 1005551 70987 1006551
rect 71015 1005551 71143 1006551
rect 71171 1005551 71299 1006551
rect 71327 1005551 71455 1006551
rect 71483 1005551 71539 1006551
rect 71659 1005551 71787 1006551
rect 71835 1005551 71963 1006551
rect 72011 1005551 72139 1006551
rect 72187 1005551 72315 1006551
rect 72363 1005551 72491 1006551
rect 72539 1005551 72667 1006551
rect 72715 1005551 72843 1006551
rect 72891 1005551 72941 1006551
rect 73007 1005551 73057 1006551
rect 73157 1005551 73285 1006551
rect 73313 1005551 73441 1006551
rect 73469 1005551 73597 1006551
rect 73625 1005551 73681 1006551
rect 73781 1005551 73909 1006551
rect 73937 1005551 74065 1006551
rect 74093 1005551 74221 1006551
rect 74249 1005551 74299 1006551
rect 74890 1005992 74943 1006142
rect 74893 1005895 74943 1005992
rect 74890 1005673 74943 1005895
rect 74893 1005542 74943 1005673
rect 75063 1005542 75119 1006142
rect 75239 1005542 75289 1006142
rect 75665 1005547 75715 1006147
rect 75835 1005547 75885 1006147
rect 110176 1005537 110226 1006137
rect 110326 1005537 110382 1006137
rect 110482 1005537 110532 1006137
rect 111216 1006053 111253 1006253
rect 111216 1005793 111253 1005993
rect 122249 1005551 122299 1006551
rect 163797 1006498 164007 1006513
rect 166113 1006498 166323 1006513
rect 163812 1006328 163992 1006498
rect 166128 1006328 166308 1006498
rect 163801 1006325 164003 1006328
rect 166117 1006325 166319 1006328
rect 163797 1006313 164007 1006325
rect 166113 1006313 166323 1006325
rect 163201 1006238 163411 1006253
rect 163437 1006238 163647 1006253
rect 163797 1006238 164007 1006253
rect 164157 1006238 164217 1006253
rect 164243 1006238 164303 1006253
rect 165817 1006238 165877 1006253
rect 165903 1006238 165963 1006253
rect 166113 1006238 166323 1006253
rect 166473 1006238 166683 1006253
rect 166709 1006238 166919 1006253
rect 122893 1005542 122943 1006142
rect 123063 1005542 123119 1006142
rect 123239 1005542 123289 1006142
rect 123665 1005547 123715 1006147
rect 123835 1005547 123885 1006147
rect 162176 1005537 162226 1006137
rect 162326 1005537 162382 1006137
rect 162482 1005537 162532 1006137
rect 163216 1006068 163396 1006238
rect 163452 1006068 163632 1006238
rect 163812 1006068 163992 1006238
rect 164172 1006068 164202 1006238
rect 164258 1006068 164288 1006238
rect 163205 1006065 163407 1006068
rect 163441 1006065 163643 1006068
rect 163801 1006065 164003 1006068
rect 164161 1006065 164213 1006068
rect 164247 1006065 164299 1006068
rect 163201 1006053 163411 1006065
rect 163437 1006053 163647 1006065
rect 163797 1006053 164007 1006065
rect 164157 1006053 164217 1006065
rect 164243 1006053 164303 1006065
rect 163201 1005978 163411 1005993
rect 163437 1005978 163647 1005993
rect 163797 1005978 164007 1005993
rect 164157 1005978 164217 1005993
rect 164243 1005978 164303 1005993
rect 163216 1005808 163396 1005978
rect 163452 1005808 163632 1005978
rect 163812 1005808 163992 1005978
rect 164172 1005808 164202 1005978
rect 164258 1005808 164288 1005978
rect 163205 1005805 163407 1005808
rect 163441 1005805 163643 1005808
rect 163801 1005805 164003 1005808
rect 164161 1005805 164213 1005808
rect 164247 1005805 164299 1005808
rect 163201 1005793 163411 1005805
rect 163437 1005793 163647 1005805
rect 163797 1005793 164007 1005805
rect 164157 1005793 164217 1005805
rect 164243 1005793 164303 1005805
rect 164449 1005803 164465 1006119
rect 165653 1005803 165671 1006119
rect 165832 1006068 165862 1006238
rect 165918 1006068 165948 1006238
rect 166128 1006068 166308 1006238
rect 166488 1006068 166668 1006238
rect 166724 1006068 166904 1006238
rect 165821 1006065 165873 1006068
rect 165907 1006065 165959 1006068
rect 166117 1006065 166319 1006068
rect 166477 1006065 166679 1006068
rect 166713 1006065 166915 1006068
rect 165817 1006053 165877 1006065
rect 165903 1006053 165963 1006065
rect 166113 1006053 166323 1006065
rect 166473 1006053 166683 1006065
rect 166709 1006053 166919 1006065
rect 165817 1005978 165877 1005993
rect 165903 1005978 165963 1005993
rect 166113 1005978 166323 1005993
rect 166473 1005978 166683 1005993
rect 166709 1005978 166919 1005993
rect 165832 1005808 165862 1005978
rect 165918 1005808 165948 1005978
rect 166128 1005808 166308 1005978
rect 166488 1005808 166668 1005978
rect 166724 1005808 166904 1005978
rect 165821 1005805 165873 1005808
rect 165907 1005805 165959 1005808
rect 166117 1005805 166319 1005808
rect 166477 1005805 166679 1005808
rect 166713 1005805 166915 1005808
rect 164449 1005777 164453 1005803
rect 165817 1005793 165877 1005805
rect 165903 1005793 165963 1005805
rect 166113 1005793 166323 1005805
rect 166473 1005793 166683 1005805
rect 166709 1005793 166919 1005805
rect 163797 1005718 164007 1005733
rect 164157 1005718 164217 1005733
rect 164243 1005718 164303 1005733
rect 163812 1005548 163992 1005718
rect 164172 1005679 164202 1005718
rect 164258 1005679 164288 1005718
rect 163801 1005545 164003 1005548
rect 163797 1005533 164007 1005545
rect 164415 1005539 164453 1005777
rect 165673 1005539 165705 1005777
rect 165817 1005718 165877 1005733
rect 165903 1005718 165963 1005733
rect 166113 1005718 166323 1005733
rect 165832 1005679 165862 1005718
rect 165918 1005679 165948 1005718
rect 166128 1005548 166308 1005718
rect 166117 1005545 166319 1005548
rect 164415 1005513 164449 1005539
rect 166113 1005533 166323 1005545
rect 167588 1005537 167638 1006137
rect 167738 1005537 167794 1006137
rect 167894 1005537 167944 1006137
rect 168441 1005551 168491 1006551
rect 168591 1005551 168647 1006551
rect 168747 1005551 168797 1006551
rect 168883 1005551 168933 1006551
rect 169033 1005551 169089 1006551
rect 169189 1005551 169245 1006551
rect 169345 1005551 169401 1006551
rect 169501 1005551 169551 1006551
rect 169617 1005551 169667 1006551
rect 169767 1005551 169895 1006551
rect 169923 1005551 170051 1006551
rect 170079 1005551 170207 1006551
rect 170235 1005551 170363 1006551
rect 170391 1005551 170519 1006551
rect 170547 1005551 170603 1006551
rect 170703 1005551 170831 1006551
rect 170859 1005551 170987 1006551
rect 171015 1005551 171143 1006551
rect 171171 1005551 171299 1006551
rect 171327 1005551 171455 1006551
rect 171483 1005551 171539 1006551
rect 171659 1005551 171787 1006551
rect 171835 1005551 171963 1006551
rect 172011 1005551 172139 1006551
rect 172187 1005551 172315 1006551
rect 172363 1005551 172491 1006551
rect 172539 1005551 172667 1006551
rect 172715 1005551 172843 1006551
rect 172891 1005551 172941 1006551
rect 173007 1005551 173057 1006551
rect 173157 1005551 173285 1006551
rect 173313 1005551 173441 1006551
rect 173469 1005551 173597 1006551
rect 173625 1005551 173681 1006551
rect 173781 1005551 173909 1006551
rect 173937 1005551 174065 1006551
rect 174093 1005551 174221 1006551
rect 174249 1005551 174299 1006551
rect 174890 1005992 174943 1006142
rect 174893 1005895 174943 1005992
rect 174890 1005673 174943 1005895
rect 174893 1005542 174943 1005673
rect 175063 1005542 175119 1006142
rect 175239 1005542 175289 1006142
rect 175665 1005547 175715 1006147
rect 175835 1005547 175885 1006147
rect 214176 1005537 214226 1006137
rect 214326 1005537 214382 1006137
rect 214482 1005537 214532 1006137
rect 215216 1006053 215253 1006253
rect 215216 1005793 215253 1005993
rect 226249 1005551 226299 1006551
rect 226893 1005542 226943 1006142
rect 227063 1005542 227119 1006142
rect 227239 1005542 227289 1006142
rect 227665 1005547 227715 1006147
rect 227835 1005547 227885 1006147
rect 274249 1005551 274299 1006551
rect 274893 1005542 274943 1006142
rect 275063 1005542 275119 1006142
rect 275239 1005542 275289 1006142
rect 275665 1005547 275715 1006147
rect 275835 1005547 275885 1006147
rect 314176 1005537 314226 1006137
rect 314326 1005537 314382 1006137
rect 314482 1005537 314532 1006137
rect 315216 1006053 315253 1006253
rect 315216 1005793 315253 1005993
rect 326249 1005551 326299 1006551
rect 367797 1006498 368007 1006513
rect 370113 1006498 370323 1006513
rect 367812 1006328 367992 1006498
rect 370128 1006328 370308 1006498
rect 367801 1006325 368003 1006328
rect 370117 1006325 370319 1006328
rect 367797 1006313 368007 1006325
rect 370113 1006313 370323 1006325
rect 367201 1006238 367411 1006253
rect 367437 1006238 367647 1006253
rect 367797 1006238 368007 1006253
rect 368157 1006238 368217 1006253
rect 368243 1006238 368303 1006253
rect 369817 1006238 369877 1006253
rect 369903 1006238 369963 1006253
rect 370113 1006238 370323 1006253
rect 370473 1006238 370683 1006253
rect 370709 1006238 370919 1006253
rect 326893 1005542 326943 1006142
rect 327063 1005542 327119 1006142
rect 327239 1005542 327289 1006142
rect 327665 1005547 327715 1006147
rect 327835 1005547 327885 1006147
rect 366176 1005537 366226 1006137
rect 366326 1005537 366382 1006137
rect 366482 1005537 366532 1006137
rect 367216 1006068 367396 1006238
rect 367452 1006068 367632 1006238
rect 367812 1006068 367992 1006238
rect 368172 1006068 368202 1006238
rect 368258 1006068 368288 1006238
rect 367205 1006065 367407 1006068
rect 367441 1006065 367643 1006068
rect 367801 1006065 368003 1006068
rect 368161 1006065 368213 1006068
rect 368247 1006065 368299 1006068
rect 367201 1006053 367411 1006065
rect 367437 1006053 367647 1006065
rect 367797 1006053 368007 1006065
rect 368157 1006053 368217 1006065
rect 368243 1006053 368303 1006065
rect 367201 1005978 367411 1005993
rect 367437 1005978 367647 1005993
rect 367797 1005978 368007 1005993
rect 368157 1005978 368217 1005993
rect 368243 1005978 368303 1005993
rect 367216 1005808 367396 1005978
rect 367452 1005808 367632 1005978
rect 367812 1005808 367992 1005978
rect 368172 1005808 368202 1005978
rect 368258 1005808 368288 1005978
rect 367205 1005805 367407 1005808
rect 367441 1005805 367643 1005808
rect 367801 1005805 368003 1005808
rect 368161 1005805 368213 1005808
rect 368247 1005805 368299 1005808
rect 367201 1005793 367411 1005805
rect 367437 1005793 367647 1005805
rect 367797 1005793 368007 1005805
rect 368157 1005793 368217 1005805
rect 368243 1005793 368303 1005805
rect 368449 1005803 368465 1006119
rect 369653 1005803 369671 1006119
rect 369832 1006068 369862 1006238
rect 369918 1006068 369948 1006238
rect 370128 1006068 370308 1006238
rect 370488 1006068 370668 1006238
rect 370724 1006068 370904 1006238
rect 369821 1006065 369873 1006068
rect 369907 1006065 369959 1006068
rect 370117 1006065 370319 1006068
rect 370477 1006065 370679 1006068
rect 370713 1006065 370915 1006068
rect 369817 1006053 369877 1006065
rect 369903 1006053 369963 1006065
rect 370113 1006053 370323 1006065
rect 370473 1006053 370683 1006065
rect 370709 1006053 370919 1006065
rect 369817 1005978 369877 1005993
rect 369903 1005978 369963 1005993
rect 370113 1005978 370323 1005993
rect 370473 1005978 370683 1005993
rect 370709 1005978 370919 1005993
rect 369832 1005808 369862 1005978
rect 369918 1005808 369948 1005978
rect 370128 1005808 370308 1005978
rect 370488 1005808 370668 1005978
rect 370724 1005808 370904 1005978
rect 369821 1005805 369873 1005808
rect 369907 1005805 369959 1005808
rect 370117 1005805 370319 1005808
rect 370477 1005805 370679 1005808
rect 370713 1005805 370915 1005808
rect 368449 1005777 368453 1005803
rect 369817 1005793 369877 1005805
rect 369903 1005793 369963 1005805
rect 370113 1005793 370323 1005805
rect 370473 1005793 370683 1005805
rect 370709 1005793 370919 1005805
rect 367797 1005718 368007 1005733
rect 368157 1005718 368217 1005733
rect 368243 1005718 368303 1005733
rect 367812 1005548 367992 1005718
rect 368172 1005679 368202 1005718
rect 368258 1005679 368288 1005718
rect 367801 1005545 368003 1005548
rect 367797 1005533 368007 1005545
rect 368415 1005539 368453 1005777
rect 369673 1005539 369705 1005777
rect 369817 1005718 369877 1005733
rect 369903 1005718 369963 1005733
rect 370113 1005718 370323 1005733
rect 369832 1005679 369862 1005718
rect 369918 1005679 369948 1005718
rect 370128 1005548 370308 1005718
rect 370117 1005545 370319 1005548
rect 368415 1005513 368449 1005539
rect 370113 1005533 370323 1005545
rect 371588 1005537 371638 1006137
rect 371738 1005537 371794 1006137
rect 371894 1005537 371944 1006137
rect 372441 1005551 372491 1006551
rect 372591 1005551 372647 1006551
rect 372747 1005551 372797 1006551
rect 372883 1005551 372933 1006551
rect 373033 1005551 373089 1006551
rect 373189 1005551 373245 1006551
rect 373345 1005551 373401 1006551
rect 373501 1005551 373551 1006551
rect 373617 1005551 373667 1006551
rect 373767 1005551 373895 1006551
rect 373923 1005551 374051 1006551
rect 374079 1005551 374207 1006551
rect 374235 1005551 374363 1006551
rect 374391 1005551 374519 1006551
rect 374547 1005551 374603 1006551
rect 374703 1005551 374831 1006551
rect 374859 1005551 374987 1006551
rect 375015 1005551 375143 1006551
rect 375171 1005551 375299 1006551
rect 375327 1005551 375455 1006551
rect 375483 1005551 375539 1006551
rect 375659 1005551 375787 1006551
rect 375835 1005551 375963 1006551
rect 376011 1005551 376139 1006551
rect 376187 1005551 376315 1006551
rect 376363 1005551 376491 1006551
rect 376539 1005551 376667 1006551
rect 376715 1005551 376843 1006551
rect 376891 1005551 376941 1006551
rect 377007 1005551 377057 1006551
rect 377157 1005551 377285 1006551
rect 377313 1005551 377441 1006551
rect 377469 1005551 377597 1006551
rect 377625 1005551 377681 1006551
rect 377781 1005551 377909 1006551
rect 377937 1005551 378065 1006551
rect 378093 1005551 378221 1006551
rect 378249 1005551 378299 1006551
rect 378890 1005992 378943 1006142
rect 378893 1005895 378943 1005992
rect 378890 1005673 378943 1005895
rect 378893 1005542 378943 1005673
rect 379063 1005542 379119 1006142
rect 379239 1005542 379289 1006142
rect 379665 1005547 379715 1006147
rect 379835 1005547 379885 1006147
rect 414176 1005537 414226 1006137
rect 414326 1005537 414382 1006137
rect 414482 1005537 414532 1006137
rect 415216 1006053 415253 1006253
rect 415216 1005793 415253 1005993
rect 426249 1005551 426299 1006551
rect 467797 1006498 468007 1006513
rect 470113 1006498 470323 1006513
rect 467812 1006328 467992 1006498
rect 470128 1006328 470308 1006498
rect 467801 1006325 468003 1006328
rect 470117 1006325 470319 1006328
rect 467797 1006313 468007 1006325
rect 470113 1006313 470323 1006325
rect 467201 1006238 467411 1006253
rect 467437 1006238 467647 1006253
rect 467797 1006238 468007 1006253
rect 468157 1006238 468217 1006253
rect 468243 1006238 468303 1006253
rect 469817 1006238 469877 1006253
rect 469903 1006238 469963 1006253
rect 470113 1006238 470323 1006253
rect 470473 1006238 470683 1006253
rect 470709 1006238 470919 1006253
rect 426893 1005542 426943 1006142
rect 427063 1005542 427119 1006142
rect 427239 1005542 427289 1006142
rect 427665 1005547 427715 1006147
rect 427835 1005547 427885 1006147
rect 466176 1005537 466226 1006137
rect 466326 1005537 466382 1006137
rect 466482 1005537 466532 1006137
rect 467216 1006068 467396 1006238
rect 467452 1006068 467632 1006238
rect 467812 1006068 467992 1006238
rect 468172 1006068 468202 1006238
rect 468258 1006068 468288 1006238
rect 467205 1006065 467407 1006068
rect 467441 1006065 467643 1006068
rect 467801 1006065 468003 1006068
rect 468161 1006065 468213 1006068
rect 468247 1006065 468299 1006068
rect 467201 1006053 467411 1006065
rect 467437 1006053 467647 1006065
rect 467797 1006053 468007 1006065
rect 468157 1006053 468217 1006065
rect 468243 1006053 468303 1006065
rect 467201 1005978 467411 1005993
rect 467437 1005978 467647 1005993
rect 467797 1005978 468007 1005993
rect 468157 1005978 468217 1005993
rect 468243 1005978 468303 1005993
rect 467216 1005808 467396 1005978
rect 467452 1005808 467632 1005978
rect 467812 1005808 467992 1005978
rect 468172 1005808 468202 1005978
rect 468258 1005808 468288 1005978
rect 467205 1005805 467407 1005808
rect 467441 1005805 467643 1005808
rect 467801 1005805 468003 1005808
rect 468161 1005805 468213 1005808
rect 468247 1005805 468299 1005808
rect 467201 1005793 467411 1005805
rect 467437 1005793 467647 1005805
rect 467797 1005793 468007 1005805
rect 468157 1005793 468217 1005805
rect 468243 1005793 468303 1005805
rect 468449 1005803 468465 1006119
rect 469653 1005803 469671 1006119
rect 469832 1006068 469862 1006238
rect 469918 1006068 469948 1006238
rect 470128 1006068 470308 1006238
rect 470488 1006068 470668 1006238
rect 470724 1006068 470904 1006238
rect 469821 1006065 469873 1006068
rect 469907 1006065 469959 1006068
rect 470117 1006065 470319 1006068
rect 470477 1006065 470679 1006068
rect 470713 1006065 470915 1006068
rect 469817 1006053 469877 1006065
rect 469903 1006053 469963 1006065
rect 470113 1006053 470323 1006065
rect 470473 1006053 470683 1006065
rect 470709 1006053 470919 1006065
rect 469817 1005978 469877 1005993
rect 469903 1005978 469963 1005993
rect 470113 1005978 470323 1005993
rect 470473 1005978 470683 1005993
rect 470709 1005978 470919 1005993
rect 469832 1005808 469862 1005978
rect 469918 1005808 469948 1005978
rect 470128 1005808 470308 1005978
rect 470488 1005808 470668 1005978
rect 470724 1005808 470904 1005978
rect 469821 1005805 469873 1005808
rect 469907 1005805 469959 1005808
rect 470117 1005805 470319 1005808
rect 470477 1005805 470679 1005808
rect 470713 1005805 470915 1005808
rect 468449 1005777 468453 1005803
rect 469817 1005793 469877 1005805
rect 469903 1005793 469963 1005805
rect 470113 1005793 470323 1005805
rect 470473 1005793 470683 1005805
rect 470709 1005793 470919 1005805
rect 467797 1005718 468007 1005733
rect 468157 1005718 468217 1005733
rect 468243 1005718 468303 1005733
rect 467812 1005548 467992 1005718
rect 468172 1005679 468202 1005718
rect 468258 1005679 468288 1005718
rect 467801 1005545 468003 1005548
rect 467797 1005533 468007 1005545
rect 468415 1005539 468453 1005777
rect 469673 1005539 469705 1005777
rect 469817 1005718 469877 1005733
rect 469903 1005718 469963 1005733
rect 470113 1005718 470323 1005733
rect 469832 1005679 469862 1005718
rect 469918 1005679 469948 1005718
rect 470128 1005548 470308 1005718
rect 470117 1005545 470319 1005548
rect 468415 1005513 468449 1005539
rect 470113 1005533 470323 1005545
rect 471588 1005537 471638 1006137
rect 471738 1005537 471794 1006137
rect 471894 1005537 471944 1006137
rect 472441 1005551 472491 1006551
rect 472591 1005551 472647 1006551
rect 472747 1005551 472797 1006551
rect 472883 1005551 472933 1006551
rect 473033 1005551 473089 1006551
rect 473189 1005551 473245 1006551
rect 473345 1005551 473401 1006551
rect 473501 1005551 473551 1006551
rect 473617 1005551 473667 1006551
rect 473767 1005551 473895 1006551
rect 473923 1005551 474051 1006551
rect 474079 1005551 474207 1006551
rect 474235 1005551 474363 1006551
rect 474391 1005551 474519 1006551
rect 474547 1005551 474603 1006551
rect 474703 1005551 474831 1006551
rect 474859 1005551 474987 1006551
rect 475015 1005551 475143 1006551
rect 475171 1005551 475299 1006551
rect 475327 1005551 475455 1006551
rect 475483 1005551 475539 1006551
rect 475659 1005551 475787 1006551
rect 475835 1005551 475963 1006551
rect 476011 1005551 476139 1006551
rect 476187 1005551 476315 1006551
rect 476363 1005551 476491 1006551
rect 476539 1005551 476667 1006551
rect 476715 1005551 476843 1006551
rect 476891 1005551 476941 1006551
rect 477007 1005551 477057 1006551
rect 477157 1005551 477285 1006551
rect 477313 1005551 477441 1006551
rect 477469 1005551 477597 1006551
rect 477625 1005551 477681 1006551
rect 477781 1005551 477909 1006551
rect 477937 1005551 478065 1006551
rect 478093 1005551 478221 1006551
rect 478249 1005551 478299 1006551
rect 478890 1005992 478943 1006142
rect 478893 1005895 478943 1005992
rect 478890 1005673 478943 1005895
rect 478893 1005542 478943 1005673
rect 479063 1005542 479119 1006142
rect 479239 1005542 479289 1006142
rect 479665 1005547 479715 1006147
rect 479835 1005547 479885 1006147
rect 518176 1005537 518226 1006137
rect 518326 1005537 518382 1006137
rect 518482 1005537 518532 1006137
rect 519216 1006053 519253 1006253
rect 519216 1005793 519253 1005993
rect 530249 1005551 530299 1006551
rect 571797 1006498 572007 1006513
rect 574113 1006498 574323 1006513
rect 571812 1006328 571992 1006498
rect 574128 1006328 574308 1006498
rect 571801 1006325 572003 1006328
rect 574117 1006325 574319 1006328
rect 571797 1006313 572007 1006325
rect 574113 1006313 574323 1006325
rect 571201 1006238 571411 1006253
rect 571437 1006238 571647 1006253
rect 571797 1006238 572007 1006253
rect 572157 1006238 572217 1006253
rect 572243 1006238 572303 1006253
rect 573817 1006238 573877 1006253
rect 573903 1006238 573963 1006253
rect 574113 1006238 574323 1006253
rect 574473 1006238 574683 1006253
rect 574709 1006238 574919 1006253
rect 530893 1005542 530943 1006142
rect 531063 1005542 531119 1006142
rect 531239 1005542 531289 1006142
rect 531665 1005547 531715 1006147
rect 531835 1005547 531885 1006147
rect 570176 1005537 570226 1006137
rect 570326 1005537 570382 1006137
rect 570482 1005537 570532 1006137
rect 571216 1006068 571396 1006238
rect 571452 1006068 571632 1006238
rect 571812 1006068 571992 1006238
rect 572172 1006068 572202 1006238
rect 572258 1006068 572288 1006238
rect 571205 1006065 571407 1006068
rect 571441 1006065 571643 1006068
rect 571801 1006065 572003 1006068
rect 572161 1006065 572213 1006068
rect 572247 1006065 572299 1006068
rect 571201 1006053 571411 1006065
rect 571437 1006053 571647 1006065
rect 571797 1006053 572007 1006065
rect 572157 1006053 572217 1006065
rect 572243 1006053 572303 1006065
rect 571201 1005978 571411 1005993
rect 571437 1005978 571647 1005993
rect 571797 1005978 572007 1005993
rect 572157 1005978 572217 1005993
rect 572243 1005978 572303 1005993
rect 571216 1005808 571396 1005978
rect 571452 1005808 571632 1005978
rect 571812 1005808 571992 1005978
rect 572172 1005808 572202 1005978
rect 572258 1005808 572288 1005978
rect 571205 1005805 571407 1005808
rect 571441 1005805 571643 1005808
rect 571801 1005805 572003 1005808
rect 572161 1005805 572213 1005808
rect 572247 1005805 572299 1005808
rect 571201 1005793 571411 1005805
rect 571437 1005793 571647 1005805
rect 571797 1005793 572007 1005805
rect 572157 1005793 572217 1005805
rect 572243 1005793 572303 1005805
rect 572449 1005803 572465 1006119
rect 573653 1005803 573671 1006119
rect 573832 1006068 573862 1006238
rect 573918 1006068 573948 1006238
rect 574128 1006068 574308 1006238
rect 574488 1006068 574668 1006238
rect 574724 1006068 574904 1006238
rect 573821 1006065 573873 1006068
rect 573907 1006065 573959 1006068
rect 574117 1006065 574319 1006068
rect 574477 1006065 574679 1006068
rect 574713 1006065 574915 1006068
rect 573817 1006053 573877 1006065
rect 573903 1006053 573963 1006065
rect 574113 1006053 574323 1006065
rect 574473 1006053 574683 1006065
rect 574709 1006053 574919 1006065
rect 573817 1005978 573877 1005993
rect 573903 1005978 573963 1005993
rect 574113 1005978 574323 1005993
rect 574473 1005978 574683 1005993
rect 574709 1005978 574919 1005993
rect 573832 1005808 573862 1005978
rect 573918 1005808 573948 1005978
rect 574128 1005808 574308 1005978
rect 574488 1005808 574668 1005978
rect 574724 1005808 574904 1005978
rect 573821 1005805 573873 1005808
rect 573907 1005805 573959 1005808
rect 574117 1005805 574319 1005808
rect 574477 1005805 574679 1005808
rect 574713 1005805 574915 1005808
rect 572449 1005777 572453 1005803
rect 573817 1005793 573877 1005805
rect 573903 1005793 573963 1005805
rect 574113 1005793 574323 1005805
rect 574473 1005793 574683 1005805
rect 574709 1005793 574919 1005805
rect 571797 1005718 572007 1005733
rect 572157 1005718 572217 1005733
rect 572243 1005718 572303 1005733
rect 571812 1005548 571992 1005718
rect 572172 1005679 572202 1005718
rect 572258 1005679 572288 1005718
rect 571801 1005545 572003 1005548
rect 571797 1005533 572007 1005545
rect 572415 1005539 572453 1005777
rect 573673 1005539 573705 1005777
rect 573817 1005718 573877 1005733
rect 573903 1005718 573963 1005733
rect 574113 1005718 574323 1005733
rect 573832 1005679 573862 1005718
rect 573918 1005679 573948 1005718
rect 574128 1005548 574308 1005718
rect 574117 1005545 574319 1005548
rect 572415 1005513 572449 1005539
rect 574113 1005533 574323 1005545
rect 575588 1005537 575638 1006137
rect 575738 1005537 575794 1006137
rect 575894 1005537 575944 1006137
rect 576441 1005551 576491 1006551
rect 576591 1005551 576647 1006551
rect 576747 1005551 576797 1006551
rect 576883 1005551 576933 1006551
rect 577033 1005551 577089 1006551
rect 577189 1005551 577245 1006551
rect 577345 1005551 577401 1006551
rect 577501 1005551 577551 1006551
rect 577617 1005551 577667 1006551
rect 577767 1005551 577895 1006551
rect 577923 1005551 578051 1006551
rect 578079 1005551 578207 1006551
rect 578235 1005551 578363 1006551
rect 578391 1005551 578519 1006551
rect 578547 1005551 578603 1006551
rect 578703 1005551 578831 1006551
rect 578859 1005551 578987 1006551
rect 579015 1005551 579143 1006551
rect 579171 1005551 579299 1006551
rect 579327 1005551 579455 1006551
rect 579483 1005551 579539 1006551
rect 579659 1005551 579787 1006551
rect 579835 1005551 579963 1006551
rect 580011 1005551 580139 1006551
rect 580187 1005551 580315 1006551
rect 580363 1005551 580491 1006551
rect 580539 1005551 580667 1006551
rect 580715 1005551 580843 1006551
rect 580891 1005551 580941 1006551
rect 581007 1005551 581057 1006551
rect 581157 1005551 581285 1006551
rect 581313 1005551 581441 1006551
rect 581469 1005551 581597 1006551
rect 581625 1005551 581681 1006551
rect 581781 1005551 581909 1006551
rect 581937 1005551 582065 1006551
rect 582093 1005551 582221 1006551
rect 582249 1005551 582299 1006551
rect 582890 1005992 582943 1006142
rect 582893 1005895 582943 1005992
rect 582890 1005673 582943 1005895
rect 582893 1005542 582943 1005673
rect 583063 1005542 583119 1006142
rect 583239 1005542 583289 1006142
rect 583665 1005547 583715 1006147
rect 583835 1005547 583885 1006147
rect 60893 1004565 60901 1004790
rect 60970 1003708 61020 1004308
rect 61120 1003708 61170 1004308
rect 62026 1004070 62076 1004670
rect 62176 1004070 62232 1004670
rect 62332 1004070 62382 1004670
rect 62554 1004004 62604 1005004
rect 62704 1004004 62760 1005004
rect 62860 1004004 62910 1005004
rect 62976 1004004 63026 1005004
rect 63126 1004004 63254 1005004
rect 63282 1004004 63410 1005004
rect 63438 1004004 63566 1005004
rect 63594 1004004 63650 1005004
rect 63750 1004004 63878 1005004
rect 63906 1004004 64034 1005004
rect 64062 1004004 64190 1005004
rect 64218 1004004 64268 1005004
rect 64420 1004004 64470 1005004
rect 64570 1004004 64698 1005004
rect 64726 1004004 64854 1005004
rect 64882 1004004 65010 1005004
rect 65038 1004004 65166 1005004
rect 65194 1004004 65322 1005004
rect 65350 1004004 65478 1005004
rect 65506 1004004 65634 1005004
rect 65662 1004004 65712 1005004
rect 65864 1004054 65914 1005054
rect 66014 1004054 66142 1005054
rect 66170 1004054 66298 1005054
rect 66326 1004054 66454 1005054
rect 66482 1004054 66610 1005054
rect 66638 1004054 66766 1005054
rect 66794 1004054 66922 1005054
rect 66950 1004054 67078 1005054
rect 67106 1004054 67156 1005054
rect 67308 1004004 67358 1005004
rect 67458 1004004 67586 1005004
rect 67614 1004004 67742 1005004
rect 67770 1004004 67898 1005004
rect 67926 1004004 68054 1005004
rect 68082 1004004 68210 1005004
rect 68238 1004004 68366 1005004
rect 68394 1004004 68522 1005004
rect 68550 1004004 68606 1005004
rect 68706 1004004 68756 1005004
rect 68908 1004404 68958 1005004
rect 69342 1004404 69392 1005004
rect 70585 1004519 70635 1005119
rect 70735 1004519 70863 1005119
rect 70891 1004519 71019 1005119
rect 71047 1004519 71097 1005119
rect 71177 1004519 71227 1005119
rect 71327 1004519 71455 1005119
rect 71483 1004519 71539 1005119
rect 71639 1004519 71767 1005119
rect 71795 1004519 71845 1005119
rect 71925 1004519 71975 1005119
rect 72075 1004519 72131 1005119
rect 72231 1004519 72281 1005119
rect 108893 1004565 108901 1004790
rect 71210 1003739 71246 1004339
rect 71570 1003739 71626 1004339
rect 71760 1003739 71810 1004339
rect 67473 1003625 67539 1003641
rect 67635 1003625 67701 1003641
rect 70043 1003571 70118 1003581
rect 70338 1003571 70413 1003581
rect 62326 1002921 62376 1003521
rect 62476 1002921 62532 1003521
rect 62632 1002921 62682 1003521
rect 62894 1002890 62944 1003490
rect 63044 1002890 63172 1003490
rect 63200 1002890 63328 1003490
rect 63356 1002890 63484 1003490
rect 63512 1002890 63562 1003490
rect 63628 1002890 63678 1003490
rect 63778 1002890 63906 1003490
rect 63934 1002890 64062 1003490
rect 64090 1002890 64218 1003490
rect 64246 1002890 64302 1003490
rect 64402 1002890 64530 1003490
rect 64558 1002890 64686 1003490
rect 64714 1002890 64842 1003490
rect 64870 1002890 64926 1003490
rect 65026 1002890 65082 1003490
rect 65182 1002890 65238 1003490
rect 65338 1002890 65388 1003490
rect 65454 1002890 65504 1003490
rect 65604 1002890 65732 1003490
rect 65760 1002890 65816 1003490
rect 65916 1002890 66044 1003490
rect 66072 1002890 66122 1003490
rect 69055 1003398 70055 1003448
rect 70118 1003398 70168 1003509
rect 70115 1003278 70168 1003398
rect 69055 1003228 70055 1003278
rect 69018 1002508 69068 1003108
rect 69188 1002508 69244 1003108
rect 69364 1002508 69414 1003108
rect 69634 1002509 69684 1003109
rect 69804 1002509 69860 1003109
rect 69980 1002509 70030 1003109
rect 70118 1002509 70168 1003278
rect 70288 1002509 70338 1003509
rect 70401 1003398 71001 1003448
rect 70401 1003298 70413 1003398
rect 72300 1003328 72350 1003928
rect 72470 1003328 72526 1003928
rect 72646 1003328 72774 1003928
rect 72822 1003328 72878 1003928
rect 72998 1003328 73054 1003928
rect 73174 1003328 73230 1003928
rect 73350 1003328 73478 1003928
rect 73526 1003328 73576 1003928
rect 108970 1003708 109020 1004308
rect 109120 1003708 109170 1004308
rect 110026 1004070 110076 1004670
rect 110176 1004070 110232 1004670
rect 110332 1004070 110382 1004670
rect 110554 1004004 110604 1005004
rect 110704 1004004 110760 1005004
rect 110860 1004004 110910 1005004
rect 110976 1004004 111026 1005004
rect 160893 1004565 160901 1004790
rect 160970 1003708 161020 1004308
rect 161120 1003708 161170 1004308
rect 162026 1004070 162076 1004670
rect 162176 1004070 162232 1004670
rect 162332 1004070 162382 1004670
rect 162554 1004004 162604 1005004
rect 162704 1004004 162760 1005004
rect 162860 1004004 162910 1005004
rect 162976 1004004 163026 1005004
rect 163126 1004004 163254 1005004
rect 163282 1004004 163410 1005004
rect 163438 1004004 163566 1005004
rect 163594 1004004 163650 1005004
rect 163750 1004004 163878 1005004
rect 163906 1004004 164034 1005004
rect 164062 1004004 164190 1005004
rect 164218 1004004 164268 1005004
rect 164420 1004004 164470 1005004
rect 164570 1004004 164698 1005004
rect 164726 1004004 164854 1005004
rect 164882 1004004 165010 1005004
rect 165038 1004004 165166 1005004
rect 165194 1004004 165322 1005004
rect 165350 1004004 165478 1005004
rect 165506 1004004 165634 1005004
rect 165662 1004004 165712 1005004
rect 165864 1004054 165914 1005054
rect 166014 1004054 166142 1005054
rect 166170 1004054 166298 1005054
rect 166326 1004054 166454 1005054
rect 166482 1004054 166610 1005054
rect 166638 1004054 166766 1005054
rect 166794 1004054 166922 1005054
rect 166950 1004054 167078 1005054
rect 167106 1004054 167156 1005054
rect 167308 1004004 167358 1005004
rect 167458 1004004 167586 1005004
rect 167614 1004004 167742 1005004
rect 167770 1004004 167898 1005004
rect 167926 1004004 168054 1005004
rect 168082 1004004 168210 1005004
rect 168238 1004004 168366 1005004
rect 168394 1004004 168522 1005004
rect 168550 1004004 168606 1005004
rect 168706 1004004 168756 1005004
rect 168908 1004404 168958 1005004
rect 169342 1004404 169392 1005004
rect 170585 1004519 170635 1005119
rect 170735 1004519 170863 1005119
rect 170891 1004519 171019 1005119
rect 171047 1004519 171097 1005119
rect 171177 1004519 171227 1005119
rect 171327 1004519 171455 1005119
rect 171483 1004519 171539 1005119
rect 171639 1004519 171767 1005119
rect 171795 1004519 171845 1005119
rect 171925 1004519 171975 1005119
rect 172075 1004519 172131 1005119
rect 172231 1004519 172281 1005119
rect 212893 1004565 212901 1004790
rect 171210 1003739 171246 1004339
rect 171570 1003739 171626 1004339
rect 171760 1003739 171810 1004339
rect 167473 1003625 167539 1003641
rect 167635 1003625 167701 1003641
rect 170043 1003571 170118 1003581
rect 170338 1003571 170413 1003581
rect 70401 1003248 71001 1003298
rect 70417 1002509 70467 1003109
rect 70587 1002509 70643 1003109
rect 70763 1002509 70813 1003109
rect 71104 1002509 71154 1003109
rect 71274 1002509 71402 1003109
rect 71450 1002509 71506 1003109
rect 71626 1002509 71754 1003109
rect 71802 1002509 71852 1003109
rect 72224 1002573 72274 1003173
rect 72394 1002573 72522 1003173
rect 72570 1002573 72698 1003173
rect 72746 1002573 72874 1003173
rect 72922 1002573 73050 1003173
rect 73098 1002573 73154 1003173
rect 73274 1002573 73402 1003173
rect 73450 1002573 73500 1003173
rect 110326 1002921 110376 1003521
rect 110476 1002921 110532 1003521
rect 110632 1002921 110682 1003521
rect 110894 1002890 110944 1003490
rect 162326 1002921 162376 1003521
rect 162476 1002921 162532 1003521
rect 162632 1002921 162682 1003521
rect 162894 1002890 162944 1003490
rect 163044 1002890 163172 1003490
rect 163200 1002890 163328 1003490
rect 163356 1002890 163484 1003490
rect 163512 1002890 163562 1003490
rect 163628 1002890 163678 1003490
rect 163778 1002890 163906 1003490
rect 163934 1002890 164062 1003490
rect 164090 1002890 164218 1003490
rect 164246 1002890 164302 1003490
rect 164402 1002890 164530 1003490
rect 164558 1002890 164686 1003490
rect 164714 1002890 164842 1003490
rect 164870 1002890 164926 1003490
rect 165026 1002890 165082 1003490
rect 165182 1002890 165238 1003490
rect 165338 1002890 165388 1003490
rect 165454 1002890 165504 1003490
rect 165604 1002890 165732 1003490
rect 165760 1002890 165816 1003490
rect 165916 1002890 166044 1003490
rect 166072 1002890 166122 1003490
rect 169055 1003398 170055 1003448
rect 170118 1003398 170168 1003509
rect 170115 1003278 170168 1003398
rect 169055 1003228 170055 1003278
rect 169018 1002508 169068 1003108
rect 169188 1002508 169244 1003108
rect 169364 1002508 169414 1003108
rect 169634 1002509 169684 1003109
rect 169804 1002509 169860 1003109
rect 169980 1002509 170030 1003109
rect 170118 1002509 170168 1003278
rect 170288 1002509 170338 1003509
rect 170401 1003398 171001 1003448
rect 170401 1003298 170413 1003398
rect 172300 1003328 172350 1003928
rect 172470 1003328 172526 1003928
rect 172646 1003328 172774 1003928
rect 172822 1003328 172878 1003928
rect 172998 1003328 173054 1003928
rect 173174 1003328 173230 1003928
rect 173350 1003328 173478 1003928
rect 173526 1003328 173576 1003928
rect 212970 1003708 213020 1004308
rect 213120 1003708 213170 1004308
rect 214026 1004070 214076 1004670
rect 214176 1004070 214232 1004670
rect 214332 1004070 214382 1004670
rect 214554 1004004 214604 1005004
rect 214704 1004004 214760 1005004
rect 214860 1004004 214910 1005004
rect 214976 1004004 215026 1005004
rect 260893 1004565 260901 1004790
rect 260970 1003708 261020 1004308
rect 261120 1003708 261170 1004308
rect 262026 1004070 262076 1004670
rect 312893 1004565 312901 1004790
rect 312970 1003708 313020 1004308
rect 313120 1003708 313170 1004308
rect 314026 1004070 314076 1004670
rect 314176 1004070 314232 1004670
rect 314332 1004070 314382 1004670
rect 314554 1004004 314604 1005004
rect 314704 1004004 314760 1005004
rect 314860 1004004 314910 1005004
rect 314976 1004004 315026 1005004
rect 364893 1004565 364901 1004790
rect 364970 1003708 365020 1004308
rect 365120 1003708 365170 1004308
rect 366026 1004070 366076 1004670
rect 366176 1004070 366232 1004670
rect 366332 1004070 366382 1004670
rect 366554 1004004 366604 1005004
rect 366704 1004004 366760 1005004
rect 366860 1004004 366910 1005004
rect 366976 1004004 367026 1005004
rect 367126 1004004 367254 1005004
rect 367282 1004004 367410 1005004
rect 367438 1004004 367566 1005004
rect 367594 1004004 367650 1005004
rect 367750 1004004 367878 1005004
rect 367906 1004004 368034 1005004
rect 368062 1004004 368190 1005004
rect 368218 1004004 368268 1005004
rect 368420 1004004 368470 1005004
rect 368570 1004004 368698 1005004
rect 368726 1004004 368854 1005004
rect 368882 1004004 369010 1005004
rect 369038 1004004 369166 1005004
rect 369194 1004004 369322 1005004
rect 369350 1004004 369478 1005004
rect 369506 1004004 369634 1005004
rect 369662 1004004 369712 1005004
rect 369864 1004054 369914 1005054
rect 370014 1004054 370142 1005054
rect 370170 1004054 370298 1005054
rect 370326 1004054 370454 1005054
rect 370482 1004054 370610 1005054
rect 370638 1004054 370766 1005054
rect 370794 1004054 370922 1005054
rect 370950 1004054 371078 1005054
rect 371106 1004054 371156 1005054
rect 371308 1004004 371358 1005004
rect 371458 1004004 371586 1005004
rect 371614 1004004 371742 1005004
rect 371770 1004004 371898 1005004
rect 371926 1004004 372054 1005004
rect 372082 1004004 372210 1005004
rect 372238 1004004 372366 1005004
rect 372394 1004004 372522 1005004
rect 372550 1004004 372606 1005004
rect 372706 1004004 372756 1005004
rect 372908 1004404 372958 1005004
rect 373342 1004404 373392 1005004
rect 374585 1004519 374635 1005119
rect 374735 1004519 374863 1005119
rect 374891 1004519 375019 1005119
rect 375047 1004519 375097 1005119
rect 375177 1004519 375227 1005119
rect 375327 1004519 375455 1005119
rect 375483 1004519 375539 1005119
rect 375639 1004519 375767 1005119
rect 375795 1004519 375845 1005119
rect 375925 1004519 375975 1005119
rect 376075 1004519 376131 1005119
rect 376231 1004519 376281 1005119
rect 412893 1004565 412901 1004790
rect 375210 1003739 375246 1004339
rect 375570 1003739 375626 1004339
rect 375760 1003739 375810 1004339
rect 371473 1003625 371539 1003641
rect 371635 1003625 371701 1003641
rect 374043 1003571 374118 1003581
rect 374338 1003571 374413 1003581
rect 170401 1003248 171001 1003298
rect 170417 1002509 170467 1003109
rect 170587 1002509 170643 1003109
rect 170763 1002509 170813 1003109
rect 171104 1002509 171154 1003109
rect 171274 1002509 171402 1003109
rect 171450 1002509 171506 1003109
rect 171626 1002509 171754 1003109
rect 171802 1002509 171852 1003109
rect 172224 1002573 172274 1003173
rect 172394 1002573 172522 1003173
rect 172570 1002573 172698 1003173
rect 172746 1002573 172874 1003173
rect 172922 1002573 173050 1003173
rect 173098 1002573 173154 1003173
rect 173274 1002573 173402 1003173
rect 173450 1002573 173500 1003173
rect 214326 1002921 214376 1003521
rect 214476 1002921 214532 1003521
rect 214632 1002921 214682 1003521
rect 214894 1002890 214944 1003490
rect 314326 1002921 314376 1003521
rect 314476 1002921 314532 1003521
rect 314632 1002921 314682 1003521
rect 314894 1002890 314944 1003490
rect 366326 1002921 366376 1003521
rect 366476 1002921 366532 1003521
rect 366632 1002921 366682 1003521
rect 366894 1002890 366944 1003490
rect 367044 1002890 367172 1003490
rect 367200 1002890 367328 1003490
rect 367356 1002890 367484 1003490
rect 367512 1002890 367562 1003490
rect 367628 1002890 367678 1003490
rect 367778 1002890 367906 1003490
rect 367934 1002890 368062 1003490
rect 368090 1002890 368218 1003490
rect 368246 1002890 368302 1003490
rect 368402 1002890 368530 1003490
rect 368558 1002890 368686 1003490
rect 368714 1002890 368842 1003490
rect 368870 1002890 368926 1003490
rect 369026 1002890 369082 1003490
rect 369182 1002890 369238 1003490
rect 369338 1002890 369388 1003490
rect 369454 1002890 369504 1003490
rect 369604 1002890 369732 1003490
rect 369760 1002890 369816 1003490
rect 369916 1002890 370044 1003490
rect 370072 1002890 370122 1003490
rect 373055 1003398 374055 1003448
rect 374118 1003398 374168 1003509
rect 374115 1003278 374168 1003398
rect 373055 1003228 374055 1003278
rect 373018 1002508 373068 1003108
rect 373188 1002508 373244 1003108
rect 373364 1002508 373414 1003108
rect 373634 1002509 373684 1003109
rect 373804 1002509 373860 1003109
rect 373980 1002509 374030 1003109
rect 374118 1002509 374168 1003278
rect 374288 1002509 374338 1003509
rect 374401 1003398 375001 1003448
rect 374401 1003298 374413 1003398
rect 376300 1003328 376350 1003928
rect 376470 1003328 376526 1003928
rect 376646 1003328 376774 1003928
rect 376822 1003328 376878 1003928
rect 376998 1003328 377054 1003928
rect 377174 1003328 377230 1003928
rect 377350 1003328 377478 1003928
rect 377526 1003328 377576 1003928
rect 412970 1003708 413020 1004308
rect 413120 1003708 413170 1004308
rect 414026 1004070 414076 1004670
rect 414176 1004070 414232 1004670
rect 414332 1004070 414382 1004670
rect 414554 1004004 414604 1005004
rect 414704 1004004 414760 1005004
rect 414860 1004004 414910 1005004
rect 414976 1004004 415026 1005004
rect 464893 1004565 464901 1004790
rect 464970 1003708 465020 1004308
rect 465120 1003708 465170 1004308
rect 466026 1004070 466076 1004670
rect 466176 1004070 466232 1004670
rect 466332 1004070 466382 1004670
rect 466554 1004004 466604 1005004
rect 466704 1004004 466760 1005004
rect 466860 1004004 466910 1005004
rect 466976 1004004 467026 1005004
rect 467126 1004004 467254 1005004
rect 467282 1004004 467410 1005004
rect 467438 1004004 467566 1005004
rect 467594 1004004 467650 1005004
rect 467750 1004004 467878 1005004
rect 467906 1004004 468034 1005004
rect 468062 1004004 468190 1005004
rect 468218 1004004 468268 1005004
rect 468420 1004004 468470 1005004
rect 468570 1004004 468698 1005004
rect 468726 1004004 468854 1005004
rect 468882 1004004 469010 1005004
rect 469038 1004004 469166 1005004
rect 469194 1004004 469322 1005004
rect 469350 1004004 469478 1005004
rect 469506 1004004 469634 1005004
rect 469662 1004004 469712 1005004
rect 469864 1004054 469914 1005054
rect 470014 1004054 470142 1005054
rect 470170 1004054 470298 1005054
rect 470326 1004054 470454 1005054
rect 470482 1004054 470610 1005054
rect 470638 1004054 470766 1005054
rect 470794 1004054 470922 1005054
rect 470950 1004054 471078 1005054
rect 471106 1004054 471156 1005054
rect 471308 1004004 471358 1005004
rect 471458 1004004 471586 1005004
rect 471614 1004004 471742 1005004
rect 471770 1004004 471898 1005004
rect 471926 1004004 472054 1005004
rect 472082 1004004 472210 1005004
rect 472238 1004004 472366 1005004
rect 472394 1004004 472522 1005004
rect 472550 1004004 472606 1005004
rect 472706 1004004 472756 1005004
rect 472908 1004404 472958 1005004
rect 473342 1004404 473392 1005004
rect 474585 1004519 474635 1005119
rect 474735 1004519 474863 1005119
rect 474891 1004519 475019 1005119
rect 475047 1004519 475097 1005119
rect 475177 1004519 475227 1005119
rect 475327 1004519 475455 1005119
rect 475483 1004519 475539 1005119
rect 475639 1004519 475767 1005119
rect 475795 1004519 475845 1005119
rect 475925 1004519 475975 1005119
rect 476075 1004519 476131 1005119
rect 476231 1004519 476281 1005119
rect 516893 1004565 516901 1004790
rect 475210 1003739 475246 1004339
rect 475570 1003739 475626 1004339
rect 475760 1003739 475810 1004339
rect 471473 1003625 471539 1003641
rect 471635 1003625 471701 1003641
rect 474043 1003571 474118 1003581
rect 474338 1003571 474413 1003581
rect 374401 1003248 375001 1003298
rect 374417 1002509 374467 1003109
rect 374587 1002509 374643 1003109
rect 374763 1002509 374813 1003109
rect 375104 1002509 375154 1003109
rect 375274 1002509 375402 1003109
rect 375450 1002509 375506 1003109
rect 375626 1002509 375754 1003109
rect 375802 1002509 375852 1003109
rect 376224 1002573 376274 1003173
rect 376394 1002573 376522 1003173
rect 376570 1002573 376698 1003173
rect 376746 1002573 376874 1003173
rect 376922 1002573 377050 1003173
rect 377098 1002573 377154 1003173
rect 377274 1002573 377402 1003173
rect 377450 1002573 377500 1003173
rect 414326 1002921 414376 1003521
rect 414476 1002921 414532 1003521
rect 414632 1002921 414682 1003521
rect 414894 1002890 414944 1003490
rect 466326 1002921 466376 1003521
rect 466476 1002921 466532 1003521
rect 466632 1002921 466682 1003521
rect 466894 1002890 466944 1003490
rect 467044 1002890 467172 1003490
rect 467200 1002890 467328 1003490
rect 467356 1002890 467484 1003490
rect 467512 1002890 467562 1003490
rect 467628 1002890 467678 1003490
rect 467778 1002890 467906 1003490
rect 467934 1002890 468062 1003490
rect 468090 1002890 468218 1003490
rect 468246 1002890 468302 1003490
rect 468402 1002890 468530 1003490
rect 468558 1002890 468686 1003490
rect 468714 1002890 468842 1003490
rect 468870 1002890 468926 1003490
rect 469026 1002890 469082 1003490
rect 469182 1002890 469238 1003490
rect 469338 1002890 469388 1003490
rect 469454 1002890 469504 1003490
rect 469604 1002890 469732 1003490
rect 469760 1002890 469816 1003490
rect 469916 1002890 470044 1003490
rect 470072 1002890 470122 1003490
rect 473055 1003398 474055 1003448
rect 474118 1003398 474168 1003509
rect 474115 1003278 474168 1003398
rect 473055 1003228 474055 1003278
rect 473018 1002508 473068 1003108
rect 473188 1002508 473244 1003108
rect 473364 1002508 473414 1003108
rect 473634 1002509 473684 1003109
rect 473804 1002509 473860 1003109
rect 473980 1002509 474030 1003109
rect 474118 1002509 474168 1003278
rect 474288 1002509 474338 1003509
rect 474401 1003398 475001 1003448
rect 474401 1003298 474413 1003398
rect 476300 1003328 476350 1003928
rect 476470 1003328 476526 1003928
rect 476646 1003328 476774 1003928
rect 476822 1003328 476878 1003928
rect 476998 1003328 477054 1003928
rect 477174 1003328 477230 1003928
rect 477350 1003328 477478 1003928
rect 477526 1003328 477576 1003928
rect 516970 1003708 517020 1004308
rect 517120 1003708 517170 1004308
rect 518026 1004070 518076 1004670
rect 518176 1004070 518232 1004670
rect 518332 1004070 518382 1004670
rect 518554 1004004 518604 1005004
rect 518704 1004004 518760 1005004
rect 518860 1004004 518910 1005004
rect 518976 1004004 519026 1005004
rect 568893 1004565 568901 1004790
rect 568970 1003708 569020 1004308
rect 569120 1003708 569170 1004308
rect 570026 1004070 570076 1004670
rect 570176 1004070 570232 1004670
rect 570332 1004070 570382 1004670
rect 570554 1004004 570604 1005004
rect 570704 1004004 570760 1005004
rect 570860 1004004 570910 1005004
rect 570976 1004004 571026 1005004
rect 571126 1004004 571254 1005004
rect 571282 1004004 571410 1005004
rect 571438 1004004 571566 1005004
rect 571594 1004004 571650 1005004
rect 571750 1004004 571878 1005004
rect 571906 1004004 572034 1005004
rect 572062 1004004 572190 1005004
rect 572218 1004004 572268 1005004
rect 572420 1004004 572470 1005004
rect 572570 1004004 572698 1005004
rect 572726 1004004 572854 1005004
rect 572882 1004004 573010 1005004
rect 573038 1004004 573166 1005004
rect 573194 1004004 573322 1005004
rect 573350 1004004 573478 1005004
rect 573506 1004004 573634 1005004
rect 573662 1004004 573712 1005004
rect 573864 1004054 573914 1005054
rect 574014 1004054 574142 1005054
rect 574170 1004054 574298 1005054
rect 574326 1004054 574454 1005054
rect 574482 1004054 574610 1005054
rect 574638 1004054 574766 1005054
rect 574794 1004054 574922 1005054
rect 574950 1004054 575078 1005054
rect 575106 1004054 575156 1005054
rect 575308 1004004 575358 1005004
rect 575458 1004004 575586 1005004
rect 575614 1004004 575742 1005004
rect 575770 1004004 575898 1005004
rect 575926 1004004 576054 1005004
rect 576082 1004004 576210 1005004
rect 576238 1004004 576366 1005004
rect 576394 1004004 576522 1005004
rect 576550 1004004 576606 1005004
rect 576706 1004004 576756 1005004
rect 576908 1004404 576958 1005004
rect 577342 1004404 577392 1005004
rect 578585 1004519 578635 1005119
rect 578735 1004519 578863 1005119
rect 578891 1004519 579019 1005119
rect 579047 1004519 579097 1005119
rect 579177 1004519 579227 1005119
rect 579327 1004519 579455 1005119
rect 579483 1004519 579539 1005119
rect 579639 1004519 579767 1005119
rect 579795 1004519 579845 1005119
rect 579925 1004519 579975 1005119
rect 580075 1004519 580131 1005119
rect 580231 1004519 580281 1005119
rect 579210 1003739 579246 1004339
rect 579570 1003739 579626 1004339
rect 579760 1003739 579810 1004339
rect 575473 1003625 575539 1003641
rect 575635 1003625 575701 1003641
rect 578043 1003571 578118 1003581
rect 578338 1003571 578413 1003581
rect 474401 1003248 475001 1003298
rect 474417 1002509 474467 1003109
rect 474587 1002509 474643 1003109
rect 474763 1002509 474813 1003109
rect 475104 1002509 475154 1003109
rect 475274 1002509 475402 1003109
rect 475450 1002509 475506 1003109
rect 475626 1002509 475754 1003109
rect 475802 1002509 475852 1003109
rect 476224 1002573 476274 1003173
rect 476394 1002573 476522 1003173
rect 476570 1002573 476698 1003173
rect 476746 1002573 476874 1003173
rect 476922 1002573 477050 1003173
rect 477098 1002573 477154 1003173
rect 477274 1002573 477402 1003173
rect 477450 1002573 477500 1003173
rect 518326 1002921 518376 1003521
rect 518476 1002921 518532 1003521
rect 518632 1002921 518682 1003521
rect 518894 1002890 518944 1003490
rect 570326 1002921 570376 1003521
rect 570476 1002921 570532 1003521
rect 570632 1002921 570682 1003521
rect 570894 1002890 570944 1003490
rect 571044 1002890 571172 1003490
rect 571200 1002890 571328 1003490
rect 571356 1002890 571484 1003490
rect 571512 1002890 571562 1003490
rect 571628 1002890 571678 1003490
rect 571778 1002890 571906 1003490
rect 571934 1002890 572062 1003490
rect 572090 1002890 572218 1003490
rect 572246 1002890 572302 1003490
rect 572402 1002890 572530 1003490
rect 572558 1002890 572686 1003490
rect 572714 1002890 572842 1003490
rect 572870 1002890 572926 1003490
rect 573026 1002890 573082 1003490
rect 573182 1002890 573238 1003490
rect 573338 1002890 573388 1003490
rect 573454 1002890 573504 1003490
rect 573604 1002890 573732 1003490
rect 573760 1002890 573816 1003490
rect 573916 1002890 574044 1003490
rect 574072 1002890 574122 1003490
rect 577055 1003398 578055 1003448
rect 578118 1003398 578168 1003509
rect 578115 1003278 578168 1003398
rect 577055 1003228 578055 1003278
rect 577018 1002508 577068 1003108
rect 577188 1002508 577244 1003108
rect 577364 1002508 577414 1003108
rect 577634 1002509 577684 1003109
rect 577804 1002509 577860 1003109
rect 577980 1002509 578030 1003109
rect 578118 1002509 578168 1003278
rect 578288 1002509 578338 1003509
rect 578401 1003398 579001 1003448
rect 578401 1003298 578413 1003398
rect 580300 1003328 580350 1003928
rect 580470 1003328 580526 1003928
rect 580646 1003328 580774 1003928
rect 580822 1003328 580878 1003928
rect 580998 1003328 581054 1003928
rect 581174 1003328 581230 1003928
rect 581350 1003328 581478 1003928
rect 581526 1003328 581576 1003928
rect 578401 1003248 579001 1003298
rect 578417 1002509 578467 1003109
rect 578587 1002509 578643 1003109
rect 578763 1002509 578813 1003109
rect 579104 1002509 579154 1003109
rect 579274 1002509 579402 1003109
rect 579450 1002509 579506 1003109
rect 579626 1002509 579754 1003109
rect 579802 1002509 579852 1003109
rect 580224 1002573 580274 1003173
rect 580394 1002573 580522 1003173
rect 580570 1002573 580698 1003173
rect 580746 1002573 580874 1003173
rect 580922 1002573 581050 1003173
rect 581098 1002573 581154 1003173
rect 581274 1002573 581402 1003173
rect 581450 1002573 581500 1003173
rect 64901 1002385 64951 1002466
rect 61234 1002054 61249 1002069
rect 61198 1002024 61249 1002054
rect 61234 1002009 61249 1002024
rect 62092 1001713 62142 1002313
rect 62262 1001713 62390 1002313
rect 62438 1001713 62494 1002313
rect 62614 1001884 62664 1002313
rect 62727 1002113 62739 1002313
rect 64898 1002113 64951 1002385
rect 62614 1001812 62667 1001884
rect 64901 1001866 64951 1002113
rect 65051 1001866 65101 1002466
rect 65167 1001866 65217 1002466
rect 65317 1001866 65445 1002466
rect 65473 1001866 65601 1002466
rect 65629 1001866 65757 1002466
rect 65835 1001866 65888 1002466
rect 62614 1001713 62664 1001812
rect 62727 1001713 62739 1001812
rect 65238 1001502 65728 1001529
rect 65838 1001466 65888 1001866
rect 65988 1001466 66116 1002466
rect 66144 1001466 66194 1002466
rect 164901 1002385 164951 1002466
rect 31303 1001420 31428 1001422
rect 66395 1001345 66407 1002345
rect 66464 1001345 66514 1002345
rect 66634 1001345 66762 1002345
rect 66810 1001345 66938 1002345
rect 66986 1001345 67042 1002345
rect 67162 1001345 67212 1002345
rect 67311 1002225 67377 1002241
rect 67797 1002225 67863 1002241
rect 67311 1001441 67377 1001457
rect 67473 1001441 67539 1001457
rect 67635 1001441 67701 1001457
rect 67797 1001441 67863 1001457
rect 67962 1001345 68012 1002345
rect 68132 1001345 68188 1002345
rect 68308 1001345 68436 1002345
rect 68484 1001345 68612 1002345
rect 68660 1001345 68710 1002345
rect 68767 1001345 68779 1002345
rect 68803 1002281 68813 1002315
rect 68803 1002213 68813 1002247
rect 68803 1002145 68813 1002179
rect 68803 1002077 68813 1002111
rect 68803 1002002 68813 1002036
rect 68803 1001934 68813 1001968
rect 68803 1001866 68813 1001900
rect 68803 1001798 68813 1001832
rect 68803 1001730 68813 1001764
rect 68803 1001662 68813 1001696
rect 68803 1001594 68813 1001628
rect 68803 1001526 68813 1001560
rect 68803 1001458 68813 1001492
rect 68803 1001390 68813 1001424
rect 68862 1001345 68912 1002345
rect 69032 1001345 69160 1002345
rect 69208 1001345 69264 1002345
rect 69384 1001345 69434 1002345
rect 69600 1001745 69650 1002345
rect 69770 1001745 69826 1002345
rect 69946 1001745 70074 1002345
rect 70122 1001745 70172 1002345
rect 70324 1001745 70374 1002345
rect 70474 1001745 70602 1002345
rect 70630 1001745 70686 1002345
rect 70786 1001745 70914 1002345
rect 70942 1001745 70992 1002345
rect 71196 1001745 71246 1002345
rect 71346 1001745 71474 1002345
rect 71502 1001745 71630 1002345
rect 71658 1001745 71714 1002345
rect 71814 1001745 71864 1002345
rect 109234 1002054 109249 1002069
rect 109198 1002024 109249 1002054
rect 109234 1002009 109249 1002024
rect 110092 1001713 110142 1002313
rect 110438 1001713 110494 1002313
rect 110614 1001713 110664 1002313
rect 161234 1002054 161249 1002069
rect 161198 1002024 161249 1002054
rect 161234 1002009 161249 1002024
rect 162092 1001713 162142 1002313
rect 162262 1001713 162390 1002313
rect 162438 1001713 162494 1002313
rect 162614 1001884 162664 1002313
rect 162727 1002113 162739 1002313
rect 164898 1002113 164951 1002385
rect 162614 1001812 162667 1001884
rect 164901 1001866 164951 1002113
rect 165051 1001866 165101 1002466
rect 165167 1001866 165217 1002466
rect 165317 1001866 165445 1002466
rect 165473 1001866 165601 1002466
rect 165629 1001866 165757 1002466
rect 165835 1001866 165888 1002466
rect 162614 1001713 162664 1001812
rect 162727 1001713 162739 1001812
rect 165238 1001502 165728 1001529
rect 165838 1001466 165888 1001866
rect 165988 1001466 166116 1002466
rect 166144 1001466 166194 1002466
rect 368901 1002385 368951 1002466
rect 166395 1001345 166407 1002345
rect 166464 1001345 166514 1002345
rect 166634 1001345 166762 1002345
rect 166810 1001345 166938 1002345
rect 166986 1001345 167042 1002345
rect 167162 1001345 167212 1002345
rect 167311 1002225 167377 1002241
rect 167797 1002225 167863 1002241
rect 167311 1001441 167377 1001457
rect 167473 1001441 167539 1001457
rect 167635 1001441 167701 1001457
rect 167797 1001441 167863 1001457
rect 167962 1001345 168012 1002345
rect 168132 1001345 168188 1002345
rect 168308 1001345 168436 1002345
rect 168484 1001345 168612 1002345
rect 168660 1001345 168710 1002345
rect 168767 1001345 168779 1002345
rect 168803 1002281 168813 1002315
rect 168803 1002213 168813 1002247
rect 168803 1002145 168813 1002179
rect 168803 1002077 168813 1002111
rect 168803 1002002 168813 1002036
rect 168803 1001934 168813 1001968
rect 168803 1001866 168813 1001900
rect 168803 1001798 168813 1001832
rect 168803 1001730 168813 1001764
rect 168803 1001662 168813 1001696
rect 168803 1001594 168813 1001628
rect 168803 1001526 168813 1001560
rect 168803 1001458 168813 1001492
rect 168803 1001390 168813 1001424
rect 168862 1001345 168912 1002345
rect 169032 1001345 169160 1002345
rect 169208 1001345 169264 1002345
rect 169384 1001345 169434 1002345
rect 169600 1001745 169650 1002345
rect 169770 1001745 169826 1002345
rect 169946 1001745 170074 1002345
rect 170122 1001745 170172 1002345
rect 170324 1001745 170374 1002345
rect 170474 1001745 170602 1002345
rect 170630 1001745 170686 1002345
rect 170786 1001745 170914 1002345
rect 170942 1001745 170992 1002345
rect 171196 1001745 171246 1002345
rect 171346 1001745 171474 1002345
rect 171502 1001745 171630 1002345
rect 171658 1001745 171714 1002345
rect 171814 1001745 171864 1002345
rect 213234 1002054 213249 1002069
rect 213198 1002024 213249 1002054
rect 213234 1002009 213249 1002024
rect 214092 1001713 214142 1002313
rect 214438 1001713 214494 1002313
rect 214614 1001713 214664 1002313
rect 261234 1002054 261249 1002069
rect 313234 1002054 313249 1002069
rect 261198 1002024 261249 1002054
rect 313198 1002024 313249 1002054
rect 261234 1002009 261249 1002024
rect 313234 1002009 313249 1002024
rect 314092 1001713 314142 1002313
rect 314438 1001713 314494 1002313
rect 314614 1001713 314664 1002313
rect 365234 1002054 365249 1002069
rect 365198 1002024 365249 1002054
rect 365234 1002009 365249 1002024
rect 366092 1001713 366142 1002313
rect 366262 1001713 366390 1002313
rect 366438 1001713 366494 1002313
rect 366614 1001884 366664 1002313
rect 366727 1002113 366739 1002313
rect 368898 1002113 368951 1002385
rect 366614 1001812 366667 1001884
rect 368901 1001866 368951 1002113
rect 369051 1001866 369101 1002466
rect 369167 1001866 369217 1002466
rect 369317 1001866 369445 1002466
rect 369473 1001866 369601 1002466
rect 369629 1001866 369757 1002466
rect 369835 1001866 369888 1002466
rect 366614 1001713 366664 1001812
rect 366727 1001713 366739 1001812
rect 369238 1001502 369728 1001529
rect 369838 1001466 369888 1001866
rect 369988 1001466 370116 1002466
rect 370144 1001466 370194 1002466
rect 468901 1002385 468951 1002466
rect 370395 1001345 370407 1002345
rect 370464 1001345 370514 1002345
rect 370634 1001345 370762 1002345
rect 370810 1001345 370938 1002345
rect 370986 1001345 371042 1002345
rect 371162 1001345 371212 1002345
rect 371311 1002225 371377 1002241
rect 371797 1002225 371863 1002241
rect 371311 1001441 371377 1001457
rect 371473 1001441 371539 1001457
rect 371635 1001441 371701 1001457
rect 371797 1001441 371863 1001457
rect 371962 1001345 372012 1002345
rect 372132 1001345 372188 1002345
rect 372308 1001345 372436 1002345
rect 372484 1001345 372612 1002345
rect 372660 1001345 372710 1002345
rect 372767 1001345 372779 1002345
rect 372803 1002281 372813 1002315
rect 372803 1002213 372813 1002247
rect 372803 1002145 372813 1002179
rect 372803 1002077 372813 1002111
rect 372803 1002002 372813 1002036
rect 372803 1001934 372813 1001968
rect 372803 1001866 372813 1001900
rect 372803 1001798 372813 1001832
rect 372803 1001730 372813 1001764
rect 372803 1001662 372813 1001696
rect 372803 1001594 372813 1001628
rect 372803 1001526 372813 1001560
rect 372803 1001458 372813 1001492
rect 372803 1001390 372813 1001424
rect 372862 1001345 372912 1002345
rect 373032 1001345 373160 1002345
rect 373208 1001345 373264 1002345
rect 373384 1001345 373434 1002345
rect 373600 1001745 373650 1002345
rect 373770 1001745 373826 1002345
rect 373946 1001745 374074 1002345
rect 374122 1001745 374172 1002345
rect 374324 1001745 374374 1002345
rect 374474 1001745 374602 1002345
rect 374630 1001745 374686 1002345
rect 374786 1001745 374914 1002345
rect 374942 1001745 374992 1002345
rect 375196 1001745 375246 1002345
rect 375346 1001745 375474 1002345
rect 375502 1001745 375630 1002345
rect 375658 1001745 375714 1002345
rect 375814 1001745 375864 1002345
rect 413234 1002054 413249 1002069
rect 413198 1002024 413249 1002054
rect 413234 1002009 413249 1002024
rect 414092 1001713 414142 1002313
rect 414438 1001713 414494 1002313
rect 414614 1001713 414664 1002313
rect 465234 1002054 465249 1002069
rect 465198 1002024 465249 1002054
rect 465234 1002009 465249 1002024
rect 466092 1001713 466142 1002313
rect 466262 1001713 466390 1002313
rect 466438 1001713 466494 1002313
rect 466614 1001884 466664 1002313
rect 466727 1002113 466739 1002313
rect 468898 1002113 468951 1002385
rect 466614 1001812 466667 1001884
rect 468901 1001866 468951 1002113
rect 469051 1001866 469101 1002466
rect 469167 1001866 469217 1002466
rect 469317 1001866 469445 1002466
rect 469473 1001866 469601 1002466
rect 469629 1001866 469757 1002466
rect 469835 1001866 469888 1002466
rect 466614 1001713 466664 1001812
rect 466727 1001713 466739 1001812
rect 469238 1001502 469728 1001529
rect 469838 1001466 469888 1001866
rect 469988 1001466 470116 1002466
rect 470144 1001466 470194 1002466
rect 572901 1002385 572951 1002466
rect 470395 1001345 470407 1002345
rect 470464 1001345 470514 1002345
rect 470634 1001345 470762 1002345
rect 470810 1001345 470938 1002345
rect 470986 1001345 471042 1002345
rect 471162 1001345 471212 1002345
rect 471311 1002225 471377 1002241
rect 471797 1002225 471863 1002241
rect 471311 1001441 471377 1001457
rect 471473 1001441 471539 1001457
rect 471635 1001441 471701 1001457
rect 471797 1001441 471863 1001457
rect 471962 1001345 472012 1002345
rect 472132 1001345 472188 1002345
rect 472308 1001345 472436 1002345
rect 472484 1001345 472612 1002345
rect 472660 1001345 472710 1002345
rect 472767 1001345 472779 1002345
rect 472803 1002281 472813 1002315
rect 472803 1002213 472813 1002247
rect 472803 1002145 472813 1002179
rect 472803 1002077 472813 1002111
rect 472803 1002002 472813 1002036
rect 472803 1001934 472813 1001968
rect 472803 1001866 472813 1001900
rect 472803 1001798 472813 1001832
rect 472803 1001730 472813 1001764
rect 472803 1001662 472813 1001696
rect 472803 1001594 472813 1001628
rect 472803 1001526 472813 1001560
rect 472803 1001458 472813 1001492
rect 472803 1001390 472813 1001424
rect 472862 1001345 472912 1002345
rect 473032 1001345 473160 1002345
rect 473208 1001345 473264 1002345
rect 473384 1001345 473434 1002345
rect 473600 1001745 473650 1002345
rect 473770 1001745 473826 1002345
rect 473946 1001745 474074 1002345
rect 474122 1001745 474172 1002345
rect 474324 1001745 474374 1002345
rect 474474 1001745 474602 1002345
rect 474630 1001745 474686 1002345
rect 474786 1001745 474914 1002345
rect 474942 1001745 474992 1002345
rect 475196 1001745 475246 1002345
rect 475346 1001745 475474 1002345
rect 475502 1001745 475630 1002345
rect 475658 1001745 475714 1002345
rect 475814 1001745 475864 1002345
rect 517234 1002054 517249 1002069
rect 517198 1002024 517249 1002054
rect 517234 1002009 517249 1002024
rect 518092 1001713 518142 1002313
rect 518438 1001713 518494 1002313
rect 518614 1001713 518664 1002313
rect 569234 1002054 569249 1002069
rect 569198 1002024 569249 1002054
rect 569234 1002009 569249 1002024
rect 570092 1001713 570142 1002313
rect 570262 1001713 570390 1002313
rect 570438 1001713 570494 1002313
rect 570614 1001884 570664 1002313
rect 570727 1002113 570739 1002313
rect 572898 1002113 572951 1002385
rect 570614 1001812 570667 1001884
rect 572901 1001866 572951 1002113
rect 573051 1001866 573101 1002466
rect 573167 1001866 573217 1002466
rect 573317 1001866 573445 1002466
rect 573473 1001866 573601 1002466
rect 573629 1001866 573757 1002466
rect 573835 1001866 573888 1002466
rect 570614 1001713 570664 1001812
rect 570727 1001713 570739 1001812
rect 573238 1001502 573728 1001529
rect 573838 1001466 573888 1001866
rect 573988 1001466 574116 1002466
rect 574144 1001466 574194 1002466
rect 574395 1001345 574407 1002345
rect 574464 1001345 574514 1002345
rect 574634 1001345 574762 1002345
rect 574810 1001345 574938 1002345
rect 574986 1001345 575042 1002345
rect 575162 1001345 575212 1002345
rect 575311 1002225 575377 1002241
rect 575797 1002225 575863 1002241
rect 575311 1001441 575377 1001457
rect 575473 1001441 575539 1001457
rect 575635 1001441 575701 1001457
rect 575797 1001441 575863 1001457
rect 575962 1001345 576012 1002345
rect 576132 1001345 576188 1002345
rect 576308 1001345 576436 1002345
rect 576484 1001345 576612 1002345
rect 576660 1001345 576710 1002345
rect 576767 1001345 576779 1002345
rect 576803 1002281 576813 1002315
rect 576803 1002213 576813 1002247
rect 576803 1002145 576813 1002179
rect 576803 1002077 576813 1002111
rect 576803 1002002 576813 1002036
rect 576803 1001934 576813 1001968
rect 576803 1001866 576813 1001900
rect 576803 1001798 576813 1001832
rect 576803 1001730 576813 1001764
rect 576803 1001662 576813 1001696
rect 576803 1001594 576813 1001628
rect 576803 1001526 576813 1001560
rect 576803 1001458 576813 1001492
rect 576803 1001390 576813 1001424
rect 576862 1001345 576912 1002345
rect 577032 1001345 577160 1002345
rect 577208 1001345 577264 1002345
rect 577384 1001345 577434 1002345
rect 577600 1001745 577650 1002345
rect 577770 1001745 577826 1002345
rect 577946 1001745 578074 1002345
rect 578122 1001745 578172 1002345
rect 578324 1001745 578374 1002345
rect 578474 1001745 578602 1002345
rect 578630 1001745 578686 1002345
rect 578786 1001745 578914 1002345
rect 578942 1001745 578992 1002345
rect 579196 1001745 579246 1002345
rect 579346 1001745 579474 1002345
rect 579502 1001745 579630 1002345
rect 579658 1001745 579714 1002345
rect 579814 1001745 579864 1002345
rect 61264 1000665 61317 1000815
rect 61267 1000215 61317 1000665
rect 61437 1000215 61493 1000815
rect 61613 1000215 61669 1000815
rect 61789 1000215 61845 1000815
rect 61965 1000215 62015 1000815
rect 62081 1000215 62131 1000815
rect 62251 1000215 62307 1000815
rect 62427 1000215 62483 1000815
rect 62603 1000215 62653 1000815
rect 62909 1000803 63119 1000815
rect 63145 1000803 63355 1000815
rect 64879 1000803 65089 1000815
rect 65115 1000803 65325 1000815
rect 62913 1000800 63115 1000803
rect 63149 1000800 63351 1000803
rect 64883 1000800 65085 1000803
rect 65119 1000800 65321 1000803
rect 62924 1000630 63104 1000800
rect 63160 1000630 63340 1000800
rect 64894 1000630 65074 1000800
rect 65130 1000630 65310 1000800
rect 62909 1000615 63119 1000630
rect 63145 1000615 63355 1000630
rect 64879 1000615 65089 1000630
rect 65115 1000615 65325 1000630
rect 63145 1000502 63355 1000517
rect 64879 1000502 65089 1000517
rect 63160 1000480 63340 1000502
rect 64894 1000480 65074 1000502
rect 65581 1000215 65631 1000815
rect 65751 1000215 65807 1000815
rect 65927 1000215 65983 1000815
rect 66103 1000215 66153 1000815
rect 66235 1000215 66285 1000815
rect 66405 1000215 66461 1000815
rect 66581 1000215 66637 1000815
rect 66757 1000215 66807 1000815
rect 67063 1000803 67273 1000815
rect 67299 1000803 67509 1000815
rect 69033 1000803 69243 1000815
rect 69269 1000803 69479 1000815
rect 67067 1000800 67269 1000803
rect 67303 1000800 67505 1000803
rect 69037 1000800 69239 1000803
rect 69273 1000800 69475 1000803
rect 67078 1000630 67258 1000800
rect 67314 1000630 67494 1000800
rect 69048 1000630 69228 1000800
rect 69284 1000630 69464 1000800
rect 67063 1000615 67273 1000630
rect 67299 1000615 67509 1000630
rect 69033 1000615 69243 1000630
rect 69269 1000615 69479 1000630
rect 67299 1000502 67509 1000517
rect 69033 1000502 69243 1000517
rect 67314 1000480 67494 1000502
rect 69048 1000480 69228 1000502
rect 69735 1000215 69785 1000815
rect 69905 1000215 69961 1000815
rect 70081 1000215 70137 1000815
rect 70257 1000215 70307 1000815
rect 70389 1000215 70439 1000815
rect 70559 1000215 70615 1000815
rect 70735 1000215 70791 1000815
rect 70911 1000215 70961 1000815
rect 71217 1000803 71427 1000815
rect 71453 1000803 71663 1000815
rect 73187 1000803 73397 1000815
rect 73423 1000803 73633 1000815
rect 71221 1000800 71423 1000803
rect 71457 1000800 71659 1000803
rect 73191 1000800 73393 1000803
rect 73427 1000800 73629 1000803
rect 71232 1000630 71412 1000800
rect 71468 1000630 71648 1000800
rect 73202 1000630 73382 1000800
rect 73438 1000630 73618 1000800
rect 71217 1000615 71427 1000630
rect 71453 1000615 71663 1000630
rect 73187 1000615 73397 1000630
rect 73423 1000615 73633 1000630
rect 71453 1000502 71663 1000517
rect 73187 1000502 73397 1000517
rect 71468 1000480 71648 1000502
rect 73202 1000480 73382 1000502
rect 73889 1000215 73939 1000815
rect 74059 1000215 74115 1000815
rect 74235 1000215 74291 1000815
rect 74411 1000215 74461 1000815
rect 109264 1000665 109317 1000815
rect 109267 1000215 109317 1000665
rect 109437 1000215 109493 1000815
rect 109613 1000215 109669 1000815
rect 109789 1000215 109845 1000815
rect 109965 1000215 110015 1000815
rect 110081 1000215 110131 1000815
rect 110251 1000215 110307 1000815
rect 110427 1000215 110483 1000815
rect 110603 1000215 110653 1000815
rect 110924 1000615 111104 1000815
rect 111160 1000615 111253 1000815
rect 111160 1000480 111253 1000517
rect 122235 1000215 122291 1000815
rect 122411 1000215 122461 1000815
rect 161264 1000665 161317 1000815
rect 161267 1000215 161317 1000665
rect 161437 1000215 161493 1000815
rect 161613 1000215 161669 1000815
rect 161789 1000215 161845 1000815
rect 161965 1000215 162015 1000815
rect 162081 1000215 162131 1000815
rect 162251 1000215 162307 1000815
rect 162427 1000215 162483 1000815
rect 162603 1000215 162653 1000815
rect 162909 1000803 163119 1000815
rect 163145 1000803 163355 1000815
rect 164879 1000803 165089 1000815
rect 165115 1000803 165325 1000815
rect 162913 1000800 163115 1000803
rect 163149 1000800 163351 1000803
rect 164883 1000800 165085 1000803
rect 165119 1000800 165321 1000803
rect 162924 1000630 163104 1000800
rect 163160 1000630 163340 1000800
rect 164894 1000630 165074 1000800
rect 165130 1000630 165310 1000800
rect 162909 1000615 163119 1000630
rect 163145 1000615 163355 1000630
rect 164879 1000615 165089 1000630
rect 165115 1000615 165325 1000630
rect 163145 1000502 163355 1000517
rect 164879 1000502 165089 1000517
rect 163160 1000480 163340 1000502
rect 164894 1000480 165074 1000502
rect 165581 1000215 165631 1000815
rect 165751 1000215 165807 1000815
rect 165927 1000215 165983 1000815
rect 166103 1000215 166153 1000815
rect 166235 1000215 166285 1000815
rect 166405 1000215 166461 1000815
rect 166581 1000215 166637 1000815
rect 166757 1000215 166807 1000815
rect 167063 1000803 167273 1000815
rect 167299 1000803 167509 1000815
rect 169033 1000803 169243 1000815
rect 169269 1000803 169479 1000815
rect 167067 1000800 167269 1000803
rect 167303 1000800 167505 1000803
rect 169037 1000800 169239 1000803
rect 169273 1000800 169475 1000803
rect 167078 1000630 167258 1000800
rect 167314 1000630 167494 1000800
rect 169048 1000630 169228 1000800
rect 169284 1000630 169464 1000800
rect 167063 1000615 167273 1000630
rect 167299 1000615 167509 1000630
rect 169033 1000615 169243 1000630
rect 169269 1000615 169479 1000630
rect 167299 1000502 167509 1000517
rect 169033 1000502 169243 1000517
rect 167314 1000480 167494 1000502
rect 169048 1000480 169228 1000502
rect 169735 1000215 169785 1000815
rect 169905 1000215 169961 1000815
rect 170081 1000215 170137 1000815
rect 170257 1000215 170307 1000815
rect 170389 1000215 170439 1000815
rect 170559 1000215 170615 1000815
rect 170735 1000215 170791 1000815
rect 170911 1000215 170961 1000815
rect 171217 1000803 171427 1000815
rect 171453 1000803 171663 1000815
rect 173187 1000803 173397 1000815
rect 173423 1000803 173633 1000815
rect 171221 1000800 171423 1000803
rect 171457 1000800 171659 1000803
rect 173191 1000800 173393 1000803
rect 173427 1000800 173629 1000803
rect 171232 1000630 171412 1000800
rect 171468 1000630 171648 1000800
rect 173202 1000630 173382 1000800
rect 173438 1000630 173618 1000800
rect 171217 1000615 171427 1000630
rect 171453 1000615 171663 1000630
rect 173187 1000615 173397 1000630
rect 173423 1000615 173633 1000630
rect 171453 1000502 171663 1000517
rect 173187 1000502 173397 1000517
rect 171468 1000480 171648 1000502
rect 173202 1000480 173382 1000502
rect 173889 1000215 173939 1000815
rect 174059 1000215 174115 1000815
rect 174235 1000215 174291 1000815
rect 174411 1000215 174461 1000815
rect 213264 1000665 213317 1000815
rect 213267 1000215 213317 1000665
rect 213437 1000215 213493 1000815
rect 213613 1000215 213669 1000815
rect 213789 1000215 213845 1000815
rect 213965 1000215 214015 1000815
rect 214081 1000215 214131 1000815
rect 214251 1000215 214307 1000815
rect 214427 1000215 214483 1000815
rect 214603 1000215 214653 1000815
rect 214924 1000615 215104 1000815
rect 215160 1000615 215253 1000815
rect 215160 1000480 215253 1000517
rect 226235 1000215 226291 1000815
rect 226411 1000215 226461 1000815
rect 261264 1000665 261317 1000815
rect 261267 1000215 261317 1000665
rect 261437 1000215 261493 1000815
rect 261613 1000215 261669 1000815
rect 261789 1000215 261845 1000815
rect 261965 1000215 262015 1000815
rect 274235 1000215 274291 1000815
rect 274411 1000215 274461 1000815
rect 313264 1000665 313317 1000815
rect 313267 1000215 313317 1000665
rect 313437 1000215 313493 1000815
rect 313613 1000215 313669 1000815
rect 313789 1000215 313845 1000815
rect 313965 1000215 314015 1000815
rect 314081 1000215 314131 1000815
rect 314251 1000215 314307 1000815
rect 314427 1000215 314483 1000815
rect 314603 1000215 314653 1000815
rect 314924 1000615 315104 1000815
rect 315160 1000615 315253 1000815
rect 315160 1000480 315253 1000517
rect 326235 1000215 326291 1000815
rect 326411 1000215 326461 1000815
rect 365264 1000665 365317 1000815
rect 365267 1000215 365317 1000665
rect 365437 1000215 365493 1000815
rect 365613 1000215 365669 1000815
rect 365789 1000215 365845 1000815
rect 365965 1000215 366015 1000815
rect 366081 1000215 366131 1000815
rect 366251 1000215 366307 1000815
rect 366427 1000215 366483 1000815
rect 366603 1000215 366653 1000815
rect 366909 1000803 367119 1000815
rect 367145 1000803 367355 1000815
rect 368879 1000803 369089 1000815
rect 369115 1000803 369325 1000815
rect 366913 1000800 367115 1000803
rect 367149 1000800 367351 1000803
rect 368883 1000800 369085 1000803
rect 369119 1000800 369321 1000803
rect 366924 1000630 367104 1000800
rect 367160 1000630 367340 1000800
rect 368894 1000630 369074 1000800
rect 369130 1000630 369310 1000800
rect 366909 1000615 367119 1000630
rect 367145 1000615 367355 1000630
rect 368879 1000615 369089 1000630
rect 369115 1000615 369325 1000630
rect 367145 1000502 367355 1000517
rect 368879 1000502 369089 1000517
rect 367160 1000480 367340 1000502
rect 368894 1000480 369074 1000502
rect 369581 1000215 369631 1000815
rect 369751 1000215 369807 1000815
rect 369927 1000215 369983 1000815
rect 370103 1000215 370153 1000815
rect 370235 1000215 370285 1000815
rect 370405 1000215 370461 1000815
rect 370581 1000215 370637 1000815
rect 370757 1000215 370807 1000815
rect 371063 1000803 371273 1000815
rect 371299 1000803 371509 1000815
rect 373033 1000803 373243 1000815
rect 373269 1000803 373479 1000815
rect 371067 1000800 371269 1000803
rect 371303 1000800 371505 1000803
rect 373037 1000800 373239 1000803
rect 373273 1000800 373475 1000803
rect 371078 1000630 371258 1000800
rect 371314 1000630 371494 1000800
rect 373048 1000630 373228 1000800
rect 373284 1000630 373464 1000800
rect 371063 1000615 371273 1000630
rect 371299 1000615 371509 1000630
rect 373033 1000615 373243 1000630
rect 373269 1000615 373479 1000630
rect 371299 1000502 371509 1000517
rect 373033 1000502 373243 1000517
rect 371314 1000480 371494 1000502
rect 373048 1000480 373228 1000502
rect 373735 1000215 373785 1000815
rect 373905 1000215 373961 1000815
rect 374081 1000215 374137 1000815
rect 374257 1000215 374307 1000815
rect 374389 1000215 374439 1000815
rect 374559 1000215 374615 1000815
rect 374735 1000215 374791 1000815
rect 374911 1000215 374961 1000815
rect 375217 1000803 375427 1000815
rect 375453 1000803 375663 1000815
rect 377187 1000803 377397 1000815
rect 377423 1000803 377633 1000815
rect 375221 1000800 375423 1000803
rect 375457 1000800 375659 1000803
rect 377191 1000800 377393 1000803
rect 377427 1000800 377629 1000803
rect 375232 1000630 375412 1000800
rect 375468 1000630 375648 1000800
rect 377202 1000630 377382 1000800
rect 377438 1000630 377618 1000800
rect 375217 1000615 375427 1000630
rect 375453 1000615 375663 1000630
rect 377187 1000615 377397 1000630
rect 377423 1000615 377633 1000630
rect 375453 1000502 375663 1000517
rect 377187 1000502 377397 1000517
rect 375468 1000480 375648 1000502
rect 377202 1000480 377382 1000502
rect 377889 1000215 377939 1000815
rect 378059 1000215 378115 1000815
rect 378235 1000215 378291 1000815
rect 378411 1000215 378461 1000815
rect 413264 1000665 413317 1000815
rect 413267 1000215 413317 1000665
rect 413437 1000215 413493 1000815
rect 413613 1000215 413669 1000815
rect 413789 1000215 413845 1000815
rect 413965 1000215 414015 1000815
rect 414081 1000215 414131 1000815
rect 414251 1000215 414307 1000815
rect 414427 1000215 414483 1000815
rect 414603 1000215 414653 1000815
rect 414924 1000615 415104 1000815
rect 415160 1000615 415253 1000815
rect 415160 1000480 415253 1000517
rect 426235 1000215 426291 1000815
rect 426411 1000215 426461 1000815
rect 465264 1000665 465317 1000815
rect 465267 1000215 465317 1000665
rect 465437 1000215 465493 1000815
rect 465613 1000215 465669 1000815
rect 465789 1000215 465845 1000815
rect 465965 1000215 466015 1000815
rect 466081 1000215 466131 1000815
rect 466251 1000215 466307 1000815
rect 466427 1000215 466483 1000815
rect 466603 1000215 466653 1000815
rect 466909 1000803 467119 1000815
rect 467145 1000803 467355 1000815
rect 468879 1000803 469089 1000815
rect 469115 1000803 469325 1000815
rect 466913 1000800 467115 1000803
rect 467149 1000800 467351 1000803
rect 468883 1000800 469085 1000803
rect 469119 1000800 469321 1000803
rect 466924 1000630 467104 1000800
rect 467160 1000630 467340 1000800
rect 468894 1000630 469074 1000800
rect 469130 1000630 469310 1000800
rect 466909 1000615 467119 1000630
rect 467145 1000615 467355 1000630
rect 468879 1000615 469089 1000630
rect 469115 1000615 469325 1000630
rect 467145 1000502 467355 1000517
rect 468879 1000502 469089 1000517
rect 467160 1000480 467340 1000502
rect 468894 1000480 469074 1000502
rect 469581 1000215 469631 1000815
rect 469751 1000215 469807 1000815
rect 469927 1000215 469983 1000815
rect 470103 1000215 470153 1000815
rect 470235 1000215 470285 1000815
rect 470405 1000215 470461 1000815
rect 470581 1000215 470637 1000815
rect 470757 1000215 470807 1000815
rect 471063 1000803 471273 1000815
rect 471299 1000803 471509 1000815
rect 473033 1000803 473243 1000815
rect 473269 1000803 473479 1000815
rect 471067 1000800 471269 1000803
rect 471303 1000800 471505 1000803
rect 473037 1000800 473239 1000803
rect 473273 1000800 473475 1000803
rect 471078 1000630 471258 1000800
rect 471314 1000630 471494 1000800
rect 473048 1000630 473228 1000800
rect 473284 1000630 473464 1000800
rect 471063 1000615 471273 1000630
rect 471299 1000615 471509 1000630
rect 473033 1000615 473243 1000630
rect 473269 1000615 473479 1000630
rect 471299 1000502 471509 1000517
rect 473033 1000502 473243 1000517
rect 471314 1000480 471494 1000502
rect 473048 1000480 473228 1000502
rect 473735 1000215 473785 1000815
rect 473905 1000215 473961 1000815
rect 474081 1000215 474137 1000815
rect 474257 1000215 474307 1000815
rect 474389 1000215 474439 1000815
rect 474559 1000215 474615 1000815
rect 474735 1000215 474791 1000815
rect 474911 1000215 474961 1000815
rect 475217 1000803 475427 1000815
rect 475453 1000803 475663 1000815
rect 477187 1000803 477397 1000815
rect 477423 1000803 477633 1000815
rect 475221 1000800 475423 1000803
rect 475457 1000800 475659 1000803
rect 477191 1000800 477393 1000803
rect 477427 1000800 477629 1000803
rect 475232 1000630 475412 1000800
rect 475468 1000630 475648 1000800
rect 477202 1000630 477382 1000800
rect 477438 1000630 477618 1000800
rect 475217 1000615 475427 1000630
rect 475453 1000615 475663 1000630
rect 477187 1000615 477397 1000630
rect 477423 1000615 477633 1000630
rect 475453 1000502 475663 1000517
rect 477187 1000502 477397 1000517
rect 475468 1000480 475648 1000502
rect 477202 1000480 477382 1000502
rect 477889 1000215 477939 1000815
rect 478059 1000215 478115 1000815
rect 478235 1000215 478291 1000815
rect 478411 1000215 478461 1000815
rect 517264 1000665 517317 1000815
rect 517267 1000215 517317 1000665
rect 517437 1000215 517493 1000815
rect 517613 1000215 517669 1000815
rect 517789 1000215 517845 1000815
rect 517965 1000215 518015 1000815
rect 518081 1000215 518131 1000815
rect 518251 1000215 518307 1000815
rect 518427 1000215 518483 1000815
rect 518603 1000215 518653 1000815
rect 518924 1000615 519104 1000815
rect 519160 1000615 519253 1000815
rect 519160 1000480 519253 1000517
rect 530235 1000215 530291 1000815
rect 530411 1000215 530461 1000815
rect 569264 1000665 569317 1000815
rect 569267 1000215 569317 1000665
rect 569437 1000215 569493 1000815
rect 569613 1000215 569669 1000815
rect 569789 1000215 569845 1000815
rect 569965 1000215 570015 1000815
rect 570081 1000215 570131 1000815
rect 570251 1000215 570307 1000815
rect 570427 1000215 570483 1000815
rect 570603 1000215 570653 1000815
rect 570909 1000803 571119 1000815
rect 571145 1000803 571355 1000815
rect 572879 1000803 573089 1000815
rect 573115 1000803 573325 1000815
rect 570913 1000800 571115 1000803
rect 571149 1000800 571351 1000803
rect 572883 1000800 573085 1000803
rect 573119 1000800 573321 1000803
rect 570924 1000630 571104 1000800
rect 571160 1000630 571340 1000800
rect 572894 1000630 573074 1000800
rect 573130 1000630 573310 1000800
rect 570909 1000615 571119 1000630
rect 571145 1000615 571355 1000630
rect 572879 1000615 573089 1000630
rect 573115 1000615 573325 1000630
rect 571145 1000502 571355 1000517
rect 572879 1000502 573089 1000517
rect 571160 1000480 571340 1000502
rect 572894 1000480 573074 1000502
rect 573581 1000215 573631 1000815
rect 573751 1000215 573807 1000815
rect 573927 1000215 573983 1000815
rect 574103 1000215 574153 1000815
rect 574235 1000215 574285 1000815
rect 574405 1000215 574461 1000815
rect 574581 1000215 574637 1000815
rect 574757 1000215 574807 1000815
rect 575063 1000803 575273 1000815
rect 575299 1000803 575509 1000815
rect 577033 1000803 577243 1000815
rect 577269 1000803 577479 1000815
rect 575067 1000800 575269 1000803
rect 575303 1000800 575505 1000803
rect 577037 1000800 577239 1000803
rect 577273 1000800 577475 1000803
rect 575078 1000630 575258 1000800
rect 575314 1000630 575494 1000800
rect 577048 1000630 577228 1000800
rect 577284 1000630 577464 1000800
rect 575063 1000615 575273 1000630
rect 575299 1000615 575509 1000630
rect 577033 1000615 577243 1000630
rect 577269 1000615 577479 1000630
rect 575299 1000502 575509 1000517
rect 577033 1000502 577243 1000517
rect 575314 1000480 575494 1000502
rect 577048 1000480 577228 1000502
rect 577735 1000215 577785 1000815
rect 577905 1000215 577961 1000815
rect 578081 1000215 578137 1000815
rect 578257 1000215 578307 1000815
rect 578389 1000215 578439 1000815
rect 578559 1000215 578615 1000815
rect 578735 1000215 578791 1000815
rect 578911 1000215 578961 1000815
rect 579217 1000803 579427 1000815
rect 579453 1000803 579663 1000815
rect 581187 1000803 581397 1000815
rect 581423 1000803 581633 1000815
rect 579221 1000800 579423 1000803
rect 579457 1000800 579659 1000803
rect 581191 1000800 581393 1000803
rect 581427 1000800 581629 1000803
rect 579232 1000630 579412 1000800
rect 579468 1000630 579648 1000800
rect 581202 1000630 581382 1000800
rect 581438 1000630 581618 1000800
rect 579217 1000615 579427 1000630
rect 579453 1000615 579663 1000630
rect 581187 1000615 581397 1000630
rect 581423 1000615 581633 1000630
rect 579453 1000502 579663 1000517
rect 581187 1000502 581397 1000517
rect 579468 1000480 579648 1000502
rect 581202 1000480 581382 1000502
rect 581889 1000215 581939 1000815
rect 582059 1000215 582115 1000815
rect 582235 1000215 582291 1000815
rect 582411 1000215 582461 1000815
rect 74642 999817 74666 999841
rect 75063 999817 75087 999841
rect 174642 999817 174666 999841
rect 175063 999817 175087 999841
rect 378642 999817 378666 999841
rect 379063 999817 379087 999841
rect 478642 999817 478666 999841
rect 479063 999817 479087 999841
rect 582642 999817 582666 999841
rect 583063 999817 583087 999841
rect 74666 999793 74690 999808
rect 75039 999793 75063 999808
rect 174666 999793 174690 999808
rect 175039 999793 175063 999808
rect 378666 999793 378690 999808
rect 379039 999793 379063 999808
rect 478666 999793 478690 999808
rect 479039 999793 479063 999808
rect 582666 999793 582690 999808
rect 583039 999793 583063 999808
rect 74470 999637 74494 999661
rect 174470 999637 174494 999661
rect 378470 999637 378494 999661
rect 478470 999637 478494 999661
rect 582470 999637 582494 999661
rect 74495 999613 74518 999637
rect 174495 999613 174518 999637
rect 378495 999613 378518 999637
rect 478495 999613 478518 999637
rect 582495 999613 582518 999637
rect 60890 998799 60940 999399
rect 61060 998799 61116 999399
rect 61236 998799 61286 999399
rect 62779 999007 62829 999607
rect 62949 999007 62999 999607
rect 63375 999002 63425 999602
rect 63545 999002 63601 999602
rect 63721 999355 63771 999602
rect 63834 999452 63846 999602
rect 64460 999452 64513 999602
rect 64463 999355 64513 999452
rect 63721 999283 63774 999355
rect 63721 999002 63771 999283
rect 63834 999133 63846 999283
rect 64460 999133 64513 999355
rect 64463 999002 64513 999133
rect 64633 999002 64689 999602
rect 64809 999002 64859 999602
rect 65235 999007 65285 999607
rect 65405 999007 65455 999607
rect 66933 999007 66983 999607
rect 67103 999007 67153 999607
rect 67529 999002 67579 999602
rect 67699 999002 67755 999602
rect 67875 999355 67925 999602
rect 67988 999452 68000 999602
rect 68614 999452 68667 999602
rect 68617 999355 68667 999452
rect 67875 999283 67928 999355
rect 67875 999002 67925 999283
rect 67988 999133 68000 999283
rect 68614 999133 68667 999355
rect 68617 999002 68667 999133
rect 68787 999002 68843 999602
rect 68963 999002 69013 999602
rect 69389 999007 69439 999607
rect 69559 999007 69609 999607
rect 71087 999007 71137 999607
rect 71257 999007 71307 999607
rect 71683 999002 71733 999602
rect 71853 999002 71909 999602
rect 72029 999355 72079 999602
rect 72142 999452 72154 999602
rect 72768 999452 72821 999602
rect 72771 999355 72821 999452
rect 72029 999283 72082 999355
rect 72029 999002 72079 999283
rect 72142 999133 72154 999283
rect 72768 999133 72821 999355
rect 72771 999002 72821 999133
rect 72941 999002 72997 999602
rect 73117 999002 73167 999602
rect 73543 999007 73593 999607
rect 73713 999007 73763 999607
rect 74690 999549 74724 999573
rect 74760 999549 74794 999573
rect 74830 999549 74864 999573
rect 74900 999549 74934 999573
rect 74970 999549 75004 999573
rect 75040 999549 75063 999573
rect 74495 999515 74518 999539
rect 74470 999491 74494 999515
rect 108890 998799 108940 999399
rect 109060 998799 109116 999399
rect 109236 998799 109286 999399
rect 110779 999007 110829 999607
rect 110949 999007 110999 999607
rect 160890 998799 160940 999399
rect 161060 998799 161116 999399
rect 161236 998799 161286 999399
rect 162779 999007 162829 999607
rect 162949 999007 162999 999607
rect 163375 999002 163425 999602
rect 163545 999002 163601 999602
rect 163721 999355 163771 999602
rect 163834 999452 163846 999602
rect 164460 999452 164513 999602
rect 164463 999355 164513 999452
rect 163721 999283 163774 999355
rect 163721 999002 163771 999283
rect 163834 999133 163846 999283
rect 164460 999133 164513 999355
rect 164463 999002 164513 999133
rect 164633 999002 164689 999602
rect 164809 999002 164859 999602
rect 165235 999007 165285 999607
rect 165405 999007 165455 999607
rect 166933 999007 166983 999607
rect 167103 999007 167153 999607
rect 167529 999002 167579 999602
rect 167699 999002 167755 999602
rect 167875 999355 167925 999602
rect 167988 999452 168000 999602
rect 168614 999452 168667 999602
rect 168617 999355 168667 999452
rect 167875 999283 167928 999355
rect 167875 999002 167925 999283
rect 167988 999133 168000 999283
rect 168614 999133 168667 999355
rect 168617 999002 168667 999133
rect 168787 999002 168843 999602
rect 168963 999002 169013 999602
rect 169389 999007 169439 999607
rect 169559 999007 169609 999607
rect 171087 999007 171137 999607
rect 171257 999007 171307 999607
rect 171683 999002 171733 999602
rect 171853 999002 171909 999602
rect 172029 999355 172079 999602
rect 172142 999452 172154 999602
rect 172768 999452 172821 999602
rect 172771 999355 172821 999452
rect 172029 999283 172082 999355
rect 172029 999002 172079 999283
rect 172142 999133 172154 999283
rect 172768 999133 172821 999355
rect 172771 999002 172821 999133
rect 172941 999002 172997 999602
rect 173117 999002 173167 999602
rect 173543 999007 173593 999607
rect 173713 999007 173763 999607
rect 174690 999549 174724 999573
rect 174760 999549 174794 999573
rect 174830 999549 174864 999573
rect 174900 999549 174934 999573
rect 174970 999549 175004 999573
rect 175040 999549 175063 999573
rect 174495 999515 174518 999539
rect 174470 999491 174494 999515
rect 212890 998799 212940 999399
rect 213060 998799 213116 999399
rect 213236 998799 213286 999399
rect 214779 999007 214829 999607
rect 214949 999007 214999 999607
rect 260890 998799 260940 999399
rect 261060 998799 261116 999399
rect 261236 998799 261286 999399
rect 312890 998799 312940 999399
rect 313060 998799 313116 999399
rect 313236 998799 313286 999399
rect 314779 999007 314829 999607
rect 314949 999007 314999 999607
rect 364890 998799 364940 999399
rect 365060 998799 365116 999399
rect 365236 998799 365286 999399
rect 366779 999007 366829 999607
rect 366949 999007 366999 999607
rect 367375 999002 367425 999602
rect 367545 999002 367601 999602
rect 367721 999355 367771 999602
rect 367834 999452 367846 999602
rect 368460 999452 368513 999602
rect 368463 999355 368513 999452
rect 367721 999283 367774 999355
rect 367721 999002 367771 999283
rect 367834 999133 367846 999283
rect 368460 999133 368513 999355
rect 368463 999002 368513 999133
rect 368633 999002 368689 999602
rect 368809 999002 368859 999602
rect 369235 999007 369285 999607
rect 369405 999007 369455 999607
rect 370933 999007 370983 999607
rect 371103 999007 371153 999607
rect 371529 999002 371579 999602
rect 371699 999002 371755 999602
rect 371875 999355 371925 999602
rect 371988 999452 372000 999602
rect 372614 999452 372667 999602
rect 372617 999355 372667 999452
rect 371875 999283 371928 999355
rect 371875 999002 371925 999283
rect 371988 999133 372000 999283
rect 372614 999133 372667 999355
rect 372617 999002 372667 999133
rect 372787 999002 372843 999602
rect 372963 999002 373013 999602
rect 373389 999007 373439 999607
rect 373559 999007 373609 999607
rect 375087 999007 375137 999607
rect 375257 999007 375307 999607
rect 375683 999002 375733 999602
rect 375853 999002 375909 999602
rect 376029 999355 376079 999602
rect 376142 999452 376154 999602
rect 376768 999452 376821 999602
rect 376771 999355 376821 999452
rect 376029 999283 376082 999355
rect 376029 999002 376079 999283
rect 376142 999133 376154 999283
rect 376768 999133 376821 999355
rect 376771 999002 376821 999133
rect 376941 999002 376997 999602
rect 377117 999002 377167 999602
rect 377543 999007 377593 999607
rect 377713 999007 377763 999607
rect 378690 999549 378724 999573
rect 378760 999549 378794 999573
rect 378830 999549 378864 999573
rect 378900 999549 378934 999573
rect 378970 999549 379004 999573
rect 379040 999549 379063 999573
rect 378495 999515 378518 999539
rect 378470 999491 378494 999515
rect 412890 998799 412940 999399
rect 413060 998799 413116 999399
rect 413236 998799 413286 999399
rect 414779 999007 414829 999607
rect 414949 999007 414999 999607
rect 464890 998799 464940 999399
rect 465060 998799 465116 999399
rect 465236 998799 465286 999399
rect 466779 999007 466829 999607
rect 466949 999007 466999 999607
rect 467375 999002 467425 999602
rect 467545 999002 467601 999602
rect 467721 999355 467771 999602
rect 467834 999452 467846 999602
rect 468460 999452 468513 999602
rect 468463 999355 468513 999452
rect 467721 999283 467774 999355
rect 467721 999002 467771 999283
rect 467834 999133 467846 999283
rect 468460 999133 468513 999355
rect 468463 999002 468513 999133
rect 468633 999002 468689 999602
rect 468809 999002 468859 999602
rect 469235 999007 469285 999607
rect 469405 999007 469455 999607
rect 470933 999007 470983 999607
rect 471103 999007 471153 999607
rect 471529 999002 471579 999602
rect 471699 999002 471755 999602
rect 471875 999355 471925 999602
rect 471988 999452 472000 999602
rect 472614 999452 472667 999602
rect 472617 999355 472667 999452
rect 471875 999283 471928 999355
rect 471875 999002 471925 999283
rect 471988 999133 472000 999283
rect 472614 999133 472667 999355
rect 472617 999002 472667 999133
rect 472787 999002 472843 999602
rect 472963 999002 473013 999602
rect 473389 999007 473439 999607
rect 473559 999007 473609 999607
rect 475087 999007 475137 999607
rect 475257 999007 475307 999607
rect 475683 999002 475733 999602
rect 475853 999002 475909 999602
rect 476029 999355 476079 999602
rect 476142 999452 476154 999602
rect 476768 999452 476821 999602
rect 476771 999355 476821 999452
rect 476029 999283 476082 999355
rect 476029 999002 476079 999283
rect 476142 999133 476154 999283
rect 476768 999133 476821 999355
rect 476771 999002 476821 999133
rect 476941 999002 476997 999602
rect 477117 999002 477167 999602
rect 477543 999007 477593 999607
rect 477713 999007 477763 999607
rect 478690 999549 478724 999573
rect 478760 999549 478794 999573
rect 478830 999549 478864 999573
rect 478900 999549 478934 999573
rect 478970 999549 479004 999573
rect 479040 999549 479063 999573
rect 478495 999515 478518 999539
rect 478470 999491 478494 999515
rect 516890 998799 516940 999399
rect 517060 998799 517116 999399
rect 517236 998799 517286 999399
rect 518779 999007 518829 999607
rect 518949 999007 518999 999607
rect 568890 998799 568940 999399
rect 569060 998799 569116 999399
rect 569236 998799 569286 999399
rect 570779 999007 570829 999607
rect 570949 999007 570999 999607
rect 571375 999002 571425 999602
rect 571545 999002 571601 999602
rect 571721 999355 571771 999602
rect 571834 999452 571846 999602
rect 572460 999452 572513 999602
rect 572463 999355 572513 999452
rect 571721 999283 571774 999355
rect 571721 999002 571771 999283
rect 571834 999133 571846 999283
rect 572460 999133 572513 999355
rect 572463 999002 572513 999133
rect 572633 999002 572689 999602
rect 572809 999002 572859 999602
rect 573235 999007 573285 999607
rect 573405 999007 573455 999607
rect 574933 999007 574983 999607
rect 575103 999007 575153 999607
rect 575529 999002 575579 999602
rect 575699 999002 575755 999602
rect 575875 999355 575925 999602
rect 575988 999452 576000 999602
rect 576614 999452 576667 999602
rect 576617 999355 576667 999452
rect 575875 999283 575928 999355
rect 575875 999002 575925 999283
rect 575988 999133 576000 999283
rect 576614 999133 576667 999355
rect 576617 999002 576667 999133
rect 576787 999002 576843 999602
rect 576963 999002 577013 999602
rect 577389 999007 577439 999607
rect 577559 999007 577609 999607
rect 579087 999007 579137 999607
rect 579257 999007 579307 999607
rect 579683 999002 579733 999602
rect 579853 999002 579909 999602
rect 580029 999355 580079 999602
rect 580142 999452 580154 999602
rect 580768 999452 580821 999602
rect 580771 999355 580821 999452
rect 580029 999283 580082 999355
rect 580029 999002 580079 999283
rect 580142 999133 580154 999283
rect 580768 999133 580821 999355
rect 580771 999002 580821 999133
rect 580941 999002 580997 999602
rect 581117 999002 581167 999602
rect 581543 999007 581593 999607
rect 581713 999007 581763 999607
rect 582690 999549 582724 999573
rect 582760 999549 582794 999573
rect 582830 999549 582864 999573
rect 582900 999549 582934 999573
rect 582970 999549 583004 999573
rect 583040 999549 583063 999573
rect 582495 999515 582518 999539
rect 582470 999491 582494 999515
rect 62318 998680 62352 998704
rect 62386 998680 62420 998704
rect 62454 998680 62488 998704
rect 62522 998680 62556 998704
rect 62590 998680 62624 998704
rect 62658 998680 62692 998704
rect 62726 998680 62760 998704
rect 62794 998680 62828 998704
rect 62862 998680 62896 998704
rect 62930 998680 62964 998704
rect 62998 998680 63032 998704
rect 63066 998680 63100 998704
rect 63134 998680 63168 998704
rect 63202 998680 63236 998704
rect 63270 998680 63304 998704
rect 63338 998680 63372 998704
rect 63406 998680 63440 998704
rect 63474 998680 63508 998704
rect 63542 998680 63576 998704
rect 63610 998680 63644 998704
rect 63678 998680 63712 998704
rect 63746 998680 63780 998704
rect 63814 998680 63848 998704
rect 63882 998680 63916 998704
rect 63950 998680 63984 998704
rect 64018 998680 64052 998704
rect 64086 998680 64120 998704
rect 64154 998680 64188 998704
rect 64222 998680 64256 998704
rect 64290 998680 64324 998704
rect 64358 998680 64392 998704
rect 64426 998680 64460 998704
rect 64494 998680 64528 998704
rect 64562 998680 64596 998704
rect 64630 998680 64664 998704
rect 64698 998680 64732 998704
rect 64766 998680 64800 998704
rect 64834 998680 64868 998704
rect 64902 998680 64936 998704
rect 64970 998680 65004 998704
rect 65038 998680 65072 998704
rect 65106 998680 65140 998704
rect 65174 998680 65208 998704
rect 65242 998680 65276 998704
rect 65310 998680 65344 998704
rect 65378 998680 65412 998704
rect 65446 998680 65480 998704
rect 65514 998680 65548 998704
rect 65582 998680 65616 998704
rect 65650 998680 65684 998704
rect 65718 998680 65752 998704
rect 65786 998680 65820 998704
rect 65854 998680 65888 998704
rect 65922 998680 65956 998704
rect 65990 998680 66024 998704
rect 66058 998680 66092 998704
rect 66126 998680 66160 998704
rect 66194 998680 66228 998704
rect 66262 998680 66296 998704
rect 66330 998680 66364 998704
rect 66398 998680 66432 998704
rect 66466 998680 66500 998704
rect 66534 998680 66568 998704
rect 66602 998680 66636 998704
rect 66670 998680 66704 998704
rect 66738 998680 66772 998704
rect 66806 998680 66840 998704
rect 66874 998680 66908 998704
rect 66942 998680 66976 998704
rect 67010 998680 67044 998704
rect 67078 998680 67112 998704
rect 67146 998680 67180 998704
rect 67214 998680 67248 998704
rect 67282 998680 67316 998704
rect 67350 998680 67384 998704
rect 67418 998680 67452 998704
rect 67486 998680 67520 998704
rect 67554 998680 67588 998704
rect 67622 998680 67656 998704
rect 67690 998680 67724 998704
rect 67758 998680 67792 998704
rect 67826 998680 67860 998704
rect 67894 998680 67928 998704
rect 67962 998680 67996 998704
rect 68030 998680 68064 998704
rect 68098 998680 68132 998704
rect 68166 998680 68200 998704
rect 68234 998680 68268 998704
rect 68302 998680 68336 998704
rect 68370 998680 68404 998704
rect 68438 998680 68472 998704
rect 68506 998680 68540 998704
rect 68574 998680 68608 998704
rect 68642 998680 68676 998704
rect 68710 998680 68744 998704
rect 68778 998680 68812 998704
rect 68846 998680 68880 998704
rect 68914 998680 68948 998704
rect 68982 998680 69016 998704
rect 69050 998680 69084 998704
rect 69118 998680 69152 998704
rect 69186 998680 69220 998704
rect 69254 998680 69288 998704
rect 69322 998680 69356 998704
rect 69390 998680 69424 998704
rect 69458 998680 69492 998704
rect 69526 998680 69560 998704
rect 69594 998680 69628 998704
rect 69662 998680 69696 998704
rect 69796 998680 69830 998704
rect 69864 998680 69898 998704
rect 69932 998680 69966 998704
rect 70000 998680 70034 998704
rect 70068 998680 70102 998704
rect 70136 998680 70170 998704
rect 70204 998680 70238 998704
rect 70272 998680 70306 998704
rect 70340 998680 70374 998704
rect 70408 998680 70442 998704
rect 70476 998680 70510 998704
rect 70544 998680 70578 998704
rect 70612 998680 70646 998704
rect 70680 998680 70714 998704
rect 70748 998680 70782 998704
rect 70816 998680 70850 998704
rect 70884 998680 70918 998704
rect 70952 998680 70986 998704
rect 71020 998680 71054 998704
rect 71088 998680 71122 998704
rect 71156 998680 71190 998704
rect 71224 998680 71258 998704
rect 71292 998680 71326 998704
rect 71360 998680 71394 998704
rect 71428 998680 71462 998704
rect 71496 998680 71530 998704
rect 71564 998680 71598 998704
rect 71632 998680 71666 998704
rect 71700 998680 71734 998704
rect 71768 998680 71802 998704
rect 71836 998680 71870 998704
rect 71904 998680 71938 998704
rect 71972 998680 72006 998704
rect 72040 998680 72074 998704
rect 72108 998680 72142 998704
rect 72176 998680 72210 998704
rect 72244 998680 72278 998704
rect 72312 998680 72346 998704
rect 72380 998680 72414 998704
rect 72448 998680 72482 998704
rect 72516 998680 72550 998704
rect 72584 998680 72618 998704
rect 72652 998680 72686 998704
rect 72720 998680 72754 998704
rect 72788 998680 72822 998704
rect 72856 998680 72890 998704
rect 162318 998680 162352 998704
rect 162386 998680 162420 998704
rect 162454 998680 162488 998704
rect 162522 998680 162556 998704
rect 162590 998680 162624 998704
rect 162658 998680 162692 998704
rect 162726 998680 162760 998704
rect 162794 998680 162828 998704
rect 162862 998680 162896 998704
rect 162930 998680 162964 998704
rect 162998 998680 163032 998704
rect 163066 998680 163100 998704
rect 163134 998680 163168 998704
rect 163202 998680 163236 998704
rect 163270 998680 163304 998704
rect 163338 998680 163372 998704
rect 163406 998680 163440 998704
rect 163474 998680 163508 998704
rect 163542 998680 163576 998704
rect 163610 998680 163644 998704
rect 163678 998680 163712 998704
rect 163746 998680 163780 998704
rect 163814 998680 163848 998704
rect 163882 998680 163916 998704
rect 163950 998680 163984 998704
rect 164018 998680 164052 998704
rect 164086 998680 164120 998704
rect 164154 998680 164188 998704
rect 164222 998680 164256 998704
rect 164290 998680 164324 998704
rect 164358 998680 164392 998704
rect 164426 998680 164460 998704
rect 164494 998680 164528 998704
rect 164562 998680 164596 998704
rect 164630 998680 164664 998704
rect 164698 998680 164732 998704
rect 164766 998680 164800 998704
rect 164834 998680 164868 998704
rect 164902 998680 164936 998704
rect 164970 998680 165004 998704
rect 165038 998680 165072 998704
rect 165106 998680 165140 998704
rect 165174 998680 165208 998704
rect 165242 998680 165276 998704
rect 165310 998680 165344 998704
rect 165378 998680 165412 998704
rect 165446 998680 165480 998704
rect 165514 998680 165548 998704
rect 165582 998680 165616 998704
rect 165650 998680 165684 998704
rect 165718 998680 165752 998704
rect 165786 998680 165820 998704
rect 165854 998680 165888 998704
rect 165922 998680 165956 998704
rect 165990 998680 166024 998704
rect 166058 998680 166092 998704
rect 166126 998680 166160 998704
rect 166194 998680 166228 998704
rect 166262 998680 166296 998704
rect 166330 998680 166364 998704
rect 166398 998680 166432 998704
rect 166466 998680 166500 998704
rect 166534 998680 166568 998704
rect 166602 998680 166636 998704
rect 166670 998680 166704 998704
rect 166738 998680 166772 998704
rect 166806 998680 166840 998704
rect 166874 998680 166908 998704
rect 166942 998680 166976 998704
rect 167010 998680 167044 998704
rect 167078 998680 167112 998704
rect 167146 998680 167180 998704
rect 167214 998680 167248 998704
rect 167282 998680 167316 998704
rect 167350 998680 167384 998704
rect 167418 998680 167452 998704
rect 167486 998680 167520 998704
rect 167554 998680 167588 998704
rect 167622 998680 167656 998704
rect 167690 998680 167724 998704
rect 167758 998680 167792 998704
rect 167826 998680 167860 998704
rect 167894 998680 167928 998704
rect 167962 998680 167996 998704
rect 168030 998680 168064 998704
rect 168098 998680 168132 998704
rect 168166 998680 168200 998704
rect 168234 998680 168268 998704
rect 168302 998680 168336 998704
rect 168370 998680 168404 998704
rect 168438 998680 168472 998704
rect 168506 998680 168540 998704
rect 168574 998680 168608 998704
rect 168642 998680 168676 998704
rect 168710 998680 168744 998704
rect 168778 998680 168812 998704
rect 168846 998680 168880 998704
rect 168914 998680 168948 998704
rect 168982 998680 169016 998704
rect 169050 998680 169084 998704
rect 169118 998680 169152 998704
rect 169186 998680 169220 998704
rect 169254 998680 169288 998704
rect 169322 998680 169356 998704
rect 169390 998680 169424 998704
rect 169458 998680 169492 998704
rect 169526 998680 169560 998704
rect 169594 998680 169628 998704
rect 169662 998680 169696 998704
rect 169796 998680 169830 998704
rect 169864 998680 169898 998704
rect 169932 998680 169966 998704
rect 170000 998680 170034 998704
rect 170068 998680 170102 998704
rect 170136 998680 170170 998704
rect 170204 998680 170238 998704
rect 170272 998680 170306 998704
rect 170340 998680 170374 998704
rect 170408 998680 170442 998704
rect 170476 998680 170510 998704
rect 170544 998680 170578 998704
rect 170612 998680 170646 998704
rect 170680 998680 170714 998704
rect 170748 998680 170782 998704
rect 170816 998680 170850 998704
rect 170884 998680 170918 998704
rect 170952 998680 170986 998704
rect 171020 998680 171054 998704
rect 171088 998680 171122 998704
rect 171156 998680 171190 998704
rect 171224 998680 171258 998704
rect 171292 998680 171326 998704
rect 171360 998680 171394 998704
rect 171428 998680 171462 998704
rect 171496 998680 171530 998704
rect 171564 998680 171598 998704
rect 171632 998680 171666 998704
rect 171700 998680 171734 998704
rect 171768 998680 171802 998704
rect 171836 998680 171870 998704
rect 171904 998680 171938 998704
rect 171972 998680 172006 998704
rect 172040 998680 172074 998704
rect 172108 998680 172142 998704
rect 172176 998680 172210 998704
rect 172244 998680 172278 998704
rect 172312 998680 172346 998704
rect 172380 998680 172414 998704
rect 172448 998680 172482 998704
rect 172516 998680 172550 998704
rect 172584 998680 172618 998704
rect 172652 998680 172686 998704
rect 172720 998680 172754 998704
rect 172788 998680 172822 998704
rect 172856 998680 172890 998704
rect 366318 998680 366352 998704
rect 366386 998680 366420 998704
rect 366454 998680 366488 998704
rect 366522 998680 366556 998704
rect 366590 998680 366624 998704
rect 366658 998680 366692 998704
rect 366726 998680 366760 998704
rect 366794 998680 366828 998704
rect 366862 998680 366896 998704
rect 366930 998680 366964 998704
rect 366998 998680 367032 998704
rect 367066 998680 367100 998704
rect 367134 998680 367168 998704
rect 367202 998680 367236 998704
rect 367270 998680 367304 998704
rect 367338 998680 367372 998704
rect 367406 998680 367440 998704
rect 367474 998680 367508 998704
rect 367542 998680 367576 998704
rect 367610 998680 367644 998704
rect 367678 998680 367712 998704
rect 367746 998680 367780 998704
rect 367814 998680 367848 998704
rect 367882 998680 367916 998704
rect 367950 998680 367984 998704
rect 368018 998680 368052 998704
rect 368086 998680 368120 998704
rect 368154 998680 368188 998704
rect 368222 998680 368256 998704
rect 368290 998680 368324 998704
rect 368358 998680 368392 998704
rect 368426 998680 368460 998704
rect 368494 998680 368528 998704
rect 368562 998680 368596 998704
rect 368630 998680 368664 998704
rect 368698 998680 368732 998704
rect 368766 998680 368800 998704
rect 368834 998680 368868 998704
rect 368902 998680 368936 998704
rect 368970 998680 369004 998704
rect 369038 998680 369072 998704
rect 369106 998680 369140 998704
rect 369174 998680 369208 998704
rect 369242 998680 369276 998704
rect 369310 998680 369344 998704
rect 369378 998680 369412 998704
rect 369446 998680 369480 998704
rect 369514 998680 369548 998704
rect 369582 998680 369616 998704
rect 369650 998680 369684 998704
rect 369718 998680 369752 998704
rect 369786 998680 369820 998704
rect 369854 998680 369888 998704
rect 369922 998680 369956 998704
rect 369990 998680 370024 998704
rect 370058 998680 370092 998704
rect 370126 998680 370160 998704
rect 370194 998680 370228 998704
rect 370262 998680 370296 998704
rect 370330 998680 370364 998704
rect 370398 998680 370432 998704
rect 370466 998680 370500 998704
rect 370534 998680 370568 998704
rect 370602 998680 370636 998704
rect 370670 998680 370704 998704
rect 370738 998680 370772 998704
rect 370806 998680 370840 998704
rect 370874 998680 370908 998704
rect 370942 998680 370976 998704
rect 371010 998680 371044 998704
rect 371078 998680 371112 998704
rect 371146 998680 371180 998704
rect 371214 998680 371248 998704
rect 371282 998680 371316 998704
rect 371350 998680 371384 998704
rect 371418 998680 371452 998704
rect 371486 998680 371520 998704
rect 371554 998680 371588 998704
rect 371622 998680 371656 998704
rect 371690 998680 371724 998704
rect 371758 998680 371792 998704
rect 371826 998680 371860 998704
rect 371894 998680 371928 998704
rect 371962 998680 371996 998704
rect 372030 998680 372064 998704
rect 372098 998680 372132 998704
rect 372166 998680 372200 998704
rect 372234 998680 372268 998704
rect 372302 998680 372336 998704
rect 372370 998680 372404 998704
rect 372438 998680 372472 998704
rect 372506 998680 372540 998704
rect 372574 998680 372608 998704
rect 372642 998680 372676 998704
rect 372710 998680 372744 998704
rect 372778 998680 372812 998704
rect 372846 998680 372880 998704
rect 372914 998680 372948 998704
rect 372982 998680 373016 998704
rect 373050 998680 373084 998704
rect 373118 998680 373152 998704
rect 373186 998680 373220 998704
rect 373254 998680 373288 998704
rect 373322 998680 373356 998704
rect 373390 998680 373424 998704
rect 373458 998680 373492 998704
rect 373526 998680 373560 998704
rect 373594 998680 373628 998704
rect 373662 998680 373696 998704
rect 373796 998680 373830 998704
rect 373864 998680 373898 998704
rect 373932 998680 373966 998704
rect 374000 998680 374034 998704
rect 374068 998680 374102 998704
rect 374136 998680 374170 998704
rect 374204 998680 374238 998704
rect 374272 998680 374306 998704
rect 374340 998680 374374 998704
rect 374408 998680 374442 998704
rect 374476 998680 374510 998704
rect 374544 998680 374578 998704
rect 374612 998680 374646 998704
rect 374680 998680 374714 998704
rect 374748 998680 374782 998704
rect 374816 998680 374850 998704
rect 374884 998680 374918 998704
rect 374952 998680 374986 998704
rect 375020 998680 375054 998704
rect 375088 998680 375122 998704
rect 375156 998680 375190 998704
rect 375224 998680 375258 998704
rect 375292 998680 375326 998704
rect 375360 998680 375394 998704
rect 375428 998680 375462 998704
rect 375496 998680 375530 998704
rect 375564 998680 375598 998704
rect 375632 998680 375666 998704
rect 375700 998680 375734 998704
rect 375768 998680 375802 998704
rect 375836 998680 375870 998704
rect 375904 998680 375938 998704
rect 375972 998680 376006 998704
rect 376040 998680 376074 998704
rect 376108 998680 376142 998704
rect 376176 998680 376210 998704
rect 376244 998680 376278 998704
rect 376312 998680 376346 998704
rect 376380 998680 376414 998704
rect 376448 998680 376482 998704
rect 376516 998680 376550 998704
rect 376584 998680 376618 998704
rect 376652 998680 376686 998704
rect 376720 998680 376754 998704
rect 376788 998680 376822 998704
rect 376856 998680 376890 998704
rect 466318 998680 466352 998704
rect 466386 998680 466420 998704
rect 466454 998680 466488 998704
rect 466522 998680 466556 998704
rect 466590 998680 466624 998704
rect 466658 998680 466692 998704
rect 466726 998680 466760 998704
rect 466794 998680 466828 998704
rect 466862 998680 466896 998704
rect 466930 998680 466964 998704
rect 466998 998680 467032 998704
rect 467066 998680 467100 998704
rect 467134 998680 467168 998704
rect 467202 998680 467236 998704
rect 467270 998680 467304 998704
rect 467338 998680 467372 998704
rect 467406 998680 467440 998704
rect 467474 998680 467508 998704
rect 467542 998680 467576 998704
rect 467610 998680 467644 998704
rect 467678 998680 467712 998704
rect 467746 998680 467780 998704
rect 467814 998680 467848 998704
rect 467882 998680 467916 998704
rect 467950 998680 467984 998704
rect 468018 998680 468052 998704
rect 468086 998680 468120 998704
rect 468154 998680 468188 998704
rect 468222 998680 468256 998704
rect 468290 998680 468324 998704
rect 468358 998680 468392 998704
rect 468426 998680 468460 998704
rect 468494 998680 468528 998704
rect 468562 998680 468596 998704
rect 468630 998680 468664 998704
rect 468698 998680 468732 998704
rect 468766 998680 468800 998704
rect 468834 998680 468868 998704
rect 468902 998680 468936 998704
rect 468970 998680 469004 998704
rect 469038 998680 469072 998704
rect 469106 998680 469140 998704
rect 469174 998680 469208 998704
rect 469242 998680 469276 998704
rect 469310 998680 469344 998704
rect 469378 998680 469412 998704
rect 469446 998680 469480 998704
rect 469514 998680 469548 998704
rect 469582 998680 469616 998704
rect 469650 998680 469684 998704
rect 469718 998680 469752 998704
rect 469786 998680 469820 998704
rect 469854 998680 469888 998704
rect 469922 998680 469956 998704
rect 469990 998680 470024 998704
rect 470058 998680 470092 998704
rect 470126 998680 470160 998704
rect 470194 998680 470228 998704
rect 470262 998680 470296 998704
rect 470330 998680 470364 998704
rect 470398 998680 470432 998704
rect 470466 998680 470500 998704
rect 470534 998680 470568 998704
rect 470602 998680 470636 998704
rect 470670 998680 470704 998704
rect 470738 998680 470772 998704
rect 470806 998680 470840 998704
rect 470874 998680 470908 998704
rect 470942 998680 470976 998704
rect 471010 998680 471044 998704
rect 471078 998680 471112 998704
rect 471146 998680 471180 998704
rect 471214 998680 471248 998704
rect 471282 998680 471316 998704
rect 471350 998680 471384 998704
rect 471418 998680 471452 998704
rect 471486 998680 471520 998704
rect 471554 998680 471588 998704
rect 471622 998680 471656 998704
rect 471690 998680 471724 998704
rect 471758 998680 471792 998704
rect 471826 998680 471860 998704
rect 471894 998680 471928 998704
rect 471962 998680 471996 998704
rect 472030 998680 472064 998704
rect 472098 998680 472132 998704
rect 472166 998680 472200 998704
rect 472234 998680 472268 998704
rect 472302 998680 472336 998704
rect 472370 998680 472404 998704
rect 472438 998680 472472 998704
rect 472506 998680 472540 998704
rect 472574 998680 472608 998704
rect 472642 998680 472676 998704
rect 472710 998680 472744 998704
rect 472778 998680 472812 998704
rect 472846 998680 472880 998704
rect 472914 998680 472948 998704
rect 472982 998680 473016 998704
rect 473050 998680 473084 998704
rect 473118 998680 473152 998704
rect 473186 998680 473220 998704
rect 473254 998680 473288 998704
rect 473322 998680 473356 998704
rect 473390 998680 473424 998704
rect 473458 998680 473492 998704
rect 473526 998680 473560 998704
rect 473594 998680 473628 998704
rect 473662 998680 473696 998704
rect 473796 998680 473830 998704
rect 473864 998680 473898 998704
rect 473932 998680 473966 998704
rect 474000 998680 474034 998704
rect 474068 998680 474102 998704
rect 474136 998680 474170 998704
rect 474204 998680 474238 998704
rect 474272 998680 474306 998704
rect 474340 998680 474374 998704
rect 474408 998680 474442 998704
rect 474476 998680 474510 998704
rect 474544 998680 474578 998704
rect 474612 998680 474646 998704
rect 474680 998680 474714 998704
rect 474748 998680 474782 998704
rect 474816 998680 474850 998704
rect 474884 998680 474918 998704
rect 474952 998680 474986 998704
rect 475020 998680 475054 998704
rect 475088 998680 475122 998704
rect 475156 998680 475190 998704
rect 475224 998680 475258 998704
rect 475292 998680 475326 998704
rect 475360 998680 475394 998704
rect 475428 998680 475462 998704
rect 475496 998680 475530 998704
rect 475564 998680 475598 998704
rect 475632 998680 475666 998704
rect 475700 998680 475734 998704
rect 475768 998680 475802 998704
rect 475836 998680 475870 998704
rect 475904 998680 475938 998704
rect 475972 998680 476006 998704
rect 476040 998680 476074 998704
rect 476108 998680 476142 998704
rect 476176 998680 476210 998704
rect 476244 998680 476278 998704
rect 476312 998680 476346 998704
rect 476380 998680 476414 998704
rect 476448 998680 476482 998704
rect 476516 998680 476550 998704
rect 476584 998680 476618 998704
rect 476652 998680 476686 998704
rect 476720 998680 476754 998704
rect 476788 998680 476822 998704
rect 476856 998680 476890 998704
rect 570318 998680 570352 998704
rect 570386 998680 570420 998704
rect 570454 998680 570488 998704
rect 570522 998680 570556 998704
rect 570590 998680 570624 998704
rect 570658 998680 570692 998704
rect 570726 998680 570760 998704
rect 570794 998680 570828 998704
rect 570862 998680 570896 998704
rect 570930 998680 570964 998704
rect 570998 998680 571032 998704
rect 571066 998680 571100 998704
rect 571134 998680 571168 998704
rect 571202 998680 571236 998704
rect 571270 998680 571304 998704
rect 571338 998680 571372 998704
rect 571406 998680 571440 998704
rect 571474 998680 571508 998704
rect 571542 998680 571576 998704
rect 571610 998680 571644 998704
rect 571678 998680 571712 998704
rect 571746 998680 571780 998704
rect 571814 998680 571848 998704
rect 571882 998680 571916 998704
rect 571950 998680 571984 998704
rect 572018 998680 572052 998704
rect 572086 998680 572120 998704
rect 572154 998680 572188 998704
rect 572222 998680 572256 998704
rect 572290 998680 572324 998704
rect 572358 998680 572392 998704
rect 572426 998680 572460 998704
rect 572494 998680 572528 998704
rect 572562 998680 572596 998704
rect 572630 998680 572664 998704
rect 572698 998680 572732 998704
rect 572766 998680 572800 998704
rect 572834 998680 572868 998704
rect 572902 998680 572936 998704
rect 572970 998680 573004 998704
rect 573038 998680 573072 998704
rect 573106 998680 573140 998704
rect 573174 998680 573208 998704
rect 573242 998680 573276 998704
rect 573310 998680 573344 998704
rect 573378 998680 573412 998704
rect 573446 998680 573480 998704
rect 573514 998680 573548 998704
rect 573582 998680 573616 998704
rect 573650 998680 573684 998704
rect 573718 998680 573752 998704
rect 573786 998680 573820 998704
rect 573854 998680 573888 998704
rect 573922 998680 573956 998704
rect 573990 998680 574024 998704
rect 574058 998680 574092 998704
rect 574126 998680 574160 998704
rect 574194 998680 574228 998704
rect 574262 998680 574296 998704
rect 574330 998680 574364 998704
rect 574398 998680 574432 998704
rect 574466 998680 574500 998704
rect 574534 998680 574568 998704
rect 574602 998680 574636 998704
rect 574670 998680 574704 998704
rect 574738 998680 574772 998704
rect 574806 998680 574840 998704
rect 574874 998680 574908 998704
rect 574942 998680 574976 998704
rect 575010 998680 575044 998704
rect 575078 998680 575112 998704
rect 575146 998680 575180 998704
rect 575214 998680 575248 998704
rect 575282 998680 575316 998704
rect 575350 998680 575384 998704
rect 575418 998680 575452 998704
rect 575486 998680 575520 998704
rect 575554 998680 575588 998704
rect 575622 998680 575656 998704
rect 575690 998680 575724 998704
rect 575758 998680 575792 998704
rect 575826 998680 575860 998704
rect 575894 998680 575928 998704
rect 575962 998680 575996 998704
rect 576030 998680 576064 998704
rect 576098 998680 576132 998704
rect 576166 998680 576200 998704
rect 576234 998680 576268 998704
rect 576302 998680 576336 998704
rect 576370 998680 576404 998704
rect 576438 998680 576472 998704
rect 576506 998680 576540 998704
rect 576574 998680 576608 998704
rect 576642 998680 576676 998704
rect 576710 998680 576744 998704
rect 576778 998680 576812 998704
rect 576846 998680 576880 998704
rect 576914 998680 576948 998704
rect 576982 998680 577016 998704
rect 577050 998680 577084 998704
rect 577118 998680 577152 998704
rect 577186 998680 577220 998704
rect 577254 998680 577288 998704
rect 577322 998680 577356 998704
rect 577390 998680 577424 998704
rect 577458 998680 577492 998704
rect 577526 998680 577560 998704
rect 577594 998680 577628 998704
rect 577662 998680 577696 998704
rect 577796 998680 577830 998704
rect 577864 998680 577898 998704
rect 577932 998680 577966 998704
rect 578000 998680 578034 998704
rect 578068 998680 578102 998704
rect 578136 998680 578170 998704
rect 578204 998680 578238 998704
rect 578272 998680 578306 998704
rect 578340 998680 578374 998704
rect 578408 998680 578442 998704
rect 578476 998680 578510 998704
rect 578544 998680 578578 998704
rect 578612 998680 578646 998704
rect 578680 998680 578714 998704
rect 578748 998680 578782 998704
rect 578816 998680 578850 998704
rect 578884 998680 578918 998704
rect 578952 998680 578986 998704
rect 579020 998680 579054 998704
rect 579088 998680 579122 998704
rect 579156 998680 579190 998704
rect 579224 998680 579258 998704
rect 579292 998680 579326 998704
rect 579360 998680 579394 998704
rect 579428 998680 579462 998704
rect 579496 998680 579530 998704
rect 579564 998680 579598 998704
rect 579632 998680 579666 998704
rect 579700 998680 579734 998704
rect 579768 998680 579802 998704
rect 579836 998680 579870 998704
rect 579904 998680 579938 998704
rect 579972 998680 580006 998704
rect 580040 998680 580074 998704
rect 580108 998680 580142 998704
rect 580176 998680 580210 998704
rect 580244 998680 580278 998704
rect 580312 998680 580346 998704
rect 580380 998680 580414 998704
rect 580448 998680 580482 998704
rect 580516 998680 580550 998704
rect 580584 998680 580618 998704
rect 580652 998680 580686 998704
rect 580720 998680 580754 998704
rect 580788 998680 580822 998704
rect 580856 998680 580890 998704
rect 69746 998654 69772 998680
rect 169746 998654 169772 998680
rect 373746 998654 373772 998680
rect 473746 998654 473772 998680
rect 577746 998654 577772 998680
rect 21000 997600 21003 997720
rect 696597 996800 696600 996920
rect 21000 981800 21003 981920
rect 282 981423 1316 981505
rect 1602 981423 2636 981505
rect 32810 981462 33035 981470
rect 38201 981393 38801 981443
rect 24572 981318 25172 981368
rect 33292 981313 33892 981363
rect 99 979374 181 981292
rect 452 981131 1146 981213
rect 381 979685 463 980991
rect 660 980928 700 980968
rect 900 980928 940 980968
rect 700 980844 740 980928
rect 860 980844 900 980928
rect 607 979881 657 980823
rect 951 979881 1001 980823
rect 1133 979685 1215 980991
rect 452 979563 1146 979645
rect 1418 979374 1500 981292
rect 1772 981131 2466 981213
rect 1703 979685 1785 980991
rect 1978 980928 2018 980968
rect 2218 980928 2258 980968
rect 2018 980844 2058 980928
rect 2178 980844 2218 980928
rect 1917 979881 1967 980823
rect 2261 979881 2311 980823
rect 2455 979685 2537 980991
rect 2737 980579 2819 981292
rect 24572 981162 25172 981290
rect 38201 981217 38801 981273
rect 33292 981163 33892 981213
rect 24572 981006 25172 981134
rect 35546 981099 35576 981135
rect 36785 981129 36935 981141
rect 35531 981084 35591 981099
rect 36785 981016 37385 981066
rect 38201 981047 38801 981097
rect 30833 980920 30857 980944
rect 30891 980920 30915 980944
rect 24572 980850 25172 980906
rect 30857 980905 30881 980907
rect 30857 980896 30887 980905
rect 30867 980883 30887 980896
rect 30891 980883 30907 980920
rect 30833 980859 30857 980883
rect 30867 980849 30911 980883
rect 14747 980665 19516 980772
rect 24572 980694 25172 980822
rect 30867 980812 30887 980849
rect 30891 980812 30907 980849
rect 36785 980840 37385 980896
rect 30867 980778 30911 980812
rect 30867 980741 30887 980778
rect 30891 980741 30907 980778
rect 30867 980707 30911 980741
rect 30867 980683 30887 980707
rect 30891 980683 30907 980707
rect 14747 980641 14844 980665
rect 13955 980617 14844 980641
rect 19390 980653 19516 980665
rect 19390 980641 19583 980653
rect 19390 980617 19605 980641
rect 19639 980617 19673 980641
rect 19707 980617 19741 980641
rect 19775 980617 19809 980641
rect 19843 980617 19877 980641
rect 19911 980617 19945 980641
rect 19979 980617 20013 980641
rect 20047 980617 20081 980641
rect 20115 980617 20149 980641
rect 20183 980617 20217 980641
rect 20251 980617 20285 980641
rect 20319 980617 20353 980641
rect 20387 980617 20421 980641
rect 20455 980617 20489 980641
rect 20523 980617 20557 980641
rect 20591 980617 20625 980641
rect 20659 980617 20693 980641
rect 2737 980511 2914 980579
rect 1772 979563 2466 979645
rect 2737 979374 2819 980511
rect 2848 980477 2955 980511
rect 19480 980340 19516 980617
rect 19547 980340 19583 980617
rect 24572 980538 25172 980666
rect 36785 980664 37385 980720
rect 36785 980488 37385 980544
rect 20809 980450 20833 980484
rect 20809 980382 20833 980416
rect 24572 980388 25172 980438
rect 20809 980340 20833 980348
rect 36785 980318 37385 980368
rect 3125 979602 3175 980202
rect 3375 979602 3425 980202
rect 282 979271 1316 979353
rect 1602 979271 2636 979353
rect 1389 979244 1392 979245
rect 1389 979243 1390 979244
rect 1391 979243 1392 979244
rect 1389 979242 1392 979243
rect 1526 979244 1529 979245
rect 1526 979243 1527 979244
rect 1528 979243 1529 979244
rect 2848 979243 2955 979277
rect 1526 979242 1529 979243
rect 5488 979080 5538 979903
rect 5658 979080 5708 979903
rect 6005 979080 6021 980299
rect 12427 980248 12493 980264
rect 24572 980258 25172 980308
rect 32930 980257 33530 980307
rect 35287 980191 35887 980241
rect 36785 980202 37385 980252
rect 24572 980108 25172 980158
rect 31463 980107 32063 980157
rect 32930 980101 33530 980157
rect 7389 980077 7406 980087
rect 7440 980077 7477 980087
rect 7511 980077 7551 980087
rect 7585 980077 7622 980087
rect 7656 980077 7696 980087
rect 7730 980077 7767 980087
rect 7801 980077 7841 980087
rect 7875 980077 7912 980087
rect 7946 980077 7986 980087
rect 8020 980077 8057 980087
rect 8091 980077 8131 980087
rect 8165 980077 8202 980087
rect 8236 980077 8296 980087
rect 8330 980077 8381 980087
rect 8996 980077 9044 980087
rect 9078 980077 9120 980087
rect 9154 980077 9197 980087
rect 9231 980077 9291 980087
rect 9325 980077 9362 980087
rect 9396 980077 9436 980087
rect 9470 980077 9507 980087
rect 9541 980077 9581 980087
rect 9615 980077 9652 980087
rect 9686 980077 9726 980087
rect 9760 980077 9797 980087
rect 9831 980077 9871 980087
rect 9905 980077 9942 980087
rect 9976 980077 9990 980087
rect 7389 980009 8389 980077
rect 8990 979983 9990 980077
rect 36785 980026 37385 980082
rect 15678 979927 16678 979977
rect 17278 979927 18278 979977
rect 31463 979951 32063 980007
rect 32930 979951 33530 980001
rect 34079 979957 34679 980007
rect 7389 979640 8389 979664
rect 15678 979660 16678 979716
rect 17278 979660 18278 979716
rect 8990 979640 9990 979641
rect 7389 979543 8389 979599
rect 8990 979543 9990 979599
rect 15678 979588 16678 979644
rect 17278 979588 18278 979644
rect 8990 979501 9990 979502
rect 15678 979086 16678 979226
rect 17278 979086 18278 979226
rect 19844 979080 19894 979851
rect 20462 979080 20512 979851
rect 31463 979801 32063 979851
rect 34079 979801 34679 979857
rect 35287 979839 35887 979895
rect 36785 979850 37385 979906
rect 32596 979729 33596 979779
rect 24573 979620 25173 979670
rect 34079 979651 34679 979701
rect 35287 979669 35887 979719
rect 36785 979680 37385 979730
rect 30171 979595 30771 979645
rect 32596 979573 33596 979629
rect 37993 979504 38593 979554
rect 30171 979419 30771 979475
rect 32596 979423 33596 979473
rect 34110 979389 34710 979439
rect 21263 979080 21313 979318
rect 22349 979080 22399 979318
rect 32596 979307 33596 979357
rect 30171 979249 30771 979299
rect 36785 979229 36985 979409
rect 37993 979334 38593 979384
rect 24573 979152 25173 979208
rect 29993 979110 30993 979160
rect 31347 979080 31547 979117
rect 31607 979080 31807 979117
rect 36785 979080 36985 979173
rect 37083 979080 37120 979173
rect 696597 977000 696600 977120
rect 692376 976783 692396 976817
rect 692463 976793 692532 976817
rect 696191 976793 696239 976817
rect 692487 976783 692532 976793
rect 696204 976783 696239 976793
rect 696340 976783 696360 976817
rect 692487 976715 692502 976739
rect 696200 976715 696215 976739
rect 692454 976691 692478 976715
rect 696224 976691 696248 976715
rect 686755 976600 687355 976650
rect 692487 976548 692505 976552
rect 692479 976518 692505 976548
rect 692487 976498 692505 976518
rect 686755 976424 687355 976480
rect 692485 976474 692505 976498
rect 692509 976474 692517 976518
rect 696215 976498 696223 976548
rect 696203 976474 696223 976498
rect 696227 976474 696245 976552
rect 692485 976440 692521 976474
rect 696203 976440 696249 976474
rect 686755 976248 687355 976304
rect 686755 976078 687355 976128
rect 685547 975902 686147 975952
rect 687155 975807 687170 975822
rect 687343 975818 687355 975822
rect 687340 975807 687355 975818
rect 685547 975732 686147 975782
rect 687155 975627 687355 975807
rect 687155 975612 687170 975627
rect 687340 975616 687355 975627
rect 687343 975612 687355 975616
rect 687042 975571 687057 975586
rect 687020 975391 687057 975571
rect 687155 975571 687170 975586
rect 687343 975582 687355 975586
rect 687340 975571 687355 975582
rect 687155 975391 687355 975571
rect 688210 975430 688260 976430
rect 688360 975540 688488 976430
rect 688516 975540 688644 976430
rect 688672 975540 688800 976430
rect 688828 975540 688956 976430
rect 688984 975540 689112 976430
rect 689140 975540 689268 976430
rect 689296 975540 689424 976430
rect 689452 975540 689580 976430
rect 689608 975540 689736 976430
rect 689764 975540 689892 976430
rect 689920 975540 690048 976430
rect 690076 975540 690204 976430
rect 690232 975540 690360 976430
rect 690388 975430 690438 976430
rect 692485 976406 692505 976440
rect 692509 976406 692517 976440
rect 696203 976406 696223 976440
rect 696227 976406 696245 976440
rect 691275 976323 691875 976373
rect 692485 976372 692521 976406
rect 696203 976372 696249 976406
rect 692485 976338 692505 976372
rect 692509 976338 692517 976372
rect 692485 976304 692521 976338
rect 692583 976328 693983 976371
rect 694719 976328 696119 976371
rect 696203 976338 696223 976372
rect 696227 976338 696245 976372
rect 696203 976304 696249 976338
rect 692485 976270 692505 976304
rect 692509 976270 692517 976304
rect 692485 976236 692521 976270
rect 691275 976173 691875 976223
rect 692485 976202 692505 976236
rect 692509 976202 692517 976236
rect 692485 976168 692521 976202
rect 692485 976134 692505 976168
rect 692509 976134 692517 976168
rect 692583 976165 693983 976293
rect 694719 976165 696119 976293
rect 696203 976270 696223 976304
rect 696227 976270 696245 976304
rect 696203 976236 696249 976270
rect 707624 976241 707658 976275
rect 707695 976241 707729 976275
rect 707769 976241 707803 976275
rect 707840 976241 707874 976275
rect 707914 976241 707948 976275
rect 707985 976241 708019 976275
rect 708059 976241 708093 976275
rect 708130 976241 708164 976275
rect 708204 976241 708238 976275
rect 708275 976241 708309 976275
rect 708369 976241 708403 976275
rect 708446 976241 708480 976275
rect 708520 976241 708554 976265
rect 708588 976241 708610 976265
rect 709211 976241 709234 976265
rect 709270 976241 709304 976275
rect 709364 976241 709398 976275
rect 709435 976241 709469 976275
rect 709509 976241 709543 976275
rect 709580 976241 709614 976275
rect 709654 976241 709688 976275
rect 709725 976241 709759 976275
rect 709799 976241 709833 976275
rect 709870 976241 709904 976275
rect 709944 976241 709978 976275
rect 710015 976241 710049 976275
rect 710089 976241 710123 976275
rect 710160 976241 710194 976275
rect 696203 976202 696223 976236
rect 696227 976202 696245 976236
rect 707610 976231 707624 976241
rect 707658 976231 707695 976241
rect 707729 976231 707769 976241
rect 707803 976231 707840 976241
rect 707874 976231 707914 976241
rect 707948 976231 707985 976241
rect 708019 976231 708059 976241
rect 708093 976231 708130 976241
rect 708164 976231 708204 976241
rect 708238 976231 708275 976241
rect 708309 976231 708369 976241
rect 708403 976231 708446 976241
rect 708480 976231 708520 976241
rect 708554 976231 708588 976241
rect 708610 976231 708634 976241
rect 709211 976231 709270 976241
rect 709304 976231 709364 976241
rect 709398 976231 709435 976241
rect 709469 976231 709509 976241
rect 709543 976231 709580 976241
rect 709614 976231 709654 976241
rect 709688 976231 709725 976241
rect 709759 976231 709799 976241
rect 709833 976231 709870 976241
rect 709904 976231 709944 976241
rect 709978 976231 710015 976241
rect 710049 976231 710089 976241
rect 710123 976231 710160 976241
rect 710194 976231 710211 976241
rect 696203 976168 696249 976202
rect 696203 976134 696223 976168
rect 696227 976134 696245 976168
rect 707610 976137 708610 976231
rect 709211 976137 710211 976231
rect 691275 976051 691875 976101
rect 692485 976100 692521 976134
rect 692485 976066 692505 976100
rect 692509 976066 692517 976100
rect 692485 976032 692521 976066
rect 692485 975998 692505 976032
rect 692509 975998 692517 976032
rect 692583 976002 693983 976130
rect 694719 976002 696119 976130
rect 696203 976100 696249 976134
rect 711579 976117 712463 976131
rect 711579 976107 711619 976117
rect 696203 976066 696223 976100
rect 696227 976066 696245 976100
rect 701730 976090 701747 976092
rect 696203 976032 696249 976066
rect 696203 975998 696223 976032
rect 696227 975998 696245 976032
rect 701692 976020 701722 976054
rect 701730 976020 701760 976090
rect 707610 976041 708610 976101
rect 709211 976041 710211 976101
rect 692485 975964 692521 975998
rect 691275 975901 691875 975951
rect 692485 975930 692505 975964
rect 692509 975930 692517 975964
rect 692485 975896 692521 975930
rect 692485 975862 692505 975896
rect 692509 975862 692517 975896
rect 692485 975828 692521 975862
rect 692583 975839 693983 975967
rect 694719 975839 696119 975967
rect 696203 975964 696249 975998
rect 696203 975930 696223 975964
rect 696227 975930 696245 975964
rect 696203 975896 696249 975930
rect 696203 975862 696223 975896
rect 696227 975862 696245 975896
rect 699322 975864 700322 975897
rect 700922 975864 701922 975897
rect 696203 975828 696249 975862
rect 707610 975844 708610 975848
rect 709211 975844 710211 975848
rect 691275 975775 691875 975825
rect 692485 975794 692505 975828
rect 692509 975794 692517 975828
rect 692485 975760 692521 975794
rect 692485 975726 692505 975760
rect 692509 975726 692517 975760
rect 692485 975692 692521 975726
rect 691275 975625 691875 975675
rect 692485 975658 692505 975692
rect 692509 975658 692517 975692
rect 692583 975676 693983 975804
rect 694719 975676 696119 975804
rect 696203 975794 696223 975828
rect 696227 975794 696245 975828
rect 707574 975794 708646 975830
rect 696203 975760 696249 975794
rect 696203 975726 696223 975760
rect 696227 975726 696245 975760
rect 707574 975753 707610 975794
rect 708610 975753 708646 975794
rect 696203 975692 696249 975726
rect 697284 975694 697350 975710
rect 707574 975697 708646 975753
rect 696203 975658 696223 975692
rect 696227 975658 696245 975692
rect 699322 975677 700322 975694
rect 700922 975677 701922 975694
rect 707574 975681 707610 975697
rect 708610 975681 708646 975697
rect 692485 975624 692521 975658
rect 692485 975590 692505 975624
rect 692509 975590 692517 975624
rect 692485 975556 692521 975590
rect 691275 975503 691875 975553
rect 692485 975540 692505 975556
rect 692509 975540 692517 975556
rect 692583 975540 693983 975641
rect 694719 975540 696119 975641
rect 696203 975624 696249 975658
rect 707574 975625 708646 975681
rect 696203 975590 696223 975624
rect 696227 975590 696245 975624
rect 696203 975556 696249 975590
rect 696203 975540 696223 975556
rect 696227 975540 696245 975556
rect 699322 975540 700322 975611
rect 700922 975540 701922 975611
rect 707574 975588 707610 975625
rect 708610 975588 708646 975625
rect 707574 975548 708646 975588
rect 709175 975794 710247 975830
rect 709175 975753 709211 975794
rect 710211 975753 710247 975794
rect 709175 975697 710247 975753
rect 709175 975681 709211 975697
rect 710211 975681 710247 975697
rect 709175 975625 710247 975681
rect 709175 975588 709211 975625
rect 710211 975588 710247 975625
rect 709175 975548 710247 975588
rect 685542 975306 686142 975356
rect 691275 975353 691875 975403
rect 685542 975130 686142 975186
rect 692583 975037 693983 975080
rect 694719 975037 696119 975080
rect 699322 975078 700322 975218
rect 700922 975078 701922 975218
rect 685542 974960 686142 975010
rect 692583 974901 693983 974944
rect 694719 974901 696119 974944
rect 680215 974478 680815 974528
rect 680215 974302 680815 974358
rect 685551 974316 686551 974366
rect 689154 974280 689204 974697
rect 689304 974280 689360 974697
rect 689460 974280 689516 974697
rect 689616 974280 689672 974697
rect 689772 974280 689828 974697
rect 689928 974280 689978 974697
rect 699322 974660 700322 974716
rect 700922 974660 701922 974716
rect 707610 974705 708610 974761
rect 709211 974705 710211 974761
rect 699322 974588 700322 974644
rect 700922 974588 701922 974644
rect 707610 974633 708610 974689
rect 709211 974633 710211 974689
rect 711579 974325 711605 976107
rect 715956 975097 716006 976097
rect 716106 975540 716234 976097
rect 716262 975097 716312 976097
rect 711579 974280 711595 974295
rect 712409 974280 712431 974285
rect 713640 974280 713641 974585
rect 713750 974572 714750 974622
rect 713750 974362 714750 974412
rect 713750 974280 714750 974296
rect 2850 895304 3850 895320
rect 2850 895188 3850 895238
rect 2850 894978 3850 895028
rect 3959 895015 3960 895320
rect 5169 895315 5191 895320
rect 6005 895305 6021 895320
rect 1288 893503 1338 894503
rect 1438 893503 1566 894060
rect 1594 893503 1644 894503
rect 5995 893493 6021 895275
rect 7389 894911 8389 894967
rect 8990 894911 9990 894967
rect 15678 894956 16678 895012
rect 17278 894956 18278 895012
rect 7389 894839 8389 894895
rect 8990 894839 9990 894895
rect 15678 894884 16678 894940
rect 17278 894884 18278 894940
rect 27622 894903 27672 895320
rect 27772 894903 27828 895320
rect 27928 894903 27984 895320
rect 28084 894903 28140 895320
rect 28240 894903 28296 895320
rect 28396 894903 28446 895320
rect 31049 895234 32049 895284
rect 36785 895242 37385 895298
rect 36785 895072 37385 895122
rect 21481 894656 22881 894699
rect 23617 894656 25017 894699
rect 31458 894590 32058 894640
rect 15678 894382 16678 894522
rect 17278 894382 18278 894522
rect 21481 894520 22881 894563
rect 23617 894520 25017 894563
rect 31458 894414 32058 894470
rect 25725 894197 26325 894247
rect 31458 894244 32058 894294
rect 7353 894016 8425 894052
rect 7353 893975 7389 894016
rect 8389 893975 8425 894016
rect 7353 893919 8425 893975
rect 7353 893903 7389 893919
rect 8389 893903 8425 893919
rect 7353 893847 8425 893903
rect 7353 893810 7389 893847
rect 8389 893810 8425 893847
rect 7353 893770 8425 893810
rect 8954 894016 10026 894052
rect 8954 893975 8990 894016
rect 9990 893975 10026 894016
rect 8954 893919 10026 893975
rect 21383 894044 21403 894060
rect 21407 894044 21415 894060
rect 21383 894010 21419 894044
rect 21481 894031 22881 894060
rect 23617 894031 25017 894060
rect 25101 894044 25121 894060
rect 25125 894044 25143 894060
rect 25725 894047 26325 894097
rect 25101 894010 25147 894044
rect 21383 893976 21403 894010
rect 21407 893976 21415 894010
rect 21383 893942 21419 893976
rect 8954 893903 8990 893919
rect 9990 893903 10026 893919
rect 15678 893906 16678 893923
rect 17278 893906 18278 893923
rect 21383 893908 21403 893942
rect 21407 893908 21415 893942
rect 8954 893847 10026 893903
rect 20250 893890 20316 893906
rect 8954 893810 8990 893847
rect 9990 893810 10026 893847
rect 8954 893770 10026 893810
rect 21383 893874 21419 893908
rect 21383 893840 21403 893874
rect 21407 893840 21415 893874
rect 21481 893868 22881 893996
rect 23617 893868 25017 893996
rect 25101 893976 25121 894010
rect 25125 893976 25143 894010
rect 25101 893942 25147 893976
rect 25101 893908 25121 893942
rect 25125 893908 25143 893942
rect 25725 893925 26325 893975
rect 25101 893874 25147 893908
rect 25101 893840 25121 893874
rect 25125 893840 25143 893874
rect 21383 893806 21419 893840
rect 21383 893772 21403 893806
rect 21407 893772 21415 893806
rect 21383 893738 21419 893772
rect 15678 893703 16678 893736
rect 17278 893703 18278 893736
rect 21383 893704 21403 893738
rect 21407 893704 21415 893738
rect 21481 893705 22881 893833
rect 23617 893705 25017 893833
rect 25101 893806 25147 893840
rect 25101 893772 25121 893806
rect 25125 893772 25143 893806
rect 25725 893775 26325 893825
rect 25101 893738 25147 893772
rect 25101 893704 25121 893738
rect 25125 893704 25143 893738
rect 21383 893670 21419 893704
rect 25101 893670 25147 893704
rect 21383 893636 21403 893670
rect 21407 893636 21415 893670
rect 7389 893559 8389 893631
rect 8990 893559 9990 893631
rect 21383 893602 21419 893636
rect 15840 893510 15870 893580
rect 15878 893546 15908 893580
rect 21383 893568 21403 893602
rect 21407 893568 21415 893602
rect 15853 893508 15870 893510
rect 21383 893534 21419 893568
rect 21481 893542 22881 893670
rect 23617 893542 25017 893670
rect 25101 893636 25121 893670
rect 25125 893636 25143 893670
rect 25725 893649 26325 893699
rect 25101 893602 25147 893636
rect 25101 893568 25121 893602
rect 25125 893568 25143 893602
rect 25101 893534 25147 893568
rect 5981 893483 6021 893493
rect 5137 893469 6021 893483
rect 21383 893500 21403 893534
rect 21407 893500 21415 893534
rect 21383 893466 21419 893500
rect 7389 893369 8389 893463
rect 7389 893359 8413 893369
rect 8990 893359 9990 893463
rect 21383 893432 21403 893466
rect 21407 893432 21415 893466
rect 21383 893398 21419 893432
rect 21383 893364 21403 893398
rect 21407 893364 21415 893398
rect 21481 893379 22881 893507
rect 23617 893379 25017 893507
rect 25101 893500 25121 893534
rect 25125 893500 25143 893534
rect 25101 893466 25147 893500
rect 25725 893499 26325 893549
rect 25101 893432 25121 893466
rect 25125 893432 25143 893466
rect 25101 893398 25147 893432
rect 25101 893364 25121 893398
rect 25125 893364 25143 893398
rect 25725 893377 26325 893427
rect 21383 893330 21419 893364
rect 25101 893330 25147 893364
rect 21383 893296 21403 893330
rect 21407 893296 21415 893330
rect 25101 893296 25121 893330
rect 25125 893296 25143 893330
rect 21383 893262 21419 893296
rect 21383 893228 21403 893262
rect 21407 893228 21415 893262
rect 21481 893229 22881 893272
rect 23617 893229 25017 893272
rect 25101 893262 25147 893296
rect 25101 893228 25121 893262
rect 25125 893228 25143 893262
rect 21383 893194 21419 893228
rect 25101 893194 25147 893228
rect 25725 893227 26325 893277
rect 21383 893160 21403 893194
rect 21407 893160 21415 893194
rect 25101 893160 25121 893194
rect 25125 893160 25143 893194
rect 27162 893170 27212 894170
rect 27312 893170 27440 894060
rect 27468 893170 27596 894060
rect 27624 893170 27752 894060
rect 27780 893170 27908 894060
rect 27936 893170 28064 894060
rect 28092 893170 28220 894060
rect 28248 893170 28376 894060
rect 28404 893170 28532 894060
rect 28560 893170 28688 894060
rect 28716 893170 28844 894060
rect 28872 893170 29000 894060
rect 29028 893170 29156 894060
rect 29184 893170 29312 894060
rect 29340 893170 29390 894170
rect 30245 894029 30445 894209
rect 30245 894018 30260 894029
rect 30245 894014 30257 894018
rect 30430 894014 30445 894029
rect 30543 894029 30580 894209
rect 30543 894014 30558 894029
rect 30245 893984 30257 893988
rect 30245 893973 30260 893984
rect 30430 893973 30445 893988
rect 30245 893793 30445 893973
rect 31453 893818 32053 893868
rect 30245 893782 30260 893793
rect 30245 893778 30257 893782
rect 30430 893778 30445 893793
rect 31453 893648 32053 893698
rect 30245 893472 30845 893522
rect 30245 893296 30845 893352
rect 21383 893126 21419 893160
rect 25101 893126 25147 893160
rect 21383 893102 21403 893126
rect 21385 893048 21403 893102
rect 21407 893082 21415 893126
rect 25101 893102 25121 893126
rect 25113 893082 25121 893102
rect 25125 893048 25143 893126
rect 30245 893120 30845 893176
rect 30245 892950 30845 893000
rect 21000 892800 21003 892920
rect 21352 892885 21376 892909
rect 25122 892885 25146 892909
rect 21385 892861 21400 892885
rect 25098 892861 25113 892885
rect 21274 892783 21294 892851
rect 21410 892817 21430 892851
rect 25068 892817 25088 892851
rect 25204 892817 25224 892851
rect 21385 892807 21430 892817
rect 25102 892807 25137 892817
rect 21361 892783 21430 892807
rect 25089 892783 25137 892807
rect 25238 892783 25258 892817
rect 680480 890427 680517 890520
rect 680615 890427 680815 890520
rect 685793 890483 685993 890520
rect 686053 890483 686253 890520
rect 686607 890440 687607 890490
rect 692427 890392 693027 890448
rect 679007 890216 679607 890266
rect 680615 890191 680815 890371
rect 686829 890301 687429 890351
rect 684004 890243 685004 890293
rect 695201 890282 695251 890520
rect 696287 890282 696337 890520
rect 682890 890161 683490 890211
rect 684004 890127 685004 890177
rect 686829 890125 687429 890181
rect 679007 890046 679607 890096
rect 684004 889971 685004 890027
rect 686829 889955 687429 890005
rect 680215 889870 680815 889920
rect 681713 889881 682313 889931
rect 682921 889899 683521 889949
rect 692427 889930 693027 889980
rect 684004 889821 685004 889871
rect 680215 889694 680815 889750
rect 681713 889705 682313 889761
rect 682921 889743 683521 889799
rect 685537 889749 686137 889799
rect 697088 889749 697138 890520
rect 697706 889749 697756 890520
rect 699322 890374 700322 890514
rect 700922 890374 701922 890514
rect 707610 890098 708610 890099
rect 699322 889956 700322 890012
rect 700922 889956 701922 890012
rect 707610 890001 708610 890057
rect 709211 890001 710211 890057
rect 707610 889959 708610 889960
rect 699322 889884 700322 889940
rect 700922 889884 701922 889940
rect 709211 889936 710211 889960
rect 682921 889593 683521 889643
rect 684070 889599 684670 889649
rect 685537 889593 686137 889649
rect 699322 889623 700322 889673
rect 700922 889623 701922 889673
rect 680215 889518 680815 889574
rect 707610 889523 708610 889617
rect 709211 889523 710211 889591
rect 707610 889513 707624 889523
rect 707658 889513 707695 889523
rect 707729 889513 707769 889523
rect 707803 889513 707840 889523
rect 707874 889513 707914 889523
rect 707948 889513 707985 889523
rect 708019 889513 708059 889523
rect 708093 889513 708130 889523
rect 708164 889513 708204 889523
rect 708238 889513 708275 889523
rect 708309 889513 708369 889523
rect 708403 889513 708446 889523
rect 708480 889513 708522 889523
rect 708556 889513 708604 889523
rect 709219 889513 709270 889523
rect 709304 889513 709364 889523
rect 709398 889513 709435 889523
rect 709469 889513 709509 889523
rect 709543 889513 709580 889523
rect 709614 889513 709654 889523
rect 709688 889513 709725 889523
rect 709759 889513 709799 889523
rect 709833 889513 709870 889523
rect 709904 889513 709944 889523
rect 709978 889513 710015 889523
rect 710049 889513 710089 889523
rect 710123 889513 710160 889523
rect 710194 889513 710211 889523
rect 684070 889443 684670 889499
rect 685537 889443 686137 889493
rect 692428 889442 693028 889492
rect 680215 889348 680815 889398
rect 681713 889359 682313 889409
rect 684070 889293 684670 889343
rect 692428 889292 693028 889342
rect 705107 889336 705173 889352
rect 711579 889301 711595 890520
rect 711892 889697 711942 890520
rect 712062 889697 712112 890520
rect 716071 890357 716074 890358
rect 714645 890323 714752 890357
rect 716071 890356 716072 890357
rect 716073 890356 716074 890357
rect 716071 890355 716074 890356
rect 716208 890357 716211 890358
rect 716208 890356 716209 890357
rect 716210 890356 716211 890357
rect 716208 890355 716211 890356
rect 714964 890247 715998 890329
rect 716284 890247 717318 890329
rect 714175 889398 714225 889998
rect 714425 889398 714475 889998
rect 680215 889232 680815 889282
rect 698017 889232 698053 889260
rect 692428 889162 693028 889212
rect 698030 889198 698077 889232
rect 698017 889164 698053 889198
rect 680215 889056 680815 889112
rect 692428 889006 693028 889134
rect 698030 889130 698077 889164
rect 698017 889096 698053 889130
rect 698030 889062 698077 889096
rect 698017 888983 698053 889062
rect 698084 888983 698120 889260
rect 714781 889191 714863 890226
rect 715134 889955 715828 890037
rect 714686 889123 714863 889191
rect 714645 889089 714863 889123
rect 680215 888880 680815 888936
rect 686719 888893 686739 888917
rect 686743 888893 686753 888917
rect 686719 888859 686757 888893
rect 686719 888822 686739 888859
rect 686743 888822 686753 888859
rect 692428 888850 693028 888978
rect 698017 888947 698210 888983
rect 698084 888935 698210 888947
rect 702756 888959 703645 888983
rect 702756 888935 702853 888959
rect 698084 888828 702853 888935
rect 686719 888788 686757 888822
rect 680215 888704 680815 888760
rect 686719 888751 686739 888788
rect 686743 888751 686753 888788
rect 686719 888741 686757 888751
rect 686699 888717 686767 888741
rect 686719 888704 686739 888717
rect 686743 888704 686753 888717
rect 686719 888695 686753 888704
rect 686719 888693 686743 888695
rect 692428 888694 693028 888750
rect 686685 888656 686709 888680
rect 686743 888656 686767 888680
rect 678799 888503 679399 888553
rect 680215 888534 680815 888584
rect 692428 888538 693028 888666
rect 680593 888531 680815 888534
rect 682009 888501 682069 888516
rect 682024 888465 682054 888501
rect 683708 888387 684308 888437
rect 678799 888327 679399 888383
rect 692428 888382 693028 888510
rect 714781 888308 714863 889089
rect 715063 888609 715145 889915
rect 715289 888777 715339 889719
rect 715633 888777 715683 889719
rect 715382 888672 715422 888756
rect 715542 888672 715582 888756
rect 715342 888632 715382 888672
rect 715582 888632 715622 888672
rect 715815 888609 715897 889915
rect 715134 888387 715828 888469
rect 716100 888308 716182 890226
rect 716454 889955 717148 890037
rect 716385 888609 716467 889915
rect 716599 888777 716649 889719
rect 716943 888777 716993 889719
rect 716700 888672 716740 888756
rect 716860 888672 716900 888756
rect 716660 888632 716700 888672
rect 716900 888632 716940 888672
rect 717137 888609 717219 889915
rect 716454 888387 717148 888469
rect 717419 888308 717501 890226
rect 683708 888237 684308 888287
rect 692428 888232 693028 888282
rect 678799 888157 679399 888207
rect 684565 888160 684790 888168
rect 696597 888000 696600 888120
rect 714964 888095 715998 888177
rect 716284 888095 717318 888177
rect 21000 861000 21003 861120
rect 282 860623 1316 860705
rect 1602 860623 2636 860705
rect 32810 860662 33035 860670
rect 38201 860593 38801 860643
rect 24572 860518 25172 860568
rect 33292 860513 33892 860563
rect 99 858574 181 860492
rect 452 860331 1146 860413
rect 381 858885 463 860191
rect 660 860128 700 860168
rect 900 860128 940 860168
rect 700 860044 740 860128
rect 860 860044 900 860128
rect 607 859081 657 860023
rect 951 859081 1001 860023
rect 1133 858885 1215 860191
rect 452 858763 1146 858845
rect 1418 858574 1500 860492
rect 1772 860331 2466 860413
rect 1703 858885 1785 860191
rect 1978 860128 2018 860168
rect 2218 860128 2258 860168
rect 2018 860044 2058 860128
rect 2178 860044 2218 860128
rect 1917 859081 1967 860023
rect 2261 859081 2311 860023
rect 2455 858885 2537 860191
rect 2737 859779 2819 860492
rect 24572 860362 25172 860490
rect 38201 860417 38801 860473
rect 33292 860363 33892 860413
rect 24572 860206 25172 860334
rect 35546 860299 35576 860335
rect 36785 860329 36935 860341
rect 35531 860284 35591 860299
rect 36785 860216 37385 860266
rect 38201 860247 38801 860297
rect 30833 860120 30857 860144
rect 30891 860120 30915 860144
rect 24572 860050 25172 860106
rect 30857 860105 30881 860107
rect 30857 860096 30887 860105
rect 30867 860083 30887 860096
rect 30891 860083 30907 860120
rect 30833 860059 30857 860083
rect 30867 860049 30911 860083
rect 14747 859865 19516 859972
rect 24572 859894 25172 860022
rect 30867 860012 30887 860049
rect 30891 860012 30907 860049
rect 36785 860040 37385 860096
rect 30867 859978 30911 860012
rect 30867 859941 30887 859978
rect 30891 859941 30907 859978
rect 30867 859907 30911 859941
rect 30867 859883 30887 859907
rect 30891 859883 30907 859907
rect 14747 859841 14844 859865
rect 13955 859817 14844 859841
rect 19390 859853 19516 859865
rect 19390 859841 19583 859853
rect 19390 859817 19605 859841
rect 19639 859817 19673 859841
rect 19707 859817 19741 859841
rect 19775 859817 19809 859841
rect 19843 859817 19877 859841
rect 19911 859817 19945 859841
rect 19979 859817 20013 859841
rect 20047 859817 20081 859841
rect 20115 859817 20149 859841
rect 20183 859817 20217 859841
rect 20251 859817 20285 859841
rect 20319 859817 20353 859841
rect 20387 859817 20421 859841
rect 20455 859817 20489 859841
rect 20523 859817 20557 859841
rect 20591 859817 20625 859841
rect 20659 859817 20693 859841
rect 2737 859711 2914 859779
rect 1772 858763 2466 858845
rect 2737 858574 2819 859711
rect 2848 859677 2955 859711
rect 19480 859540 19516 859817
rect 19547 859540 19583 859817
rect 24572 859738 25172 859866
rect 36785 859864 37385 859920
rect 36785 859688 37385 859744
rect 20809 859650 20833 859684
rect 20809 859582 20833 859616
rect 24572 859588 25172 859638
rect 20809 859540 20833 859548
rect 36785 859518 37385 859568
rect 3125 858802 3175 859402
rect 3375 858802 3425 859402
rect 282 858471 1316 858553
rect 1602 858471 2636 858553
rect 1389 858444 1392 858445
rect 1389 858443 1390 858444
rect 1391 858443 1392 858444
rect 1389 858442 1392 858443
rect 1526 858444 1529 858445
rect 1526 858443 1527 858444
rect 1528 858443 1529 858444
rect 2848 858443 2955 858477
rect 1526 858442 1529 858443
rect 5488 858280 5538 859103
rect 5658 858280 5708 859103
rect 6005 858280 6021 859499
rect 12427 859448 12493 859464
rect 24572 859458 25172 859508
rect 32930 859457 33530 859507
rect 35287 859391 35887 859441
rect 36785 859402 37385 859452
rect 24572 859308 25172 859358
rect 31463 859307 32063 859357
rect 32930 859301 33530 859357
rect 7389 859277 7406 859287
rect 7440 859277 7477 859287
rect 7511 859277 7551 859287
rect 7585 859277 7622 859287
rect 7656 859277 7696 859287
rect 7730 859277 7767 859287
rect 7801 859277 7841 859287
rect 7875 859277 7912 859287
rect 7946 859277 7986 859287
rect 8020 859277 8057 859287
rect 8091 859277 8131 859287
rect 8165 859277 8202 859287
rect 8236 859277 8296 859287
rect 8330 859277 8381 859287
rect 8996 859277 9044 859287
rect 9078 859277 9120 859287
rect 9154 859277 9197 859287
rect 9231 859277 9291 859287
rect 9325 859277 9362 859287
rect 9396 859277 9436 859287
rect 9470 859277 9507 859287
rect 9541 859277 9581 859287
rect 9615 859277 9652 859287
rect 9686 859277 9726 859287
rect 9760 859277 9797 859287
rect 9831 859277 9871 859287
rect 9905 859277 9942 859287
rect 9976 859277 9990 859287
rect 7389 859209 8389 859277
rect 8990 859183 9990 859277
rect 36785 859226 37385 859282
rect 15678 859127 16678 859177
rect 17278 859127 18278 859177
rect 31463 859151 32063 859207
rect 32930 859151 33530 859201
rect 34079 859157 34679 859207
rect 7389 858840 8389 858864
rect 15678 858860 16678 858916
rect 17278 858860 18278 858916
rect 8990 858840 9990 858841
rect 7389 858743 8389 858799
rect 8990 858743 9990 858799
rect 15678 858788 16678 858844
rect 17278 858788 18278 858844
rect 8990 858701 9990 858702
rect 15678 858286 16678 858426
rect 17278 858286 18278 858426
rect 19844 858280 19894 859051
rect 20462 858280 20512 859051
rect 31463 859001 32063 859051
rect 34079 859001 34679 859057
rect 35287 859039 35887 859095
rect 36785 859050 37385 859106
rect 32596 858929 33596 858979
rect 24573 858820 25173 858870
rect 34079 858851 34679 858901
rect 35287 858869 35887 858919
rect 36785 858880 37385 858930
rect 30171 858795 30771 858845
rect 32596 858773 33596 858829
rect 37993 858704 38593 858754
rect 30171 858619 30771 858675
rect 32596 858623 33596 858673
rect 34110 858589 34710 858639
rect 21263 858280 21313 858518
rect 22349 858280 22399 858518
rect 32596 858507 33596 858557
rect 30171 858449 30771 858499
rect 36785 858429 36985 858609
rect 37993 858534 38593 858584
rect 24573 858352 25173 858408
rect 29993 858310 30993 858360
rect 31347 858280 31547 858317
rect 31607 858280 31807 858317
rect 36785 858280 36985 858373
rect 37083 858280 37120 858373
rect 696597 856200 696600 856320
rect 692376 855983 692396 856017
rect 692463 855993 692532 856017
rect 696191 855993 696239 856017
rect 692487 855983 692532 855993
rect 696204 855983 696239 855993
rect 696340 855983 696360 856017
rect 692487 855915 692502 855939
rect 696200 855915 696215 855939
rect 692454 855891 692478 855915
rect 696224 855891 696248 855915
rect 686755 855800 687355 855850
rect 692487 855748 692505 855752
rect 692479 855718 692505 855748
rect 692487 855698 692505 855718
rect 686755 855624 687355 855680
rect 692485 855674 692505 855698
rect 692509 855674 692517 855718
rect 696215 855698 696223 855748
rect 696203 855674 696223 855698
rect 696227 855674 696245 855752
rect 692485 855640 692521 855674
rect 696203 855640 696249 855674
rect 686755 855448 687355 855504
rect 686755 855278 687355 855328
rect 685547 855102 686147 855152
rect 687155 855007 687170 855022
rect 687343 855018 687355 855022
rect 687340 855007 687355 855018
rect 685547 854932 686147 854982
rect 687155 854827 687355 855007
rect 687155 854812 687170 854827
rect 687340 854816 687355 854827
rect 687343 854812 687355 854816
rect 687042 854771 687057 854786
rect 687020 854591 687057 854771
rect 687155 854771 687170 854786
rect 687343 854782 687355 854786
rect 687340 854771 687355 854782
rect 687155 854591 687355 854771
rect 688210 854630 688260 855630
rect 688360 854740 688488 855630
rect 688516 854740 688644 855630
rect 688672 854740 688800 855630
rect 688828 854740 688956 855630
rect 688984 854740 689112 855630
rect 689140 854740 689268 855630
rect 689296 854740 689424 855630
rect 689452 854740 689580 855630
rect 689608 854740 689736 855630
rect 689764 854740 689892 855630
rect 689920 854740 690048 855630
rect 690076 854740 690204 855630
rect 690232 854740 690360 855630
rect 690388 854630 690438 855630
rect 692485 855606 692505 855640
rect 692509 855606 692517 855640
rect 696203 855606 696223 855640
rect 696227 855606 696245 855640
rect 691275 855523 691875 855573
rect 692485 855572 692521 855606
rect 696203 855572 696249 855606
rect 692485 855538 692505 855572
rect 692509 855538 692517 855572
rect 692485 855504 692521 855538
rect 692583 855528 693983 855571
rect 694719 855528 696119 855571
rect 696203 855538 696223 855572
rect 696227 855538 696245 855572
rect 696203 855504 696249 855538
rect 692485 855470 692505 855504
rect 692509 855470 692517 855504
rect 692485 855436 692521 855470
rect 691275 855373 691875 855423
rect 692485 855402 692505 855436
rect 692509 855402 692517 855436
rect 692485 855368 692521 855402
rect 692485 855334 692505 855368
rect 692509 855334 692517 855368
rect 692583 855365 693983 855493
rect 694719 855365 696119 855493
rect 696203 855470 696223 855504
rect 696227 855470 696245 855504
rect 696203 855436 696249 855470
rect 707624 855441 707658 855475
rect 707695 855441 707729 855475
rect 707769 855441 707803 855475
rect 707840 855441 707874 855475
rect 707914 855441 707948 855475
rect 707985 855441 708019 855475
rect 708059 855441 708093 855475
rect 708130 855441 708164 855475
rect 708204 855441 708238 855475
rect 708275 855441 708309 855475
rect 708369 855441 708403 855475
rect 708446 855441 708480 855475
rect 708520 855441 708554 855465
rect 708588 855441 708610 855465
rect 709211 855441 709234 855465
rect 709270 855441 709304 855475
rect 709364 855441 709398 855475
rect 709435 855441 709469 855475
rect 709509 855441 709543 855475
rect 709580 855441 709614 855475
rect 709654 855441 709688 855475
rect 709725 855441 709759 855475
rect 709799 855441 709833 855475
rect 709870 855441 709904 855475
rect 709944 855441 709978 855475
rect 710015 855441 710049 855475
rect 710089 855441 710123 855475
rect 710160 855441 710194 855475
rect 696203 855402 696223 855436
rect 696227 855402 696245 855436
rect 707610 855431 707624 855441
rect 707658 855431 707695 855441
rect 707729 855431 707769 855441
rect 707803 855431 707840 855441
rect 707874 855431 707914 855441
rect 707948 855431 707985 855441
rect 708019 855431 708059 855441
rect 708093 855431 708130 855441
rect 708164 855431 708204 855441
rect 708238 855431 708275 855441
rect 708309 855431 708369 855441
rect 708403 855431 708446 855441
rect 708480 855431 708520 855441
rect 708554 855431 708588 855441
rect 708610 855431 708634 855441
rect 709211 855431 709270 855441
rect 709304 855431 709364 855441
rect 709398 855431 709435 855441
rect 709469 855431 709509 855441
rect 709543 855431 709580 855441
rect 709614 855431 709654 855441
rect 709688 855431 709725 855441
rect 709759 855431 709799 855441
rect 709833 855431 709870 855441
rect 709904 855431 709944 855441
rect 709978 855431 710015 855441
rect 710049 855431 710089 855441
rect 710123 855431 710160 855441
rect 710194 855431 710211 855441
rect 696203 855368 696249 855402
rect 696203 855334 696223 855368
rect 696227 855334 696245 855368
rect 707610 855337 708610 855431
rect 709211 855337 710211 855431
rect 691275 855251 691875 855301
rect 692485 855300 692521 855334
rect 692485 855266 692505 855300
rect 692509 855266 692517 855300
rect 692485 855232 692521 855266
rect 692485 855198 692505 855232
rect 692509 855198 692517 855232
rect 692583 855202 693983 855330
rect 694719 855202 696119 855330
rect 696203 855300 696249 855334
rect 711579 855317 712463 855331
rect 711579 855307 711619 855317
rect 696203 855266 696223 855300
rect 696227 855266 696245 855300
rect 701730 855290 701747 855292
rect 696203 855232 696249 855266
rect 696203 855198 696223 855232
rect 696227 855198 696245 855232
rect 701692 855220 701722 855254
rect 701730 855220 701760 855290
rect 707610 855241 708610 855301
rect 709211 855241 710211 855301
rect 692485 855164 692521 855198
rect 691275 855101 691875 855151
rect 692485 855130 692505 855164
rect 692509 855130 692517 855164
rect 692485 855096 692521 855130
rect 692485 855062 692505 855096
rect 692509 855062 692517 855096
rect 692485 855028 692521 855062
rect 692583 855039 693983 855167
rect 694719 855039 696119 855167
rect 696203 855164 696249 855198
rect 696203 855130 696223 855164
rect 696227 855130 696245 855164
rect 696203 855096 696249 855130
rect 696203 855062 696223 855096
rect 696227 855062 696245 855096
rect 699322 855064 700322 855097
rect 700922 855064 701922 855097
rect 696203 855028 696249 855062
rect 707610 855044 708610 855048
rect 709211 855044 710211 855048
rect 691275 854975 691875 855025
rect 692485 854994 692505 855028
rect 692509 854994 692517 855028
rect 692485 854960 692521 854994
rect 692485 854926 692505 854960
rect 692509 854926 692517 854960
rect 692485 854892 692521 854926
rect 691275 854825 691875 854875
rect 692485 854858 692505 854892
rect 692509 854858 692517 854892
rect 692583 854876 693983 855004
rect 694719 854876 696119 855004
rect 696203 854994 696223 855028
rect 696227 854994 696245 855028
rect 707574 854994 708646 855030
rect 696203 854960 696249 854994
rect 696203 854926 696223 854960
rect 696227 854926 696245 854960
rect 707574 854953 707610 854994
rect 708610 854953 708646 854994
rect 696203 854892 696249 854926
rect 697284 854894 697350 854910
rect 707574 854897 708646 854953
rect 696203 854858 696223 854892
rect 696227 854858 696245 854892
rect 699322 854877 700322 854894
rect 700922 854877 701922 854894
rect 707574 854881 707610 854897
rect 708610 854881 708646 854897
rect 692485 854824 692521 854858
rect 692485 854790 692505 854824
rect 692509 854790 692517 854824
rect 692485 854756 692521 854790
rect 691275 854703 691875 854753
rect 692485 854740 692505 854756
rect 692509 854740 692517 854756
rect 692583 854740 693983 854841
rect 694719 854740 696119 854841
rect 696203 854824 696249 854858
rect 707574 854825 708646 854881
rect 696203 854790 696223 854824
rect 696227 854790 696245 854824
rect 696203 854756 696249 854790
rect 696203 854740 696223 854756
rect 696227 854740 696245 854756
rect 699322 854740 700322 854811
rect 700922 854740 701922 854811
rect 707574 854788 707610 854825
rect 708610 854788 708646 854825
rect 707574 854748 708646 854788
rect 709175 854994 710247 855030
rect 709175 854953 709211 854994
rect 710211 854953 710247 854994
rect 709175 854897 710247 854953
rect 709175 854881 709211 854897
rect 710211 854881 710247 854897
rect 709175 854825 710247 854881
rect 709175 854788 709211 854825
rect 710211 854788 710247 854825
rect 709175 854748 710247 854788
rect 685542 854506 686142 854556
rect 691275 854553 691875 854603
rect 685542 854330 686142 854386
rect 692583 854237 693983 854280
rect 694719 854237 696119 854280
rect 699322 854278 700322 854418
rect 700922 854278 701922 854418
rect 685542 854160 686142 854210
rect 692583 854101 693983 854144
rect 694719 854101 696119 854144
rect 680215 853678 680815 853728
rect 680215 853502 680815 853558
rect 685551 853516 686551 853566
rect 689154 853480 689204 853897
rect 689304 853480 689360 853897
rect 689460 853480 689516 853897
rect 689616 853480 689672 853897
rect 689772 853480 689828 853897
rect 689928 853480 689978 853897
rect 699322 853860 700322 853916
rect 700922 853860 701922 853916
rect 707610 853905 708610 853961
rect 709211 853905 710211 853961
rect 699322 853788 700322 853844
rect 700922 853788 701922 853844
rect 707610 853833 708610 853889
rect 709211 853833 710211 853889
rect 711579 853525 711605 855307
rect 715956 854297 716006 855297
rect 716106 854740 716234 855297
rect 716262 854297 716312 855297
rect 711579 853480 711595 853495
rect 712409 853480 712431 853485
rect 713640 853480 713641 853785
rect 713750 853772 714750 853822
rect 713750 853562 714750 853612
rect 713750 853480 714750 853496
rect 2850 847304 3850 847320
rect 2850 847188 3850 847238
rect 2850 846978 3850 847028
rect 3959 847015 3960 847320
rect 5169 847315 5191 847320
rect 6005 847305 6021 847320
rect 1288 845503 1338 846503
rect 1438 845503 1566 846060
rect 1594 845503 1644 846503
rect 5995 845493 6021 847275
rect 7389 846911 8389 846967
rect 8990 846911 9990 846967
rect 15678 846956 16678 847012
rect 17278 846956 18278 847012
rect 7389 846839 8389 846895
rect 8990 846839 9990 846895
rect 15678 846884 16678 846940
rect 17278 846884 18278 846940
rect 27622 846903 27672 847320
rect 27772 846903 27828 847320
rect 27928 846903 27984 847320
rect 28084 846903 28140 847320
rect 28240 846903 28296 847320
rect 28396 846903 28446 847320
rect 31049 847234 32049 847284
rect 36785 847242 37385 847298
rect 36785 847072 37385 847122
rect 21481 846656 22881 846699
rect 23617 846656 25017 846699
rect 31458 846590 32058 846640
rect 15678 846382 16678 846522
rect 17278 846382 18278 846522
rect 21481 846520 22881 846563
rect 23617 846520 25017 846563
rect 31458 846414 32058 846470
rect 25725 846197 26325 846247
rect 31458 846244 32058 846294
rect 7353 846016 8425 846052
rect 7353 845975 7389 846016
rect 8389 845975 8425 846016
rect 7353 845919 8425 845975
rect 7353 845903 7389 845919
rect 8389 845903 8425 845919
rect 7353 845847 8425 845903
rect 7353 845810 7389 845847
rect 8389 845810 8425 845847
rect 7353 845770 8425 845810
rect 8954 846016 10026 846052
rect 8954 845975 8990 846016
rect 9990 845975 10026 846016
rect 8954 845919 10026 845975
rect 21383 846044 21403 846060
rect 21407 846044 21415 846060
rect 21383 846010 21419 846044
rect 21481 846031 22881 846060
rect 23617 846031 25017 846060
rect 25101 846044 25121 846060
rect 25125 846044 25143 846060
rect 25725 846047 26325 846097
rect 25101 846010 25147 846044
rect 21383 845976 21403 846010
rect 21407 845976 21415 846010
rect 21383 845942 21419 845976
rect 8954 845903 8990 845919
rect 9990 845903 10026 845919
rect 15678 845906 16678 845923
rect 17278 845906 18278 845923
rect 21383 845908 21403 845942
rect 21407 845908 21415 845942
rect 8954 845847 10026 845903
rect 20250 845890 20316 845906
rect 8954 845810 8990 845847
rect 9990 845810 10026 845847
rect 8954 845770 10026 845810
rect 21383 845874 21419 845908
rect 21383 845840 21403 845874
rect 21407 845840 21415 845874
rect 21481 845868 22881 845996
rect 23617 845868 25017 845996
rect 25101 845976 25121 846010
rect 25125 845976 25143 846010
rect 25101 845942 25147 845976
rect 25101 845908 25121 845942
rect 25125 845908 25143 845942
rect 25725 845925 26325 845975
rect 25101 845874 25147 845908
rect 25101 845840 25121 845874
rect 25125 845840 25143 845874
rect 21383 845806 21419 845840
rect 21383 845772 21403 845806
rect 21407 845772 21415 845806
rect 21383 845738 21419 845772
rect 15678 845703 16678 845736
rect 17278 845703 18278 845736
rect 21383 845704 21403 845738
rect 21407 845704 21415 845738
rect 21481 845705 22881 845833
rect 23617 845705 25017 845833
rect 25101 845806 25147 845840
rect 25101 845772 25121 845806
rect 25125 845772 25143 845806
rect 25725 845775 26325 845825
rect 25101 845738 25147 845772
rect 25101 845704 25121 845738
rect 25125 845704 25143 845738
rect 21383 845670 21419 845704
rect 25101 845670 25147 845704
rect 21383 845636 21403 845670
rect 21407 845636 21415 845670
rect 7389 845559 8389 845631
rect 8990 845559 9990 845631
rect 21383 845602 21419 845636
rect 15840 845510 15870 845580
rect 15878 845546 15908 845580
rect 21383 845568 21403 845602
rect 21407 845568 21415 845602
rect 15853 845508 15870 845510
rect 21383 845534 21419 845568
rect 21481 845542 22881 845670
rect 23617 845542 25017 845670
rect 25101 845636 25121 845670
rect 25125 845636 25143 845670
rect 25725 845649 26325 845699
rect 25101 845602 25147 845636
rect 25101 845568 25121 845602
rect 25125 845568 25143 845602
rect 25101 845534 25147 845568
rect 5981 845483 6021 845493
rect 5137 845469 6021 845483
rect 21383 845500 21403 845534
rect 21407 845500 21415 845534
rect 21383 845466 21419 845500
rect 7389 845369 8389 845463
rect 7389 845359 8413 845369
rect 8990 845359 9990 845463
rect 21383 845432 21403 845466
rect 21407 845432 21415 845466
rect 21383 845398 21419 845432
rect 21383 845364 21403 845398
rect 21407 845364 21415 845398
rect 21481 845379 22881 845507
rect 23617 845379 25017 845507
rect 25101 845500 25121 845534
rect 25125 845500 25143 845534
rect 25101 845466 25147 845500
rect 25725 845499 26325 845549
rect 25101 845432 25121 845466
rect 25125 845432 25143 845466
rect 25101 845398 25147 845432
rect 25101 845364 25121 845398
rect 25125 845364 25143 845398
rect 25725 845377 26325 845427
rect 21383 845330 21419 845364
rect 25101 845330 25147 845364
rect 21383 845296 21403 845330
rect 21407 845296 21415 845330
rect 25101 845296 25121 845330
rect 25125 845296 25143 845330
rect 21383 845262 21419 845296
rect 21383 845228 21403 845262
rect 21407 845228 21415 845262
rect 21481 845229 22881 845272
rect 23617 845229 25017 845272
rect 25101 845262 25147 845296
rect 25101 845228 25121 845262
rect 25125 845228 25143 845262
rect 21383 845194 21419 845228
rect 25101 845194 25147 845228
rect 25725 845227 26325 845277
rect 21383 845160 21403 845194
rect 21407 845160 21415 845194
rect 25101 845160 25121 845194
rect 25125 845160 25143 845194
rect 27162 845170 27212 846170
rect 27312 845170 27440 846060
rect 27468 845170 27596 846060
rect 27624 845170 27752 846060
rect 27780 845170 27908 846060
rect 27936 845170 28064 846060
rect 28092 845170 28220 846060
rect 28248 845170 28376 846060
rect 28404 845170 28532 846060
rect 28560 845170 28688 846060
rect 28716 845170 28844 846060
rect 28872 845170 29000 846060
rect 29028 845170 29156 846060
rect 29184 845170 29312 846060
rect 29340 845170 29390 846170
rect 30245 846029 30445 846209
rect 30245 846018 30260 846029
rect 30245 846014 30257 846018
rect 30430 846014 30445 846029
rect 30543 846029 30580 846209
rect 30543 846014 30558 846029
rect 30245 845984 30257 845988
rect 30245 845973 30260 845984
rect 30430 845973 30445 845988
rect 30245 845793 30445 845973
rect 31453 845818 32053 845868
rect 30245 845782 30260 845793
rect 30245 845778 30257 845782
rect 30430 845778 30445 845793
rect 31453 845648 32053 845698
rect 30245 845472 30845 845522
rect 30245 845296 30845 845352
rect 21383 845126 21419 845160
rect 25101 845126 25147 845160
rect 21383 845102 21403 845126
rect 21385 845048 21403 845102
rect 21407 845082 21415 845126
rect 25101 845102 25121 845126
rect 25113 845082 25121 845102
rect 25125 845048 25143 845126
rect 30245 845120 30845 845176
rect 30245 844950 30845 845000
rect 21000 844800 21003 844920
rect 21352 844885 21376 844909
rect 25122 844885 25146 844909
rect 21385 844861 21400 844885
rect 25098 844861 25113 844885
rect 21274 844783 21294 844851
rect 21410 844817 21430 844851
rect 25068 844817 25088 844851
rect 25204 844817 25224 844851
rect 21385 844807 21430 844817
rect 25102 844807 25137 844817
rect 21361 844783 21430 844807
rect 25089 844783 25137 844807
rect 25238 844783 25258 844817
rect 680480 842427 680517 842520
rect 680615 842427 680815 842520
rect 685793 842483 685993 842520
rect 686053 842483 686253 842520
rect 686607 842440 687607 842490
rect 692427 842392 693027 842448
rect 679007 842216 679607 842266
rect 680615 842191 680815 842371
rect 686829 842301 687429 842351
rect 684004 842243 685004 842293
rect 695201 842282 695251 842520
rect 696287 842282 696337 842520
rect 682890 842161 683490 842211
rect 684004 842127 685004 842177
rect 686829 842125 687429 842181
rect 679007 842046 679607 842096
rect 684004 841971 685004 842027
rect 686829 841955 687429 842005
rect 680215 841870 680815 841920
rect 681713 841881 682313 841931
rect 682921 841899 683521 841949
rect 692427 841930 693027 841980
rect 684004 841821 685004 841871
rect 680215 841694 680815 841750
rect 681713 841705 682313 841761
rect 682921 841743 683521 841799
rect 685537 841749 686137 841799
rect 697088 841749 697138 842520
rect 697706 841749 697756 842520
rect 699322 842374 700322 842514
rect 700922 842374 701922 842514
rect 707610 842098 708610 842099
rect 699322 841956 700322 842012
rect 700922 841956 701922 842012
rect 707610 842001 708610 842057
rect 709211 842001 710211 842057
rect 707610 841959 708610 841960
rect 699322 841884 700322 841940
rect 700922 841884 701922 841940
rect 709211 841936 710211 841960
rect 682921 841593 683521 841643
rect 684070 841599 684670 841649
rect 685537 841593 686137 841649
rect 699322 841623 700322 841673
rect 700922 841623 701922 841673
rect 680215 841518 680815 841574
rect 707610 841523 708610 841617
rect 709211 841523 710211 841591
rect 707610 841513 707624 841523
rect 707658 841513 707695 841523
rect 707729 841513 707769 841523
rect 707803 841513 707840 841523
rect 707874 841513 707914 841523
rect 707948 841513 707985 841523
rect 708019 841513 708059 841523
rect 708093 841513 708130 841523
rect 708164 841513 708204 841523
rect 708238 841513 708275 841523
rect 708309 841513 708369 841523
rect 708403 841513 708446 841523
rect 708480 841513 708522 841523
rect 708556 841513 708604 841523
rect 709219 841513 709270 841523
rect 709304 841513 709364 841523
rect 709398 841513 709435 841523
rect 709469 841513 709509 841523
rect 709543 841513 709580 841523
rect 709614 841513 709654 841523
rect 709688 841513 709725 841523
rect 709759 841513 709799 841523
rect 709833 841513 709870 841523
rect 709904 841513 709944 841523
rect 709978 841513 710015 841523
rect 710049 841513 710089 841523
rect 710123 841513 710160 841523
rect 710194 841513 710211 841523
rect 684070 841443 684670 841499
rect 685537 841443 686137 841493
rect 692428 841442 693028 841492
rect 680215 841348 680815 841398
rect 681713 841359 682313 841409
rect 684070 841293 684670 841343
rect 692428 841292 693028 841342
rect 705107 841336 705173 841352
rect 711579 841301 711595 842520
rect 711892 841697 711942 842520
rect 712062 841697 712112 842520
rect 716071 842357 716074 842358
rect 714645 842323 714752 842357
rect 716071 842356 716072 842357
rect 716073 842356 716074 842357
rect 716071 842355 716074 842356
rect 716208 842357 716211 842358
rect 716208 842356 716209 842357
rect 716210 842356 716211 842357
rect 716208 842355 716211 842356
rect 714964 842247 715998 842329
rect 716284 842247 717318 842329
rect 714175 841398 714225 841998
rect 714425 841398 714475 841998
rect 680215 841232 680815 841282
rect 698017 841232 698053 841260
rect 692428 841162 693028 841212
rect 698030 841198 698077 841232
rect 698017 841164 698053 841198
rect 680215 841056 680815 841112
rect 692428 841006 693028 841134
rect 698030 841130 698077 841164
rect 698017 841096 698053 841130
rect 698030 841062 698077 841096
rect 698017 840983 698053 841062
rect 698084 840983 698120 841260
rect 714781 841191 714863 842226
rect 715134 841955 715828 842037
rect 714686 841123 714863 841191
rect 714645 841089 714863 841123
rect 680215 840880 680815 840936
rect 686719 840893 686739 840917
rect 686743 840893 686753 840917
rect 686719 840859 686757 840893
rect 686719 840822 686739 840859
rect 686743 840822 686753 840859
rect 692428 840850 693028 840978
rect 698017 840947 698210 840983
rect 698084 840935 698210 840947
rect 702756 840959 703645 840983
rect 702756 840935 702853 840959
rect 698084 840828 702853 840935
rect 686719 840788 686757 840822
rect 680215 840704 680815 840760
rect 686719 840751 686739 840788
rect 686743 840751 686753 840788
rect 686719 840741 686757 840751
rect 686699 840717 686767 840741
rect 686719 840704 686739 840717
rect 686743 840704 686753 840717
rect 686719 840695 686753 840704
rect 686719 840693 686743 840695
rect 692428 840694 693028 840750
rect 686685 840656 686709 840680
rect 686743 840656 686767 840680
rect 678799 840503 679399 840553
rect 680215 840534 680815 840584
rect 692428 840538 693028 840666
rect 680593 840531 680815 840534
rect 682009 840501 682069 840516
rect 682024 840465 682054 840501
rect 683708 840387 684308 840437
rect 678799 840327 679399 840383
rect 692428 840382 693028 840510
rect 714781 840308 714863 841089
rect 715063 840609 715145 841915
rect 715289 840777 715339 841719
rect 715633 840777 715683 841719
rect 715382 840672 715422 840756
rect 715542 840672 715582 840756
rect 715342 840632 715382 840672
rect 715582 840632 715622 840672
rect 715815 840609 715897 841915
rect 715134 840387 715828 840469
rect 716100 840308 716182 842226
rect 716454 841955 717148 842037
rect 716385 840609 716467 841915
rect 716599 840777 716649 841719
rect 716943 840777 716993 841719
rect 716700 840672 716740 840756
rect 716860 840672 716900 840756
rect 716660 840632 716700 840672
rect 716900 840632 716940 840672
rect 717137 840609 717219 841915
rect 716454 840387 717148 840469
rect 717419 840308 717501 842226
rect 683708 840237 684308 840287
rect 692428 840232 693028 840282
rect 678799 840157 679399 840207
rect 684565 840160 684790 840168
rect 696597 840000 696600 840120
rect 714964 840095 715998 840177
rect 716284 840095 717318 840177
rect 21000 813000 21003 813120
rect 282 812623 1316 812705
rect 1602 812623 2636 812705
rect 32810 812662 33035 812670
rect 38201 812593 38801 812643
rect 24572 812518 25172 812568
rect 33292 812513 33892 812563
rect 99 810574 181 812492
rect 452 812331 1146 812413
rect 381 810885 463 812191
rect 660 812128 700 812168
rect 900 812128 940 812168
rect 700 812044 740 812128
rect 860 812044 900 812128
rect 607 811081 657 812023
rect 951 811081 1001 812023
rect 1133 810885 1215 812191
rect 452 810763 1146 810845
rect 1418 810574 1500 812492
rect 1772 812331 2466 812413
rect 1703 810885 1785 812191
rect 1978 812128 2018 812168
rect 2218 812128 2258 812168
rect 2018 812044 2058 812128
rect 2178 812044 2218 812128
rect 1917 811081 1967 812023
rect 2261 811081 2311 812023
rect 2455 810885 2537 812191
rect 2737 811779 2819 812492
rect 24572 812362 25172 812490
rect 38201 812417 38801 812473
rect 33292 812363 33892 812413
rect 24572 812206 25172 812334
rect 35546 812299 35576 812335
rect 36785 812329 36935 812341
rect 35531 812284 35591 812299
rect 36785 812216 37385 812266
rect 38201 812247 38801 812297
rect 30833 812120 30857 812144
rect 30891 812120 30915 812144
rect 24572 812050 25172 812106
rect 30857 812105 30881 812107
rect 30857 812096 30887 812105
rect 30867 812083 30887 812096
rect 30891 812083 30907 812120
rect 30833 812059 30857 812083
rect 30867 812049 30911 812083
rect 14747 811865 19516 811972
rect 24572 811894 25172 812022
rect 30867 812012 30887 812049
rect 30891 812012 30907 812049
rect 36785 812040 37385 812096
rect 30867 811978 30911 812012
rect 30867 811941 30887 811978
rect 30891 811941 30907 811978
rect 30867 811907 30911 811941
rect 30867 811883 30887 811907
rect 30891 811883 30907 811907
rect 14747 811841 14844 811865
rect 13955 811817 14844 811841
rect 19390 811853 19516 811865
rect 19390 811841 19583 811853
rect 19390 811817 19605 811841
rect 19639 811817 19673 811841
rect 19707 811817 19741 811841
rect 19775 811817 19809 811841
rect 19843 811817 19877 811841
rect 19911 811817 19945 811841
rect 19979 811817 20013 811841
rect 20047 811817 20081 811841
rect 20115 811817 20149 811841
rect 20183 811817 20217 811841
rect 20251 811817 20285 811841
rect 20319 811817 20353 811841
rect 20387 811817 20421 811841
rect 20455 811817 20489 811841
rect 20523 811817 20557 811841
rect 20591 811817 20625 811841
rect 20659 811817 20693 811841
rect 2737 811711 2914 811779
rect 1772 810763 2466 810845
rect 2737 810574 2819 811711
rect 2848 811677 2955 811711
rect 19480 811540 19516 811817
rect 19547 811540 19583 811817
rect 24572 811738 25172 811866
rect 36785 811864 37385 811920
rect 36785 811688 37385 811744
rect 20809 811650 20833 811684
rect 20809 811582 20833 811616
rect 24572 811588 25172 811638
rect 20809 811540 20833 811548
rect 36785 811518 37385 811568
rect 3125 810802 3175 811402
rect 3375 810802 3425 811402
rect 282 810471 1316 810553
rect 1602 810471 2636 810553
rect 1389 810444 1392 810445
rect 1389 810443 1390 810444
rect 1391 810443 1392 810444
rect 1389 810442 1392 810443
rect 1526 810444 1529 810445
rect 1526 810443 1527 810444
rect 1528 810443 1529 810444
rect 2848 810443 2955 810477
rect 1526 810442 1529 810443
rect 5488 810280 5538 811103
rect 5658 810280 5708 811103
rect 6005 810280 6021 811499
rect 12427 811448 12493 811464
rect 24572 811458 25172 811508
rect 32930 811457 33530 811507
rect 35287 811391 35887 811441
rect 36785 811402 37385 811452
rect 24572 811308 25172 811358
rect 31463 811307 32063 811357
rect 32930 811301 33530 811357
rect 7389 811277 7406 811287
rect 7440 811277 7477 811287
rect 7511 811277 7551 811287
rect 7585 811277 7622 811287
rect 7656 811277 7696 811287
rect 7730 811277 7767 811287
rect 7801 811277 7841 811287
rect 7875 811277 7912 811287
rect 7946 811277 7986 811287
rect 8020 811277 8057 811287
rect 8091 811277 8131 811287
rect 8165 811277 8202 811287
rect 8236 811277 8296 811287
rect 8330 811277 8381 811287
rect 8996 811277 9044 811287
rect 9078 811277 9120 811287
rect 9154 811277 9197 811287
rect 9231 811277 9291 811287
rect 9325 811277 9362 811287
rect 9396 811277 9436 811287
rect 9470 811277 9507 811287
rect 9541 811277 9581 811287
rect 9615 811277 9652 811287
rect 9686 811277 9726 811287
rect 9760 811277 9797 811287
rect 9831 811277 9871 811287
rect 9905 811277 9942 811287
rect 9976 811277 9990 811287
rect 7389 811209 8389 811277
rect 8990 811183 9990 811277
rect 36785 811226 37385 811282
rect 15678 811127 16678 811177
rect 17278 811127 18278 811177
rect 31463 811151 32063 811207
rect 32930 811151 33530 811201
rect 34079 811157 34679 811207
rect 7389 810840 8389 810864
rect 15678 810860 16678 810916
rect 17278 810860 18278 810916
rect 8990 810840 9990 810841
rect 7389 810743 8389 810799
rect 8990 810743 9990 810799
rect 15678 810788 16678 810844
rect 17278 810788 18278 810844
rect 8990 810701 9990 810702
rect 15678 810286 16678 810426
rect 17278 810286 18278 810426
rect 19844 810280 19894 811051
rect 20462 810280 20512 811051
rect 31463 811001 32063 811051
rect 34079 811001 34679 811057
rect 35287 811039 35887 811095
rect 36785 811050 37385 811106
rect 32596 810929 33596 810979
rect 24573 810820 25173 810870
rect 34079 810851 34679 810901
rect 35287 810869 35887 810919
rect 36785 810880 37385 810930
rect 30171 810795 30771 810845
rect 32596 810773 33596 810829
rect 37993 810704 38593 810754
rect 30171 810619 30771 810675
rect 32596 810623 33596 810673
rect 34110 810589 34710 810639
rect 21263 810280 21313 810518
rect 22349 810280 22399 810518
rect 32596 810507 33596 810557
rect 30171 810449 30771 810499
rect 36785 810429 36985 810609
rect 37993 810534 38593 810584
rect 24573 810352 25173 810408
rect 29993 810310 30993 810360
rect 31347 810280 31547 810317
rect 31607 810280 31807 810317
rect 36785 810280 36985 810373
rect 37083 810280 37120 810373
rect 696597 804200 696600 804320
rect 692376 803983 692396 804017
rect 692463 803993 692532 804017
rect 696191 803993 696239 804017
rect 692487 803983 692532 803993
rect 696204 803983 696239 803993
rect 696340 803983 696360 804017
rect 692487 803915 692502 803939
rect 696200 803915 696215 803939
rect 692454 803891 692478 803915
rect 696224 803891 696248 803915
rect 686755 803800 687355 803850
rect 692487 803748 692505 803752
rect 692479 803718 692505 803748
rect 692487 803698 692505 803718
rect 686755 803624 687355 803680
rect 692485 803674 692505 803698
rect 692509 803674 692517 803718
rect 696215 803698 696223 803748
rect 696203 803674 696223 803698
rect 696227 803674 696245 803752
rect 692485 803640 692521 803674
rect 696203 803640 696249 803674
rect 686755 803448 687355 803504
rect 686755 803278 687355 803328
rect 685547 803102 686147 803152
rect 687155 803007 687170 803022
rect 687343 803018 687355 803022
rect 687340 803007 687355 803018
rect 685547 802932 686147 802982
rect 687155 802827 687355 803007
rect 687155 802812 687170 802827
rect 687340 802816 687355 802827
rect 687343 802812 687355 802816
rect 687042 802771 687057 802786
rect 687020 802591 687057 802771
rect 687042 802576 687057 802591
rect 687155 802771 687170 802786
rect 687343 802782 687355 802786
rect 687340 802771 687355 802782
rect 687155 802591 687355 802771
rect 688210 802630 688260 803630
rect 688360 802630 688488 803630
rect 688516 802630 688644 803630
rect 688672 802630 688800 803630
rect 688828 802630 688956 803630
rect 688984 802630 689112 803630
rect 689140 802630 689268 803630
rect 689296 802630 689424 803630
rect 689452 802630 689580 803630
rect 689608 802630 689736 803630
rect 689764 802630 689892 803630
rect 689920 802630 690048 803630
rect 690076 802630 690204 803630
rect 690232 802630 690360 803630
rect 690388 802630 690438 803630
rect 692485 803606 692505 803640
rect 692509 803606 692517 803640
rect 696203 803606 696223 803640
rect 696227 803606 696245 803640
rect 691275 803523 691875 803573
rect 692485 803572 692521 803606
rect 696203 803572 696249 803606
rect 692485 803538 692505 803572
rect 692509 803538 692517 803572
rect 692485 803504 692521 803538
rect 692583 803528 693983 803571
rect 694719 803528 696119 803571
rect 696203 803538 696223 803572
rect 696227 803538 696245 803572
rect 696203 803504 696249 803538
rect 692485 803470 692505 803504
rect 692509 803470 692517 803504
rect 692485 803436 692521 803470
rect 691275 803373 691875 803423
rect 692485 803402 692505 803436
rect 692509 803402 692517 803436
rect 692485 803368 692521 803402
rect 692485 803334 692505 803368
rect 692509 803334 692517 803368
rect 692583 803365 693983 803493
rect 694719 803365 696119 803493
rect 696203 803470 696223 803504
rect 696227 803470 696245 803504
rect 696203 803436 696249 803470
rect 707624 803441 707658 803475
rect 707695 803441 707729 803475
rect 707769 803441 707803 803475
rect 707840 803441 707874 803475
rect 707914 803441 707948 803475
rect 707985 803441 708019 803475
rect 708059 803441 708093 803475
rect 708130 803441 708164 803475
rect 708204 803441 708238 803475
rect 708275 803441 708309 803475
rect 708369 803441 708403 803475
rect 708446 803441 708480 803475
rect 708520 803441 708554 803465
rect 708588 803441 708610 803465
rect 709211 803441 709234 803465
rect 709270 803441 709304 803475
rect 709364 803441 709398 803475
rect 709435 803441 709469 803475
rect 709509 803441 709543 803475
rect 709580 803441 709614 803475
rect 709654 803441 709688 803475
rect 709725 803441 709759 803475
rect 709799 803441 709833 803475
rect 709870 803441 709904 803475
rect 709944 803441 709978 803475
rect 710015 803441 710049 803475
rect 710089 803441 710123 803475
rect 710160 803441 710194 803475
rect 696203 803402 696223 803436
rect 696227 803402 696245 803436
rect 707610 803431 707624 803441
rect 707658 803431 707695 803441
rect 707729 803431 707769 803441
rect 707803 803431 707840 803441
rect 707874 803431 707914 803441
rect 707948 803431 707985 803441
rect 708019 803431 708059 803441
rect 708093 803431 708130 803441
rect 708164 803431 708204 803441
rect 708238 803431 708275 803441
rect 708309 803431 708369 803441
rect 708403 803431 708446 803441
rect 708480 803431 708520 803441
rect 708554 803431 708588 803441
rect 708610 803431 708634 803441
rect 709211 803431 709270 803441
rect 709304 803431 709364 803441
rect 709398 803431 709435 803441
rect 709469 803431 709509 803441
rect 709543 803431 709580 803441
rect 709614 803431 709654 803441
rect 709688 803431 709725 803441
rect 709759 803431 709799 803441
rect 709833 803431 709870 803441
rect 709904 803431 709944 803441
rect 709978 803431 710015 803441
rect 710049 803431 710089 803441
rect 710123 803431 710160 803441
rect 710194 803431 710211 803441
rect 696203 803368 696249 803402
rect 696203 803334 696223 803368
rect 696227 803334 696245 803368
rect 707610 803337 708610 803431
rect 709211 803337 710211 803431
rect 691275 803251 691875 803301
rect 692485 803300 692521 803334
rect 692485 803266 692505 803300
rect 692509 803266 692517 803300
rect 692485 803232 692521 803266
rect 692485 803198 692505 803232
rect 692509 803198 692517 803232
rect 692583 803202 693983 803330
rect 694719 803202 696119 803330
rect 696203 803300 696249 803334
rect 711579 803317 712463 803331
rect 711579 803307 711619 803317
rect 696203 803266 696223 803300
rect 696227 803266 696245 803300
rect 701730 803290 701747 803292
rect 696203 803232 696249 803266
rect 696203 803198 696223 803232
rect 696227 803198 696245 803232
rect 701692 803220 701722 803254
rect 701730 803220 701760 803290
rect 707610 803241 708610 803301
rect 709211 803241 710211 803301
rect 692485 803164 692521 803198
rect 691275 803101 691875 803151
rect 692485 803130 692505 803164
rect 692509 803130 692517 803164
rect 692485 803096 692521 803130
rect 692485 803062 692505 803096
rect 692509 803062 692517 803096
rect 692485 803028 692521 803062
rect 692583 803039 693983 803167
rect 694719 803039 696119 803167
rect 696203 803164 696249 803198
rect 696203 803130 696223 803164
rect 696227 803130 696245 803164
rect 696203 803096 696249 803130
rect 696203 803062 696223 803096
rect 696227 803062 696245 803096
rect 699322 803064 700322 803097
rect 700922 803064 701922 803097
rect 696203 803028 696249 803062
rect 707610 803044 708610 803048
rect 709211 803044 710211 803048
rect 691275 802975 691875 803025
rect 692485 802994 692505 803028
rect 692509 802994 692517 803028
rect 692485 802960 692521 802994
rect 692485 802926 692505 802960
rect 692509 802926 692517 802960
rect 692485 802892 692521 802926
rect 691275 802825 691875 802875
rect 692485 802858 692505 802892
rect 692509 802858 692517 802892
rect 692583 802876 693983 803004
rect 694719 802876 696119 803004
rect 696203 802994 696223 803028
rect 696227 802994 696245 803028
rect 707574 802994 708646 803030
rect 696203 802960 696249 802994
rect 696203 802926 696223 802960
rect 696227 802926 696245 802960
rect 707574 802953 707610 802994
rect 708610 802953 708646 802994
rect 696203 802892 696249 802926
rect 697284 802894 697350 802910
rect 707574 802897 708646 802953
rect 696203 802858 696223 802892
rect 696227 802858 696245 802892
rect 699322 802877 700322 802894
rect 700922 802877 701922 802894
rect 707574 802881 707610 802897
rect 708610 802881 708646 802897
rect 692485 802824 692521 802858
rect 692485 802790 692505 802824
rect 692509 802790 692517 802824
rect 692485 802756 692521 802790
rect 691275 802703 691875 802753
rect 692485 802722 692505 802756
rect 692509 802722 692517 802756
rect 692485 802688 692521 802722
rect 692583 802713 693983 802841
rect 694719 802713 696119 802841
rect 696203 802824 696249 802858
rect 707574 802825 708646 802881
rect 696203 802790 696223 802824
rect 696227 802790 696245 802824
rect 696203 802756 696249 802790
rect 696203 802722 696223 802756
rect 696227 802722 696245 802756
rect 699322 802739 700322 802811
rect 700922 802739 701922 802811
rect 707574 802788 707610 802825
rect 708610 802788 708646 802825
rect 707574 802748 708646 802788
rect 709175 802994 710247 803030
rect 709175 802953 709211 802994
rect 710211 802953 710247 802994
rect 709175 802897 710247 802953
rect 709175 802881 709211 802897
rect 710211 802881 710247 802897
rect 709175 802825 710247 802881
rect 709175 802788 709211 802825
rect 710211 802788 710247 802825
rect 709175 802748 710247 802788
rect 696203 802688 696249 802722
rect 692485 802654 692505 802688
rect 692509 802654 692517 802688
rect 692485 802620 692521 802654
rect 687155 802576 687170 802591
rect 687340 802580 687355 802591
rect 687343 802576 687355 802580
rect 685542 802506 686142 802556
rect 691275 802553 691875 802603
rect 692485 802586 692505 802620
rect 692509 802586 692517 802620
rect 692485 802552 692521 802586
rect 692485 802518 692505 802552
rect 692509 802518 692517 802552
rect 692583 802550 693983 802678
rect 694719 802550 696119 802678
rect 696203 802654 696223 802688
rect 696227 802654 696245 802688
rect 696203 802620 696249 802654
rect 696203 802586 696223 802620
rect 696227 802586 696245 802620
rect 696203 802552 696249 802586
rect 696203 802518 696223 802552
rect 696227 802518 696245 802552
rect 692485 802484 692521 802518
rect 692485 802450 692505 802484
rect 692509 802450 692517 802484
rect 692485 802416 692521 802450
rect 679817 802330 679841 802354
rect 685542 802330 686142 802386
rect 692485 802382 692505 802416
rect 692509 802382 692517 802416
rect 692583 802387 693983 802515
rect 694719 802387 696119 802515
rect 696203 802484 696249 802518
rect 696203 802450 696223 802484
rect 696227 802450 696245 802484
rect 699322 802478 700322 802550
rect 700922 802478 701922 802550
rect 707610 802523 708610 802595
rect 709211 802523 710211 802595
rect 699392 802467 699426 802478
rect 699460 802467 699494 802478
rect 699528 802467 699562 802478
rect 699596 802467 699630 802478
rect 699664 802467 699698 802478
rect 699732 802467 699766 802478
rect 699800 802467 699834 802478
rect 699868 802467 699902 802478
rect 699936 802467 699970 802478
rect 700004 802467 700038 802478
rect 700072 802467 700106 802478
rect 700140 802467 700174 802478
rect 700208 802467 700242 802478
rect 700276 802467 700310 802478
rect 700934 802467 700968 802478
rect 701002 802467 701036 802478
rect 701070 802467 701104 802478
rect 701138 802467 701172 802478
rect 701206 802467 701240 802478
rect 701274 802467 701308 802478
rect 701342 802467 701376 802478
rect 701410 802467 701444 802478
rect 701478 802467 701512 802478
rect 701546 802467 701580 802478
rect 701614 802467 701648 802478
rect 701682 802467 701716 802478
rect 701750 802467 701784 802478
rect 701818 802467 701852 802478
rect 699392 802457 699450 802467
rect 699460 802457 699518 802467
rect 699528 802457 699586 802467
rect 699596 802457 699654 802467
rect 699664 802457 699722 802467
rect 699732 802457 699790 802467
rect 699800 802457 699858 802467
rect 699868 802457 699926 802467
rect 699936 802457 699994 802467
rect 700004 802457 700062 802467
rect 700072 802457 700130 802467
rect 700140 802457 700198 802467
rect 700208 802457 700266 802467
rect 700276 802457 700334 802467
rect 700934 802457 700992 802467
rect 701002 802457 701060 802467
rect 701070 802457 701128 802467
rect 701138 802457 701196 802467
rect 701206 802457 701264 802467
rect 701274 802457 701332 802467
rect 701342 802457 701400 802467
rect 701410 802457 701468 802467
rect 701478 802457 701536 802467
rect 701546 802457 701604 802467
rect 701614 802457 701672 802467
rect 701682 802457 701740 802467
rect 701750 802457 701808 802467
rect 701818 802457 701876 802467
rect 696203 802416 696249 802450
rect 699368 802433 700334 802457
rect 700910 802433 701876 802457
rect 699392 802418 699416 802433
rect 699460 802418 699484 802433
rect 699528 802418 699552 802433
rect 699596 802418 699620 802433
rect 699664 802418 699688 802433
rect 699732 802418 699756 802433
rect 699800 802418 699824 802433
rect 699868 802418 699892 802433
rect 699936 802418 699960 802433
rect 700004 802418 700028 802433
rect 700072 802418 700096 802433
rect 700140 802418 700164 802433
rect 700208 802418 700232 802433
rect 700276 802418 700300 802433
rect 700934 802418 700958 802433
rect 701002 802418 701026 802433
rect 701070 802418 701094 802433
rect 701138 802418 701162 802433
rect 701206 802418 701230 802433
rect 701274 802418 701298 802433
rect 701342 802418 701366 802433
rect 701410 802418 701434 802433
rect 701478 802418 701502 802433
rect 701546 802418 701570 802433
rect 701614 802418 701638 802433
rect 701682 802418 701706 802433
rect 701750 802418 701774 802433
rect 701818 802418 701842 802433
rect 696203 802382 696223 802416
rect 696227 802382 696245 802416
rect 692485 802348 692521 802382
rect 696203 802348 696249 802382
rect 679549 802307 679573 802330
rect 679793 802306 679808 802330
rect 692485 802314 692505 802348
rect 692509 802314 692517 802348
rect 696203 802314 696223 802348
rect 696227 802314 696245 802348
rect 692485 802280 692521 802314
rect 696203 802280 696249 802314
rect 679549 802237 679573 802271
rect 692485 802246 692505 802280
rect 692509 802246 692517 802280
rect 692485 802212 692521 802246
rect 692583 802237 693983 802280
rect 694719 802237 696119 802280
rect 696203 802246 696223 802280
rect 696227 802246 696245 802280
rect 699322 802263 700322 802418
rect 696203 802212 696249 802246
rect 699322 802229 700334 802263
rect 700922 802253 701922 802418
rect 700910 802229 701922 802253
rect 699322 802218 700322 802229
rect 700922 802218 701922 802229
rect 707574 802263 708646 802299
rect 707574 802226 707610 802263
rect 708610 802226 708646 802263
rect 679549 802167 679573 802201
rect 685542 802160 686142 802210
rect 685601 802157 685895 802160
rect 685920 802157 686142 802160
rect 692485 802178 692505 802212
rect 692509 802178 692517 802212
rect 696203 802178 696223 802212
rect 696227 802178 696245 802212
rect 699392 802205 699416 802218
rect 699460 802205 699484 802218
rect 699528 802205 699552 802218
rect 699596 802205 699620 802218
rect 699664 802205 699688 802218
rect 699732 802205 699756 802218
rect 699800 802205 699824 802218
rect 699868 802205 699892 802218
rect 699936 802205 699960 802218
rect 700004 802205 700028 802218
rect 700072 802205 700096 802218
rect 700140 802205 700164 802218
rect 700208 802205 700232 802218
rect 700276 802205 700300 802218
rect 700934 802205 700958 802218
rect 701002 802205 701026 802218
rect 701070 802205 701094 802218
rect 701138 802205 701162 802218
rect 701206 802205 701230 802218
rect 701274 802205 701298 802218
rect 701342 802205 701366 802218
rect 701410 802205 701434 802218
rect 701478 802205 701502 802218
rect 701546 802205 701570 802218
rect 701614 802205 701638 802218
rect 701682 802205 701706 802218
rect 701750 802205 701774 802218
rect 701818 802205 701842 802218
rect 707574 802186 708646 802226
rect 709175 802263 710247 802299
rect 709175 802226 709211 802263
rect 710211 802226 710247 802263
rect 709175 802186 710247 802226
rect 692485 802144 692521 802178
rect 696203 802144 696249 802178
rect 679549 802097 679573 802131
rect 692485 802110 692505 802144
rect 692509 802110 692517 802144
rect 692485 802076 692521 802110
rect 692583 802101 693983 802144
rect 694719 802101 696119 802144
rect 696203 802110 696223 802144
rect 696227 802110 696245 802144
rect 696203 802076 696249 802110
rect 679549 802027 679573 802061
rect 692485 802042 692505 802076
rect 692509 802042 692517 802076
rect 692485 802008 692521 802042
rect 679549 801957 679573 801991
rect 692485 801974 692505 802008
rect 692509 801974 692517 802008
rect 679793 801933 679808 801957
rect 692485 801940 692521 801974
rect 679817 801909 679841 801933
rect 692485 801906 692505 801940
rect 692509 801906 692517 801940
rect 692583 801938 693983 802066
rect 694719 801938 696119 802066
rect 696203 802042 696223 802076
rect 696227 802042 696245 802076
rect 696203 802008 696249 802042
rect 696203 801974 696223 802008
rect 696227 801974 696245 802008
rect 696203 801940 696249 801974
rect 696203 801906 696223 801940
rect 696227 801906 696245 801940
rect 687685 801838 687709 801862
rect 687661 801814 687675 801838
rect 687669 801797 687675 801814
rect 679515 801762 679539 801785
rect 679613 801762 679637 801785
rect 679491 801737 679515 801761
rect 679637 801737 679661 801761
rect 680215 801678 680815 801728
rect 680215 801502 680815 801558
rect 685551 801516 686551 801566
rect 680215 801326 680815 801382
rect 685551 801360 686551 801488
rect 689154 801439 689204 801897
rect 689151 801355 689204 801439
rect 680215 801156 680815 801206
rect 685551 801204 686551 801332
rect 685551 801048 686551 801176
rect 686865 801116 687465 801166
rect 679007 800980 679607 801030
rect 680615 800885 680630 800900
rect 680803 800896 680815 800900
rect 680800 800885 680815 800896
rect 685551 800892 686551 800948
rect 686865 800940 687465 801068
rect 679007 800810 679607 800860
rect 680615 800705 680815 800885
rect 683328 800793 683928 800843
rect 682573 800717 683173 800767
rect 680615 800690 680630 800705
rect 680800 800694 680815 800705
rect 680803 800690 680815 800694
rect 680502 800649 680517 800664
rect 680480 800469 680517 800649
rect 680502 800454 680517 800469
rect 680615 800649 680630 800664
rect 680803 800660 680815 800664
rect 680800 800649 680815 800660
rect 680615 800469 680815 800649
rect 682573 800541 683173 800669
rect 683328 800617 683928 800745
rect 685551 800736 686551 800864
rect 686865 800764 687465 800820
rect 685551 800580 686551 800708
rect 686865 800588 687465 800716
rect 680615 800454 680630 800469
rect 680800 800458 680815 800469
rect 680803 800454 680815 800458
rect 683328 800441 683928 800497
rect 679002 800384 679602 800434
rect 685551 800424 686551 800552
rect 682573 800365 683173 800421
rect 686865 800412 687465 800468
rect 679002 800208 679602 800264
rect 682573 800189 683173 800317
rect 683328 800265 683928 800321
rect 685551 800274 686551 800324
rect 686865 800236 687465 800364
rect 685551 800158 686551 800208
rect 678680 800123 678704 800157
rect 678680 800055 678704 800089
rect 679002 800038 679602 800088
rect 679061 800035 679355 800038
rect 679380 800035 679602 800038
rect 678680 799987 678704 800021
rect 682573 800013 683173 800141
rect 683328 800089 683928 800145
rect 678680 799919 678704 799953
rect 678680 799851 678704 799885
rect 682573 799837 683173 799965
rect 683328 799913 683928 800041
rect 685551 799982 686551 800110
rect 686865 800060 687465 800116
rect 678680 799783 678704 799817
rect 685551 799806 686551 799934
rect 686865 799884 687465 800012
rect 678680 799715 678704 799749
rect 678680 799647 678704 799681
rect 682573 799661 683173 799789
rect 683328 799737 683928 799793
rect 685551 799630 686551 799758
rect 686865 799708 687465 799836
rect 678680 799579 678704 799613
rect 683328 799567 683928 799617
rect 678680 799511 678704 799545
rect 682573 799491 683173 799541
rect 684519 799498 685119 799548
rect 678680 799443 678704 799477
rect 685551 799454 686551 799582
rect 686865 799532 687465 799660
rect 679133 799409 679283 799421
rect 679452 799409 679602 799421
rect 678680 799375 678704 799409
rect 2850 799304 3850 799320
rect 2850 799188 3850 799238
rect 2850 798978 3850 799028
rect 3959 799015 3960 799320
rect 5169 799315 5191 799320
rect 6005 799305 6021 799320
rect 1288 797503 1338 798503
rect 1438 797503 1566 798060
rect 1594 797503 1644 798503
rect 5995 797493 6021 799275
rect 7389 798911 8389 798967
rect 8990 798911 9990 798967
rect 15678 798956 16678 799012
rect 17278 798956 18278 799012
rect 7389 798839 8389 798895
rect 8990 798839 9990 798895
rect 15678 798884 16678 798940
rect 17278 798884 18278 798940
rect 27622 798903 27672 799320
rect 27772 798903 27828 799320
rect 27928 798903 27984 799320
rect 28084 798903 28140 799320
rect 28240 798903 28296 799320
rect 28396 798903 28446 799320
rect 678680 799307 678704 799341
rect 31049 799234 32049 799284
rect 36785 799242 37385 799298
rect 679002 799296 679602 799346
rect 684519 799342 685119 799398
rect 685551 799278 686551 799406
rect 686865 799356 687465 799484
rect 678680 799239 678704 799273
rect 678680 799171 678704 799205
rect 684519 799192 685119 799242
rect 36785 799072 37385 799122
rect 678680 799103 678704 799137
rect 679002 799120 679602 799176
rect 681745 799081 682345 799131
rect 682509 799069 683109 799119
rect 678680 799035 678704 799069
rect 683739 799027 684339 799077
rect 684519 799062 685119 799112
rect 685551 799102 686551 799230
rect 686865 799180 687465 799308
rect 678680 798967 678704 799001
rect 679002 798950 679602 799000
rect 678680 798899 678704 798933
rect 680502 798915 680517 798930
rect 678680 798831 678704 798865
rect 678680 798763 678704 798797
rect 680480 798735 680517 798915
rect 21481 798656 22881 798699
rect 23617 798656 25017 798699
rect 678680 798695 678704 798729
rect 680502 798720 680517 798735
rect 680615 798915 680630 798930
rect 680803 798926 680815 798930
rect 680800 798915 680815 798926
rect 681745 798925 682345 798981
rect 680615 798735 680815 798915
rect 681745 798769 682345 798897
rect 682509 798893 683109 799021
rect 684519 798906 685119 799034
rect 685551 798926 686551 799054
rect 686865 799004 687465 799060
rect 683739 798837 684339 798893
rect 686865 798828 687465 798956
rect 680615 798720 680630 798735
rect 680800 798724 680815 798735
rect 680803 798720 680815 798724
rect 680615 798679 680630 798694
rect 680803 798690 680815 798694
rect 680800 798679 680815 798690
rect 31458 798590 32058 798640
rect 678680 798627 678704 798661
rect 15678 798382 16678 798522
rect 17278 798382 18278 798522
rect 21481 798520 22881 798563
rect 23617 798520 25017 798563
rect 678680 798559 678704 798593
rect 678680 798491 678704 798525
rect 679007 798524 679607 798574
rect 680615 798499 680815 798679
rect 681745 798613 682345 798741
rect 682509 798717 683109 798773
rect 684519 798750 685119 798806
rect 685551 798750 686551 798806
rect 682509 798541 683109 798669
rect 684519 798594 685119 798722
rect 685551 798594 686551 798722
rect 686865 798652 687465 798780
rect 680615 798484 680630 798499
rect 680800 798488 680815 798499
rect 680803 798484 680815 798488
rect 31458 798414 32058 798470
rect 681745 798463 682345 798513
rect 683739 798477 684339 798513
rect 678680 798423 678704 798457
rect 684519 798444 685119 798494
rect 685551 798438 686551 798566
rect 686865 798476 687465 798604
rect 678680 798355 678704 798389
rect 679007 798354 679607 798404
rect 682509 798371 683109 798421
rect 25725 798197 26325 798247
rect 31458 798244 32058 798294
rect 678680 798287 678704 798321
rect 684519 798314 685119 798364
rect 678680 798219 678704 798253
rect 7353 798016 8425 798052
rect 7353 797975 7389 798016
rect 8389 797975 8425 798016
rect 7353 797919 8425 797975
rect 7353 797903 7389 797919
rect 8389 797903 8425 797919
rect 7353 797847 8425 797903
rect 7353 797810 7389 797847
rect 8389 797810 8425 797847
rect 7353 797770 8425 797810
rect 8954 798016 10026 798052
rect 8954 797975 8990 798016
rect 9990 797975 10026 798016
rect 8954 797919 10026 797975
rect 21383 798044 21403 798060
rect 21407 798044 21415 798060
rect 21383 798010 21419 798044
rect 21481 798031 22881 798060
rect 23617 798031 25017 798060
rect 25101 798044 25121 798060
rect 25125 798044 25143 798060
rect 25725 798047 26325 798097
rect 25101 798010 25147 798044
rect 21383 797976 21403 798010
rect 21407 797976 21415 798010
rect 21383 797942 21419 797976
rect 8954 797903 8990 797919
rect 9990 797903 10026 797919
rect 15678 797906 16678 797923
rect 17278 797906 18278 797923
rect 21383 797908 21403 797942
rect 21407 797908 21415 797942
rect 8954 797847 10026 797903
rect 20250 797890 20316 797906
rect 8954 797810 8990 797847
rect 9990 797810 10026 797847
rect 8954 797770 10026 797810
rect 21383 797874 21419 797908
rect 21383 797840 21403 797874
rect 21407 797840 21415 797874
rect 21481 797868 22881 797996
rect 23617 797868 25017 797996
rect 25101 797976 25121 798010
rect 25125 797976 25143 798010
rect 25101 797942 25147 797976
rect 25101 797908 25121 797942
rect 25125 797908 25143 797942
rect 25725 797925 26325 797975
rect 25101 797874 25147 797908
rect 25101 797840 25121 797874
rect 25125 797840 25143 797874
rect 21383 797806 21419 797840
rect 21383 797772 21403 797806
rect 21407 797772 21415 797806
rect 21383 797738 21419 797772
rect 15678 797703 16678 797736
rect 17278 797703 18278 797736
rect 21383 797704 21403 797738
rect 21407 797704 21415 797738
rect 21481 797705 22881 797833
rect 23617 797705 25017 797833
rect 25101 797806 25147 797840
rect 25101 797772 25121 797806
rect 25125 797772 25143 797806
rect 25725 797775 26325 797825
rect 25101 797738 25147 797772
rect 25101 797704 25121 797738
rect 25125 797704 25143 797738
rect 21383 797670 21419 797704
rect 25101 797670 25147 797704
rect 21383 797636 21403 797670
rect 21407 797636 21415 797670
rect 7389 797559 8389 797631
rect 8990 797559 9990 797631
rect 21383 797602 21419 797636
rect 15840 797510 15870 797580
rect 15878 797546 15908 797580
rect 21383 797568 21403 797602
rect 21407 797568 21415 797602
rect 15853 797508 15870 797510
rect 21383 797534 21419 797568
rect 21481 797542 22881 797670
rect 23617 797542 25017 797670
rect 25101 797636 25121 797670
rect 25125 797636 25143 797670
rect 25725 797649 26325 797699
rect 25101 797602 25147 797636
rect 25101 797568 25121 797602
rect 25125 797568 25143 797602
rect 25101 797534 25147 797568
rect 5981 797483 6021 797493
rect 5137 797469 6021 797483
rect 21383 797500 21403 797534
rect 21407 797500 21415 797534
rect 21383 797466 21419 797500
rect 7389 797369 8389 797463
rect 7389 797359 8413 797369
rect 8990 797359 9990 797463
rect 21383 797432 21403 797466
rect 21407 797432 21415 797466
rect 21383 797398 21419 797432
rect 21383 797364 21403 797398
rect 21407 797364 21415 797398
rect 21481 797379 22881 797507
rect 23617 797379 25017 797507
rect 25101 797500 25121 797534
rect 25125 797500 25143 797534
rect 25101 797466 25147 797500
rect 25725 797499 26325 797549
rect 25101 797432 25121 797466
rect 25125 797432 25143 797466
rect 25101 797398 25147 797432
rect 25101 797364 25121 797398
rect 25125 797364 25143 797398
rect 25725 797377 26325 797427
rect 21383 797330 21419 797364
rect 25101 797330 25147 797364
rect 21383 797296 21403 797330
rect 21407 797296 21415 797330
rect 25101 797296 25121 797330
rect 25125 797296 25143 797330
rect 21383 797262 21419 797296
rect 21383 797228 21403 797262
rect 21407 797228 21415 797262
rect 21481 797229 22881 797272
rect 23617 797229 25017 797272
rect 25101 797262 25147 797296
rect 25101 797228 25121 797262
rect 25125 797228 25143 797262
rect 21383 797194 21419 797228
rect 25101 797194 25147 797228
rect 25725 797227 26325 797277
rect 21383 797160 21403 797194
rect 21407 797160 21415 797194
rect 25101 797160 25121 797194
rect 25125 797160 25143 797194
rect 27162 797170 27212 798170
rect 27312 797170 27440 798060
rect 27468 797170 27596 798060
rect 27624 797170 27752 798060
rect 27780 797170 27908 798060
rect 27936 797170 28064 798060
rect 28092 797170 28220 798060
rect 28248 797170 28376 798060
rect 28404 797170 28532 798060
rect 28560 797170 28688 798060
rect 28716 797170 28844 798060
rect 28872 797170 29000 798060
rect 29028 797170 29156 798060
rect 29184 797170 29312 798060
rect 29340 797170 29390 798170
rect 30245 798029 30445 798209
rect 30245 798018 30260 798029
rect 30245 798014 30257 798018
rect 30430 798014 30445 798029
rect 30543 798029 30580 798209
rect 678680 798151 678704 798185
rect 680215 798178 680815 798228
rect 681745 798209 682345 798259
rect 678680 798083 678704 798117
rect 30543 798014 30558 798029
rect 678680 798015 678704 798049
rect 680215 798002 680815 798058
rect 681745 798053 682345 798181
rect 682509 798030 683109 798080
rect 30245 797984 30257 797988
rect 30245 797973 30260 797984
rect 30430 797973 30445 797988
rect 30245 797793 30445 797973
rect 678680 797947 678704 797981
rect 678680 797879 678704 797913
rect 681745 797897 682345 797953
rect 31453 797818 32053 797868
rect 678680 797811 678704 797845
rect 680215 797826 680815 797882
rect 30245 797782 30260 797793
rect 30245 797778 30257 797782
rect 30430 797778 30445 797793
rect 678680 797743 678704 797777
rect 681745 797741 682345 797869
rect 682509 797854 683109 797910
rect 31453 797648 32053 797698
rect 678680 797675 678704 797709
rect 680215 797656 680815 797706
rect 682509 797684 683109 797734
rect 683248 797680 683298 798268
rect 683398 797680 683448 798268
rect 684519 798158 685119 798286
rect 685551 798282 686551 798410
rect 686865 798300 687465 798428
rect 684519 798002 685119 798130
rect 685551 798126 686551 798254
rect 686865 798124 687465 798252
rect 685551 797970 686551 798098
rect 686865 797954 687465 798004
rect 684519 797852 685119 797902
rect 685551 797814 686551 797870
rect 686865 797838 687465 797888
rect 683248 797668 683448 797680
rect 685551 797658 686551 797786
rect 686865 797662 687465 797790
rect 678680 797607 678704 797641
rect 681745 797591 682345 797641
rect 683571 797605 683581 797646
rect 678680 797539 678704 797573
rect 680215 797524 680815 797574
rect 682509 797555 683509 797605
rect 30245 797472 30845 797522
rect 678680 797471 678704 797505
rect 685551 797502 686551 797630
rect 686865 797486 687465 797542
rect 678680 797403 678704 797437
rect 30245 797296 30845 797352
rect 678680 797335 678704 797369
rect 680215 797348 680815 797404
rect 681745 797389 682345 797439
rect 682509 797385 683509 797435
rect 683278 797382 683398 797385
rect 683571 797382 683581 797385
rect 685551 797346 686551 797474
rect 678680 797267 678704 797301
rect 678680 797199 678704 797233
rect 21383 797126 21419 797160
rect 25101 797126 25147 797160
rect 21383 797102 21403 797126
rect 21385 797048 21403 797102
rect 21407 797082 21415 797126
rect 25101 797102 25121 797126
rect 25113 797082 25121 797102
rect 25125 797048 25143 797126
rect 30245 797120 30845 797176
rect 680215 797172 680815 797228
rect 681745 797213 682345 797341
rect 682509 797247 683109 797297
rect 678680 797131 678704 797165
rect 678680 797063 678704 797097
rect 678654 797013 678680 797039
rect 680215 797002 680815 797052
rect 681745 797037 682345 797093
rect 682509 797071 683109 797127
rect 30245 796950 30845 797000
rect 678680 796929 678704 796963
rect 21000 796800 21003 796920
rect 21352 796885 21376 796909
rect 25122 796885 25146 796909
rect 21385 796861 21400 796885
rect 25098 796861 25113 796885
rect 678680 796861 678704 796895
rect 21274 796783 21294 796851
rect 21410 796817 21430 796851
rect 25068 796817 25088 796851
rect 25204 796817 25224 796851
rect 21385 796807 21430 796817
rect 25102 796807 25137 796817
rect 21361 796783 21430 796807
rect 25089 796783 25137 796807
rect 25238 796783 25258 796817
rect 678680 796793 678704 796827
rect 679007 796826 679607 796876
rect 681745 796867 682345 796917
rect 682509 796901 683109 796951
rect 678680 796725 678704 796759
rect 680615 796731 680630 796746
rect 680803 796742 680815 796746
rect 680800 796731 680815 796742
rect 678680 796657 678704 796691
rect 679007 796656 679607 796706
rect 678680 796589 678704 796623
rect 678680 796521 678704 796555
rect 680615 796551 680815 796731
rect 681345 796651 682345 796701
rect 682508 796631 683108 796681
rect 680615 796536 680630 796551
rect 680800 796540 680815 796551
rect 680803 796536 680815 796540
rect 680502 796495 680517 796510
rect 678680 796453 678704 796487
rect 678680 796385 678704 796419
rect 678680 796317 678704 796351
rect 680480 796315 680517 796495
rect 680502 796300 680517 796315
rect 680615 796495 680630 796510
rect 680803 796506 680815 796510
rect 680800 796495 680815 796506
rect 680615 796315 680815 796495
rect 681345 796475 682345 796531
rect 682508 796455 683108 796511
rect 680615 796300 680630 796315
rect 680800 796304 680815 796315
rect 680803 796300 680815 796304
rect 681345 796299 682345 796427
rect 682508 796285 683108 796335
rect 683228 796322 683278 797322
rect 683398 796322 683448 797322
rect 685551 797190 686551 797318
rect 686865 797310 687465 797438
rect 685551 797034 686551 797162
rect 686865 797140 687465 797190
rect 686865 797024 687465 797074
rect 685551 796884 686551 796934
rect 686865 796848 687465 796976
rect 685551 796768 686551 796818
rect 686865 796672 687465 796800
rect 684404 796609 685004 796659
rect 685551 796612 686551 796668
rect 685551 796456 686551 796512
rect 686865 796496 687465 796624
rect 685551 796300 686551 796356
rect 686865 796320 687465 796376
rect 678680 796249 678704 796283
rect 679002 796230 679602 796280
rect 678680 796181 678704 796215
rect 678680 796113 678704 796147
rect 681345 796129 682345 796179
rect 684404 796175 685004 796225
rect 685551 796150 686551 796200
rect 686865 796150 687465 796200
rect 678680 796045 678704 796079
rect 679002 796054 679602 796110
rect 681390 796070 681424 796080
rect 681458 796070 681492 796080
rect 681526 796070 681560 796080
rect 681594 796070 681628 796080
rect 681662 796070 681696 796080
rect 681730 796070 681764 796080
rect 681798 796070 681832 796080
rect 681866 796070 681900 796080
rect 681934 796070 681968 796080
rect 682002 796070 682036 796080
rect 682077 796070 682111 796080
rect 682145 796070 682179 796080
rect 682213 796070 682247 796080
rect 682281 796070 682315 796080
rect 681345 796034 682345 796046
rect 678680 795977 678704 796011
rect 678680 795909 678704 795943
rect 679002 795884 679602 795934
rect 681345 795927 682345 795977
rect 684004 795973 685004 796023
rect 685551 796014 686551 796064
rect 686865 796034 687465 796084
rect 679061 795881 679355 795884
rect 679380 795881 679602 795884
rect 678680 795841 678704 795875
rect 678680 795773 678704 795807
rect 681345 795751 682345 795879
rect 684004 795817 685004 795873
rect 685551 795858 686551 795914
rect 686865 795858 687465 795914
rect 686686 795812 686714 795840
rect 678680 795705 678704 795739
rect 678680 795637 678704 795671
rect 678680 795569 678704 795603
rect 681345 795575 682345 795703
rect 684004 795661 685004 795789
rect 685551 795708 686551 795758
rect 686865 795688 687465 795738
rect 678680 795501 678704 795535
rect 684004 795505 685004 795633
rect 687573 795554 687585 801277
rect 689154 801107 689204 801355
rect 689151 801023 689204 801107
rect 689154 800897 689204 801023
rect 689304 800897 689360 801897
rect 689460 800897 689516 801897
rect 689616 800897 689672 801897
rect 689772 800897 689828 801897
rect 689928 800897 689978 801897
rect 692485 801872 692521 801906
rect 692485 801838 692505 801872
rect 692509 801838 692517 801872
rect 690952 801509 691122 801815
rect 692485 801804 692521 801838
rect 692485 801770 692505 801804
rect 692509 801770 692517 801804
rect 692583 801775 693983 801903
rect 694719 801775 696119 801903
rect 696203 801872 696249 801906
rect 696203 801838 696223 801872
rect 696227 801838 696245 801872
rect 699322 801860 700322 801916
rect 700922 801860 701922 801916
rect 707610 801905 708610 801961
rect 709211 801905 710211 801961
rect 696203 801804 696249 801838
rect 696203 801770 696223 801804
rect 696227 801770 696245 801804
rect 699322 801788 700322 801844
rect 700922 801788 701922 801844
rect 707610 801833 708610 801889
rect 709211 801833 710211 801889
rect 692485 801736 692521 801770
rect 692485 801702 692505 801736
rect 692509 801702 692517 801736
rect 692485 801668 692521 801702
rect 692485 801634 692505 801668
rect 692509 801634 692517 801668
rect 692485 801600 692521 801634
rect 692583 801612 693983 801740
rect 694719 801612 696119 801740
rect 696203 801736 696249 801770
rect 696203 801702 696223 801736
rect 696227 801702 696245 801736
rect 696203 801668 696249 801702
rect 696203 801634 696223 801668
rect 696227 801634 696245 801668
rect 696203 801600 696249 801634
rect 692485 801566 692505 801600
rect 692509 801566 692517 801600
rect 692485 801532 692521 801566
rect 692485 801498 692505 801532
rect 692509 801498 692517 801532
rect 692485 801464 692521 801498
rect 692485 801430 692505 801464
rect 692509 801430 692517 801464
rect 692583 801449 693983 801577
rect 694719 801449 696119 801577
rect 696203 801566 696223 801600
rect 696227 801566 696245 801600
rect 696203 801532 696249 801566
rect 696203 801498 696223 801532
rect 696227 801498 696245 801532
rect 696203 801464 696249 801498
rect 699322 801486 700322 801558
rect 700922 801486 701922 801558
rect 707610 801531 708610 801603
rect 709211 801531 710211 801603
rect 711579 801553 711605 803307
rect 715956 802297 716006 803297
rect 716106 802297 716234 803297
rect 716262 802297 716312 803297
rect 699392 801475 699426 801486
rect 699460 801475 699494 801486
rect 699528 801475 699562 801486
rect 699596 801475 699630 801486
rect 699664 801475 699698 801486
rect 699732 801475 699766 801486
rect 699800 801475 699834 801486
rect 699868 801475 699902 801486
rect 699936 801475 699970 801486
rect 700004 801475 700038 801486
rect 700072 801475 700106 801486
rect 700140 801475 700174 801486
rect 700208 801475 700242 801486
rect 700276 801475 700310 801486
rect 700934 801475 700968 801486
rect 701002 801475 701036 801486
rect 701070 801475 701104 801486
rect 701138 801475 701172 801486
rect 701206 801475 701240 801486
rect 701274 801475 701308 801486
rect 701342 801475 701376 801486
rect 701410 801475 701444 801486
rect 701478 801475 701512 801486
rect 701546 801475 701580 801486
rect 701614 801475 701648 801486
rect 701682 801475 701716 801486
rect 701750 801475 701784 801486
rect 701818 801475 701852 801486
rect 711511 801485 711663 801553
rect 712447 801501 712557 801511
rect 711579 801482 711663 801485
rect 699392 801465 699450 801475
rect 699460 801465 699518 801475
rect 699528 801465 699586 801475
rect 699596 801465 699654 801475
rect 699664 801465 699722 801475
rect 699732 801465 699790 801475
rect 699800 801465 699858 801475
rect 699868 801465 699926 801475
rect 699936 801465 699994 801475
rect 700004 801465 700062 801475
rect 700072 801465 700130 801475
rect 700140 801465 700198 801475
rect 700208 801465 700266 801475
rect 700276 801465 700334 801475
rect 700934 801465 700992 801475
rect 701002 801465 701060 801475
rect 701070 801465 701128 801475
rect 701138 801465 701196 801475
rect 701206 801465 701264 801475
rect 701274 801465 701332 801475
rect 701342 801465 701400 801475
rect 701410 801465 701468 801475
rect 701478 801465 701536 801475
rect 701546 801465 701604 801475
rect 701614 801465 701672 801475
rect 701682 801465 701740 801475
rect 701750 801465 701808 801475
rect 701818 801465 701876 801475
rect 696203 801430 696223 801464
rect 696227 801430 696245 801464
rect 699368 801441 700334 801465
rect 700910 801441 701876 801465
rect 711541 801461 711633 801482
rect 692485 801396 692521 801430
rect 692485 801362 692505 801396
rect 692509 801362 692517 801396
rect 692485 801328 692521 801362
rect 692485 801294 692505 801328
rect 692509 801294 692517 801328
rect 692485 801260 692521 801294
rect 692583 801286 693983 801414
rect 694719 801286 696119 801414
rect 696203 801396 696249 801430
rect 699392 801426 699416 801441
rect 699460 801426 699484 801441
rect 699528 801426 699552 801441
rect 699596 801426 699620 801441
rect 699664 801426 699688 801441
rect 699732 801426 699756 801441
rect 699800 801426 699824 801441
rect 699868 801426 699892 801441
rect 699936 801426 699960 801441
rect 700004 801426 700028 801441
rect 700072 801426 700096 801441
rect 700140 801426 700164 801441
rect 700208 801426 700232 801441
rect 700276 801426 700300 801441
rect 700934 801426 700958 801441
rect 701002 801426 701026 801441
rect 701070 801426 701094 801441
rect 701138 801426 701162 801441
rect 701206 801426 701230 801441
rect 701274 801426 701298 801441
rect 701342 801426 701366 801441
rect 701410 801426 701434 801441
rect 701478 801426 701502 801441
rect 701546 801426 701570 801441
rect 701614 801426 701638 801441
rect 701682 801426 701706 801441
rect 701750 801426 701774 801441
rect 701818 801426 701842 801441
rect 696203 801362 696223 801396
rect 696227 801362 696245 801396
rect 696203 801328 696249 801362
rect 696203 801294 696223 801328
rect 696227 801294 696245 801328
rect 696203 801260 696249 801294
rect 699322 801271 700322 801426
rect 692485 801226 692505 801260
rect 692509 801226 692517 801260
rect 692485 801192 692521 801226
rect 692485 801158 692505 801192
rect 692509 801158 692517 801192
rect 692485 801124 692521 801158
rect 692485 801090 692505 801124
rect 692509 801090 692517 801124
rect 692583 801123 693983 801251
rect 694719 801123 696119 801251
rect 696203 801226 696223 801260
rect 696227 801226 696245 801260
rect 699322 801237 700334 801271
rect 700922 801261 701922 801426
rect 707610 801271 708610 801331
rect 709211 801271 710211 801331
rect 700910 801237 701922 801261
rect 699322 801226 700322 801237
rect 700922 801226 701922 801237
rect 696203 801192 696249 801226
rect 699392 801213 699416 801226
rect 699460 801213 699484 801226
rect 699528 801213 699552 801226
rect 699596 801213 699620 801226
rect 699664 801213 699688 801226
rect 699732 801213 699756 801226
rect 699800 801213 699824 801226
rect 699868 801213 699892 801226
rect 699936 801213 699960 801226
rect 700004 801213 700028 801226
rect 700072 801213 700096 801226
rect 700140 801213 700164 801226
rect 700208 801213 700232 801226
rect 700276 801213 700300 801226
rect 700934 801213 700958 801226
rect 701002 801213 701026 801226
rect 701070 801213 701094 801226
rect 701138 801213 701162 801226
rect 701206 801213 701230 801226
rect 701274 801213 701298 801226
rect 701342 801213 701366 801226
rect 701410 801213 701434 801226
rect 701478 801213 701502 801226
rect 701546 801213 701570 801226
rect 701614 801213 701638 801226
rect 701682 801213 701706 801226
rect 701750 801213 701774 801226
rect 701818 801213 701842 801226
rect 696203 801158 696223 801192
rect 696227 801158 696245 801192
rect 696203 801124 696249 801158
rect 696203 801090 696223 801124
rect 696227 801090 696245 801124
rect 692485 801056 692521 801090
rect 696203 801056 696249 801090
rect 692485 801022 692505 801056
rect 692509 801022 692517 801056
rect 696203 801022 696223 801056
rect 696227 801022 696245 801056
rect 692485 800988 692521 801022
rect 692485 800954 692505 800988
rect 692509 800954 692517 800988
rect 692583 800966 693983 801016
rect 694719 800966 696119 801016
rect 696203 800988 696249 801022
rect 696203 800954 696223 800988
rect 696227 800954 696245 800988
rect 692485 800920 692521 800954
rect 696203 800920 696249 800954
rect 692485 800896 692505 800920
rect 692487 800852 692505 800896
rect 692509 800886 692517 800920
rect 696203 800896 696223 800920
rect 696215 800886 696223 800896
rect 696227 800852 696245 800920
rect 697284 800870 697350 800886
rect 699322 800868 700322 800924
rect 700922 800868 701922 800924
rect 707610 800913 708610 800969
rect 709211 800913 710211 800969
rect 692174 800787 692186 800811
rect 692288 800787 692312 800811
rect 696390 800787 696414 800811
rect 696516 800787 696528 800811
rect 699322 800796 700322 800852
rect 700922 800796 701922 800852
rect 707610 800841 708610 800897
rect 709211 800841 710211 800897
rect 692264 800763 692288 800777
rect 696414 800763 696438 800777
rect 692288 800729 692312 800753
rect 696390 800729 696414 800753
rect 688940 800475 688990 800675
rect 689110 800475 689238 800675
rect 689286 800475 689342 800675
rect 689462 800475 689590 800675
rect 689638 800559 689688 800675
rect 692736 800597 695966 800699
rect 689638 800475 689691 800559
rect 699322 800494 700322 800566
rect 700922 800494 701922 800566
rect 707610 800539 708610 800611
rect 709211 800539 710211 800611
rect 699392 800483 699426 800494
rect 699460 800483 699494 800494
rect 699528 800483 699562 800494
rect 699596 800483 699630 800494
rect 699664 800483 699698 800494
rect 699732 800483 699766 800494
rect 699800 800483 699834 800494
rect 699868 800483 699902 800494
rect 699936 800483 699970 800494
rect 700004 800483 700038 800494
rect 700072 800483 700106 800494
rect 700140 800483 700174 800494
rect 700208 800483 700242 800494
rect 700276 800483 700310 800494
rect 700934 800483 700968 800494
rect 701002 800483 701036 800494
rect 701070 800483 701104 800494
rect 701138 800483 701172 800494
rect 701206 800483 701240 800494
rect 701274 800483 701308 800494
rect 701342 800483 701376 800494
rect 701410 800483 701444 800494
rect 701478 800483 701512 800494
rect 701546 800483 701580 800494
rect 701614 800483 701648 800494
rect 701682 800483 701716 800494
rect 701750 800483 701784 800494
rect 701818 800483 701852 800494
rect 689649 800471 689683 800475
rect 699392 800473 699450 800483
rect 699460 800473 699518 800483
rect 699528 800473 699586 800483
rect 699596 800473 699654 800483
rect 699664 800473 699722 800483
rect 699732 800473 699790 800483
rect 699800 800473 699858 800483
rect 699868 800473 699926 800483
rect 699936 800473 699994 800483
rect 700004 800473 700062 800483
rect 700072 800473 700130 800483
rect 700140 800473 700198 800483
rect 700208 800473 700266 800483
rect 700276 800473 700334 800483
rect 700934 800473 700992 800483
rect 701002 800473 701060 800483
rect 701070 800473 701128 800483
rect 701138 800473 701196 800483
rect 701206 800473 701264 800483
rect 701274 800473 701332 800483
rect 701342 800473 701400 800483
rect 701410 800473 701468 800483
rect 701478 800473 701536 800483
rect 701546 800473 701604 800483
rect 701614 800473 701672 800483
rect 701682 800473 701740 800483
rect 701750 800473 701808 800483
rect 701818 800473 701876 800483
rect 692451 800444 692475 800468
rect 692509 800444 692533 800468
rect 696169 800444 696193 800468
rect 696227 800444 696251 800468
rect 699368 800449 700334 800473
rect 700910 800449 701876 800473
rect 692485 800410 692499 800444
rect 696203 800410 696217 800444
rect 699392 800434 699416 800449
rect 699460 800434 699484 800449
rect 699528 800434 699552 800449
rect 699596 800434 699620 800449
rect 699664 800434 699688 800449
rect 699732 800434 699756 800449
rect 699800 800434 699824 800449
rect 699868 800434 699892 800449
rect 699936 800434 699960 800449
rect 700004 800434 700028 800449
rect 700072 800434 700096 800449
rect 700140 800434 700164 800449
rect 700208 800434 700232 800449
rect 700276 800434 700300 800449
rect 700934 800434 700958 800449
rect 701002 800434 701026 800449
rect 701070 800434 701094 800449
rect 701138 800434 701162 800449
rect 701206 800434 701230 800449
rect 701274 800434 701298 800449
rect 701342 800434 701366 800449
rect 701410 800434 701434 800449
rect 701478 800434 701502 800449
rect 701546 800434 701570 800449
rect 701614 800434 701638 800449
rect 701682 800434 701706 800449
rect 701750 800434 701774 800449
rect 701818 800434 701842 800449
rect 692451 800386 692475 800410
rect 692509 800386 692533 800410
rect 696169 800386 696193 800410
rect 696227 800386 696251 800410
rect 690664 800318 691664 800368
rect 692515 800280 693915 800330
rect 694787 800280 696187 800330
rect 699322 800279 700322 800434
rect 699322 800245 700334 800279
rect 700922 800269 701922 800434
rect 703539 800286 703699 800290
rect 707610 800279 708610 800339
rect 709211 800279 710211 800339
rect 700910 800245 701922 800269
rect 690242 800219 690326 800222
rect 690242 800214 690442 800219
rect 690238 800180 690442 800214
rect 690242 800169 690442 800180
rect 690664 800162 691664 800218
rect 687686 800128 687720 800162
rect 687686 800104 687710 800128
rect 689649 800127 689683 800131
rect 688940 799927 688990 800127
rect 689110 799927 689238 800127
rect 689286 799927 689342 800127
rect 689462 799927 689590 800127
rect 689638 800043 689691 800127
rect 689638 799927 689688 800043
rect 690242 799993 690442 800121
rect 692515 800117 693915 800245
rect 694787 800117 696187 800245
rect 699322 800234 700322 800245
rect 700922 800234 701922 800245
rect 699392 800221 699416 800234
rect 699460 800221 699484 800234
rect 699528 800221 699552 800234
rect 699596 800221 699620 800234
rect 699664 800221 699688 800234
rect 699732 800221 699756 800234
rect 699800 800221 699824 800234
rect 699868 800221 699892 800234
rect 699936 800221 699960 800234
rect 700004 800221 700028 800234
rect 700072 800221 700096 800234
rect 700140 800221 700164 800234
rect 700208 800221 700232 800234
rect 700276 800221 700300 800234
rect 700934 800221 700958 800234
rect 701002 800221 701026 800234
rect 701070 800221 701094 800234
rect 701138 800221 701162 800234
rect 701206 800221 701230 800234
rect 701274 800221 701298 800234
rect 701342 800221 701366 800234
rect 701410 800221 701434 800234
rect 701478 800221 701502 800234
rect 701546 800221 701570 800234
rect 701614 800221 701638 800234
rect 701682 800221 701706 800234
rect 701750 800221 701774 800234
rect 701818 800221 701842 800234
rect 703541 800140 703701 800144
rect 690664 800006 691664 800062
rect 692515 799954 693915 800082
rect 694787 799954 696187 800082
rect 690242 799817 690442 799873
rect 690664 799850 691664 799906
rect 692515 799791 693915 799919
rect 694787 799791 696187 799919
rect 699322 799876 700322 799932
rect 700922 799876 701922 799932
rect 707610 799921 708610 799977
rect 709211 799921 710211 799977
rect 699322 799804 700322 799860
rect 700922 799804 701922 799860
rect 707610 799849 708610 799905
rect 709211 799849 710211 799905
rect 689154 799579 689204 799705
rect 687686 799501 687720 799535
rect 687798 799515 687822 799539
rect 687774 799491 687798 799504
rect 689151 799495 689204 799579
rect 687798 799456 687822 799480
rect 689154 799247 689204 799495
rect 689151 799163 689204 799247
rect 689154 798705 689204 799163
rect 689304 798705 689360 799705
rect 689460 798705 689516 799705
rect 689616 798705 689672 799705
rect 689772 798705 689828 799705
rect 689928 798705 689978 799705
rect 690242 799641 690442 799769
rect 690664 799700 691664 799750
rect 690790 799697 690874 799700
rect 691123 799697 691207 799700
rect 692515 799628 693915 799756
rect 694787 799628 696187 799756
rect 704735 799731 705041 799833
rect 704719 799715 705057 799731
rect 690242 799465 690442 799521
rect 692515 799465 693915 799593
rect 694787 799465 696187 799593
rect 699322 799502 700322 799574
rect 700922 799502 701922 799574
rect 707610 799547 708610 799619
rect 709211 799547 710211 799619
rect 699392 799491 699426 799502
rect 699460 799491 699494 799502
rect 699528 799491 699562 799502
rect 699596 799491 699630 799502
rect 699664 799491 699698 799502
rect 699732 799491 699766 799502
rect 699800 799491 699834 799502
rect 699868 799491 699902 799502
rect 699936 799491 699970 799502
rect 700004 799491 700038 799502
rect 700072 799491 700106 799502
rect 700140 799491 700174 799502
rect 700208 799491 700242 799502
rect 700276 799491 700310 799502
rect 700934 799491 700968 799502
rect 701002 799491 701036 799502
rect 701070 799491 701104 799502
rect 701138 799491 701172 799502
rect 701206 799491 701240 799502
rect 701274 799491 701308 799502
rect 701342 799491 701376 799502
rect 701410 799491 701444 799502
rect 701478 799491 701512 799502
rect 701546 799491 701580 799502
rect 701614 799491 701648 799502
rect 701682 799491 701716 799502
rect 701750 799491 701784 799502
rect 701818 799491 701852 799502
rect 699392 799481 699450 799491
rect 699460 799481 699518 799491
rect 699528 799481 699586 799491
rect 699596 799481 699654 799491
rect 699664 799481 699722 799491
rect 699732 799481 699790 799491
rect 699800 799481 699858 799491
rect 699868 799481 699926 799491
rect 699936 799481 699994 799491
rect 700004 799481 700062 799491
rect 700072 799481 700130 799491
rect 700140 799481 700198 799491
rect 700208 799481 700266 799491
rect 700276 799481 700334 799491
rect 700934 799481 700992 799491
rect 701002 799481 701060 799491
rect 701070 799481 701128 799491
rect 701138 799481 701196 799491
rect 701206 799481 701264 799491
rect 701274 799481 701332 799491
rect 701342 799481 701400 799491
rect 701410 799481 701468 799491
rect 701478 799481 701536 799491
rect 701546 799481 701604 799491
rect 701614 799481 701672 799491
rect 701682 799481 701740 799491
rect 701750 799481 701808 799491
rect 701818 799481 701876 799491
rect 699368 799457 700334 799481
rect 700910 799457 701876 799481
rect 699392 799442 699416 799457
rect 699460 799442 699484 799457
rect 699528 799442 699552 799457
rect 699596 799442 699620 799457
rect 699664 799442 699688 799457
rect 699732 799442 699756 799457
rect 699800 799442 699824 799457
rect 699868 799442 699892 799457
rect 699936 799442 699960 799457
rect 700004 799442 700028 799457
rect 700072 799442 700096 799457
rect 700140 799442 700164 799457
rect 700208 799442 700232 799457
rect 700276 799442 700300 799457
rect 700934 799442 700958 799457
rect 701002 799442 701026 799457
rect 701070 799442 701094 799457
rect 701138 799442 701162 799457
rect 701206 799442 701230 799457
rect 701274 799442 701298 799457
rect 701342 799442 701366 799457
rect 701410 799442 701434 799457
rect 701478 799442 701502 799457
rect 701546 799442 701570 799457
rect 701614 799442 701638 799457
rect 701682 799442 701706 799457
rect 701750 799442 701774 799457
rect 701818 799442 701842 799457
rect 690242 799289 690442 799417
rect 692515 799302 693915 799430
rect 694787 799302 696187 799430
rect 690790 799286 690874 799289
rect 691123 799286 691207 799289
rect 699322 799287 700322 799442
rect 690664 799236 691664 799286
rect 699322 799253 700334 799287
rect 700922 799277 701922 799442
rect 707610 799287 708610 799347
rect 709211 799287 710211 799347
rect 700910 799253 701922 799277
rect 699322 799242 700322 799253
rect 700922 799242 701922 799253
rect 699392 799229 699416 799242
rect 699460 799229 699484 799242
rect 699528 799229 699552 799242
rect 699596 799229 699620 799242
rect 699664 799229 699688 799242
rect 699732 799229 699756 799242
rect 699800 799229 699824 799242
rect 699868 799229 699892 799242
rect 699936 799229 699960 799242
rect 700004 799229 700028 799242
rect 700072 799229 700096 799242
rect 700140 799229 700164 799242
rect 700208 799229 700232 799242
rect 700276 799229 700300 799242
rect 700934 799229 700958 799242
rect 701002 799229 701026 799242
rect 701070 799229 701094 799242
rect 701138 799229 701162 799242
rect 701206 799229 701230 799242
rect 701274 799229 701298 799242
rect 701342 799229 701366 799242
rect 701410 799229 701434 799242
rect 701478 799229 701502 799242
rect 701546 799229 701570 799242
rect 701614 799229 701638 799242
rect 701682 799229 701706 799242
rect 701750 799229 701774 799242
rect 701818 799229 701842 799242
rect 690242 799113 690442 799169
rect 692515 799152 693915 799195
rect 694787 799152 696187 799195
rect 690664 799080 691664 799136
rect 690242 798937 690442 799065
rect 692515 799016 693915 799059
rect 694787 799016 696187 799059
rect 690664 798924 691664 798980
rect 692515 798853 693915 798981
rect 694787 798853 696187 798981
rect 703541 798944 703701 798948
rect 699322 798884 700322 798940
rect 700922 798884 701922 798940
rect 707610 798929 708610 798985
rect 709211 798929 710211 798985
rect 690242 798806 690442 798817
rect 690238 798772 690442 798806
rect 690242 798767 690442 798772
rect 690664 798768 691664 798824
rect 690242 798764 690326 798767
rect 692515 798690 693915 798818
rect 694787 798690 696187 798818
rect 699322 798812 700322 798868
rect 700922 798812 701922 798868
rect 707610 798857 708610 798913
rect 709211 798857 710211 798913
rect 703541 798798 703701 798802
rect 690664 798618 691664 798668
rect 692515 798527 693915 798655
rect 694787 798527 696187 798655
rect 699322 798510 700322 798582
rect 700922 798510 701922 798582
rect 707610 798555 708610 798627
rect 709211 798555 710211 798627
rect 699392 798499 699426 798510
rect 699460 798499 699494 798510
rect 699528 798499 699562 798510
rect 699596 798499 699630 798510
rect 699664 798499 699698 798510
rect 699732 798499 699766 798510
rect 699800 798499 699834 798510
rect 699868 798499 699902 798510
rect 699936 798499 699970 798510
rect 700004 798499 700038 798510
rect 700072 798499 700106 798510
rect 700140 798499 700174 798510
rect 700208 798499 700242 798510
rect 700276 798499 700310 798510
rect 700934 798499 700968 798510
rect 701002 798499 701036 798510
rect 701070 798499 701104 798510
rect 701138 798499 701172 798510
rect 701206 798499 701240 798510
rect 701274 798499 701308 798510
rect 701342 798499 701376 798510
rect 701410 798499 701444 798510
rect 701478 798499 701512 798510
rect 701546 798499 701580 798510
rect 701614 798499 701648 798510
rect 701682 798499 701716 798510
rect 701750 798499 701784 798510
rect 701818 798499 701852 798510
rect 692515 798364 693915 798492
rect 694787 798364 696187 798492
rect 699392 798489 699450 798499
rect 699460 798489 699518 798499
rect 699528 798489 699586 798499
rect 699596 798489 699654 798499
rect 699664 798489 699722 798499
rect 699732 798489 699790 798499
rect 699800 798489 699858 798499
rect 699868 798489 699926 798499
rect 699936 798489 699994 798499
rect 700004 798489 700062 798499
rect 700072 798489 700130 798499
rect 700140 798489 700198 798499
rect 700208 798489 700266 798499
rect 700276 798489 700334 798499
rect 700934 798489 700992 798499
rect 701002 798489 701060 798499
rect 701070 798489 701128 798499
rect 701138 798489 701196 798499
rect 701206 798489 701264 798499
rect 701274 798489 701332 798499
rect 701342 798489 701400 798499
rect 701410 798489 701468 798499
rect 701478 798489 701536 798499
rect 701546 798489 701604 798499
rect 701614 798489 701672 798499
rect 701682 798489 701740 798499
rect 701750 798489 701808 798499
rect 701818 798489 701876 798499
rect 699368 798465 700334 798489
rect 700910 798465 701876 798489
rect 699392 798450 699416 798465
rect 699460 798450 699484 798465
rect 699528 798450 699552 798465
rect 699596 798450 699620 798465
rect 699664 798450 699688 798465
rect 699732 798450 699756 798465
rect 699800 798450 699824 798465
rect 699868 798450 699892 798465
rect 699936 798450 699960 798465
rect 700004 798450 700028 798465
rect 700072 798450 700096 798465
rect 700140 798450 700164 798465
rect 700208 798450 700232 798465
rect 700276 798450 700300 798465
rect 700934 798450 700958 798465
rect 701002 798450 701026 798465
rect 701070 798450 701094 798465
rect 701138 798450 701162 798465
rect 701206 798450 701230 798465
rect 701274 798450 701298 798465
rect 701342 798450 701366 798465
rect 701410 798450 701434 798465
rect 701478 798450 701502 798465
rect 701546 798450 701570 798465
rect 701614 798450 701638 798465
rect 701682 798450 701706 798465
rect 701750 798450 701774 798465
rect 701818 798450 701842 798465
rect 692515 798201 693915 798329
rect 694787 798201 696187 798329
rect 699322 798295 700322 798450
rect 699322 798261 700334 798295
rect 700922 798285 701922 798450
rect 707610 798295 708610 798355
rect 709211 798295 710211 798355
rect 700910 798261 701922 798285
rect 699322 798250 700322 798261
rect 700922 798250 701922 798261
rect 699392 798237 699416 798250
rect 699460 798237 699484 798250
rect 699528 798237 699552 798250
rect 699596 798237 699620 798250
rect 699664 798237 699688 798250
rect 699732 798237 699756 798250
rect 699800 798237 699824 798250
rect 699868 798237 699892 798250
rect 699936 798237 699960 798250
rect 700004 798237 700028 798250
rect 700072 798237 700096 798250
rect 700140 798237 700164 798250
rect 700208 798237 700232 798250
rect 700276 798237 700300 798250
rect 700934 798237 700958 798250
rect 701002 798237 701026 798250
rect 701070 798237 701094 798250
rect 701138 798237 701162 798250
rect 701206 798237 701230 798250
rect 701274 798237 701298 798250
rect 701342 798237 701366 798250
rect 701410 798237 701434 798250
rect 701478 798237 701502 798250
rect 701546 798237 701570 798250
rect 701614 798237 701638 798250
rect 701682 798237 701706 798250
rect 701750 798237 701774 798250
rect 701818 798237 701842 798250
rect 692515 798038 693915 798166
rect 694787 798038 696187 798166
rect 692047 797468 696655 798004
rect 699322 797892 700322 797948
rect 700922 797892 701922 797948
rect 707610 797937 708610 797993
rect 709211 797937 710211 797993
rect 699322 797820 700322 797876
rect 700922 797820 701922 797876
rect 707610 797865 708610 797921
rect 709211 797865 710211 797921
rect 697314 797582 697620 797752
rect 699322 797518 700322 797590
rect 700922 797518 701922 797590
rect 707610 797563 708610 797635
rect 709211 797563 710211 797635
rect 704719 797527 705057 797543
rect 699392 797507 699426 797518
rect 699460 797507 699494 797518
rect 699528 797507 699562 797518
rect 699596 797507 699630 797518
rect 699664 797507 699698 797518
rect 699732 797507 699766 797518
rect 699800 797507 699834 797518
rect 699868 797507 699902 797518
rect 699936 797507 699970 797518
rect 700004 797507 700038 797518
rect 700072 797507 700106 797518
rect 700140 797507 700174 797518
rect 700208 797507 700242 797518
rect 700276 797507 700310 797518
rect 700934 797507 700968 797518
rect 701002 797507 701036 797518
rect 701070 797507 701104 797518
rect 701138 797507 701172 797518
rect 701206 797507 701240 797518
rect 701274 797507 701308 797518
rect 701342 797507 701376 797518
rect 701410 797507 701444 797518
rect 701478 797507 701512 797518
rect 701546 797507 701580 797518
rect 701614 797507 701648 797518
rect 701682 797507 701716 797518
rect 701750 797507 701784 797518
rect 701818 797507 701852 797518
rect 699392 797497 699450 797507
rect 699460 797497 699518 797507
rect 699528 797497 699586 797507
rect 699596 797497 699654 797507
rect 699664 797497 699722 797507
rect 699732 797497 699790 797507
rect 699800 797497 699858 797507
rect 699868 797497 699926 797507
rect 699936 797497 699994 797507
rect 700004 797497 700062 797507
rect 700072 797497 700130 797507
rect 700140 797497 700198 797507
rect 700208 797497 700266 797507
rect 700276 797497 700334 797507
rect 700934 797497 700992 797507
rect 701002 797497 701060 797507
rect 701070 797497 701128 797507
rect 701138 797497 701196 797507
rect 701206 797497 701264 797507
rect 701274 797497 701332 797507
rect 701342 797497 701400 797507
rect 701410 797497 701468 797507
rect 701478 797497 701536 797507
rect 701546 797497 701604 797507
rect 701614 797497 701672 797507
rect 701682 797497 701740 797507
rect 701750 797497 701808 797507
rect 701818 797497 701876 797507
rect 699368 797473 700334 797497
rect 700910 797473 701876 797497
rect 699392 797458 699416 797473
rect 699460 797458 699484 797473
rect 699528 797458 699552 797473
rect 699596 797458 699620 797473
rect 699664 797458 699688 797473
rect 699732 797458 699756 797473
rect 699800 797458 699824 797473
rect 699868 797458 699892 797473
rect 699936 797458 699960 797473
rect 700004 797458 700028 797473
rect 700072 797458 700096 797473
rect 700140 797458 700164 797473
rect 700208 797458 700232 797473
rect 700276 797458 700300 797473
rect 700934 797458 700958 797473
rect 701002 797458 701026 797473
rect 701070 797458 701094 797473
rect 701138 797458 701162 797473
rect 701206 797458 701230 797473
rect 701274 797458 701298 797473
rect 701342 797458 701366 797473
rect 701410 797458 701434 797473
rect 701478 797458 701502 797473
rect 701546 797458 701570 797473
rect 701614 797458 701638 797473
rect 701682 797458 701706 797473
rect 701750 797458 701774 797473
rect 701818 797458 701842 797473
rect 699322 797303 700322 797458
rect 692463 797268 692511 797292
rect 696191 797268 696239 797292
rect 692487 797214 692511 797268
rect 696215 797214 696239 797268
rect 699322 797269 700334 797303
rect 700922 797293 701922 797458
rect 704735 797425 705041 797527
rect 707610 797303 708610 797363
rect 709211 797303 710211 797363
rect 700910 797269 701922 797293
rect 699322 797258 700322 797269
rect 700922 797258 701922 797269
rect 699392 797245 699416 797258
rect 699460 797245 699484 797258
rect 699528 797245 699552 797258
rect 699596 797245 699620 797258
rect 699664 797245 699688 797258
rect 699732 797245 699756 797258
rect 699800 797245 699824 797258
rect 699868 797245 699892 797258
rect 699936 797245 699960 797258
rect 700004 797245 700028 797258
rect 700072 797245 700096 797258
rect 700140 797245 700164 797258
rect 700208 797245 700232 797258
rect 700276 797245 700300 797258
rect 700934 797245 700958 797258
rect 701002 797245 701026 797258
rect 701070 797245 701094 797258
rect 701138 797245 701162 797258
rect 701206 797245 701230 797258
rect 701274 797245 701298 797258
rect 701342 797245 701366 797258
rect 701410 797245 701434 797258
rect 701478 797245 701502 797258
rect 701546 797245 701570 797258
rect 701614 797245 701638 797258
rect 701682 797245 701706 797258
rect 701750 797245 701774 797258
rect 701818 797245 701842 797258
rect 692463 797190 692511 797214
rect 696191 797190 696239 797214
rect 687686 797119 687720 797153
rect 687798 797141 687822 797165
rect 687686 797095 687710 797119
rect 687774 797117 687798 797129
rect 687798 797081 687822 797105
rect 692450 797037 692474 797061
rect 692508 797037 692532 797061
rect 696170 797037 696194 797061
rect 696228 797037 696252 797061
rect 692484 797013 692498 797037
rect 696204 797013 696218 797037
rect 692484 796935 692487 796959
rect 696215 796935 696218 796959
rect 692508 796911 692532 796935
rect 696170 796911 696194 796935
rect 699322 796900 700322 796956
rect 700922 796900 701922 796956
rect 707610 796945 708610 797001
rect 709211 796945 710211 797001
rect 692515 796805 693915 796848
rect 694787 796805 696187 796848
rect 699322 796828 700322 796884
rect 700922 796828 701922 796884
rect 707610 796873 708610 796929
rect 709211 796873 710211 796929
rect 692515 796642 693915 796770
rect 694787 796642 696187 796770
rect 688883 796473 688918 796502
rect 692515 796479 693915 796607
rect 694787 796479 696187 796607
rect 699322 796526 700322 796598
rect 700922 796526 701922 796598
rect 707610 796571 708610 796643
rect 709211 796571 710211 796643
rect 699392 796515 699426 796526
rect 699460 796515 699494 796526
rect 699528 796515 699562 796526
rect 699596 796515 699630 796526
rect 699664 796515 699698 796526
rect 699732 796515 699766 796526
rect 699800 796515 699834 796526
rect 699868 796515 699902 796526
rect 699936 796515 699970 796526
rect 700004 796515 700038 796526
rect 700072 796515 700106 796526
rect 700140 796515 700174 796526
rect 700208 796515 700242 796526
rect 700276 796515 700310 796526
rect 700934 796515 700968 796526
rect 701002 796515 701036 796526
rect 701070 796515 701104 796526
rect 701138 796515 701172 796526
rect 701206 796515 701240 796526
rect 701274 796515 701308 796526
rect 701342 796515 701376 796526
rect 701410 796515 701444 796526
rect 701478 796515 701512 796526
rect 701546 796515 701580 796526
rect 701614 796515 701648 796526
rect 701682 796515 701716 796526
rect 701750 796515 701784 796526
rect 701818 796515 701852 796526
rect 699392 796505 699450 796515
rect 699460 796505 699518 796515
rect 699528 796505 699586 796515
rect 699596 796505 699654 796515
rect 699664 796505 699722 796515
rect 699732 796505 699790 796515
rect 699800 796505 699858 796515
rect 699868 796505 699926 796515
rect 699936 796505 699994 796515
rect 700004 796505 700062 796515
rect 700072 796505 700130 796515
rect 700140 796505 700198 796515
rect 700208 796505 700266 796515
rect 700276 796505 700334 796515
rect 700934 796505 700992 796515
rect 701002 796505 701060 796515
rect 701070 796505 701128 796515
rect 701138 796505 701196 796515
rect 701206 796505 701264 796515
rect 701274 796505 701332 796515
rect 701342 796505 701400 796515
rect 701410 796505 701468 796515
rect 701478 796505 701536 796515
rect 701546 796505 701604 796515
rect 701614 796505 701672 796515
rect 701682 796505 701740 796515
rect 701750 796505 701808 796515
rect 701818 796505 701876 796515
rect 699368 796481 700334 796505
rect 700910 796481 701876 796505
rect 688883 796468 688884 796473
rect 688917 796468 688918 796473
rect 688917 796439 688951 796468
rect 699392 796466 699416 796481
rect 699460 796466 699484 796481
rect 699528 796466 699552 796481
rect 699596 796466 699620 796481
rect 699664 796466 699688 796481
rect 699732 796466 699756 796481
rect 699800 796466 699824 796481
rect 699868 796466 699892 796481
rect 699936 796466 699960 796481
rect 700004 796466 700028 796481
rect 700072 796466 700096 796481
rect 700140 796466 700164 796481
rect 700208 796466 700232 796481
rect 700276 796466 700300 796481
rect 700934 796466 700958 796481
rect 701002 796466 701026 796481
rect 701070 796466 701094 796481
rect 701138 796466 701162 796481
rect 701206 796466 701230 796481
rect 701274 796466 701298 796481
rect 701342 796466 701366 796481
rect 701410 796466 701434 796481
rect 701478 796466 701502 796481
rect 701546 796466 701570 796481
rect 701614 796466 701638 796481
rect 701682 796466 701706 796481
rect 701750 796466 701774 796481
rect 701818 796466 701842 796481
rect 688917 796370 688951 796404
rect 688917 796301 688951 796335
rect 692515 796316 693915 796444
rect 694787 796316 696187 796444
rect 699322 796311 700322 796466
rect 688917 796232 688951 796266
rect 688917 796163 688951 796197
rect 692515 796153 693915 796281
rect 694787 796153 696187 796281
rect 699322 796277 700334 796311
rect 700922 796301 701922 796466
rect 707610 796311 708610 796371
rect 709211 796311 710211 796371
rect 700910 796277 701922 796301
rect 699322 796266 700322 796277
rect 700922 796266 701922 796277
rect 699392 796253 699416 796266
rect 699460 796253 699484 796266
rect 699528 796253 699552 796266
rect 699596 796253 699620 796266
rect 699664 796253 699688 796266
rect 699732 796253 699756 796266
rect 699800 796253 699824 796266
rect 699868 796253 699892 796266
rect 699936 796253 699960 796266
rect 700004 796253 700028 796266
rect 700072 796253 700096 796266
rect 700140 796253 700164 796266
rect 700208 796253 700232 796266
rect 700276 796253 700300 796266
rect 700934 796253 700958 796266
rect 701002 796253 701026 796266
rect 701070 796253 701094 796266
rect 701138 796253 701162 796266
rect 701206 796253 701230 796266
rect 701274 796253 701298 796266
rect 701342 796253 701366 796266
rect 701410 796253 701434 796266
rect 701478 796253 701502 796266
rect 701546 796253 701570 796266
rect 701614 796253 701638 796266
rect 701682 796253 701706 796266
rect 701750 796253 701774 796266
rect 701818 796253 701842 796266
rect 688917 796094 688951 796128
rect 688917 796025 688951 796059
rect 692515 795996 693915 796046
rect 694787 795996 696187 796046
rect 688917 795956 688951 795990
rect 698017 795933 698120 795969
rect 688917 795887 688951 795921
rect 692463 795885 692511 795909
rect 696191 795885 696239 795909
rect 688917 795818 688951 795852
rect 692487 795831 692511 795885
rect 696215 795831 696239 795885
rect 698017 795858 698053 795933
rect 692463 795807 692511 795831
rect 696191 795807 696239 795831
rect 698030 795824 698077 795858
rect 698017 795790 698053 795824
rect 688917 795749 688951 795783
rect 698030 795756 698077 795790
rect 698017 795722 698053 795756
rect 688917 795680 688951 795714
rect 698030 795688 698077 795722
rect 698017 795654 698053 795688
rect 688917 795611 688951 795645
rect 692463 795629 692521 795653
rect 696191 795629 696249 795653
rect 692487 795619 692521 795629
rect 696215 795619 696249 795629
rect 698030 795620 698077 795654
rect 698017 795586 698053 795620
rect 686879 795544 687585 795554
rect 686882 795528 687585 795544
rect 688917 795542 688951 795576
rect 692487 795547 692521 795581
rect 696215 795547 696249 795581
rect 678680 795433 678704 795467
rect 681345 795399 682345 795455
rect 678680 795365 678704 795399
rect 684004 795349 685004 795477
rect 688917 795473 688951 795507
rect 692487 795475 692521 795509
rect 696215 795475 696249 795509
rect 688917 795404 688951 795438
rect 692487 795427 692521 795437
rect 696215 795427 696249 795437
rect 692463 795403 692521 795427
rect 696191 795403 696249 795427
rect 688917 795335 688951 795369
rect 678680 795297 678704 795331
rect 678680 795229 678704 795263
rect 679133 795255 679283 795267
rect 679452 795255 679602 795267
rect 681345 795229 682345 795279
rect 678680 795161 678704 795195
rect 684004 795193 685004 795321
rect 688917 795266 688951 795300
rect 679002 795142 679602 795192
rect 678680 795093 678704 795127
rect 681441 795064 681457 795130
rect 682225 795064 682241 795130
rect 678680 795025 678704 795059
rect 684004 795037 685004 795165
rect 685537 795161 686137 795211
rect 688917 795197 688951 795231
rect 692463 795214 692521 795248
rect 696191 795214 696249 795248
rect 688917 795128 688951 795162
rect 678680 794957 678704 794991
rect 679002 794966 679602 795022
rect 678680 794889 678704 794923
rect 681441 794902 681457 794968
rect 683625 794902 683641 794968
rect 684004 794881 685004 795009
rect 685537 795005 686137 795061
rect 688917 795059 688951 795093
rect 692515 795084 693915 795127
rect 694787 795084 696187 795127
rect 688917 794990 688951 795024
rect 688917 794921 688951 794955
rect 692515 794921 693915 795049
rect 694787 794921 696187 795049
rect 685537 794855 686137 794905
rect 678680 794821 678704 794855
rect 679002 794796 679602 794846
rect 678680 794753 678704 794787
rect 680502 794761 680517 794776
rect 678680 794685 678704 794719
rect 678680 794617 678704 794651
rect 678680 794549 678704 794583
rect 680480 794581 680517 794761
rect 680502 794566 680517 794581
rect 680615 794761 680630 794776
rect 680803 794772 680815 794776
rect 680800 794761 680815 794772
rect 680615 794581 680815 794761
rect 681441 794740 681457 794806
rect 683625 794740 683641 794806
rect 684004 794725 685004 794853
rect 688917 794852 688951 794886
rect 688917 794783 688951 794817
rect 692515 794758 693915 794886
rect 694787 794758 696187 794886
rect 688917 794714 688951 794748
rect 686829 794649 687429 794699
rect 688917 794645 688951 794679
rect 680615 794566 680630 794581
rect 680800 794570 680815 794581
rect 681441 794578 681457 794644
rect 682225 794578 682241 794644
rect 684004 794575 685004 794625
rect 688917 794576 688951 794610
rect 692515 794595 693915 794723
rect 694787 794595 696187 794723
rect 680803 794566 680815 794570
rect 680615 794525 680630 794540
rect 680803 794536 680815 794540
rect 680800 794525 680815 794536
rect 678680 794481 678704 794515
rect 678680 794413 678704 794447
rect 678680 794345 678704 794379
rect 679007 794370 679607 794420
rect 680615 794345 680815 794525
rect 681345 794429 682345 794479
rect 686829 794473 687429 794529
rect 688917 794507 688951 794541
rect 688917 794438 688951 794472
rect 692515 794432 693915 794560
rect 694787 794432 696187 794560
rect 684054 794373 685054 794423
rect 688917 794393 688951 794403
rect 688893 794369 688951 794393
rect 680615 794330 680630 794345
rect 680800 794334 680815 794345
rect 680803 794330 680815 794334
rect 678680 794277 678704 794311
rect 681345 794253 682345 794309
rect 678680 794209 678704 794243
rect 679007 794200 679607 794250
rect 684054 794217 685054 794345
rect 686829 794303 687429 794353
rect 692515 794269 693915 794397
rect 694787 794269 696187 794397
rect 678680 794141 678704 794175
rect 678680 794073 678704 794107
rect 681345 794077 682345 794205
rect 678680 794005 678704 794039
rect 680215 794024 680815 794074
rect 684054 794061 685054 794189
rect 685793 794182 685805 794186
rect 685793 794171 685808 794182
rect 685978 794171 685993 794186
rect 678680 793937 678704 793971
rect 678680 793869 678704 793903
rect 680215 793848 680815 793904
rect 681345 793901 682345 794029
rect 684054 793905 685054 794033
rect 685793 793991 685993 794171
rect 685793 793980 685808 793991
rect 685793 793976 685805 793980
rect 685978 793976 685993 793991
rect 686053 794182 686065 794186
rect 686053 794171 686068 794182
rect 686238 794171 686253 794186
rect 686053 793991 686253 794171
rect 686607 794164 687607 794214
rect 697088 794171 697138 795571
rect 697238 794171 697366 795571
rect 697394 794171 697522 795571
rect 697550 794171 697678 795571
rect 697706 794171 697756 795571
rect 698030 795552 698077 795586
rect 698017 795518 698053 795552
rect 698030 795484 698077 795518
rect 698017 795450 698053 795484
rect 698030 795416 698077 795450
rect 698017 795382 698053 795416
rect 698030 795348 698077 795382
rect 698017 795314 698053 795348
rect 698030 795280 698077 795314
rect 698017 795246 698053 795280
rect 698030 795212 698077 795246
rect 698017 795178 698053 795212
rect 698030 795144 698077 795178
rect 698017 795110 698053 795144
rect 698030 795076 698077 795110
rect 698017 795042 698053 795076
rect 698030 795008 698077 795042
rect 698017 794974 698053 795008
rect 698030 794940 698077 794974
rect 698017 794906 698053 794940
rect 698030 794872 698077 794906
rect 698017 794838 698053 794872
rect 698030 794804 698077 794838
rect 698017 794770 698053 794804
rect 698030 794736 698077 794770
rect 698017 794702 698053 794736
rect 698030 794668 698077 794702
rect 698017 794634 698053 794668
rect 698030 794600 698077 794634
rect 698017 794566 698053 794600
rect 698030 794532 698077 794566
rect 698017 794498 698053 794532
rect 698030 794464 698077 794498
rect 698017 794430 698053 794464
rect 698030 794396 698077 794430
rect 698017 794362 698053 794396
rect 698030 794328 698077 794362
rect 698017 794294 698053 794328
rect 698030 794260 698077 794294
rect 698017 794226 698053 794260
rect 698030 794192 698077 794226
rect 692515 794119 693915 794162
rect 694787 794119 696187 794162
rect 698017 794158 698053 794192
rect 698030 794124 698077 794158
rect 698017 794090 698053 794124
rect 686607 794014 687607 794064
rect 698030 794056 698077 794090
rect 686053 793980 686068 793991
rect 686053 793976 686065 793980
rect 686238 793976 686253 793991
rect 685793 793946 685805 793950
rect 685793 793935 685808 793946
rect 685978 793935 685993 793950
rect 678680 793801 678704 793835
rect 678680 793733 678704 793767
rect 681345 793731 682345 793781
rect 684054 793749 685054 793877
rect 685793 793755 685993 793935
rect 685793 793744 685808 793755
rect 685793 793740 685805 793744
rect 685978 793740 685993 793755
rect 686053 793946 686065 793950
rect 686053 793935 686068 793946
rect 686238 793935 686253 793950
rect 686053 793755 686253 793935
rect 686607 793855 687607 793905
rect 692463 793809 692511 793833
rect 696191 793809 696239 793833
rect 686053 793744 686068 793755
rect 686053 793740 686065 793744
rect 686238 793740 686253 793755
rect 678680 793665 678704 793699
rect 680215 793672 680815 793728
rect 681345 793662 682345 793674
rect 678680 793597 678704 793631
rect 684054 793593 685054 793721
rect 686607 793705 687607 793755
rect 692487 793731 692511 793809
rect 696215 793755 696239 793809
rect 696191 793731 696239 793755
rect 696617 793772 696651 793773
rect 696617 793749 696626 793772
rect 696617 793731 696675 793749
rect 696651 793715 696675 793731
rect 696651 793647 696675 793681
rect 685533 793586 685545 793590
rect 685533 793575 685548 793586
rect 685718 793575 685733 793590
rect 678680 793529 678704 793563
rect 680215 793502 680815 793552
rect 678680 793461 678704 793495
rect 678680 793393 678704 793427
rect 680215 793370 680815 793420
rect 681466 793411 682466 793461
rect 684054 793437 685054 793565
rect 678680 793325 678704 793359
rect 678680 793257 678704 793291
rect 681466 793255 682466 793383
rect 682890 793339 683490 793389
rect 678680 793189 678704 793223
rect 680215 793194 680815 793250
rect 682890 793183 683490 793311
rect 684054 793281 685054 793409
rect 685533 793395 685733 793575
rect 685533 793384 685548 793395
rect 685533 793380 685545 793384
rect 685718 793380 685733 793395
rect 685793 793586 685805 793590
rect 685793 793575 685808 793586
rect 685978 793575 685993 793590
rect 685793 793395 685993 793575
rect 685793 793384 685808 793395
rect 685793 793380 685805 793384
rect 685978 793380 685993 793395
rect 686053 793586 686065 793590
rect 686053 793575 686068 793586
rect 686238 793575 686253 793590
rect 686053 793395 686253 793575
rect 686053 793384 686068 793395
rect 686053 793380 686065 793384
rect 686238 793380 686253 793395
rect 686313 793586 686325 793590
rect 686313 793575 686328 793586
rect 686498 793575 686513 793590
rect 686313 793395 686513 793575
rect 686313 793384 686328 793395
rect 686313 793380 686325 793384
rect 686498 793380 686513 793395
rect 686627 793586 686639 793590
rect 686627 793575 686642 793586
rect 686812 793575 686827 793590
rect 686627 793395 686827 793575
rect 686627 793384 686642 793395
rect 686627 793380 686639 793384
rect 686812 793380 686827 793395
rect 686887 793586 686899 793590
rect 686887 793575 686902 793586
rect 687072 793575 687087 793590
rect 686887 793395 687087 793575
rect 686887 793384 686902 793395
rect 686887 793380 686899 793384
rect 687072 793380 687087 793395
rect 687147 793586 687159 793590
rect 687147 793575 687162 793586
rect 687332 793575 687347 793590
rect 696651 793579 696675 793613
rect 687147 793395 687347 793575
rect 696651 793511 696675 793545
rect 696651 793443 696675 793477
rect 687147 793384 687162 793395
rect 687147 793380 687159 793384
rect 687332 793380 687347 793395
rect 696651 793375 696675 793409
rect 696651 793307 696675 793341
rect 685718 793215 685733 793230
rect 685679 793185 685733 793215
rect 678680 793121 678704 793155
rect 681466 793105 682466 793155
rect 684054 793131 685054 793181
rect 685718 793170 685733 793185
rect 685793 793226 685805 793230
rect 685793 793215 685808 793226
rect 685978 793215 685993 793230
rect 685793 793185 685993 793215
rect 685793 793174 685808 793185
rect 685793 793170 685805 793174
rect 685978 793170 685993 793185
rect 686053 793226 686065 793230
rect 686053 793215 686068 793226
rect 686238 793215 686253 793230
rect 686812 793215 686827 793230
rect 686053 793185 686253 793215
rect 686807 793185 686827 793215
rect 686053 793174 686068 793185
rect 686053 793170 686065 793174
rect 686238 793170 686253 793185
rect 686812 793170 686827 793185
rect 686887 793226 686899 793230
rect 686887 793215 686902 793226
rect 687072 793215 687087 793230
rect 686887 793185 687087 793215
rect 686887 793174 686902 793185
rect 686887 793170 686899 793174
rect 687072 793170 687087 793185
rect 687147 793226 687159 793230
rect 687147 793215 687162 793226
rect 687332 793215 687347 793230
rect 687147 793185 687347 793215
rect 687147 793174 687162 793185
rect 687147 793170 687159 793174
rect 687332 793170 687347 793185
rect 685718 793129 685733 793144
rect 681794 793102 682466 793105
rect 685679 793099 685733 793129
rect 678680 793053 678704 793087
rect 685718 793084 685733 793099
rect 685793 793140 685805 793144
rect 685793 793129 685808 793140
rect 685978 793129 685993 793144
rect 685793 793099 685993 793129
rect 685793 793088 685808 793099
rect 685793 793084 685805 793088
rect 685978 793084 685993 793099
rect 686053 793140 686065 793144
rect 686053 793129 686068 793140
rect 686238 793129 686253 793144
rect 686812 793129 686827 793144
rect 686053 793099 686253 793129
rect 686807 793099 686827 793129
rect 686053 793088 686068 793099
rect 686053 793084 686065 793088
rect 686238 793084 686253 793099
rect 686812 793084 686827 793099
rect 686887 793140 686899 793144
rect 686887 793129 686902 793140
rect 687072 793129 687087 793144
rect 686887 793099 687087 793129
rect 686887 793088 686902 793099
rect 686887 793084 686899 793088
rect 687072 793084 687087 793099
rect 687147 793140 687159 793144
rect 687147 793129 687162 793140
rect 687332 793129 687347 793144
rect 687147 793099 687347 793129
rect 687147 793088 687162 793099
rect 687147 793084 687159 793088
rect 687332 793084 687347 793099
rect 678680 792985 678704 793019
rect 680215 793018 680815 793074
rect 682890 793027 683490 793083
rect 678680 792917 678704 792951
rect 678680 792849 678704 792883
rect 680215 792848 680815 792898
rect 678680 792781 678704 792815
rect 678680 792713 678704 792747
rect 678680 792645 678704 792679
rect 679007 792672 679607 792722
rect 678680 792577 678704 792611
rect 680615 792577 680630 792592
rect 680803 792588 680815 792592
rect 680800 792577 680815 792588
rect 678680 792509 678704 792543
rect 679007 792502 679607 792552
rect 678680 792441 678704 792475
rect 678680 792373 678704 792407
rect 680615 792397 680815 792577
rect 681502 792505 681529 792995
rect 681866 792896 682466 793024
rect 682890 792871 683490 792999
rect 684004 792929 685004 792979
rect 685539 792940 685777 792972
rect 685803 792920 686119 792938
rect 681866 792740 682466 792868
rect 684004 792773 685004 792901
rect 682890 792721 683490 792771
rect 681866 792584 682466 792712
rect 682890 792605 683490 792655
rect 684004 792617 685004 792745
rect 681866 792434 682466 792484
rect 682890 792449 683490 792505
rect 684004 792461 685004 792589
rect 692427 792522 693027 792572
rect 680615 792382 680630 792397
rect 680800 792386 680815 792397
rect 680803 792382 680815 792386
rect 680502 792341 680517 792356
rect 678680 792305 678704 792339
rect 678680 792237 678704 792271
rect 678680 792169 678704 792203
rect 680480 792161 680517 792341
rect 680502 792146 680517 792161
rect 680615 792341 680630 792356
rect 680803 792352 680815 792356
rect 680800 792341 680815 792352
rect 680615 792161 680815 792341
rect 681866 792318 682466 792368
rect 682890 792293 683490 792349
rect 684004 792305 685004 792433
rect 692427 792366 693027 792494
rect 693888 792375 694194 792545
rect 694388 792375 694694 792545
rect 689309 792278 689909 792328
rect 681866 792168 682466 792218
rect 682041 792165 682385 792168
rect 680615 792146 680630 792161
rect 680800 792150 680815 792161
rect 680803 792146 680815 792150
rect 682890 792137 683490 792193
rect 684004 792149 685004 792277
rect 678680 792101 678704 792135
rect 679002 792076 679602 792126
rect 689309 792122 689909 792250
rect 692427 792210 693027 792338
rect 678680 792033 678704 792067
rect 678680 791965 678704 791999
rect 682890 791981 683490 792109
rect 684004 791993 685004 792121
rect 689309 791966 689909 792094
rect 692427 792054 693027 792110
rect 678680 791897 678704 791931
rect 679002 791900 679602 791956
rect 678680 791829 678704 791863
rect 682890 791825 683490 791953
rect 684004 791837 685004 791965
rect 692427 791898 693027 792026
rect 689309 791810 689909 791866
rect 678680 791761 678704 791795
rect 679002 791730 679602 791780
rect 679061 791727 679355 791730
rect 679380 791727 679602 791730
rect 678680 791693 678704 791727
rect 682890 791669 683490 791797
rect 684004 791687 685004 791737
rect 685803 791720 686119 791732
rect 685539 791716 686119 791720
rect 685513 791682 685537 791716
rect 685539 791682 685777 791716
rect 678680 791625 678704 791659
rect 689309 791654 689909 791782
rect 690910 791754 691110 791765
rect 692427 791742 693027 791870
rect 690910 791640 691110 791690
rect 678680 791557 678704 791591
rect 678680 791489 678704 791523
rect 682890 791513 683490 791569
rect 685718 791555 685733 791570
rect 684004 791485 685004 791535
rect 685679 791525 685733 791555
rect 685718 791510 685733 791525
rect 685793 791566 685805 791570
rect 685793 791555 685808 791566
rect 685978 791555 685993 791570
rect 685793 791525 685993 791555
rect 685793 791514 685808 791525
rect 685793 791510 685805 791514
rect 685978 791510 685993 791525
rect 686053 791566 686065 791570
rect 686053 791555 686068 791566
rect 686238 791555 686253 791570
rect 686812 791555 686827 791570
rect 686053 791525 686253 791555
rect 686807 791525 686827 791555
rect 686053 791514 686068 791525
rect 686053 791510 686065 791514
rect 686238 791510 686253 791525
rect 686812 791510 686827 791525
rect 686887 791566 686899 791570
rect 686887 791555 686902 791566
rect 687072 791555 687087 791570
rect 686887 791525 687087 791555
rect 686887 791514 686902 791525
rect 686887 791510 686899 791514
rect 687072 791510 687087 791525
rect 687147 791566 687159 791570
rect 687147 791555 687162 791566
rect 687332 791555 687347 791570
rect 687147 791525 687347 791555
rect 687147 791514 687162 791525
rect 687147 791510 687159 791514
rect 687332 791510 687347 791525
rect 689309 791498 689909 791626
rect 692427 791592 693027 791642
rect 693888 791575 694194 791745
rect 694388 791575 694694 791745
rect 678680 791421 678704 791455
rect 678680 791353 678704 791387
rect 682890 791357 683490 791485
rect 690910 791484 691110 791540
rect 685718 791469 685733 791484
rect 684004 791329 685004 791457
rect 685679 791439 685733 791469
rect 685718 791424 685733 791439
rect 685793 791480 685805 791484
rect 685793 791469 685808 791480
rect 685978 791469 685993 791484
rect 685793 791439 685993 791469
rect 685793 791428 685808 791439
rect 685793 791424 685805 791428
rect 685978 791424 685993 791439
rect 686053 791480 686065 791484
rect 686053 791469 686068 791480
rect 686238 791469 686253 791484
rect 686812 791469 686827 791484
rect 686053 791439 686253 791469
rect 686807 791439 686827 791469
rect 686053 791428 686068 791439
rect 686053 791424 686065 791428
rect 686238 791424 686253 791439
rect 686812 791424 686827 791439
rect 686887 791480 686899 791484
rect 686887 791469 686902 791480
rect 687072 791469 687087 791484
rect 686887 791439 687087 791469
rect 686887 791428 686902 791439
rect 686887 791424 686899 791428
rect 687072 791424 687087 791439
rect 687147 791480 687159 791484
rect 687147 791469 687162 791480
rect 687332 791469 687347 791484
rect 687147 791439 687347 791469
rect 692427 791462 693027 791512
rect 687147 791428 687162 791439
rect 687147 791424 687159 791428
rect 687332 791424 687347 791439
rect 689309 791348 689909 791398
rect 690910 791334 691110 791384
rect 678680 791285 678704 791319
rect 678680 791217 678704 791251
rect 682890 791201 683490 791329
rect 692427 791312 693027 791362
rect 678680 791149 678704 791183
rect 684004 791173 685004 791301
rect 685533 791270 685545 791274
rect 685533 791259 685548 791270
rect 685718 791259 685733 791274
rect 678680 791081 678704 791115
rect 679133 791101 679283 791113
rect 679452 791101 679602 791113
rect 678680 791013 678704 791047
rect 682890 791045 683490 791173
rect 679002 790988 679602 791038
rect 684004 791017 685004 791145
rect 685533 791079 685733 791259
rect 685533 791068 685548 791079
rect 685533 791064 685545 791068
rect 685718 791064 685733 791079
rect 685793 791270 685805 791274
rect 685793 791259 685808 791270
rect 685978 791259 685993 791274
rect 685793 791079 685993 791259
rect 685793 791068 685808 791079
rect 685793 791064 685805 791068
rect 685978 791064 685993 791079
rect 686053 791270 686065 791274
rect 686053 791259 686068 791270
rect 686238 791259 686253 791274
rect 686053 791079 686253 791259
rect 686053 791068 686068 791079
rect 686053 791064 686065 791068
rect 686238 791064 686253 791079
rect 686313 791270 686325 791274
rect 686313 791259 686328 791270
rect 686498 791259 686513 791274
rect 686313 791079 686513 791259
rect 686313 791068 686328 791079
rect 686313 791064 686325 791068
rect 686498 791064 686513 791079
rect 686627 791270 686639 791274
rect 686627 791259 686642 791270
rect 686812 791259 686827 791274
rect 686627 791079 686827 791259
rect 686627 791068 686642 791079
rect 686627 791064 686639 791068
rect 686812 791064 686827 791079
rect 686887 791270 686899 791274
rect 686887 791259 686902 791270
rect 687072 791259 687087 791274
rect 686887 791079 687087 791259
rect 686887 791068 686902 791079
rect 686887 791064 686899 791068
rect 687072 791064 687087 791079
rect 687147 791270 687159 791274
rect 687147 791259 687162 791270
rect 687332 791259 687347 791274
rect 687147 791079 687347 791259
rect 689309 791218 689909 791268
rect 692427 791140 693027 791190
rect 687147 791068 687162 791079
rect 687147 791064 687159 791068
rect 687332 791064 687347 791079
rect 689309 791068 689909 791118
rect 692427 790990 693027 791040
rect 678680 790945 678704 790979
rect 678680 790877 678704 790911
rect 682890 790895 683490 790945
rect 678680 790809 678704 790843
rect 679002 790812 679602 790868
rect 684004 790861 685004 790917
rect 685793 790910 685805 790914
rect 685793 790899 685808 790910
rect 685978 790899 685993 790914
rect 682890 790779 683490 790829
rect 678680 790741 678704 790775
rect 678680 790673 678704 790707
rect 679002 790642 679602 790692
rect 678680 790605 678704 790639
rect 682890 790623 683490 790751
rect 684004 790705 685004 790833
rect 685793 790719 685993 790899
rect 685793 790708 685808 790719
rect 685793 790704 685805 790708
rect 685978 790704 685993 790719
rect 686053 790910 686065 790914
rect 686053 790899 686068 790910
rect 686238 790899 686253 790914
rect 686607 790899 687607 790949
rect 690910 790934 691110 790984
rect 686053 790719 686253 790899
rect 692427 790860 693027 790910
rect 686607 790749 687607 790799
rect 690910 790778 691110 790834
rect 686053 790708 686068 790719
rect 686053 790704 686065 790708
rect 686238 790704 686253 790719
rect 692427 790704 693027 790832
rect 693888 790775 694194 790945
rect 694388 790775 694694 790945
rect 680502 790607 680517 790622
rect 678680 790537 678704 790571
rect 678680 790469 678704 790503
rect 678680 790401 678704 790435
rect 680480 790427 680517 790607
rect 680502 790412 680517 790427
rect 680615 790607 680630 790622
rect 680803 790618 680815 790622
rect 680800 790607 680815 790618
rect 680615 790427 680815 790607
rect 682890 790467 683490 790595
rect 684004 790549 685004 790677
rect 685793 790674 685805 790678
rect 685793 790663 685808 790674
rect 685978 790663 685993 790678
rect 680615 790412 680630 790427
rect 680800 790416 680815 790427
rect 680803 790412 680815 790416
rect 680615 790371 680630 790386
rect 680803 790382 680815 790386
rect 680800 790371 680815 790382
rect 678680 790333 678704 790367
rect 678680 790265 678704 790299
rect 678680 790197 678704 790231
rect 679007 790216 679607 790266
rect 680615 790191 680815 790371
rect 682890 790311 683490 790439
rect 684004 790393 685004 790521
rect 685793 790483 685993 790663
rect 685793 790472 685808 790483
rect 685793 790468 685805 790472
rect 685978 790468 685993 790483
rect 686053 790674 686065 790678
rect 686053 790663 686068 790674
rect 686238 790663 686253 790678
rect 686053 790483 686253 790663
rect 686607 790590 687607 790640
rect 690910 790628 691110 790678
rect 692427 790548 693027 790676
rect 686053 790472 686068 790483
rect 686053 790468 686065 790472
rect 686238 790468 686253 790483
rect 686607 790440 687607 790490
rect 692427 790392 693027 790448
rect 686829 790301 687429 790351
rect 684004 790243 685004 790293
rect 692427 790236 693027 790364
rect 695201 790282 695251 793282
rect 695351 790282 695479 793282
rect 695507 790282 695635 793282
rect 695663 790282 695791 793282
rect 695819 790282 695947 793282
rect 695975 790282 696103 793282
rect 696131 790282 696259 793282
rect 696287 790282 696337 793282
rect 696651 793239 696675 793273
rect 696651 793171 696675 793205
rect 696651 793103 696675 793137
rect 696651 793035 696675 793069
rect 696651 792967 696675 793001
rect 696651 792899 696675 792933
rect 696651 792831 696675 792865
rect 696651 792763 696675 792797
rect 696651 792695 696675 792729
rect 696651 792627 696675 792661
rect 697088 792641 697138 794041
rect 697238 792641 697366 794041
rect 697394 792641 697522 794041
rect 697550 792641 697678 794041
rect 697706 792641 697756 794041
rect 698017 794022 698053 794056
rect 698030 793988 698077 794022
rect 698017 793954 698053 793988
rect 698030 793920 698077 793954
rect 698017 793886 698053 793920
rect 698030 793852 698077 793886
rect 698017 793818 698053 793852
rect 698030 793784 698077 793818
rect 698017 793750 698053 793784
rect 698030 793716 698077 793750
rect 698017 793682 698053 793716
rect 698030 793648 698077 793682
rect 698017 793614 698053 793648
rect 698030 793580 698077 793614
rect 698017 793546 698053 793580
rect 698030 793512 698077 793546
rect 698017 793478 698053 793512
rect 698030 793444 698077 793478
rect 698017 793410 698053 793444
rect 698030 793376 698077 793410
rect 698017 793342 698053 793376
rect 698030 793308 698077 793342
rect 698017 793274 698053 793308
rect 698030 793240 698077 793274
rect 698017 793206 698053 793240
rect 698030 793172 698077 793206
rect 698017 793138 698053 793172
rect 698030 793104 698077 793138
rect 698017 793070 698053 793104
rect 698030 793036 698077 793070
rect 698017 793002 698053 793036
rect 698030 792968 698077 793002
rect 698017 792934 698053 792968
rect 698030 792900 698077 792934
rect 698017 792866 698053 792900
rect 698030 792832 698077 792866
rect 698017 792798 698053 792832
rect 698030 792764 698077 792798
rect 698017 792730 698053 792764
rect 698030 792696 698077 792730
rect 698017 792662 698053 792696
rect 698030 792628 698077 792662
rect 698017 792594 698053 792628
rect 696651 792559 696675 792593
rect 698030 792560 698077 792594
rect 698017 792526 698053 792560
rect 696651 792491 696675 792525
rect 698030 792492 698077 792526
rect 696651 792423 696675 792457
rect 698017 792428 698053 792492
rect 698030 792394 698077 792428
rect 696651 792355 696675 792389
rect 698017 792360 698053 792394
rect 698030 792326 698077 792360
rect 696651 792287 696675 792321
rect 698017 792292 698053 792326
rect 696651 792219 696675 792253
rect 696651 792151 696675 792185
rect 696651 792083 696675 792117
rect 696651 792015 696675 792049
rect 696651 791947 696675 791981
rect 696651 791879 696675 791913
rect 696651 791811 696675 791845
rect 696651 791743 696675 791777
rect 696651 791675 696675 791709
rect 696651 791607 696675 791641
rect 696651 791539 696675 791573
rect 696651 791471 696675 791505
rect 696651 791403 696675 791437
rect 696651 791335 696675 791369
rect 696651 791267 696675 791301
rect 696651 791199 696675 791233
rect 696651 791131 696675 791165
rect 696651 791063 696675 791097
rect 696651 790995 696675 791029
rect 696651 790927 696675 790961
rect 696651 790859 696675 790893
rect 697088 790879 697138 792279
rect 697238 790879 697366 792279
rect 697394 790879 697522 792279
rect 697550 790879 697678 792279
rect 697706 790879 697756 792279
rect 698030 792258 698077 792292
rect 698017 792224 698053 792258
rect 698030 792190 698077 792224
rect 698017 792156 698053 792190
rect 698030 792122 698077 792156
rect 698017 792088 698053 792122
rect 698030 792054 698077 792088
rect 698017 792020 698053 792054
rect 698030 791986 698077 792020
rect 698017 791952 698053 791986
rect 698030 791918 698077 791952
rect 698017 791884 698053 791918
rect 698030 791850 698077 791884
rect 698017 791816 698053 791850
rect 698030 791782 698077 791816
rect 698017 791748 698053 791782
rect 698030 791714 698077 791748
rect 698017 791680 698053 791714
rect 698030 791646 698077 791680
rect 698017 791612 698053 791646
rect 698030 791578 698077 791612
rect 698017 791544 698053 791578
rect 698030 791510 698077 791544
rect 698017 791476 698053 791510
rect 698030 791442 698077 791476
rect 698017 791408 698053 791442
rect 698030 791374 698077 791408
rect 698017 791340 698053 791374
rect 698030 791306 698077 791340
rect 698017 791272 698053 791306
rect 698030 791238 698077 791272
rect 698017 791204 698053 791238
rect 698030 791170 698077 791204
rect 698017 791136 698053 791170
rect 698030 791102 698077 791136
rect 698017 791068 698053 791102
rect 698030 791034 698077 791068
rect 698017 791000 698053 791034
rect 698030 790966 698077 791000
rect 698017 790932 698053 790966
rect 698030 790898 698077 790932
rect 698017 790864 698053 790898
rect 698030 790830 698077 790864
rect 696651 790791 696675 790825
rect 698017 790796 698053 790830
rect 698030 790762 698077 790796
rect 696651 790723 696675 790757
rect 696651 790655 696675 790689
rect 696651 790587 696675 790621
rect 696651 790519 696675 790553
rect 696651 790451 696675 790485
rect 696651 790383 696675 790417
rect 696651 790315 696675 790349
rect 696651 790247 696675 790281
rect 680615 790176 680630 790191
rect 680800 790180 680815 790191
rect 680803 790176 680815 790180
rect 678680 790129 678704 790163
rect 682890 790161 683490 790211
rect 684004 790127 685004 790177
rect 686829 790125 687429 790181
rect 678680 790061 678704 790095
rect 679007 790046 679607 790096
rect 692427 790080 693027 790208
rect 696651 790179 696675 790213
rect 696651 790111 696675 790145
rect 696651 790043 696675 790077
rect 678680 789993 678704 790027
rect 681664 790002 681812 790006
rect 681641 789994 681812 790002
rect 682113 789994 682313 790006
rect 684004 789971 685004 790027
rect 678680 789925 678704 789959
rect 686829 789955 687429 790005
rect 678680 789857 678704 789891
rect 680215 789870 680815 789920
rect 681713 789881 682313 789931
rect 682921 789899 683521 789949
rect 692427 789930 693027 789980
rect 696651 789975 696675 790009
rect 696651 789907 696675 789941
rect 678680 789789 678704 789823
rect 684004 789821 685004 789871
rect 678680 789721 678704 789755
rect 680215 789694 680815 789750
rect 681713 789705 682313 789761
rect 682921 789743 683521 789799
rect 685537 789749 686137 789799
rect 697088 789749 697138 790749
rect 697238 789749 697366 790749
rect 697394 789749 697522 790749
rect 697550 789749 697678 790749
rect 697706 789749 697756 790749
rect 698017 790728 698053 790762
rect 698030 790694 698077 790728
rect 698017 790660 698053 790694
rect 698030 790626 698077 790660
rect 698017 790592 698053 790626
rect 698030 790558 698077 790592
rect 698017 790524 698053 790558
rect 698030 790490 698077 790524
rect 698017 790456 698053 790490
rect 698030 790422 698077 790456
rect 698017 790388 698053 790422
rect 698030 790354 698077 790388
rect 698017 790320 698053 790354
rect 698030 790286 698077 790320
rect 698017 790252 698053 790286
rect 698030 790218 698077 790252
rect 698017 790184 698053 790218
rect 698030 790150 698077 790184
rect 698017 790116 698053 790150
rect 698030 790082 698077 790116
rect 698017 790048 698053 790082
rect 698030 790014 698077 790048
rect 698017 789980 698053 790014
rect 698030 789946 698077 789980
rect 698017 789912 698053 789946
rect 698030 789878 698077 789912
rect 698017 789844 698053 789878
rect 698030 789810 698077 789844
rect 698017 789776 698053 789810
rect 698030 789742 698077 789776
rect 698017 789708 698053 789742
rect 678680 789653 678704 789687
rect 698030 789674 698077 789708
rect 678680 789585 678704 789619
rect 680215 789518 680815 789574
rect 681713 789529 682313 789657
rect 682921 789593 683521 789643
rect 684070 789599 684670 789649
rect 685537 789593 686137 789649
rect 698017 789640 698053 789674
rect 698030 789606 698077 789640
rect 698017 789572 698053 789606
rect 698030 789538 698077 789572
rect 698017 789504 698053 789538
rect 684070 789443 684670 789499
rect 685537 789443 686137 789493
rect 692428 789442 693028 789492
rect 698030 789470 698077 789504
rect 698017 789436 698053 789470
rect 680215 789348 680815 789398
rect 681713 789359 682313 789409
rect 698030 789402 698077 789436
rect 698017 789368 698053 789402
rect 684070 789293 684670 789343
rect 692428 789292 693028 789342
rect 698030 789334 698077 789368
rect 698017 789300 698053 789334
rect 680215 789232 680815 789282
rect 698030 789266 698077 789300
rect 698017 789232 698053 789266
rect 692428 789162 693028 789212
rect 698030 789198 698077 789232
rect 698017 789164 698053 789198
rect 680215 789056 680815 789112
rect 692428 789006 693028 789134
rect 698030 789130 698077 789164
rect 698017 789096 698053 789130
rect 698030 789062 698077 789096
rect 698017 788983 698053 789062
rect 698084 788983 698120 795933
rect 699322 795908 700322 795964
rect 700922 795908 701922 795964
rect 707610 795953 708610 796009
rect 709211 795953 710211 796009
rect 699322 795836 700322 795892
rect 700922 795836 701922 795892
rect 707610 795881 708610 795937
rect 709211 795881 710211 795937
rect 699322 795534 700322 795606
rect 700922 795534 701922 795606
rect 707610 795579 708610 795651
rect 709211 795579 710211 795651
rect 699392 795523 699426 795534
rect 699460 795523 699494 795534
rect 699528 795523 699562 795534
rect 699596 795523 699630 795534
rect 699664 795523 699698 795534
rect 699732 795523 699766 795534
rect 699800 795523 699834 795534
rect 699868 795523 699902 795534
rect 699936 795523 699970 795534
rect 700004 795523 700038 795534
rect 700072 795523 700106 795534
rect 700140 795523 700174 795534
rect 700208 795523 700242 795534
rect 700276 795523 700310 795534
rect 700934 795523 700968 795534
rect 701002 795523 701036 795534
rect 701070 795523 701104 795534
rect 701138 795523 701172 795534
rect 701206 795523 701240 795534
rect 701274 795523 701308 795534
rect 701342 795523 701376 795534
rect 701410 795523 701444 795534
rect 701478 795523 701512 795534
rect 701546 795523 701580 795534
rect 701614 795523 701648 795534
rect 701682 795523 701716 795534
rect 701750 795523 701784 795534
rect 701818 795523 701852 795534
rect 699392 795513 699450 795523
rect 699460 795513 699518 795523
rect 699528 795513 699586 795523
rect 699596 795513 699654 795523
rect 699664 795513 699722 795523
rect 699732 795513 699790 795523
rect 699800 795513 699858 795523
rect 699868 795513 699926 795523
rect 699936 795513 699994 795523
rect 700004 795513 700062 795523
rect 700072 795513 700130 795523
rect 700140 795513 700198 795523
rect 700208 795513 700266 795523
rect 700276 795513 700334 795523
rect 700934 795513 700992 795523
rect 701002 795513 701060 795523
rect 701070 795513 701128 795523
rect 701138 795513 701196 795523
rect 701206 795513 701264 795523
rect 701274 795513 701332 795523
rect 701342 795513 701400 795523
rect 701410 795513 701468 795523
rect 701478 795513 701536 795523
rect 701546 795513 701604 795523
rect 701614 795513 701672 795523
rect 701682 795513 701740 795523
rect 701750 795513 701808 795523
rect 701818 795513 701876 795523
rect 699368 795489 700334 795513
rect 700910 795489 701876 795513
rect 699392 795474 699416 795489
rect 699460 795474 699484 795489
rect 699528 795474 699552 795489
rect 699596 795474 699620 795489
rect 699664 795474 699688 795489
rect 699732 795474 699756 795489
rect 699800 795474 699824 795489
rect 699868 795474 699892 795489
rect 699936 795474 699960 795489
rect 700004 795474 700028 795489
rect 700072 795474 700096 795489
rect 700140 795474 700164 795489
rect 700208 795474 700232 795489
rect 700276 795474 700300 795489
rect 700934 795474 700958 795489
rect 701002 795474 701026 795489
rect 701070 795474 701094 795489
rect 701138 795474 701162 795489
rect 701206 795474 701230 795489
rect 701274 795474 701298 795489
rect 701342 795474 701366 795489
rect 701410 795474 701434 795489
rect 701478 795474 701502 795489
rect 701546 795474 701570 795489
rect 701614 795474 701638 795489
rect 701682 795474 701706 795489
rect 701750 795474 701774 795489
rect 701818 795474 701842 795489
rect 699322 795319 700322 795474
rect 699322 795285 700334 795319
rect 700922 795309 701922 795474
rect 707610 795319 708610 795379
rect 709211 795319 710211 795379
rect 700910 795285 701922 795309
rect 699322 795274 700322 795285
rect 700922 795274 701922 795285
rect 699392 795261 699416 795274
rect 699460 795261 699484 795274
rect 699528 795261 699552 795274
rect 699596 795261 699620 795274
rect 699664 795261 699688 795274
rect 699732 795261 699756 795274
rect 699800 795261 699824 795274
rect 699868 795261 699892 795274
rect 699936 795261 699960 795274
rect 700004 795261 700028 795274
rect 700072 795261 700096 795274
rect 700140 795261 700164 795274
rect 700208 795261 700232 795274
rect 700276 795261 700300 795274
rect 700934 795261 700958 795274
rect 701002 795261 701026 795274
rect 701070 795261 701094 795274
rect 701138 795261 701162 795274
rect 701206 795261 701230 795274
rect 701274 795261 701298 795274
rect 701342 795261 701366 795274
rect 701410 795261 701434 795274
rect 701478 795261 701502 795274
rect 701546 795261 701570 795274
rect 701614 795261 701638 795274
rect 701682 795261 701706 795274
rect 701750 795261 701774 795274
rect 701818 795261 701842 795274
rect 699322 794916 700322 794972
rect 700922 794916 701922 794972
rect 707610 794961 708610 795017
rect 709211 794961 710211 795017
rect 699322 794844 700322 794900
rect 700922 794844 701922 794900
rect 707610 794889 708610 794945
rect 709211 794889 710211 794945
rect 699322 794542 700322 794614
rect 700922 794542 701922 794614
rect 707610 794587 708610 794659
rect 709211 794587 710211 794659
rect 699392 794531 699426 794542
rect 699460 794531 699494 794542
rect 699528 794531 699562 794542
rect 699596 794531 699630 794542
rect 699664 794531 699698 794542
rect 699732 794531 699766 794542
rect 699800 794531 699834 794542
rect 699868 794531 699902 794542
rect 699936 794531 699970 794542
rect 700004 794531 700038 794542
rect 700072 794531 700106 794542
rect 700140 794531 700174 794542
rect 700208 794531 700242 794542
rect 700276 794531 700310 794542
rect 700934 794531 700968 794542
rect 701002 794531 701036 794542
rect 701070 794531 701104 794542
rect 701138 794531 701172 794542
rect 701206 794531 701240 794542
rect 701274 794531 701308 794542
rect 701342 794531 701376 794542
rect 701410 794531 701444 794542
rect 701478 794531 701512 794542
rect 701546 794531 701580 794542
rect 701614 794531 701648 794542
rect 701682 794531 701716 794542
rect 701750 794531 701784 794542
rect 701818 794531 701852 794542
rect 699392 794521 699450 794531
rect 699460 794521 699518 794531
rect 699528 794521 699586 794531
rect 699596 794521 699654 794531
rect 699664 794521 699722 794531
rect 699732 794521 699790 794531
rect 699800 794521 699858 794531
rect 699868 794521 699926 794531
rect 699936 794521 699994 794531
rect 700004 794521 700062 794531
rect 700072 794521 700130 794531
rect 700140 794521 700198 794531
rect 700208 794521 700266 794531
rect 700276 794521 700334 794531
rect 700934 794521 700992 794531
rect 701002 794521 701060 794531
rect 701070 794521 701128 794531
rect 701138 794521 701196 794531
rect 701206 794521 701264 794531
rect 701274 794521 701332 794531
rect 701342 794521 701400 794531
rect 701410 794521 701468 794531
rect 701478 794521 701536 794531
rect 701546 794521 701604 794531
rect 701614 794521 701672 794531
rect 701682 794521 701740 794531
rect 701750 794521 701808 794531
rect 701818 794521 701876 794531
rect 699368 794497 700334 794521
rect 700910 794497 701876 794521
rect 699392 794482 699416 794497
rect 699460 794482 699484 794497
rect 699528 794482 699552 794497
rect 699596 794482 699620 794497
rect 699664 794482 699688 794497
rect 699732 794482 699756 794497
rect 699800 794482 699824 794497
rect 699868 794482 699892 794497
rect 699936 794482 699960 794497
rect 700004 794482 700028 794497
rect 700072 794482 700096 794497
rect 700140 794482 700164 794497
rect 700208 794482 700232 794497
rect 700276 794482 700300 794497
rect 700934 794482 700958 794497
rect 701002 794482 701026 794497
rect 701070 794482 701094 794497
rect 701138 794482 701162 794497
rect 701206 794482 701230 794497
rect 701274 794482 701298 794497
rect 701342 794482 701366 794497
rect 701410 794482 701434 794497
rect 701478 794482 701502 794497
rect 701546 794482 701570 794497
rect 701614 794482 701638 794497
rect 701682 794482 701706 794497
rect 701750 794482 701774 794497
rect 701818 794482 701842 794497
rect 699322 794327 700322 794482
rect 699322 794293 700334 794327
rect 700922 794317 701922 794482
rect 707610 794327 708610 794387
rect 709211 794327 710211 794387
rect 711541 794345 711629 801461
rect 711892 800200 711942 801200
rect 712062 800200 712112 801200
rect 711892 799079 711942 800079
rect 712062 799079 712112 800079
rect 711892 797958 711942 798958
rect 712062 797958 712112 798958
rect 711892 796848 711942 797848
rect 712062 796848 712112 797848
rect 711892 795727 711942 796727
rect 712062 795727 712112 796727
rect 711892 794606 711942 795606
rect 712062 794606 712112 795606
rect 712409 794371 712431 801485
rect 712469 801459 712487 801501
rect 712499 801459 712505 801467
rect 712499 801455 712511 801459
rect 712539 801455 712557 801501
rect 713640 799461 713674 801785
rect 713750 801772 714750 801822
rect 717367 801820 717413 801853
rect 717367 801819 717379 801820
rect 717401 801819 717413 801820
rect 717401 801809 717600 801819
rect 717401 801786 717413 801809
rect 713750 801562 714750 801612
rect 713750 801446 714750 801496
rect 713750 801230 714750 801358
rect 713750 801014 714750 801070
rect 713750 800798 714750 800926
rect 713750 800588 714750 800638
rect 714478 800585 714750 800588
rect 715486 799931 715536 800931
rect 715696 799931 715824 800931
rect 715912 799931 715962 800931
rect 713641 799345 713663 799461
rect 713640 799309 713674 799345
rect 713750 799314 714750 799364
rect 713750 799158 714750 799214
rect 713750 799002 714750 799130
rect 713750 798846 714750 798974
rect 713750 798690 714750 798746
rect 716425 798709 716725 798721
rect 713750 798534 714750 798662
rect 716425 798596 717425 798646
rect 713750 798378 714750 798506
rect 716425 798440 717425 798568
rect 713750 798222 714750 798350
rect 716425 798284 717425 798340
rect 713750 798072 714750 798122
rect 713750 797956 714750 798006
rect 713750 797800 714750 797928
rect 713750 797644 714750 797772
rect 713750 797488 714750 797616
rect 715354 797587 715404 798187
rect 715504 797587 715560 798187
rect 715660 797587 715716 798187
rect 715816 797587 715872 798187
rect 715972 797587 716022 798187
rect 716425 798128 717425 798256
rect 716425 797978 717425 798028
rect 716425 797862 717425 797912
rect 716425 797706 717425 797834
rect 716425 797550 717425 797606
rect 716425 797394 717425 797522
rect 713750 797332 714750 797388
rect 713750 797176 714750 797304
rect 716425 797244 717425 797294
rect 713750 797020 714750 797148
rect 713750 796870 714750 796920
rect 713750 796742 714750 796792
rect 713750 796586 714750 796642
rect 713750 796436 714750 796486
rect 713750 796320 714350 796370
rect 713750 796164 714350 796292
rect 715510 796191 715560 797191
rect 715660 796191 715788 797191
rect 715816 796191 715944 797191
rect 715972 796191 716022 797191
rect 716425 797128 717425 797178
rect 716425 796972 717425 797028
rect 716425 796822 717425 796872
rect 716425 796706 717425 796756
rect 716425 796550 717425 796678
rect 716425 796394 717425 796522
rect 716425 796238 717425 796366
rect 716425 796082 717425 796210
rect 713750 796008 714350 796064
rect 713750 795852 714350 795980
rect 716425 795932 717425 795982
rect 713750 795696 714350 795752
rect 713750 795446 714350 795496
rect 714565 795443 714765 795455
rect 713750 795330 714750 795380
rect 713750 795120 714750 795170
rect 716413 795092 716447 795150
rect 713750 795004 714750 795054
rect 713750 794794 714750 794844
rect 713750 794678 714750 794728
rect 713750 794468 714750 794518
rect 713750 794352 714750 794402
rect 700910 794293 701922 794317
rect 699322 794282 700322 794293
rect 700922 794282 701922 794293
rect 711541 794311 711633 794345
rect 699392 794269 699416 794282
rect 699460 794269 699484 794282
rect 699528 794269 699552 794282
rect 699596 794269 699620 794282
rect 699664 794269 699688 794282
rect 699732 794269 699756 794282
rect 699800 794269 699824 794282
rect 699868 794269 699892 794282
rect 699936 794269 699960 794282
rect 700004 794269 700028 794282
rect 700072 794269 700096 794282
rect 700140 794269 700164 794282
rect 700208 794269 700232 794282
rect 700276 794269 700300 794282
rect 700934 794269 700958 794282
rect 701002 794269 701026 794282
rect 701070 794269 701094 794282
rect 701138 794269 701162 794282
rect 701206 794269 701230 794282
rect 701274 794269 701298 794282
rect 701342 794269 701366 794282
rect 701410 794269 701434 794282
rect 701478 794269 701502 794282
rect 701546 794269 701570 794282
rect 701614 794269 701638 794282
rect 701682 794269 701706 794282
rect 701750 794269 701774 794282
rect 701818 794269 701842 794282
rect 699322 793924 700322 793980
rect 700922 793924 701922 793980
rect 707610 793969 708610 794025
rect 709211 793969 710211 794025
rect 699322 793852 700322 793908
rect 700922 793852 701922 793908
rect 707610 793897 708610 793953
rect 709211 793897 710211 793953
rect 699322 793550 700322 793622
rect 700922 793550 701922 793622
rect 707610 793595 708610 793667
rect 709211 793595 710211 793667
rect 699392 793539 699426 793550
rect 699460 793539 699494 793550
rect 699528 793539 699562 793550
rect 699596 793539 699630 793550
rect 699664 793539 699698 793550
rect 699732 793539 699766 793550
rect 699800 793539 699834 793550
rect 699868 793539 699902 793550
rect 699936 793539 699970 793550
rect 700004 793539 700038 793550
rect 700072 793539 700106 793550
rect 700140 793539 700174 793550
rect 700208 793539 700242 793550
rect 700276 793539 700310 793550
rect 700934 793539 700968 793550
rect 701002 793539 701036 793550
rect 701070 793539 701104 793550
rect 701138 793539 701172 793550
rect 701206 793539 701240 793550
rect 701274 793539 701308 793550
rect 701342 793539 701376 793550
rect 701410 793539 701444 793550
rect 701478 793539 701512 793550
rect 701546 793539 701580 793550
rect 701614 793539 701648 793550
rect 701682 793539 701716 793550
rect 701750 793539 701784 793550
rect 701818 793539 701852 793550
rect 699392 793529 699450 793539
rect 699460 793529 699518 793539
rect 699528 793529 699586 793539
rect 699596 793529 699654 793539
rect 699664 793529 699722 793539
rect 699732 793529 699790 793539
rect 699800 793529 699858 793539
rect 699868 793529 699926 793539
rect 699936 793529 699994 793539
rect 700004 793529 700062 793539
rect 700072 793529 700130 793539
rect 700140 793529 700198 793539
rect 700208 793529 700266 793539
rect 700276 793529 700334 793539
rect 700934 793529 700992 793539
rect 701002 793529 701060 793539
rect 701070 793529 701128 793539
rect 701138 793529 701196 793539
rect 701206 793529 701264 793539
rect 701274 793529 701332 793539
rect 701342 793529 701400 793539
rect 701410 793529 701468 793539
rect 701478 793529 701536 793539
rect 701546 793529 701604 793539
rect 701614 793529 701672 793539
rect 701682 793529 701740 793539
rect 701750 793529 701808 793539
rect 701818 793529 701876 793539
rect 699368 793505 700334 793529
rect 700910 793505 701876 793529
rect 699392 793490 699416 793505
rect 699460 793490 699484 793505
rect 699528 793490 699552 793505
rect 699596 793490 699620 793505
rect 699664 793490 699688 793505
rect 699732 793490 699756 793505
rect 699800 793490 699824 793505
rect 699868 793490 699892 793505
rect 699936 793490 699960 793505
rect 700004 793490 700028 793505
rect 700072 793490 700096 793505
rect 700140 793490 700164 793505
rect 700208 793490 700232 793505
rect 700276 793490 700300 793505
rect 700934 793490 700958 793505
rect 701002 793490 701026 793505
rect 701070 793490 701094 793505
rect 701138 793490 701162 793505
rect 701206 793490 701230 793505
rect 701274 793490 701298 793505
rect 701342 793490 701366 793505
rect 701410 793490 701434 793505
rect 701478 793490 701502 793505
rect 701546 793490 701570 793505
rect 701614 793490 701638 793505
rect 701682 793490 701706 793505
rect 701750 793490 701774 793505
rect 701818 793490 701842 793505
rect 699322 793335 700322 793490
rect 699322 793301 700334 793335
rect 700922 793325 701922 793490
rect 707610 793335 708610 793395
rect 709211 793335 710211 793395
rect 700910 793301 701922 793325
rect 699322 793290 700322 793301
rect 700922 793290 701922 793301
rect 699392 793277 699416 793290
rect 699460 793277 699484 793290
rect 699528 793277 699552 793290
rect 699596 793277 699620 793290
rect 699664 793277 699688 793290
rect 699732 793277 699756 793290
rect 699800 793277 699824 793290
rect 699868 793277 699892 793290
rect 699936 793277 699960 793290
rect 700004 793277 700028 793290
rect 700072 793277 700096 793290
rect 700140 793277 700164 793290
rect 700208 793277 700232 793290
rect 700276 793277 700300 793290
rect 700934 793277 700958 793290
rect 701002 793277 701026 793290
rect 701070 793277 701094 793290
rect 701138 793277 701162 793290
rect 701206 793277 701230 793290
rect 701274 793277 701298 793290
rect 701342 793277 701366 793290
rect 701410 793277 701434 793290
rect 701478 793277 701502 793290
rect 701546 793277 701570 793290
rect 701614 793277 701638 793290
rect 701682 793277 701706 793290
rect 701750 793277 701774 793290
rect 701818 793277 701842 793290
rect 699322 792932 700322 792988
rect 700922 792932 701922 792988
rect 707610 792977 708610 793033
rect 709211 792977 710211 793033
rect 699322 792860 700322 792916
rect 700922 792860 701922 792916
rect 707610 792905 708610 792961
rect 709211 792905 710211 792961
rect 699322 792558 700322 792630
rect 700922 792558 701922 792630
rect 707610 792603 708610 792675
rect 709211 792603 710211 792675
rect 699392 792547 699426 792558
rect 699460 792547 699494 792558
rect 699528 792547 699562 792558
rect 699596 792547 699630 792558
rect 699664 792547 699698 792558
rect 699732 792547 699766 792558
rect 699800 792547 699834 792558
rect 699868 792547 699902 792558
rect 699936 792547 699970 792558
rect 700004 792547 700038 792558
rect 700072 792547 700106 792558
rect 700140 792547 700174 792558
rect 700208 792547 700242 792558
rect 700276 792547 700310 792558
rect 700934 792547 700968 792558
rect 701002 792547 701036 792558
rect 701070 792547 701104 792558
rect 701138 792547 701172 792558
rect 701206 792547 701240 792558
rect 701274 792547 701308 792558
rect 701342 792547 701376 792558
rect 701410 792547 701444 792558
rect 701478 792547 701512 792558
rect 701546 792547 701580 792558
rect 701614 792547 701648 792558
rect 701682 792547 701716 792558
rect 701750 792547 701784 792558
rect 701818 792547 701852 792558
rect 699392 792537 699450 792547
rect 699460 792537 699518 792547
rect 699528 792537 699586 792547
rect 699596 792537 699654 792547
rect 699664 792537 699722 792547
rect 699732 792537 699790 792547
rect 699800 792537 699858 792547
rect 699868 792537 699926 792547
rect 699936 792537 699994 792547
rect 700004 792537 700062 792547
rect 700072 792537 700130 792547
rect 700140 792537 700198 792547
rect 700208 792537 700266 792547
rect 700276 792537 700334 792547
rect 700934 792537 700992 792547
rect 701002 792537 701060 792547
rect 701070 792537 701128 792547
rect 701138 792537 701196 792547
rect 701206 792537 701264 792547
rect 701274 792537 701332 792547
rect 701342 792537 701400 792547
rect 701410 792537 701468 792547
rect 701478 792537 701536 792547
rect 701546 792537 701604 792547
rect 701614 792537 701672 792547
rect 701682 792537 701740 792547
rect 701750 792537 701808 792547
rect 701818 792537 701876 792547
rect 699368 792513 700334 792537
rect 700910 792513 701876 792537
rect 699392 792498 699416 792513
rect 699460 792498 699484 792513
rect 699528 792498 699552 792513
rect 699596 792498 699620 792513
rect 699664 792498 699688 792513
rect 699732 792498 699756 792513
rect 699800 792498 699824 792513
rect 699868 792498 699892 792513
rect 699936 792498 699960 792513
rect 700004 792498 700028 792513
rect 700072 792498 700096 792513
rect 700140 792498 700164 792513
rect 700208 792498 700232 792513
rect 700276 792498 700300 792513
rect 700934 792498 700958 792513
rect 701002 792498 701026 792513
rect 701070 792498 701094 792513
rect 701138 792498 701162 792513
rect 701206 792498 701230 792513
rect 701274 792498 701298 792513
rect 701342 792498 701366 792513
rect 701410 792498 701434 792513
rect 701478 792498 701502 792513
rect 701546 792498 701570 792513
rect 701614 792498 701638 792513
rect 701682 792498 701706 792513
rect 701750 792498 701774 792513
rect 701818 792498 701842 792513
rect 699322 792343 700322 792498
rect 699322 792309 700334 792343
rect 700922 792333 701922 792498
rect 707610 792343 708610 792403
rect 709211 792343 710211 792403
rect 700910 792309 701922 792333
rect 699322 792298 700322 792309
rect 700922 792298 701922 792309
rect 699392 792285 699416 792298
rect 699460 792285 699484 792298
rect 699528 792285 699552 792298
rect 699596 792285 699620 792298
rect 699664 792285 699688 792298
rect 699732 792285 699756 792298
rect 699800 792285 699824 792298
rect 699868 792285 699892 792298
rect 699936 792285 699960 792298
rect 700004 792285 700028 792298
rect 700072 792285 700096 792298
rect 700140 792285 700164 792298
rect 700208 792285 700232 792298
rect 700276 792285 700300 792298
rect 700934 792285 700958 792298
rect 701002 792285 701026 792298
rect 701070 792285 701094 792298
rect 701138 792285 701162 792298
rect 701206 792285 701230 792298
rect 701274 792285 701298 792298
rect 701342 792285 701366 792298
rect 701410 792285 701434 792298
rect 701478 792285 701502 792298
rect 701546 792285 701570 792298
rect 701614 792285 701638 792298
rect 701682 792285 701706 792298
rect 701750 792285 701774 792298
rect 701818 792285 701842 792298
rect 699322 791940 700322 791996
rect 700922 791940 701922 791996
rect 707610 791985 708610 792041
rect 709211 791985 710211 792041
rect 699322 791868 700322 791924
rect 700922 791868 701922 791924
rect 707610 791913 708610 791969
rect 709211 791913 710211 791969
rect 699322 791566 700322 791638
rect 700922 791566 701922 791638
rect 707610 791611 708610 791683
rect 709211 791611 710211 791683
rect 699392 791555 699426 791566
rect 699460 791555 699494 791566
rect 699528 791555 699562 791566
rect 699596 791555 699630 791566
rect 699664 791555 699698 791566
rect 699732 791555 699766 791566
rect 699800 791555 699834 791566
rect 699868 791555 699902 791566
rect 699936 791555 699970 791566
rect 700004 791555 700038 791566
rect 700072 791555 700106 791566
rect 700140 791555 700174 791566
rect 700208 791555 700242 791566
rect 700276 791555 700310 791566
rect 700934 791555 700968 791566
rect 701002 791555 701036 791566
rect 701070 791555 701104 791566
rect 701138 791555 701172 791566
rect 701206 791555 701240 791566
rect 701274 791555 701308 791566
rect 701342 791555 701376 791566
rect 701410 791555 701444 791566
rect 701478 791555 701512 791566
rect 701546 791555 701580 791566
rect 701614 791555 701648 791566
rect 701682 791555 701716 791566
rect 701750 791555 701784 791566
rect 701818 791555 701852 791566
rect 699392 791545 699450 791555
rect 699460 791545 699518 791555
rect 699528 791545 699586 791555
rect 699596 791545 699654 791555
rect 699664 791545 699722 791555
rect 699732 791545 699790 791555
rect 699800 791545 699858 791555
rect 699868 791545 699926 791555
rect 699936 791545 699994 791555
rect 700004 791545 700062 791555
rect 700072 791545 700130 791555
rect 700140 791545 700198 791555
rect 700208 791545 700266 791555
rect 700276 791545 700334 791555
rect 700934 791545 700992 791555
rect 701002 791545 701060 791555
rect 701070 791545 701128 791555
rect 701138 791545 701196 791555
rect 701206 791545 701264 791555
rect 701274 791545 701332 791555
rect 701342 791545 701400 791555
rect 701410 791545 701468 791555
rect 701478 791545 701536 791555
rect 701546 791545 701604 791555
rect 701614 791545 701672 791555
rect 701682 791545 701740 791555
rect 701750 791545 701808 791555
rect 701818 791545 701876 791555
rect 699368 791521 700334 791545
rect 700910 791521 701876 791545
rect 699392 791506 699416 791521
rect 699460 791506 699484 791521
rect 699528 791506 699552 791521
rect 699596 791506 699620 791521
rect 699664 791506 699688 791521
rect 699732 791506 699756 791521
rect 699800 791506 699824 791521
rect 699868 791506 699892 791521
rect 699936 791506 699960 791521
rect 700004 791506 700028 791521
rect 700072 791506 700096 791521
rect 700140 791506 700164 791521
rect 700208 791506 700232 791521
rect 700276 791506 700300 791521
rect 700934 791506 700958 791521
rect 701002 791506 701026 791521
rect 701070 791506 701094 791521
rect 701138 791506 701162 791521
rect 701206 791506 701230 791521
rect 701274 791506 701298 791521
rect 701342 791506 701366 791521
rect 701410 791506 701434 791521
rect 701478 791506 701502 791521
rect 701546 791506 701570 791521
rect 701614 791506 701638 791521
rect 701682 791506 701706 791521
rect 701750 791506 701774 791521
rect 701818 791506 701842 791521
rect 699322 791351 700322 791506
rect 699322 791317 700334 791351
rect 700922 791341 701922 791506
rect 705107 791360 705173 791376
rect 707610 791351 708610 791411
rect 709211 791351 710211 791411
rect 700910 791317 701922 791341
rect 699322 791306 700322 791317
rect 700922 791306 701922 791317
rect 699392 791293 699416 791306
rect 699460 791293 699484 791306
rect 699528 791293 699552 791306
rect 699596 791293 699620 791306
rect 699664 791293 699688 791306
rect 699732 791293 699756 791306
rect 699800 791293 699824 791306
rect 699868 791293 699892 791306
rect 699936 791293 699960 791306
rect 700004 791293 700028 791306
rect 700072 791293 700096 791306
rect 700140 791293 700164 791306
rect 700208 791293 700232 791306
rect 700276 791293 700300 791306
rect 700934 791293 700958 791306
rect 701002 791293 701026 791306
rect 701070 791293 701094 791306
rect 701138 791293 701162 791306
rect 701206 791293 701230 791306
rect 701274 791293 701298 791306
rect 701342 791293 701366 791306
rect 701410 791293 701434 791306
rect 701478 791293 701502 791306
rect 701546 791293 701570 791306
rect 701614 791293 701638 791306
rect 701682 791293 701706 791306
rect 701750 791293 701774 791306
rect 701818 791293 701842 791306
rect 699322 790948 700322 791004
rect 700922 790948 701922 791004
rect 707610 790993 708610 791049
rect 709211 790993 710211 791049
rect 699322 790876 700322 790932
rect 700922 790876 701922 790932
rect 707610 790921 708610 790977
rect 709211 790921 710211 790977
rect 699322 790574 700322 790646
rect 700922 790574 701922 790646
rect 707610 790619 708610 790691
rect 709211 790619 710211 790691
rect 699392 790563 699426 790574
rect 699460 790563 699494 790574
rect 699528 790563 699562 790574
rect 699596 790563 699630 790574
rect 699664 790563 699698 790574
rect 699732 790563 699766 790574
rect 699800 790563 699834 790574
rect 699868 790563 699902 790574
rect 699936 790563 699970 790574
rect 700004 790563 700038 790574
rect 700072 790563 700106 790574
rect 700140 790563 700174 790574
rect 700208 790563 700242 790574
rect 700276 790563 700310 790574
rect 700934 790563 700968 790574
rect 701002 790563 701036 790574
rect 701070 790563 701104 790574
rect 701138 790563 701172 790574
rect 701206 790563 701240 790574
rect 701274 790563 701308 790574
rect 701342 790563 701376 790574
rect 701410 790563 701444 790574
rect 701478 790563 701512 790574
rect 701546 790563 701580 790574
rect 701614 790563 701648 790574
rect 701682 790563 701716 790574
rect 701750 790563 701784 790574
rect 701818 790563 701852 790574
rect 699392 790553 699450 790563
rect 699460 790553 699518 790563
rect 699528 790553 699586 790563
rect 699596 790553 699654 790563
rect 699664 790553 699722 790563
rect 699732 790553 699790 790563
rect 699800 790553 699858 790563
rect 699868 790553 699926 790563
rect 699936 790553 699994 790563
rect 700004 790553 700062 790563
rect 700072 790553 700130 790563
rect 700140 790553 700198 790563
rect 700208 790553 700266 790563
rect 700276 790553 700334 790563
rect 700934 790553 700992 790563
rect 701002 790553 701060 790563
rect 701070 790553 701128 790563
rect 701138 790553 701196 790563
rect 701206 790553 701264 790563
rect 701274 790553 701332 790563
rect 701342 790553 701400 790563
rect 701410 790553 701468 790563
rect 701478 790553 701536 790563
rect 701546 790553 701604 790563
rect 701614 790553 701672 790563
rect 701682 790553 701740 790563
rect 701750 790553 701808 790563
rect 701818 790553 701876 790563
rect 699368 790529 700334 790553
rect 700910 790529 701876 790553
rect 699392 790514 699416 790529
rect 699460 790514 699484 790529
rect 699528 790514 699552 790529
rect 699596 790514 699620 790529
rect 699664 790514 699688 790529
rect 699732 790514 699756 790529
rect 699800 790514 699824 790529
rect 699868 790514 699892 790529
rect 699936 790514 699960 790529
rect 700004 790514 700028 790529
rect 700072 790514 700096 790529
rect 700140 790514 700164 790529
rect 700208 790514 700232 790529
rect 700276 790514 700300 790529
rect 700934 790514 700958 790529
rect 701002 790514 701026 790529
rect 701070 790514 701094 790529
rect 701138 790514 701162 790529
rect 701206 790514 701230 790529
rect 701274 790514 701298 790529
rect 701342 790514 701366 790529
rect 701410 790514 701434 790529
rect 701478 790514 701502 790529
rect 701546 790514 701570 790529
rect 701614 790514 701638 790529
rect 701682 790514 701706 790529
rect 701750 790514 701774 790529
rect 701818 790514 701842 790529
rect 699322 790359 700322 790514
rect 699322 790325 700334 790359
rect 700922 790349 701922 790514
rect 707610 790359 708610 790419
rect 709211 790359 710211 790419
rect 700910 790325 701922 790349
rect 699322 790314 700322 790325
rect 700922 790314 701922 790325
rect 699392 790301 699416 790314
rect 699460 790301 699484 790314
rect 699528 790301 699552 790314
rect 699596 790301 699620 790314
rect 699664 790301 699688 790314
rect 699732 790301 699756 790314
rect 699800 790301 699824 790314
rect 699868 790301 699892 790314
rect 699936 790301 699960 790314
rect 700004 790301 700028 790314
rect 700072 790301 700096 790314
rect 700140 790301 700164 790314
rect 700208 790301 700232 790314
rect 700276 790301 700300 790314
rect 700934 790301 700958 790314
rect 701002 790301 701026 790314
rect 701070 790301 701094 790314
rect 701138 790301 701162 790314
rect 701206 790301 701230 790314
rect 701274 790301 701298 790314
rect 701342 790301 701366 790314
rect 701410 790301 701434 790314
rect 701478 790301 701502 790314
rect 701546 790301 701570 790314
rect 701614 790301 701638 790314
rect 701682 790301 701706 790314
rect 701750 790301 701774 790314
rect 701818 790301 701842 790314
rect 709211 790148 710211 790152
rect 707574 790099 707610 790134
rect 708610 790099 708646 790134
rect 707574 790098 708646 790099
rect 707574 790057 707610 790098
rect 708610 790057 708646 790098
rect 699322 789956 700322 790012
rect 700922 789956 701922 790012
rect 707574 790001 708646 790057
rect 707574 789964 707610 790001
rect 708610 789964 708646 790001
rect 707574 789959 708646 789964
rect 699322 789884 700322 789940
rect 700922 789884 701922 789940
rect 707574 789924 707610 789959
rect 708610 789924 708646 789959
rect 709175 790098 710247 790134
rect 709175 790057 709211 790098
rect 710211 790057 710247 790098
rect 709175 790001 710247 790057
rect 709175 789964 709211 790001
rect 710211 789964 710247 790001
rect 709175 789936 710247 789964
rect 709175 789924 709211 789936
rect 710211 789924 710247 789936
rect 707610 789713 708610 789785
rect 709211 789713 710211 789785
rect 699322 789623 700322 789673
rect 700922 789623 701922 789673
rect 707610 789523 708610 789617
rect 707610 789513 708644 789523
rect 709211 789513 710211 789591
rect 711541 789437 711629 794311
rect 713750 794136 714750 794264
rect 716417 794152 717417 794202
rect 711892 793049 711942 794049
rect 712062 793049 712112 794049
rect 713750 793920 714750 794048
rect 716417 793996 717417 794052
rect 716417 793846 717417 793896
rect 713750 793704 714750 793832
rect 716417 793730 717017 793780
rect 716417 793580 717017 793630
rect 713750 793488 714750 793544
rect 716417 793464 717417 793514
rect 713750 793272 714750 793400
rect 716417 793308 717417 793364
rect 713750 793056 714750 793184
rect 716417 793152 717417 793280
rect 716417 792996 717417 793052
rect 711892 791928 711942 792928
rect 712062 791928 712112 792928
rect 713750 792840 714750 792968
rect 716417 792840 717417 792968
rect 713750 792624 714750 792752
rect 716417 792684 717417 792740
rect 716417 792474 717417 792524
rect 713750 792408 714750 792464
rect 716417 792308 717417 792358
rect 713750 792192 714750 792248
rect 716417 792152 717417 792280
rect 713750 791976 714750 792104
rect 716417 791996 717417 792052
rect 711892 790807 711942 791807
rect 712062 790807 712112 791807
rect 713750 791760 714750 791888
rect 716417 791780 717417 791836
rect 713750 791544 714750 791672
rect 716417 791570 717417 791620
rect 713750 791328 714750 791456
rect 716417 791454 717417 791504
rect 716417 791298 717417 791426
rect 713750 791118 714750 791168
rect 716417 791148 717417 791198
rect 711892 789697 711942 790697
rect 712062 789697 712112 790697
rect 714686 790357 714794 790424
rect 714645 790323 714794 790357
rect 716071 790357 716074 790358
rect 716071 790356 716072 790357
rect 716073 790356 716074 790357
rect 716071 790355 716074 790356
rect 716208 790357 716211 790358
rect 716208 790356 716209 790357
rect 716210 790356 716211 790357
rect 716208 790355 716211 790356
rect 714964 790247 715998 790329
rect 716284 790247 717318 790329
rect 705107 789336 705173 789352
rect 711541 789302 711633 789437
rect 714175 789398 714225 789998
rect 714425 789398 714475 789998
rect 711579 789301 711595 789302
rect 714781 789191 714863 790226
rect 715134 789955 715828 790037
rect 714686 789123 714863 789191
rect 714645 789089 714863 789123
rect 680215 788880 680815 788936
rect 686719 788893 686739 788917
rect 686743 788893 686753 788917
rect 686719 788859 686757 788893
rect 686719 788822 686739 788859
rect 686743 788822 686753 788859
rect 692428 788850 693028 788978
rect 698017 788947 698210 788983
rect 698084 788935 698210 788947
rect 702756 788959 703645 788983
rect 702756 788935 702853 788959
rect 698084 788828 702853 788935
rect 686719 788788 686757 788822
rect 680215 788704 680815 788760
rect 686719 788751 686739 788788
rect 686743 788751 686753 788788
rect 686719 788741 686757 788751
rect 686699 788717 686767 788741
rect 686719 788704 686739 788717
rect 686743 788704 686753 788717
rect 686719 788695 686753 788704
rect 686719 788693 686743 788695
rect 692428 788694 693028 788750
rect 686685 788656 686709 788680
rect 686743 788656 686767 788680
rect 678799 788503 679399 788553
rect 680215 788534 680815 788584
rect 692428 788538 693028 788666
rect 680593 788531 680815 788534
rect 682009 788501 682069 788516
rect 682024 788465 682054 788501
rect 683708 788387 684308 788437
rect 678799 788327 679399 788383
rect 692428 788382 693028 788510
rect 714781 788308 714863 789089
rect 715063 788609 715145 789915
rect 715342 789752 715382 789792
rect 715582 789752 715622 789792
rect 715289 788777 715339 789719
rect 715382 789668 715422 789752
rect 715542 789668 715582 789752
rect 715633 788777 715683 789719
rect 715382 788672 715422 788756
rect 715542 788672 715582 788756
rect 715342 788632 715382 788672
rect 715582 788632 715622 788672
rect 715815 788609 715897 789915
rect 715134 788387 715828 788469
rect 716100 788308 716182 790226
rect 716454 789955 717148 790037
rect 716385 788609 716467 789915
rect 716660 789752 716700 789792
rect 716900 789752 716940 789792
rect 716599 788777 716649 789719
rect 716700 789668 716740 789752
rect 716860 789668 716900 789752
rect 716943 788777 716993 789719
rect 716700 788672 716740 788756
rect 716860 788672 716900 788756
rect 716660 788632 716700 788672
rect 716900 788632 716940 788672
rect 717137 788609 717219 789915
rect 716454 788387 717148 788469
rect 717419 788308 717501 790226
rect 683708 788237 684308 788287
rect 692428 788232 693028 788282
rect 678799 788157 679399 788207
rect 684565 788160 684790 788168
rect 696597 788000 696600 788120
rect 714964 788095 715998 788177
rect 716284 788095 717318 788177
rect 21000 765000 21003 765120
rect 282 764623 1316 764705
rect 1602 764623 2636 764705
rect 32810 764662 33035 764670
rect 38201 764593 38801 764643
rect 24572 764518 25172 764568
rect 33292 764513 33892 764563
rect 99 762574 181 764492
rect 452 764331 1146 764413
rect 381 762885 463 764191
rect 660 764128 700 764168
rect 900 764128 940 764168
rect 700 764044 740 764128
rect 860 764044 900 764128
rect 607 763081 657 764023
rect 700 763048 740 763132
rect 860 763048 900 763132
rect 951 763081 1001 764023
rect 660 763008 700 763048
rect 900 763008 940 763048
rect 1133 762885 1215 764191
rect 452 762763 1146 762845
rect 1418 762574 1500 764492
rect 1772 764331 2466 764413
rect 1703 762885 1785 764191
rect 1978 764128 2018 764168
rect 2218 764128 2258 764168
rect 2018 764044 2058 764128
rect 2178 764044 2218 764128
rect 1917 763081 1967 764023
rect 2018 763048 2058 763132
rect 2178 763048 2218 763132
rect 2261 763081 2311 764023
rect 1978 763008 2018 763048
rect 2218 763008 2258 763048
rect 2455 762885 2537 764191
rect 2737 763779 2819 764492
rect 24572 764362 25172 764490
rect 38201 764417 38801 764473
rect 33292 764363 33892 764413
rect 24572 764206 25172 764334
rect 35546 764299 35576 764335
rect 36785 764329 36935 764341
rect 35531 764284 35591 764299
rect 36785 764216 37385 764266
rect 38201 764247 38801 764297
rect 30833 764120 30857 764144
rect 30891 764120 30915 764144
rect 24572 764050 25172 764106
rect 30857 764105 30881 764107
rect 30857 764096 30887 764105
rect 30867 764083 30887 764096
rect 30891 764083 30907 764120
rect 30833 764059 30857 764083
rect 30867 764049 30911 764083
rect 14747 763865 19516 763972
rect 24572 763894 25172 764022
rect 30867 764012 30887 764049
rect 30891 764012 30907 764049
rect 36785 764040 37385 764096
rect 30867 763978 30911 764012
rect 30867 763941 30887 763978
rect 30891 763941 30907 763978
rect 30867 763907 30911 763941
rect 30867 763883 30887 763907
rect 30891 763883 30907 763907
rect 14747 763841 14844 763865
rect 13955 763817 14844 763841
rect 19390 763853 19516 763865
rect 19390 763841 19583 763853
rect 19390 763817 19605 763841
rect 19639 763817 19673 763841
rect 19707 763817 19741 763841
rect 19775 763817 19809 763841
rect 19843 763817 19877 763841
rect 19911 763817 19945 763841
rect 19979 763817 20013 763841
rect 20047 763817 20081 763841
rect 20115 763817 20149 763841
rect 20183 763817 20217 763841
rect 20251 763817 20285 763841
rect 20319 763817 20353 763841
rect 20387 763817 20421 763841
rect 20455 763817 20489 763841
rect 20523 763817 20557 763841
rect 20591 763817 20625 763841
rect 20659 763817 20693 763841
rect 2737 763711 2914 763779
rect 1772 762763 2466 762845
rect 2737 762574 2819 763711
rect 2848 763677 2955 763711
rect 6005 763498 6021 763499
rect 3125 762802 3175 763402
rect 3375 762802 3425 763402
rect 5967 763363 6059 763498
rect 12427 763448 12493 763464
rect 282 762471 1316 762553
rect 1602 762471 2636 762553
rect 2806 762477 2914 762545
rect 1389 762444 1392 762445
rect 1389 762443 1390 762444
rect 1391 762443 1392 762444
rect 1389 762442 1392 762443
rect 1526 762444 1529 762445
rect 1526 762443 1527 762444
rect 1528 762443 1529 762444
rect 2848 762443 2955 762477
rect 1526 762442 1529 762443
rect 5488 762103 5538 763103
rect 5658 762103 5708 763103
rect 183 761602 1183 761652
rect 2850 761632 3850 761682
rect 183 761446 1183 761574
rect 2850 761416 3850 761544
rect 183 761296 1183 761346
rect 183 761180 1183 761230
rect 2850 761200 3850 761328
rect 183 760964 1183 761020
rect 2850 760984 3850 761112
rect 5488 760993 5538 761993
rect 5658 760993 5708 761993
rect 183 760748 1183 760804
rect 2850 760768 3850 760896
rect 183 760592 1183 760720
rect 2850 760552 3850 760608
rect 183 760442 1183 760492
rect 2850 760336 3850 760392
rect 183 760276 1183 760326
rect 2850 760120 3850 760248
rect 183 760060 1183 760116
rect 183 759904 1183 760032
rect 2850 759904 3850 760032
rect 5488 759872 5538 760872
rect 5658 759872 5708 760872
rect 183 759748 1183 759804
rect 183 759592 1183 759720
rect 2850 759688 3850 759816
rect 183 759436 1183 759492
rect 2850 759472 3850 759600
rect 183 759286 1183 759336
rect 2850 759256 3850 759312
rect 583 759170 1183 759220
rect 583 759020 1183 759070
rect 2850 759040 3850 759168
rect 183 758904 1183 758954
rect 2850 758824 3850 758952
rect 183 758748 1183 758804
rect 5488 758751 5538 759751
rect 5658 758751 5708 759751
rect 183 758598 1183 758648
rect 2850 758608 3850 758736
rect 5971 758489 6059 763363
rect 7406 763287 7440 763321
rect 7477 763287 7511 763321
rect 7551 763287 7585 763321
rect 7622 763287 7656 763321
rect 7696 763287 7730 763321
rect 7767 763287 7801 763321
rect 7841 763287 7875 763321
rect 7912 763287 7946 763321
rect 7986 763287 8020 763321
rect 8057 763287 8091 763321
rect 8131 763287 8165 763321
rect 8202 763287 8236 763321
rect 8296 763287 8330 763321
rect 8381 763311 8423 763321
rect 8381 763287 8389 763311
rect 8415 763287 8423 763311
rect 8956 763311 8996 763321
rect 8956 763287 8962 763311
rect 8990 763287 8996 763311
rect 9044 763287 9078 763321
rect 9120 763287 9154 763321
rect 9197 763287 9231 763321
rect 9291 763287 9325 763321
rect 9362 763287 9396 763321
rect 9436 763287 9470 763321
rect 9507 763287 9541 763321
rect 9581 763287 9615 763321
rect 9652 763287 9686 763321
rect 9726 763287 9760 763321
rect 9797 763287 9831 763321
rect 9871 763287 9905 763321
rect 9942 763287 9976 763321
rect 7389 763277 7406 763287
rect 7440 763277 7477 763287
rect 7511 763277 7551 763287
rect 7585 763277 7622 763287
rect 7656 763277 7696 763287
rect 7730 763277 7767 763287
rect 7801 763277 7841 763287
rect 7875 763277 7912 763287
rect 7946 763277 7986 763287
rect 8020 763277 8057 763287
rect 8091 763277 8131 763287
rect 8165 763277 8202 763287
rect 8236 763277 8296 763287
rect 8330 763277 8381 763287
rect 8389 763277 8423 763287
rect 8990 763277 9044 763287
rect 9078 763277 9120 763287
rect 9154 763277 9197 763287
rect 9231 763277 9291 763287
rect 9325 763277 9362 763287
rect 9396 763277 9436 763287
rect 9470 763277 9507 763287
rect 9541 763277 9581 763287
rect 9615 763277 9652 763287
rect 9686 763277 9726 763287
rect 9760 763277 9797 763287
rect 9831 763277 9871 763287
rect 9905 763277 9942 763287
rect 9976 763277 9990 763287
rect 7389 763209 8389 763277
rect 8990 763183 9990 763277
rect 7389 763087 8389 763147
rect 8990 763087 9990 763147
rect 15678 763127 16678 763177
rect 17278 763127 18278 763177
rect 7353 762864 7389 762876
rect 8389 762864 8425 762876
rect 7353 762840 8425 762864
rect 7353 762799 7389 762840
rect 8389 762799 8425 762840
rect 7353 762743 8425 762799
rect 7353 762706 7389 762743
rect 8389 762706 8425 762743
rect 7353 762666 8425 762706
rect 8954 762841 8990 762876
rect 9990 762841 10026 762876
rect 15678 762860 16678 762916
rect 17278 762860 18278 762916
rect 8954 762840 10026 762841
rect 8954 762799 8990 762840
rect 9990 762799 10026 762840
rect 8954 762743 10026 762799
rect 15678 762788 16678 762844
rect 17278 762788 18278 762844
rect 8954 762706 8990 762743
rect 9990 762706 10026 762743
rect 8954 762701 10026 762706
rect 8954 762666 8990 762701
rect 9990 762666 10026 762701
rect 7389 762441 8389 762513
rect 8990 762441 9990 762513
rect 15678 762486 16678 762558
rect 17278 762486 18278 762558
rect 15748 762475 15782 762486
rect 15816 762475 15850 762486
rect 15884 762475 15918 762486
rect 15952 762475 15986 762486
rect 16020 762475 16054 762486
rect 16088 762475 16122 762486
rect 16156 762475 16190 762486
rect 16224 762475 16258 762486
rect 16292 762475 16326 762486
rect 16360 762475 16394 762486
rect 16428 762475 16462 762486
rect 16496 762475 16530 762486
rect 16564 762475 16598 762486
rect 16632 762475 16666 762486
rect 17290 762475 17324 762486
rect 17358 762475 17392 762486
rect 17426 762475 17460 762486
rect 17494 762475 17528 762486
rect 17562 762475 17596 762486
rect 17630 762475 17664 762486
rect 17698 762475 17732 762486
rect 17766 762475 17800 762486
rect 17834 762475 17868 762486
rect 17902 762475 17936 762486
rect 17970 762475 18004 762486
rect 18038 762475 18072 762486
rect 18106 762475 18140 762486
rect 18174 762475 18208 762486
rect 15748 762465 15806 762475
rect 15816 762465 15874 762475
rect 15884 762465 15942 762475
rect 15952 762465 16010 762475
rect 16020 762465 16078 762475
rect 16088 762465 16146 762475
rect 16156 762465 16214 762475
rect 16224 762465 16282 762475
rect 16292 762465 16350 762475
rect 16360 762465 16418 762475
rect 16428 762465 16486 762475
rect 16496 762465 16554 762475
rect 16564 762465 16622 762475
rect 16632 762465 16690 762475
rect 17290 762465 17348 762475
rect 17358 762465 17416 762475
rect 17426 762465 17484 762475
rect 17494 762465 17552 762475
rect 17562 762465 17620 762475
rect 17630 762465 17688 762475
rect 17698 762465 17756 762475
rect 17766 762465 17824 762475
rect 17834 762465 17892 762475
rect 17902 762465 17960 762475
rect 17970 762465 18028 762475
rect 18038 762465 18096 762475
rect 18106 762465 18164 762475
rect 18174 762465 18232 762475
rect 15724 762441 16690 762465
rect 17266 762441 18232 762465
rect 15748 762426 15772 762441
rect 15816 762426 15840 762441
rect 15884 762426 15908 762441
rect 15952 762426 15976 762441
rect 16020 762426 16044 762441
rect 16088 762426 16112 762441
rect 16156 762426 16180 762441
rect 16224 762426 16248 762441
rect 16292 762426 16316 762441
rect 16360 762426 16384 762441
rect 16428 762426 16452 762441
rect 16496 762426 16520 762441
rect 16564 762426 16588 762441
rect 16632 762426 16656 762441
rect 17290 762426 17314 762441
rect 17358 762426 17382 762441
rect 17426 762426 17450 762441
rect 17494 762426 17518 762441
rect 17562 762426 17586 762441
rect 17630 762426 17654 762441
rect 17698 762426 17722 762441
rect 17766 762426 17790 762441
rect 17834 762426 17858 762441
rect 17902 762426 17926 762441
rect 17970 762426 17994 762441
rect 18038 762426 18062 762441
rect 18106 762426 18130 762441
rect 18174 762426 18198 762441
rect 15678 762271 16678 762426
rect 7389 762181 8389 762241
rect 8990 762181 9990 762241
rect 15678 762237 16690 762271
rect 17278 762261 18278 762426
rect 17266 762237 18278 762261
rect 15678 762226 16678 762237
rect 17278 762226 18278 762237
rect 15748 762213 15772 762226
rect 15816 762213 15840 762226
rect 15884 762213 15908 762226
rect 15952 762213 15976 762226
rect 16020 762213 16044 762226
rect 16088 762213 16112 762226
rect 16156 762213 16180 762226
rect 16224 762213 16248 762226
rect 16292 762213 16316 762226
rect 16360 762213 16384 762226
rect 16428 762213 16452 762226
rect 16496 762213 16520 762226
rect 16564 762213 16588 762226
rect 16632 762213 16656 762226
rect 17290 762213 17314 762226
rect 17358 762213 17382 762226
rect 17426 762213 17450 762226
rect 17494 762213 17518 762226
rect 17562 762213 17586 762226
rect 17630 762213 17654 762226
rect 17698 762213 17722 762226
rect 17766 762213 17790 762226
rect 17834 762213 17858 762226
rect 17902 762213 17926 762226
rect 17970 762213 17994 762226
rect 18038 762213 18062 762226
rect 18106 762213 18130 762226
rect 18174 762213 18198 762226
rect 7389 761823 8389 761879
rect 8990 761823 9990 761879
rect 15678 761868 16678 761924
rect 17278 761868 18278 761924
rect 7389 761751 8389 761807
rect 8990 761751 9990 761807
rect 15678 761796 16678 761852
rect 17278 761796 18278 761852
rect 7389 761449 8389 761521
rect 8990 761449 9990 761521
rect 15678 761494 16678 761566
rect 17278 761494 18278 761566
rect 15748 761483 15782 761494
rect 15816 761483 15850 761494
rect 15884 761483 15918 761494
rect 15952 761483 15986 761494
rect 16020 761483 16054 761494
rect 16088 761483 16122 761494
rect 16156 761483 16190 761494
rect 16224 761483 16258 761494
rect 16292 761483 16326 761494
rect 16360 761483 16394 761494
rect 16428 761483 16462 761494
rect 16496 761483 16530 761494
rect 16564 761483 16598 761494
rect 16632 761483 16666 761494
rect 17290 761483 17324 761494
rect 17358 761483 17392 761494
rect 17426 761483 17460 761494
rect 17494 761483 17528 761494
rect 17562 761483 17596 761494
rect 17630 761483 17664 761494
rect 17698 761483 17732 761494
rect 17766 761483 17800 761494
rect 17834 761483 17868 761494
rect 17902 761483 17936 761494
rect 17970 761483 18004 761494
rect 18038 761483 18072 761494
rect 18106 761483 18140 761494
rect 18174 761483 18208 761494
rect 15748 761473 15806 761483
rect 15816 761473 15874 761483
rect 15884 761473 15942 761483
rect 15952 761473 16010 761483
rect 16020 761473 16078 761483
rect 16088 761473 16146 761483
rect 16156 761473 16214 761483
rect 16224 761473 16282 761483
rect 16292 761473 16350 761483
rect 16360 761473 16418 761483
rect 16428 761473 16486 761483
rect 16496 761473 16554 761483
rect 16564 761473 16622 761483
rect 16632 761473 16690 761483
rect 17290 761473 17348 761483
rect 17358 761473 17416 761483
rect 17426 761473 17484 761483
rect 17494 761473 17552 761483
rect 17562 761473 17620 761483
rect 17630 761473 17688 761483
rect 17698 761473 17756 761483
rect 17766 761473 17824 761483
rect 17834 761473 17892 761483
rect 17902 761473 17960 761483
rect 17970 761473 18028 761483
rect 18038 761473 18096 761483
rect 18106 761473 18164 761483
rect 18174 761473 18232 761483
rect 15724 761449 16690 761473
rect 17266 761449 18232 761473
rect 12427 761424 12493 761440
rect 15748 761434 15772 761449
rect 15816 761434 15840 761449
rect 15884 761434 15908 761449
rect 15952 761434 15976 761449
rect 16020 761434 16044 761449
rect 16088 761434 16112 761449
rect 16156 761434 16180 761449
rect 16224 761434 16248 761449
rect 16292 761434 16316 761449
rect 16360 761434 16384 761449
rect 16428 761434 16452 761449
rect 16496 761434 16520 761449
rect 16564 761434 16588 761449
rect 16632 761434 16656 761449
rect 17290 761434 17314 761449
rect 17358 761434 17382 761449
rect 17426 761434 17450 761449
rect 17494 761434 17518 761449
rect 17562 761434 17586 761449
rect 17630 761434 17654 761449
rect 17698 761434 17722 761449
rect 17766 761434 17790 761449
rect 17834 761434 17858 761449
rect 17902 761434 17926 761449
rect 17970 761434 17994 761449
rect 18038 761434 18062 761449
rect 18106 761434 18130 761449
rect 18174 761434 18198 761449
rect 15678 761279 16678 761434
rect 7389 761189 8389 761249
rect 8990 761189 9990 761249
rect 15678 761245 16690 761279
rect 17278 761269 18278 761434
rect 17266 761245 18278 761269
rect 15678 761234 16678 761245
rect 17278 761234 18278 761245
rect 15748 761221 15772 761234
rect 15816 761221 15840 761234
rect 15884 761221 15908 761234
rect 15952 761221 15976 761234
rect 16020 761221 16044 761234
rect 16088 761221 16112 761234
rect 16156 761221 16180 761234
rect 16224 761221 16248 761234
rect 16292 761221 16316 761234
rect 16360 761221 16384 761234
rect 16428 761221 16452 761234
rect 16496 761221 16520 761234
rect 16564 761221 16588 761234
rect 16632 761221 16656 761234
rect 17290 761221 17314 761234
rect 17358 761221 17382 761234
rect 17426 761221 17450 761234
rect 17494 761221 17518 761234
rect 17562 761221 17586 761234
rect 17630 761221 17654 761234
rect 17698 761221 17722 761234
rect 17766 761221 17790 761234
rect 17834 761221 17858 761234
rect 17902 761221 17926 761234
rect 17970 761221 17994 761234
rect 18038 761221 18062 761234
rect 18106 761221 18130 761234
rect 18174 761221 18198 761234
rect 7389 760831 8389 760887
rect 8990 760831 9990 760887
rect 15678 760876 16678 760932
rect 17278 760876 18278 760932
rect 7389 760759 8389 760815
rect 8990 760759 9990 760815
rect 15678 760804 16678 760860
rect 17278 760804 18278 760860
rect 7389 760457 8389 760529
rect 8990 760457 9990 760529
rect 15678 760502 16678 760574
rect 17278 760502 18278 760574
rect 15748 760491 15782 760502
rect 15816 760491 15850 760502
rect 15884 760491 15918 760502
rect 15952 760491 15986 760502
rect 16020 760491 16054 760502
rect 16088 760491 16122 760502
rect 16156 760491 16190 760502
rect 16224 760491 16258 760502
rect 16292 760491 16326 760502
rect 16360 760491 16394 760502
rect 16428 760491 16462 760502
rect 16496 760491 16530 760502
rect 16564 760491 16598 760502
rect 16632 760491 16666 760502
rect 17290 760491 17324 760502
rect 17358 760491 17392 760502
rect 17426 760491 17460 760502
rect 17494 760491 17528 760502
rect 17562 760491 17596 760502
rect 17630 760491 17664 760502
rect 17698 760491 17732 760502
rect 17766 760491 17800 760502
rect 17834 760491 17868 760502
rect 17902 760491 17936 760502
rect 17970 760491 18004 760502
rect 18038 760491 18072 760502
rect 18106 760491 18140 760502
rect 18174 760491 18208 760502
rect 15748 760481 15806 760491
rect 15816 760481 15874 760491
rect 15884 760481 15942 760491
rect 15952 760481 16010 760491
rect 16020 760481 16078 760491
rect 16088 760481 16146 760491
rect 16156 760481 16214 760491
rect 16224 760481 16282 760491
rect 16292 760481 16350 760491
rect 16360 760481 16418 760491
rect 16428 760481 16486 760491
rect 16496 760481 16554 760491
rect 16564 760481 16622 760491
rect 16632 760481 16690 760491
rect 17290 760481 17348 760491
rect 17358 760481 17416 760491
rect 17426 760481 17484 760491
rect 17494 760481 17552 760491
rect 17562 760481 17620 760491
rect 17630 760481 17688 760491
rect 17698 760481 17756 760491
rect 17766 760481 17824 760491
rect 17834 760481 17892 760491
rect 17902 760481 17960 760491
rect 17970 760481 18028 760491
rect 18038 760481 18096 760491
rect 18106 760481 18164 760491
rect 18174 760481 18232 760491
rect 15724 760457 16690 760481
rect 17266 760457 18232 760481
rect 15748 760442 15772 760457
rect 15816 760442 15840 760457
rect 15884 760442 15908 760457
rect 15952 760442 15976 760457
rect 16020 760442 16044 760457
rect 16088 760442 16112 760457
rect 16156 760442 16180 760457
rect 16224 760442 16248 760457
rect 16292 760442 16316 760457
rect 16360 760442 16384 760457
rect 16428 760442 16452 760457
rect 16496 760442 16520 760457
rect 16564 760442 16588 760457
rect 16632 760442 16656 760457
rect 17290 760442 17314 760457
rect 17358 760442 17382 760457
rect 17426 760442 17450 760457
rect 17494 760442 17518 760457
rect 17562 760442 17586 760457
rect 17630 760442 17654 760457
rect 17698 760442 17722 760457
rect 17766 760442 17790 760457
rect 17834 760442 17858 760457
rect 17902 760442 17926 760457
rect 17970 760442 17994 760457
rect 18038 760442 18062 760457
rect 18106 760442 18130 760457
rect 18174 760442 18198 760457
rect 15678 760287 16678 760442
rect 7389 760197 8389 760257
rect 8990 760197 9990 760257
rect 15678 760253 16690 760287
rect 17278 760277 18278 760442
rect 17266 760253 18278 760277
rect 15678 760242 16678 760253
rect 17278 760242 18278 760253
rect 15748 760229 15772 760242
rect 15816 760229 15840 760242
rect 15884 760229 15908 760242
rect 15952 760229 15976 760242
rect 16020 760229 16044 760242
rect 16088 760229 16112 760242
rect 16156 760229 16180 760242
rect 16224 760229 16248 760242
rect 16292 760229 16316 760242
rect 16360 760229 16384 760242
rect 16428 760229 16452 760242
rect 16496 760229 16520 760242
rect 16564 760229 16588 760242
rect 16632 760229 16656 760242
rect 17290 760229 17314 760242
rect 17358 760229 17382 760242
rect 17426 760229 17450 760242
rect 17494 760229 17518 760242
rect 17562 760229 17586 760242
rect 17630 760229 17654 760242
rect 17698 760229 17722 760242
rect 17766 760229 17790 760242
rect 17834 760229 17858 760242
rect 17902 760229 17926 760242
rect 17970 760229 17994 760242
rect 18038 760229 18062 760242
rect 18106 760229 18130 760242
rect 18174 760229 18198 760242
rect 7389 759839 8389 759895
rect 8990 759839 9990 759895
rect 15678 759884 16678 759940
rect 17278 759884 18278 759940
rect 7389 759767 8389 759823
rect 8990 759767 9990 759823
rect 15678 759812 16678 759868
rect 17278 759812 18278 759868
rect 7389 759465 8389 759537
rect 8990 759465 9990 759537
rect 15678 759510 16678 759582
rect 17278 759510 18278 759582
rect 15748 759499 15782 759510
rect 15816 759499 15850 759510
rect 15884 759499 15918 759510
rect 15952 759499 15986 759510
rect 16020 759499 16054 759510
rect 16088 759499 16122 759510
rect 16156 759499 16190 759510
rect 16224 759499 16258 759510
rect 16292 759499 16326 759510
rect 16360 759499 16394 759510
rect 16428 759499 16462 759510
rect 16496 759499 16530 759510
rect 16564 759499 16598 759510
rect 16632 759499 16666 759510
rect 17290 759499 17324 759510
rect 17358 759499 17392 759510
rect 17426 759499 17460 759510
rect 17494 759499 17528 759510
rect 17562 759499 17596 759510
rect 17630 759499 17664 759510
rect 17698 759499 17732 759510
rect 17766 759499 17800 759510
rect 17834 759499 17868 759510
rect 17902 759499 17936 759510
rect 17970 759499 18004 759510
rect 18038 759499 18072 759510
rect 18106 759499 18140 759510
rect 18174 759499 18208 759510
rect 15748 759489 15806 759499
rect 15816 759489 15874 759499
rect 15884 759489 15942 759499
rect 15952 759489 16010 759499
rect 16020 759489 16078 759499
rect 16088 759489 16146 759499
rect 16156 759489 16214 759499
rect 16224 759489 16282 759499
rect 16292 759489 16350 759499
rect 16360 759489 16418 759499
rect 16428 759489 16486 759499
rect 16496 759489 16554 759499
rect 16564 759489 16622 759499
rect 16632 759489 16690 759499
rect 17290 759489 17348 759499
rect 17358 759489 17416 759499
rect 17426 759489 17484 759499
rect 17494 759489 17552 759499
rect 17562 759489 17620 759499
rect 17630 759489 17688 759499
rect 17698 759489 17756 759499
rect 17766 759489 17824 759499
rect 17834 759489 17892 759499
rect 17902 759489 17960 759499
rect 17970 759489 18028 759499
rect 18038 759489 18096 759499
rect 18106 759489 18164 759499
rect 18174 759489 18232 759499
rect 15724 759465 16690 759489
rect 17266 759465 18232 759489
rect 15748 759450 15772 759465
rect 15816 759450 15840 759465
rect 15884 759450 15908 759465
rect 15952 759450 15976 759465
rect 16020 759450 16044 759465
rect 16088 759450 16112 759465
rect 16156 759450 16180 759465
rect 16224 759450 16248 759465
rect 16292 759450 16316 759465
rect 16360 759450 16384 759465
rect 16428 759450 16452 759465
rect 16496 759450 16520 759465
rect 16564 759450 16588 759465
rect 16632 759450 16656 759465
rect 17290 759450 17314 759465
rect 17358 759450 17382 759465
rect 17426 759450 17450 759465
rect 17494 759450 17518 759465
rect 17562 759450 17586 759465
rect 17630 759450 17654 759465
rect 17698 759450 17722 759465
rect 17766 759450 17790 759465
rect 17834 759450 17858 759465
rect 17902 759450 17926 759465
rect 17970 759450 17994 759465
rect 18038 759450 18062 759465
rect 18106 759450 18130 759465
rect 18174 759450 18198 759465
rect 15678 759295 16678 759450
rect 7389 759205 8389 759265
rect 8990 759205 9990 759265
rect 15678 759261 16690 759295
rect 17278 759285 18278 759450
rect 17266 759261 18278 759285
rect 15678 759250 16678 759261
rect 17278 759250 18278 759261
rect 15748 759237 15772 759250
rect 15816 759237 15840 759250
rect 15884 759237 15908 759250
rect 15952 759237 15976 759250
rect 16020 759237 16044 759250
rect 16088 759237 16112 759250
rect 16156 759237 16180 759250
rect 16224 759237 16248 759250
rect 16292 759237 16316 759250
rect 16360 759237 16384 759250
rect 16428 759237 16452 759250
rect 16496 759237 16520 759250
rect 16564 759237 16588 759250
rect 16632 759237 16656 759250
rect 17290 759237 17314 759250
rect 17358 759237 17382 759250
rect 17426 759237 17450 759250
rect 17494 759237 17518 759250
rect 17562 759237 17586 759250
rect 17630 759237 17654 759250
rect 17698 759237 17722 759250
rect 17766 759237 17790 759250
rect 17834 759237 17858 759250
rect 17902 759237 17926 759250
rect 17970 759237 17994 759250
rect 18038 759237 18062 759250
rect 18106 759237 18130 759250
rect 18174 759237 18198 759250
rect 7389 758847 8389 758903
rect 8990 758847 9990 758903
rect 15678 758892 16678 758948
rect 17278 758892 18278 758948
rect 7389 758775 8389 758831
rect 8990 758775 9990 758831
rect 15678 758820 16678 758876
rect 17278 758820 18278 758876
rect 5967 758455 6059 758489
rect 7389 758473 8389 758545
rect 8990 758473 9990 758545
rect 15678 758518 16678 758590
rect 17278 758518 18278 758590
rect 15748 758507 15782 758518
rect 15816 758507 15850 758518
rect 15884 758507 15918 758518
rect 15952 758507 15986 758518
rect 16020 758507 16054 758518
rect 16088 758507 16122 758518
rect 16156 758507 16190 758518
rect 16224 758507 16258 758518
rect 16292 758507 16326 758518
rect 16360 758507 16394 758518
rect 16428 758507 16462 758518
rect 16496 758507 16530 758518
rect 16564 758507 16598 758518
rect 16632 758507 16666 758518
rect 17290 758507 17324 758518
rect 17358 758507 17392 758518
rect 17426 758507 17460 758518
rect 17494 758507 17528 758518
rect 17562 758507 17596 758518
rect 17630 758507 17664 758518
rect 17698 758507 17732 758518
rect 17766 758507 17800 758518
rect 17834 758507 17868 758518
rect 17902 758507 17936 758518
rect 17970 758507 18004 758518
rect 18038 758507 18072 758518
rect 18106 758507 18140 758518
rect 18174 758507 18208 758518
rect 15748 758497 15806 758507
rect 15816 758497 15874 758507
rect 15884 758497 15942 758507
rect 15952 758497 16010 758507
rect 16020 758497 16078 758507
rect 16088 758497 16146 758507
rect 16156 758497 16214 758507
rect 16224 758497 16282 758507
rect 16292 758497 16350 758507
rect 16360 758497 16418 758507
rect 16428 758497 16486 758507
rect 16496 758497 16554 758507
rect 16564 758497 16622 758507
rect 16632 758497 16690 758507
rect 17290 758497 17348 758507
rect 17358 758497 17416 758507
rect 17426 758497 17484 758507
rect 17494 758497 17552 758507
rect 17562 758497 17620 758507
rect 17630 758497 17688 758507
rect 17698 758497 17756 758507
rect 17766 758497 17824 758507
rect 17834 758497 17892 758507
rect 17902 758497 17960 758507
rect 17970 758497 18028 758507
rect 18038 758497 18096 758507
rect 18106 758497 18164 758507
rect 18174 758497 18232 758507
rect 15724 758473 16690 758497
rect 17266 758473 18232 758497
rect 15748 758458 15772 758473
rect 15816 758458 15840 758473
rect 15884 758458 15908 758473
rect 15952 758458 15976 758473
rect 16020 758458 16044 758473
rect 16088 758458 16112 758473
rect 16156 758458 16180 758473
rect 16224 758458 16248 758473
rect 16292 758458 16316 758473
rect 16360 758458 16384 758473
rect 16428 758458 16452 758473
rect 16496 758458 16520 758473
rect 16564 758458 16588 758473
rect 16632 758458 16656 758473
rect 17290 758458 17314 758473
rect 17358 758458 17382 758473
rect 17426 758458 17450 758473
rect 17494 758458 17518 758473
rect 17562 758458 17586 758473
rect 17630 758458 17654 758473
rect 17698 758458 17722 758473
rect 17766 758458 17790 758473
rect 17834 758458 17858 758473
rect 17902 758458 17926 758473
rect 17970 758458 17994 758473
rect 18038 758458 18062 758473
rect 18106 758458 18130 758473
rect 18174 758458 18198 758473
rect 2850 758398 3850 758448
rect 2850 758282 3850 758332
rect 2850 758072 3850 758122
rect 2850 757956 3850 758006
rect 2850 757746 3850 757796
rect 1153 757660 1187 757718
rect 2850 757630 3850 757680
rect 2850 757420 3850 757470
rect 2850 757417 3107 757420
rect 3250 757304 3850 757354
rect 3250 757048 3850 757104
rect 3250 756892 3850 757020
rect 175 756818 1175 756868
rect 175 756662 1175 756790
rect 3250 756736 3850 756792
rect 175 756506 1175 756634
rect 175 756350 1175 756478
rect 175 756194 1175 756322
rect 175 756044 1175 756094
rect 175 755928 1175 755978
rect 175 755772 1175 755828
rect 175 755622 1175 755672
rect 1578 755609 1628 756609
rect 1728 755609 1856 756609
rect 1884 755609 2012 756609
rect 2040 755609 2090 756609
rect 3250 756580 3850 756708
rect 3250 756430 3850 756480
rect 2850 756314 3850 756364
rect 2850 756158 3850 756214
rect 2850 756008 3850 756058
rect 2850 755880 3850 755930
rect 2850 755724 3850 755852
rect 2850 755568 3850 755696
rect 175 755506 1175 755556
rect 175 755350 1175 755478
rect 2850 755412 3850 755468
rect 2850 755256 3850 755384
rect 175 755194 1175 755250
rect 175 755038 1175 755166
rect 175 754888 1175 754938
rect 175 754772 1175 754822
rect 175 754616 1175 754744
rect 1578 754613 1628 755213
rect 1728 754613 1784 755213
rect 1884 754613 1940 755213
rect 2040 754613 2096 755213
rect 2196 754613 2246 755213
rect 2850 755100 3850 755228
rect 2850 754944 3850 755072
rect 2850 754794 3850 754844
rect 2850 754678 3850 754728
rect 2850 754522 3850 754650
rect 175 754460 1175 754516
rect 175 754304 1175 754432
rect 2850 754366 3850 754494
rect 2850 754210 3850 754338
rect 175 754154 1175 754204
rect 803 754151 1175 754154
rect 2850 754054 3850 754110
rect 2850 753898 3850 754026
rect 2850 753742 3850 753870
rect 2850 753586 3850 753642
rect 2850 753436 3850 753486
rect 3926 753455 3960 753491
rect 3967 753339 3989 753455
rect 1638 751869 1688 752869
rect 1848 751869 1976 752869
rect 2064 751869 2114 752869
rect 2850 752275 3050 752287
rect 2850 752162 3850 752212
rect 2850 751946 3850 752074
rect 2850 751730 3850 751786
rect 2850 751514 3850 751642
rect 2850 751304 3850 751354
rect 2850 751188 3850 751238
rect 2850 750978 3850 751028
rect 3926 751015 3960 753339
rect 5169 751315 5191 758429
rect 5488 757194 5538 758194
rect 5658 757194 5708 758194
rect 5488 756073 5538 757073
rect 5658 756073 5708 757073
rect 5488 754952 5538 755952
rect 5658 754952 5708 755952
rect 5488 753842 5538 754842
rect 5658 753842 5708 754842
rect 5488 752721 5538 753721
rect 5658 752721 5708 753721
rect 5488 751600 5538 752600
rect 5658 751600 5708 752600
rect 5971 751386 6059 758455
rect 15678 758303 16678 758458
rect 7389 758213 8389 758273
rect 8990 758213 9990 758273
rect 15678 758269 16690 758303
rect 17278 758293 18278 758458
rect 17266 758269 18278 758293
rect 15678 758258 16678 758269
rect 17278 758258 18278 758269
rect 15748 758245 15772 758258
rect 15816 758245 15840 758258
rect 15884 758245 15908 758258
rect 15952 758245 15976 758258
rect 16020 758245 16044 758258
rect 16088 758245 16112 758258
rect 16156 758245 16180 758258
rect 16224 758245 16248 758258
rect 16292 758245 16316 758258
rect 16360 758245 16384 758258
rect 16428 758245 16452 758258
rect 16496 758245 16520 758258
rect 16564 758245 16588 758258
rect 16632 758245 16656 758258
rect 17290 758245 17314 758258
rect 17358 758245 17382 758258
rect 17426 758245 17450 758258
rect 17494 758245 17518 758258
rect 17562 758245 17586 758258
rect 17630 758245 17654 758258
rect 17698 758245 17722 758258
rect 17766 758245 17790 758258
rect 17834 758245 17858 758258
rect 17902 758245 17926 758258
rect 17970 758245 17994 758258
rect 18038 758245 18062 758258
rect 18106 758245 18130 758258
rect 18174 758245 18198 758258
rect 7389 757855 8389 757911
rect 8990 757855 9990 757911
rect 15678 757900 16678 757956
rect 17278 757900 18278 757956
rect 7389 757783 8389 757839
rect 8990 757783 9990 757839
rect 15678 757828 16678 757884
rect 17278 757828 18278 757884
rect 7389 757481 8389 757553
rect 8990 757481 9990 757553
rect 15678 757526 16678 757598
rect 17278 757526 18278 757598
rect 15748 757515 15782 757526
rect 15816 757515 15850 757526
rect 15884 757515 15918 757526
rect 15952 757515 15986 757526
rect 16020 757515 16054 757526
rect 16088 757515 16122 757526
rect 16156 757515 16190 757526
rect 16224 757515 16258 757526
rect 16292 757515 16326 757526
rect 16360 757515 16394 757526
rect 16428 757515 16462 757526
rect 16496 757515 16530 757526
rect 16564 757515 16598 757526
rect 16632 757515 16666 757526
rect 17290 757515 17324 757526
rect 17358 757515 17392 757526
rect 17426 757515 17460 757526
rect 17494 757515 17528 757526
rect 17562 757515 17596 757526
rect 17630 757515 17664 757526
rect 17698 757515 17732 757526
rect 17766 757515 17800 757526
rect 17834 757515 17868 757526
rect 17902 757515 17936 757526
rect 17970 757515 18004 757526
rect 18038 757515 18072 757526
rect 18106 757515 18140 757526
rect 18174 757515 18208 757526
rect 15748 757505 15806 757515
rect 15816 757505 15874 757515
rect 15884 757505 15942 757515
rect 15952 757505 16010 757515
rect 16020 757505 16078 757515
rect 16088 757505 16146 757515
rect 16156 757505 16214 757515
rect 16224 757505 16282 757515
rect 16292 757505 16350 757515
rect 16360 757505 16418 757515
rect 16428 757505 16486 757515
rect 16496 757505 16554 757515
rect 16564 757505 16622 757515
rect 16632 757505 16690 757515
rect 17290 757505 17348 757515
rect 17358 757505 17416 757515
rect 17426 757505 17484 757515
rect 17494 757505 17552 757515
rect 17562 757505 17620 757515
rect 17630 757505 17688 757515
rect 17698 757505 17756 757515
rect 17766 757505 17824 757515
rect 17834 757505 17892 757515
rect 17902 757505 17960 757515
rect 17970 757505 18028 757515
rect 18038 757505 18096 757515
rect 18106 757505 18164 757515
rect 18174 757505 18232 757515
rect 15724 757481 16690 757505
rect 17266 757481 18232 757505
rect 15748 757466 15772 757481
rect 15816 757466 15840 757481
rect 15884 757466 15908 757481
rect 15952 757466 15976 757481
rect 16020 757466 16044 757481
rect 16088 757466 16112 757481
rect 16156 757466 16180 757481
rect 16224 757466 16248 757481
rect 16292 757466 16316 757481
rect 16360 757466 16384 757481
rect 16428 757466 16452 757481
rect 16496 757466 16520 757481
rect 16564 757466 16588 757481
rect 16632 757466 16656 757481
rect 17290 757466 17314 757481
rect 17358 757466 17382 757481
rect 17426 757466 17450 757481
rect 17494 757466 17518 757481
rect 17562 757466 17586 757481
rect 17630 757466 17654 757481
rect 17698 757466 17722 757481
rect 17766 757466 17790 757481
rect 17834 757466 17858 757481
rect 17902 757466 17926 757481
rect 17970 757466 17994 757481
rect 18038 757466 18062 757481
rect 18106 757466 18130 757481
rect 18174 757466 18198 757481
rect 15678 757311 16678 757466
rect 7389 757221 8389 757281
rect 8990 757221 9990 757281
rect 15678 757277 16690 757311
rect 17278 757301 18278 757466
rect 17266 757277 18278 757301
rect 15678 757266 16678 757277
rect 17278 757266 18278 757277
rect 15748 757253 15772 757266
rect 15816 757253 15840 757266
rect 15884 757253 15908 757266
rect 15952 757253 15976 757266
rect 16020 757253 16044 757266
rect 16088 757253 16112 757266
rect 16156 757253 16180 757266
rect 16224 757253 16248 757266
rect 16292 757253 16316 757266
rect 16360 757253 16384 757266
rect 16428 757253 16452 757266
rect 16496 757253 16520 757266
rect 16564 757253 16588 757266
rect 16632 757253 16656 757266
rect 17290 757253 17314 757266
rect 17358 757253 17382 757266
rect 17426 757253 17450 757266
rect 17494 757253 17518 757266
rect 17562 757253 17586 757266
rect 17630 757253 17654 757266
rect 17698 757253 17722 757266
rect 17766 757253 17790 757266
rect 17834 757253 17858 757266
rect 17902 757253 17926 757266
rect 17970 757253 17994 757266
rect 18038 757253 18062 757266
rect 18106 757253 18130 757266
rect 18174 757253 18198 757266
rect 7389 756863 8389 756919
rect 8990 756863 9990 756919
rect 15678 756908 16678 756964
rect 17278 756908 18278 756964
rect 7389 756791 8389 756847
rect 8990 756791 9990 756847
rect 15678 756836 16678 756892
rect 17278 756836 18278 756892
rect 19480 756867 19516 763817
rect 19547 756867 19583 763817
rect 24572 763738 25172 763866
rect 36785 763864 37385 763920
rect 36785 763688 37385 763744
rect 20809 763650 20833 763684
rect 20809 763582 20833 763616
rect 24572 763588 25172 763638
rect 20809 763514 20833 763548
rect 36785 763518 37385 763568
rect 20809 763446 20833 763480
rect 24572 763458 25172 763508
rect 32930 763457 33530 763507
rect 20809 763378 20833 763412
rect 35287 763391 35887 763441
rect 36785 763402 37385 763452
rect 20809 763310 20833 763344
rect 24572 763308 25172 763358
rect 31463 763307 32063 763357
rect 32930 763301 33530 763357
rect 20809 763242 20833 763276
rect 35287 763215 35887 763343
rect 36785 763226 37385 763282
rect 20809 763174 20833 763208
rect 31463 763151 32063 763207
rect 32930 763151 33530 763201
rect 34079 763157 34679 763207
rect 20809 763106 20833 763140
rect 19844 762051 19894 763051
rect 19994 762051 20122 763051
rect 20150 762051 20278 763051
rect 20306 762051 20434 763051
rect 20462 762051 20512 763051
rect 20809 763038 20833 763072
rect 20809 762970 20833 763004
rect 20973 763000 21007 763024
rect 21041 763000 21075 763024
rect 21109 763000 21143 763024
rect 21177 763000 21211 763024
rect 21245 763000 21279 763024
rect 21313 763000 21347 763024
rect 21381 763000 21415 763024
rect 21449 763000 21483 763024
rect 21517 763000 21551 763024
rect 21585 763000 21619 763024
rect 21653 763000 21687 763024
rect 21721 763000 21755 763024
rect 21789 763000 21823 763024
rect 21857 763000 21891 763024
rect 21925 763000 21959 763024
rect 21993 763000 22027 763024
rect 22061 763000 22095 763024
rect 22129 763000 22163 763024
rect 22197 763000 22210 763024
rect 31463 763001 32063 763051
rect 34079 763001 34679 763057
rect 35287 763039 35887 763095
rect 36785 763050 37385 763106
rect 20809 762902 20833 762936
rect 32596 762929 33596 762979
rect 20809 762834 20833 762868
rect 24573 762820 25173 762870
rect 34079 762851 34679 762901
rect 35287 762869 35887 762919
rect 36785 762880 37385 762930
rect 35287 762866 35559 762869
rect 35716 762866 35887 762869
rect 20809 762766 20833 762800
rect 30171 762795 30771 762845
rect 20809 762698 20833 762732
rect 24573 762664 25173 762792
rect 32596 762773 33596 762829
rect 37993 762704 38593 762754
rect 19844 760521 19894 761921
rect 19994 760521 20122 761921
rect 20150 760521 20278 761921
rect 20306 760521 20434 761921
rect 20462 760521 20512 761921
rect 20809 760219 20833 760253
rect 19844 758759 19894 760159
rect 19994 758759 20122 760159
rect 20150 758759 20278 760159
rect 20306 758759 20434 760159
rect 20462 758759 20512 760159
rect 20809 760151 20833 760185
rect 20809 760083 20833 760117
rect 20809 760015 20833 760049
rect 20809 759947 20833 759981
rect 20809 759879 20833 759913
rect 20809 759811 20833 759845
rect 20809 759743 20833 759777
rect 20809 759675 20833 759709
rect 20809 759607 20833 759641
rect 20809 759539 20833 759573
rect 21263 759518 21313 762518
rect 21413 759518 21541 762518
rect 21569 759518 21697 762518
rect 21725 759518 21853 762518
rect 21881 759518 22009 762518
rect 22037 759518 22165 762518
rect 22193 759518 22321 762518
rect 22349 759518 22399 762518
rect 24573 762508 25173 762636
rect 30171 762619 30771 762675
rect 32596 762623 33596 762673
rect 34110 762589 34710 762639
rect 36785 762620 36797 762624
rect 36785 762609 36800 762620
rect 36970 762609 36985 762624
rect 26348 762530 26372 762564
rect 32596 762507 33596 762557
rect 26348 762461 26372 762495
rect 30171 762449 30771 762499
rect 24573 762352 25173 762408
rect 24573 762196 25173 762324
rect 29993 762310 30993 762360
rect 32596 762351 33596 762479
rect 34110 762433 34710 762561
rect 36785 762429 36985 762609
rect 37993 762534 38593 762584
rect 36785 762418 36800 762429
rect 36785 762414 36797 762418
rect 36970 762414 36985 762429
rect 31347 762317 31362 762332
rect 31535 762328 31547 762332
rect 31532 762317 31547 762328
rect 24573 762040 25173 762168
rect 26490 762122 26690 762172
rect 29993 762160 30993 762210
rect 31347 762137 31547 762317
rect 31347 762122 31362 762137
rect 31532 762126 31547 762137
rect 31535 762122 31547 762126
rect 31607 762317 31622 762332
rect 31795 762328 31807 762332
rect 31792 762317 31807 762328
rect 31607 762137 31807 762317
rect 32596 762195 33596 762323
rect 34110 762277 34710 762405
rect 36785 762384 36797 762388
rect 36785 762373 36800 762384
rect 36970 762373 36985 762388
rect 31607 762122 31622 762137
rect 31792 762126 31807 762137
rect 31795 762122 31807 762126
rect 31347 762081 31362 762096
rect 31535 762092 31547 762096
rect 31532 762081 31547 762092
rect 22906 761855 23212 762025
rect 23406 761855 23712 762025
rect 26490 761966 26690 762022
rect 29993 762001 30993 762051
rect 24573 761890 25173 761940
rect 31347 761901 31547 762081
rect 26490 761816 26690 761866
rect 29993 761851 30993 761901
rect 31347 761886 31362 761901
rect 31532 761890 31547 761901
rect 31535 761886 31547 761890
rect 31607 762081 31622 762096
rect 31795 762092 31807 762096
rect 31792 762081 31807 762092
rect 31607 761901 31807 762081
rect 32596 762039 33596 762167
rect 34110 762121 34710 762249
rect 36785 762193 36985 762373
rect 36785 762182 36800 762193
rect 36785 762178 36797 762182
rect 36970 762178 36985 762193
rect 37083 762373 37098 762388
rect 37083 762193 37120 762373
rect 37083 762178 37098 762193
rect 37998 762108 38598 762158
rect 34110 761971 34710 762021
rect 31607 761886 31622 761901
rect 31792 761890 31807 761901
rect 31795 761886 31807 761890
rect 32596 761883 33596 761939
rect 37998 761932 38598 761988
rect 34110 761855 34710 761905
rect 24573 761760 25173 761810
rect 27691 761682 28291 761732
rect 30253 761721 30268 761736
rect 30441 761732 30453 761736
rect 30438 761721 30453 761732
rect 24573 761610 25173 761660
rect 27691 761532 28291 761582
rect 30253 761541 30453 761721
rect 30253 761526 30268 761541
rect 30438 761530 30453 761541
rect 30441 761526 30453 761530
rect 30513 761721 30528 761736
rect 30701 761732 30713 761736
rect 30698 761721 30713 761732
rect 30513 761541 30713 761721
rect 30513 761526 30528 761541
rect 30698 761530 30713 761541
rect 30701 761526 30713 761530
rect 30773 761721 30788 761736
rect 30961 761732 30973 761736
rect 30958 761721 30973 761732
rect 30773 761541 30973 761721
rect 30773 761526 30788 761541
rect 30958 761530 30973 761541
rect 30961 761526 30973 761530
rect 31087 761721 31102 761736
rect 31275 761732 31287 761736
rect 31272 761721 31287 761732
rect 31087 761541 31287 761721
rect 31087 761526 31102 761541
rect 31272 761530 31287 761541
rect 31275 761526 31287 761530
rect 31347 761721 31362 761736
rect 31535 761732 31547 761736
rect 31532 761721 31547 761732
rect 31347 761541 31547 761721
rect 31347 761526 31362 761541
rect 31532 761530 31547 761541
rect 31535 761526 31547 761530
rect 31607 761721 31622 761736
rect 31795 761732 31807 761736
rect 31792 761721 31807 761732
rect 31607 761541 31807 761721
rect 31607 761526 31622 761541
rect 31792 761530 31807 761541
rect 31795 761526 31807 761530
rect 31867 761721 31882 761736
rect 32055 761732 32067 761736
rect 32052 761721 32067 761732
rect 32596 761727 33596 761855
rect 31867 761541 32067 761721
rect 34110 761699 34710 761827
rect 37998 761762 38598 761812
rect 37998 761759 38220 761762
rect 38245 761759 38539 761762
rect 32596 761571 33596 761699
rect 34110 761543 34710 761671
rect 31867 761526 31882 761541
rect 32052 761530 32067 761541
rect 32055 761526 32067 761530
rect 22619 761446 22647 761474
rect 24573 761438 25173 761488
rect 26490 761416 26690 761466
rect 27691 761402 28291 761452
rect 32596 761415 33596 761543
rect 34110 761387 34710 761515
rect 24573 761288 25173 761338
rect 26490 761260 26690 761316
rect 27691 761246 28291 761374
rect 30253 761361 30268 761376
rect 30441 761372 30453 761376
rect 30438 761361 30453 761372
rect 30253 761331 30453 761361
rect 30253 761316 30268 761331
rect 30438 761320 30453 761331
rect 30441 761316 30453 761320
rect 30513 761361 30528 761376
rect 30701 761372 30713 761376
rect 30698 761361 30713 761372
rect 30513 761331 30713 761361
rect 30513 761316 30528 761331
rect 30698 761320 30713 761331
rect 30701 761316 30713 761320
rect 30773 761361 30788 761376
rect 31347 761361 31362 761376
rect 31535 761372 31547 761376
rect 31532 761361 31547 761372
rect 30773 761331 30793 761361
rect 31347 761331 31547 761361
rect 30773 761316 30788 761331
rect 31347 761316 31362 761331
rect 31532 761320 31547 761331
rect 31535 761316 31547 761320
rect 31607 761361 31622 761376
rect 31795 761372 31807 761376
rect 31792 761361 31807 761372
rect 31607 761331 31807 761361
rect 31607 761316 31622 761331
rect 31792 761320 31807 761331
rect 31795 761316 31807 761320
rect 31867 761361 31882 761376
rect 31867 761331 31921 761361
rect 31867 761316 31882 761331
rect 30253 761275 30268 761290
rect 30441 761286 30453 761290
rect 30438 761275 30453 761286
rect 30253 761245 30453 761275
rect 30253 761230 30268 761245
rect 30438 761234 30453 761245
rect 30441 761230 30453 761234
rect 30513 761275 30528 761290
rect 30701 761286 30713 761290
rect 30698 761275 30713 761286
rect 30513 761245 30713 761275
rect 30513 761230 30528 761245
rect 30698 761234 30713 761245
rect 30701 761230 30713 761234
rect 30773 761275 30788 761290
rect 31347 761275 31362 761290
rect 31535 761286 31547 761290
rect 31532 761275 31547 761286
rect 30773 761245 30793 761275
rect 31347 761245 31547 761275
rect 30773 761230 30788 761245
rect 31347 761230 31362 761245
rect 31532 761234 31547 761245
rect 31535 761230 31547 761234
rect 31607 761275 31622 761290
rect 31795 761286 31807 761290
rect 31792 761275 31807 761286
rect 31607 761245 31807 761275
rect 31607 761230 31622 761245
rect 31792 761234 31807 761245
rect 31795 761230 31807 761234
rect 31867 761275 31882 761290
rect 31867 761245 31921 761275
rect 32596 761265 33596 761315
rect 31867 761230 31882 761245
rect 34110 761231 34710 761287
rect 22906 761055 23212 761225
rect 23406 761055 23712 761225
rect 24573 761158 25173 761208
rect 24573 761002 25173 761130
rect 26490 761107 26690 761160
rect 27691 761090 28291 761218
rect 31823 761084 32061 761118
rect 31481 761080 32061 761084
rect 31481 761068 31797 761080
rect 32596 761063 33596 761113
rect 34110 761075 34710 761203
rect 37998 761133 38148 761145
rect 38317 761133 38467 761145
rect 24573 760846 25173 760974
rect 27691 760934 28291 760990
rect 32596 760907 33596 761035
rect 34110 760919 34710 761047
rect 37998 761020 38598 761070
rect 27691 760778 28291 760906
rect 25286 760758 25310 760762
rect 32596 760751 33596 760879
rect 34110 760763 34710 760891
rect 37998 760844 38598 760900
rect 24573 760690 25173 760746
rect 25286 760687 25310 760721
rect 24573 760534 25173 760662
rect 25286 760615 25310 760649
rect 27691 760622 28291 760750
rect 32596 760595 33596 760723
rect 35287 760695 35487 760707
rect 37998 760674 38598 760724
rect 34110 760607 34710 760663
rect 36785 760650 36797 760654
rect 36785 760639 36800 760650
rect 36970 760639 36985 760654
rect 35134 760582 35734 760632
rect 25286 760543 25310 760577
rect 22906 760255 23212 760425
rect 23406 760255 23712 760425
rect 24573 760378 25173 760506
rect 25286 760471 25310 760505
rect 27691 760472 28291 760522
rect 32596 760439 33596 760567
rect 34110 760451 34710 760507
rect 35134 760432 35734 760482
rect 36785 760459 36985 760639
rect 36785 760448 36800 760459
rect 36785 760444 36797 760448
rect 36970 760444 36985 760459
rect 37083 760639 37098 760654
rect 37083 760459 37120 760639
rect 37083 760444 37098 760459
rect 36785 760414 36797 760418
rect 32596 760283 33596 760411
rect 36785 760403 36800 760414
rect 36970 760403 36985 760418
rect 34110 760295 34710 760351
rect 35134 760316 35734 760366
rect 24573 760228 25173 760278
rect 32596 760127 33596 760255
rect 34110 760145 34710 760195
rect 35134 760160 35734 760288
rect 32596 759971 33596 760099
rect 34110 760029 34710 760079
rect 35134 760004 35734 760132
rect 31481 759862 31797 759880
rect 34110 759873 34710 760001
rect 31823 759828 32061 759860
rect 32596 759821 33596 759871
rect 35134 759848 35734 759976
rect 36071 759805 36098 760295
rect 36785 760223 36985 760403
rect 37993 760248 38593 760298
rect 36785 760212 36800 760223
rect 36785 760208 36797 760212
rect 36970 760208 36985 760223
rect 37993 760078 38593 760128
rect 36785 759902 37385 759952
rect 34110 759717 34710 759773
rect 30253 759701 30268 759716
rect 30441 759712 30453 759716
rect 30438 759701 30453 759712
rect 30253 759671 30453 759701
rect 30253 759656 30268 759671
rect 30438 759660 30453 759671
rect 30441 759656 30453 759660
rect 30513 759701 30528 759716
rect 30701 759712 30713 759716
rect 30698 759701 30713 759712
rect 30513 759671 30713 759701
rect 30513 759656 30528 759671
rect 30698 759660 30713 759671
rect 30701 759656 30713 759660
rect 30773 759701 30788 759716
rect 31347 759701 31362 759716
rect 31535 759712 31547 759716
rect 31532 759701 31547 759712
rect 30773 759671 30793 759701
rect 31347 759671 31547 759701
rect 30773 759656 30788 759671
rect 31347 759656 31362 759671
rect 31532 759660 31547 759671
rect 31535 759656 31547 759660
rect 31607 759701 31622 759716
rect 31795 759712 31807 759716
rect 31792 759701 31807 759712
rect 31607 759671 31807 759701
rect 31607 759656 31622 759671
rect 31792 759660 31807 759671
rect 31795 759656 31807 759660
rect 31867 759701 31882 759716
rect 31867 759671 31921 759701
rect 35134 759698 35734 759770
rect 36785 759726 37385 759782
rect 31867 759656 31882 759671
rect 30253 759615 30268 759630
rect 30441 759626 30453 759630
rect 30438 759615 30453 759626
rect 30253 759585 30453 759615
rect 30253 759570 30268 759585
rect 30438 759574 30453 759585
rect 30441 759570 30453 759574
rect 30513 759615 30528 759630
rect 30701 759626 30713 759630
rect 30698 759615 30713 759626
rect 30513 759585 30713 759615
rect 30513 759570 30528 759585
rect 30698 759574 30713 759585
rect 30701 759570 30713 759574
rect 30773 759615 30788 759630
rect 31347 759615 31362 759630
rect 31535 759626 31547 759630
rect 31532 759615 31547 759626
rect 30773 759585 30793 759615
rect 31347 759585 31547 759615
rect 30773 759570 30788 759585
rect 31347 759570 31362 759585
rect 31532 759574 31547 759585
rect 31535 759570 31547 759574
rect 31607 759615 31622 759630
rect 31795 759626 31807 759630
rect 31792 759615 31807 759626
rect 31607 759585 31807 759615
rect 31607 759570 31622 759585
rect 31792 759574 31807 759585
rect 31795 759570 31807 759574
rect 31867 759615 31882 759630
rect 32546 759619 33546 759669
rect 31867 759585 31921 759615
rect 31867 759570 31882 759585
rect 20809 759471 20833 759505
rect 32546 759463 33546 759591
rect 34110 759561 34710 759689
rect 35134 759645 36134 759695
rect 35134 759489 36134 759617
rect 36785 759550 37385 759606
rect 20809 759403 20833 759437
rect 30253 759405 30268 759420
rect 30441 759416 30453 759420
rect 30438 759405 30453 759416
rect 20809 759335 20833 759369
rect 20809 759267 20833 759301
rect 20809 759199 20833 759233
rect 30253 759225 30453 759405
rect 30253 759210 30268 759225
rect 30438 759214 30453 759225
rect 30441 759210 30453 759214
rect 30513 759405 30528 759420
rect 30701 759416 30713 759420
rect 30698 759405 30713 759416
rect 30513 759225 30713 759405
rect 30513 759210 30528 759225
rect 30698 759214 30713 759225
rect 30701 759210 30713 759214
rect 30773 759405 30788 759420
rect 30961 759416 30973 759420
rect 30958 759405 30973 759416
rect 30773 759225 30973 759405
rect 30773 759210 30788 759225
rect 30958 759214 30973 759225
rect 30961 759210 30973 759214
rect 31087 759405 31102 759420
rect 31275 759416 31287 759420
rect 31272 759405 31287 759416
rect 31087 759225 31287 759405
rect 31087 759210 31102 759225
rect 31272 759214 31287 759225
rect 31275 759210 31287 759214
rect 31347 759405 31362 759420
rect 31535 759416 31547 759420
rect 31532 759405 31547 759416
rect 31347 759225 31547 759405
rect 31347 759210 31362 759225
rect 31532 759214 31547 759225
rect 31535 759210 31547 759214
rect 31607 759405 31622 759420
rect 31795 759416 31807 759420
rect 31792 759405 31807 759416
rect 31607 759225 31807 759405
rect 31607 759210 31622 759225
rect 31792 759214 31807 759225
rect 31795 759210 31807 759214
rect 31867 759405 31882 759420
rect 32055 759416 32067 759420
rect 32052 759405 32067 759416
rect 31867 759225 32067 759405
rect 32546 759307 33546 759435
rect 34110 759411 34710 759461
rect 35134 759339 36134 759389
rect 36785 759380 37385 759430
rect 31867 759210 31882 759225
rect 32052 759214 32067 759225
rect 32055 759210 32067 759214
rect 20809 759131 20833 759165
rect 32546 759151 33546 759279
rect 36785 759248 37385 759298
rect 35285 759162 35319 759172
rect 35353 759162 35387 759172
rect 35421 759162 35455 759172
rect 35489 759162 35523 759172
rect 35564 759162 35598 759172
rect 35632 759162 35666 759172
rect 35700 759162 35734 759172
rect 35768 759162 35802 759172
rect 35836 759162 35870 759172
rect 35904 759162 35938 759172
rect 35972 759162 36006 759172
rect 36040 759162 36074 759172
rect 36108 759162 36142 759172
rect 36176 759162 36210 759172
rect 35255 759126 36255 759138
rect 20809 759063 20833 759097
rect 20940 759085 20983 759103
rect 20940 759069 20949 759085
rect 20974 759069 20983 759085
rect 25113 759069 25349 759093
rect 25383 759069 25417 759093
rect 20974 759051 21008 759069
rect 20809 758995 20833 759029
rect 20974 759028 21003 759051
rect 21361 759045 21409 759069
rect 20949 759027 20983 759028
rect 21385 758991 21409 759045
rect 25113 758991 25137 759069
rect 29993 759045 30993 759095
rect 31347 759045 31362 759060
rect 31535 759056 31547 759060
rect 31532 759045 31547 759056
rect 21361 758967 21409 758991
rect 25089 758967 25137 758991
rect 20809 758927 20833 758961
rect 20809 758859 20833 758893
rect 20809 758791 20833 758825
rect 20809 758723 20833 758757
rect 20809 758655 20833 758689
rect 21413 758638 22813 758681
rect 23685 758638 25085 758681
rect 19844 757229 19894 758629
rect 19994 757229 20122 758629
rect 20150 757229 20278 758629
rect 20306 757229 20434 758629
rect 20462 757229 20512 758629
rect 20809 758587 20833 758621
rect 20809 758519 20833 758553
rect 20809 758451 20833 758485
rect 21413 758475 22813 758603
rect 23685 758475 25085 758603
rect 20809 758383 20833 758417
rect 20809 758315 20833 758349
rect 21413 758312 22813 758440
rect 23685 758312 25085 758440
rect 20809 758247 20833 758281
rect 20809 758179 20833 758213
rect 21413 758149 22813 758277
rect 23685 758149 25085 758277
rect 20809 758111 20833 758145
rect 20809 758043 20833 758077
rect 20809 757975 20833 758009
rect 21413 757986 22813 758114
rect 23685 757986 25085 758114
rect 20809 757907 20833 757941
rect 20809 757839 20833 757873
rect 21413 757823 22813 757951
rect 23685 757823 25085 757951
rect 20809 757771 20833 757805
rect 20809 757703 20833 757737
rect 21413 757673 22813 757716
rect 23685 757673 25085 757716
rect 20809 757635 20833 757669
rect 20809 757567 20833 757601
rect 21361 757552 21419 757586
rect 25089 757552 25147 757586
rect 20809 757499 20833 757533
rect 20809 757431 20833 757465
rect 20809 757363 20833 757397
rect 21361 757373 21419 757397
rect 25089 757373 25147 757397
rect 21385 757363 21419 757373
rect 25113 757363 25147 757373
rect 20809 757295 20833 757329
rect 21385 757291 21419 757325
rect 25113 757291 25147 757325
rect 20809 757227 20833 757261
rect 21385 757219 21419 757253
rect 25113 757219 25147 757253
rect 20809 757159 20833 757193
rect 21385 757171 21419 757181
rect 25113 757171 25147 757181
rect 21361 757147 21419 757171
rect 25089 757147 25147 757171
rect 20809 757091 20833 757125
rect 20809 757023 20833 757057
rect 20809 756955 20833 756989
rect 21361 756969 21409 756993
rect 25089 756969 25137 756993
rect 20809 756887 20833 756921
rect 21385 756915 21409 756969
rect 25113 756915 25137 756969
rect 21361 756891 21409 756915
rect 25089 756891 25137 756915
rect 19480 756831 19583 756867
rect 21413 756754 22813 756804
rect 23685 756754 25085 756804
rect 7389 756489 8389 756561
rect 8990 756489 9990 756561
rect 15678 756534 16678 756606
rect 17278 756534 18278 756606
rect 21413 756591 22813 756719
rect 23685 756591 25085 756719
rect 15748 756523 15782 756534
rect 15816 756523 15850 756534
rect 15884 756523 15918 756534
rect 15952 756523 15986 756534
rect 16020 756523 16054 756534
rect 16088 756523 16122 756534
rect 16156 756523 16190 756534
rect 16224 756523 16258 756534
rect 16292 756523 16326 756534
rect 16360 756523 16394 756534
rect 16428 756523 16462 756534
rect 16496 756523 16530 756534
rect 16564 756523 16598 756534
rect 16632 756523 16666 756534
rect 17290 756523 17324 756534
rect 17358 756523 17392 756534
rect 17426 756523 17460 756534
rect 17494 756523 17528 756534
rect 17562 756523 17596 756534
rect 17630 756523 17664 756534
rect 17698 756523 17732 756534
rect 17766 756523 17800 756534
rect 17834 756523 17868 756534
rect 17902 756523 17936 756534
rect 17970 756523 18004 756534
rect 18038 756523 18072 756534
rect 18106 756523 18140 756534
rect 18174 756523 18208 756534
rect 15748 756513 15806 756523
rect 15816 756513 15874 756523
rect 15884 756513 15942 756523
rect 15952 756513 16010 756523
rect 16020 756513 16078 756523
rect 16088 756513 16146 756523
rect 16156 756513 16214 756523
rect 16224 756513 16282 756523
rect 16292 756513 16350 756523
rect 16360 756513 16418 756523
rect 16428 756513 16486 756523
rect 16496 756513 16554 756523
rect 16564 756513 16622 756523
rect 16632 756513 16690 756523
rect 17290 756513 17348 756523
rect 17358 756513 17416 756523
rect 17426 756513 17484 756523
rect 17494 756513 17552 756523
rect 17562 756513 17620 756523
rect 17630 756513 17688 756523
rect 17698 756513 17756 756523
rect 17766 756513 17824 756523
rect 17834 756513 17892 756523
rect 17902 756513 17960 756523
rect 17970 756513 18028 756523
rect 18038 756513 18096 756523
rect 18106 756513 18164 756523
rect 18174 756513 18232 756523
rect 15724 756489 16690 756513
rect 17266 756489 18232 756513
rect 15748 756474 15772 756489
rect 15816 756474 15840 756489
rect 15884 756474 15908 756489
rect 15952 756474 15976 756489
rect 16020 756474 16044 756489
rect 16088 756474 16112 756489
rect 16156 756474 16180 756489
rect 16224 756474 16248 756489
rect 16292 756474 16316 756489
rect 16360 756474 16384 756489
rect 16428 756474 16452 756489
rect 16496 756474 16520 756489
rect 16564 756474 16588 756489
rect 16632 756474 16656 756489
rect 17290 756474 17314 756489
rect 17358 756474 17382 756489
rect 17426 756474 17450 756489
rect 17494 756474 17518 756489
rect 17562 756474 17586 756489
rect 17630 756474 17654 756489
rect 17698 756474 17722 756489
rect 17766 756474 17790 756489
rect 17834 756474 17858 756489
rect 17902 756474 17926 756489
rect 17970 756474 17994 756489
rect 18038 756474 18062 756489
rect 18106 756474 18130 756489
rect 18174 756474 18198 756489
rect 15678 756319 16678 756474
rect 7389 756229 8389 756289
rect 8990 756229 9990 756289
rect 15678 756285 16690 756319
rect 17278 756309 18278 756474
rect 21413 756428 22813 756556
rect 23685 756428 25085 756556
rect 17266 756285 18278 756309
rect 15678 756274 16678 756285
rect 17278 756274 18278 756285
rect 15748 756261 15772 756274
rect 15816 756261 15840 756274
rect 15884 756261 15908 756274
rect 15952 756261 15976 756274
rect 16020 756261 16044 756274
rect 16088 756261 16112 756274
rect 16156 756261 16180 756274
rect 16224 756261 16248 756274
rect 16292 756261 16316 756274
rect 16360 756261 16384 756274
rect 16428 756261 16452 756274
rect 16496 756261 16520 756274
rect 16564 756261 16588 756274
rect 16632 756261 16656 756274
rect 17290 756261 17314 756274
rect 17358 756261 17382 756274
rect 17426 756261 17450 756274
rect 17494 756261 17518 756274
rect 17562 756261 17586 756274
rect 17630 756261 17654 756274
rect 17698 756261 17722 756274
rect 17766 756261 17790 756274
rect 17834 756261 17858 756274
rect 17902 756261 17926 756274
rect 17970 756261 17994 756274
rect 18038 756261 18062 756274
rect 18106 756261 18130 756274
rect 18174 756261 18198 756274
rect 21413 756265 22813 756393
rect 23685 756265 25085 756393
rect 21413 756102 22813 756230
rect 23685 756102 25085 756230
rect 7389 755871 8389 755927
rect 8990 755871 9990 755927
rect 15678 755916 16678 755972
rect 17278 755916 18278 755972
rect 21413 755952 22813 755995
rect 23685 755952 25085 755995
rect 7389 755799 8389 755855
rect 8990 755799 9990 755855
rect 15678 755844 16678 755900
rect 17278 755844 18278 755900
rect 21406 755865 21430 755889
rect 25068 755865 25092 755889
rect 21382 755841 21385 755865
rect 25113 755841 25116 755865
rect 21382 755763 21396 755787
rect 25102 755763 25116 755787
rect 21348 755739 21372 755763
rect 21406 755739 21430 755763
rect 25068 755739 25092 755763
rect 25126 755739 25150 755763
rect 25524 755703 25548 759001
rect 29993 758895 30993 758945
rect 31347 758865 31547 759045
rect 31347 758850 31362 758865
rect 31532 758854 31547 758865
rect 31535 758850 31547 758854
rect 31607 759045 31622 759060
rect 31795 759056 31807 759060
rect 31792 759045 31807 759056
rect 31607 758865 31807 759045
rect 32546 758995 33546 759123
rect 36785 759072 37385 759128
rect 35255 759019 36255 759069
rect 31607 758850 31622 758865
rect 31792 758854 31807 758865
rect 31795 758850 31807 758854
rect 32546 758839 33546 758967
rect 35255 758843 36255 758971
rect 36785 758896 37385 758952
rect 31347 758809 31362 758824
rect 31535 758820 31547 758824
rect 31532 758809 31547 758820
rect 29993 758736 30993 758786
rect 29993 758586 30993 758636
rect 31347 758629 31547 758809
rect 31347 758614 31362 758629
rect 31532 758618 31547 758629
rect 31535 758614 31547 758618
rect 31607 758809 31622 758824
rect 31795 758820 31807 758824
rect 31792 758809 31807 758820
rect 31607 758629 31807 758809
rect 32546 758683 33546 758811
rect 35255 758667 36255 758795
rect 36785 758726 37385 758776
rect 31607 758614 31622 758629
rect 31792 758618 31807 758629
rect 31795 758614 31807 758618
rect 32546 758527 33546 758655
rect 37993 758550 38593 758600
rect 28647 758450 28671 758477
rect 30171 758447 30771 758497
rect 35255 758491 36255 758547
rect 36785 758466 36797 758470
rect 36785 758455 36800 758466
rect 36970 758455 36985 758470
rect 28683 758397 28717 758431
rect 32546 758377 33546 758427
rect 28683 758328 28717 758362
rect 28683 758259 28717 758293
rect 30171 758271 30771 758327
rect 35255 758321 36255 758371
rect 36785 758275 36985 758455
rect 37993 758380 38593 758430
rect 36785 758264 36800 758275
rect 36785 758260 36797 758264
rect 36970 758260 36985 758275
rect 36785 758230 36797 758234
rect 28683 758190 28717 758224
rect 32596 758175 33596 758225
rect 35359 758156 35375 758222
rect 36143 758156 36159 758222
rect 36785 758219 36800 758230
rect 36970 758219 36985 758234
rect 28683 758121 28717 758155
rect 30171 758101 30771 758151
rect 28683 758052 28717 758086
rect 32596 758019 33596 758147
rect 28683 757983 28717 758017
rect 33959 757994 33975 758060
rect 36143 757994 36159 758060
rect 36785 758039 36985 758219
rect 36785 758028 36800 758039
rect 36785 758024 36797 758028
rect 36970 758024 36985 758039
rect 37083 758219 37098 758234
rect 37083 758039 37120 758219
rect 37083 758024 37098 758039
rect 28683 757914 28717 757948
rect 31463 757895 32063 757945
rect 28683 757845 28717 757879
rect 32596 757863 33596 757991
rect 37998 757954 38598 758004
rect 28683 757776 28717 757810
rect 28683 757707 28717 757741
rect 31463 757739 32063 757795
rect 32596 757707 33596 757835
rect 33959 757832 33975 757898
rect 36143 757832 36159 757898
rect 37998 757778 38598 757834
rect 28683 757638 28717 757672
rect 28683 757569 28717 757603
rect 31463 757589 32063 757639
rect 32596 757551 33596 757679
rect 35359 757670 35375 757736
rect 36143 757670 36159 757736
rect 37998 757608 38598 757658
rect 37998 757605 38220 757608
rect 38245 757605 38539 757608
rect 28683 757500 28717 757534
rect 28683 757431 28717 757465
rect 28683 757362 28717 757396
rect 32596 757395 33596 757523
rect 35255 757521 36255 757571
rect 28683 757293 28717 757327
rect 28683 757224 28717 757258
rect 30015 757256 30718 757272
rect 30015 757246 30721 757256
rect 28683 757155 28717 757189
rect 28683 757086 28717 757120
rect 28683 757017 28717 757051
rect 28683 756948 28717 756982
rect 28683 756879 28717 756913
rect 28683 756810 28717 756844
rect 28683 756741 28717 756775
rect 28683 756672 28717 756706
rect 28683 756603 28717 756637
rect 28683 756534 28717 756568
rect 28683 756465 28717 756499
rect 28683 756396 28717 756430
rect 28682 756361 28683 756366
rect 28682 756332 28717 756361
rect 28647 756303 28671 756332
rect 28647 756234 28671 756268
rect 28647 756165 28671 756199
rect 28647 756096 28671 756130
rect 28647 756027 28671 756061
rect 28647 755958 28671 755992
rect 28647 755889 28671 755923
rect 28647 755820 28671 755854
rect 28647 755751 28671 755785
rect 28647 755682 28671 755716
rect 29778 755695 29802 755719
rect 29802 755671 29826 755683
rect 29880 755681 29914 755715
rect 25524 755635 25548 755669
rect 7389 755497 8389 755569
rect 8990 755497 9990 755569
rect 15678 755542 16678 755614
rect 17278 755542 18278 755614
rect 28647 755613 28671 755647
rect 29778 755635 29802 755659
rect 21361 755586 21409 755610
rect 25089 755586 25137 755610
rect 15748 755531 15782 755542
rect 15816 755531 15850 755542
rect 15884 755531 15918 755542
rect 15952 755531 15986 755542
rect 16020 755531 16054 755542
rect 16088 755531 16122 755542
rect 16156 755531 16190 755542
rect 16224 755531 16258 755542
rect 16292 755531 16326 755542
rect 16360 755531 16394 755542
rect 16428 755531 16462 755542
rect 16496 755531 16530 755542
rect 16564 755531 16598 755542
rect 16632 755531 16666 755542
rect 17290 755531 17324 755542
rect 17358 755531 17392 755542
rect 17426 755531 17460 755542
rect 17494 755531 17528 755542
rect 17562 755531 17596 755542
rect 17630 755531 17664 755542
rect 17698 755531 17732 755542
rect 17766 755531 17800 755542
rect 17834 755531 17868 755542
rect 17902 755531 17936 755542
rect 17970 755531 18004 755542
rect 18038 755531 18072 755542
rect 18106 755531 18140 755542
rect 18174 755531 18208 755542
rect 21385 755532 21409 755586
rect 25113 755532 25137 755586
rect 28647 755544 28671 755578
rect 15748 755521 15806 755531
rect 15816 755521 15874 755531
rect 15884 755521 15942 755531
rect 15952 755521 16010 755531
rect 16020 755521 16078 755531
rect 16088 755521 16146 755531
rect 16156 755521 16214 755531
rect 16224 755521 16282 755531
rect 16292 755521 16350 755531
rect 16360 755521 16418 755531
rect 16428 755521 16486 755531
rect 16496 755521 16554 755531
rect 16564 755521 16622 755531
rect 16632 755521 16690 755531
rect 17290 755521 17348 755531
rect 17358 755521 17416 755531
rect 17426 755521 17484 755531
rect 17494 755521 17552 755531
rect 17562 755521 17620 755531
rect 17630 755521 17688 755531
rect 17698 755521 17756 755531
rect 17766 755521 17824 755531
rect 17834 755521 17892 755531
rect 17902 755521 17960 755531
rect 17970 755521 18028 755531
rect 18038 755521 18096 755531
rect 18106 755521 18164 755531
rect 18174 755521 18232 755531
rect 15724 755497 16690 755521
rect 17266 755497 18232 755521
rect 21361 755508 21409 755532
rect 25089 755508 25137 755532
rect 15748 755482 15772 755497
rect 15816 755482 15840 755497
rect 15884 755482 15908 755497
rect 15952 755482 15976 755497
rect 16020 755482 16044 755497
rect 16088 755482 16112 755497
rect 16156 755482 16180 755497
rect 16224 755482 16248 755497
rect 16292 755482 16316 755497
rect 16360 755482 16384 755497
rect 16428 755482 16452 755497
rect 16496 755482 16520 755497
rect 16564 755482 16588 755497
rect 16632 755482 16656 755497
rect 17290 755482 17314 755497
rect 17358 755482 17382 755497
rect 17426 755482 17450 755497
rect 17494 755482 17518 755497
rect 17562 755482 17586 755497
rect 17630 755482 17654 755497
rect 17698 755482 17722 755497
rect 17766 755482 17790 755497
rect 17834 755482 17858 755497
rect 17902 755482 17926 755497
rect 17970 755482 17994 755497
rect 18038 755482 18062 755497
rect 18106 755482 18130 755497
rect 18174 755482 18198 755497
rect 7389 755237 8389 755297
rect 8990 755237 9990 755297
rect 12559 755273 12865 755375
rect 15678 755327 16678 755482
rect 15678 755293 16690 755327
rect 17278 755317 18278 755482
rect 28647 755475 28671 755509
rect 28647 755406 28671 755440
rect 28647 755337 28671 755371
rect 17266 755293 18278 755317
rect 15678 755282 16678 755293
rect 17278 755282 18278 755293
rect 12543 755257 12881 755273
rect 15748 755269 15772 755282
rect 15816 755269 15840 755282
rect 15884 755269 15908 755282
rect 15952 755269 15976 755282
rect 16020 755269 16044 755282
rect 16088 755269 16112 755282
rect 16156 755269 16180 755282
rect 16224 755269 16248 755282
rect 16292 755269 16316 755282
rect 16360 755269 16384 755282
rect 16428 755269 16452 755282
rect 16496 755269 16520 755282
rect 16564 755269 16588 755282
rect 16632 755269 16656 755282
rect 17290 755269 17314 755282
rect 17358 755269 17382 755282
rect 17426 755269 17450 755282
rect 17494 755269 17518 755282
rect 17562 755269 17586 755282
rect 17630 755269 17654 755282
rect 17698 755269 17722 755282
rect 17766 755269 17790 755282
rect 17834 755269 17858 755282
rect 17902 755269 17926 755282
rect 17970 755269 17994 755282
rect 18038 755269 18062 755282
rect 18106 755269 18130 755282
rect 18174 755269 18198 755282
rect 19980 755048 20286 755218
rect 7389 754879 8389 754935
rect 8990 754879 9990 754935
rect 15678 754924 16678 754980
rect 17278 754924 18278 754980
rect 7389 754807 8389 754863
rect 8990 754807 9990 754863
rect 15678 754852 16678 754908
rect 17278 754852 18278 754908
rect 20945 754796 25553 755332
rect 28647 755268 28671 755302
rect 28647 755199 28671 755233
rect 28647 755154 28671 755164
rect 21413 754706 22813 754796
rect 23685 754706 25085 754796
rect 7389 754505 8389 754577
rect 8990 754505 9990 754577
rect 15678 754550 16678 754622
rect 17278 754550 18278 754622
rect 15748 754539 15782 754550
rect 15816 754539 15850 754550
rect 15884 754539 15918 754550
rect 15952 754539 15986 754550
rect 16020 754539 16054 754550
rect 16088 754539 16122 754550
rect 16156 754539 16190 754550
rect 16224 754539 16258 754550
rect 16292 754539 16326 754550
rect 16360 754539 16394 754550
rect 16428 754539 16462 754550
rect 16496 754539 16530 754550
rect 16564 754539 16598 754550
rect 16632 754539 16666 754550
rect 17290 754539 17324 754550
rect 17358 754539 17392 754550
rect 17426 754539 17460 754550
rect 17494 754539 17528 754550
rect 17562 754539 17596 754550
rect 17630 754539 17664 754550
rect 17698 754539 17732 754550
rect 17766 754539 17800 754550
rect 17834 754539 17868 754550
rect 17902 754539 17936 754550
rect 17970 754539 18004 754550
rect 18038 754539 18072 754550
rect 18106 754539 18140 754550
rect 18174 754539 18208 754550
rect 21413 754543 22813 754671
rect 23685 754543 25085 754671
rect 15748 754529 15806 754539
rect 15816 754529 15874 754539
rect 15884 754529 15942 754539
rect 15952 754529 16010 754539
rect 16020 754529 16078 754539
rect 16088 754529 16146 754539
rect 16156 754529 16214 754539
rect 16224 754529 16282 754539
rect 16292 754529 16350 754539
rect 16360 754529 16418 754539
rect 16428 754529 16486 754539
rect 16496 754529 16554 754539
rect 16564 754529 16622 754539
rect 16632 754529 16690 754539
rect 17290 754529 17348 754539
rect 17358 754529 17416 754539
rect 17426 754529 17484 754539
rect 17494 754529 17552 754539
rect 17562 754529 17620 754539
rect 17630 754529 17688 754539
rect 17698 754529 17756 754539
rect 17766 754529 17824 754539
rect 17834 754529 17892 754539
rect 17902 754529 17960 754539
rect 17970 754529 18028 754539
rect 18038 754529 18096 754539
rect 18106 754529 18164 754539
rect 18174 754529 18232 754539
rect 15724 754505 16690 754529
rect 17266 754505 18232 754529
rect 15748 754490 15772 754505
rect 15816 754490 15840 754505
rect 15884 754490 15908 754505
rect 15952 754490 15976 754505
rect 16020 754490 16044 754505
rect 16088 754490 16112 754505
rect 16156 754490 16180 754505
rect 16224 754490 16248 754505
rect 16292 754490 16316 754505
rect 16360 754490 16384 754505
rect 16428 754490 16452 754505
rect 16496 754490 16520 754505
rect 16564 754490 16588 754505
rect 16632 754490 16656 754505
rect 17290 754490 17314 754505
rect 17358 754490 17382 754505
rect 17426 754490 17450 754505
rect 17494 754490 17518 754505
rect 17562 754490 17586 754505
rect 17630 754490 17654 754505
rect 17698 754490 17722 754505
rect 17766 754490 17790 754505
rect 17834 754490 17858 754505
rect 17902 754490 17926 754505
rect 17970 754490 17994 754505
rect 18038 754490 18062 754505
rect 18106 754490 18130 754505
rect 18174 754490 18198 754505
rect 15678 754335 16678 754490
rect 7389 754245 8389 754305
rect 8990 754245 9990 754305
rect 15678 754301 16690 754335
rect 17278 754325 18278 754490
rect 21413 754380 22813 754508
rect 23685 754380 25085 754508
rect 17266 754301 18278 754325
rect 15678 754290 16678 754301
rect 17278 754290 18278 754301
rect 15748 754277 15772 754290
rect 15816 754277 15840 754290
rect 15884 754277 15908 754290
rect 15952 754277 15976 754290
rect 16020 754277 16044 754290
rect 16088 754277 16112 754290
rect 16156 754277 16180 754290
rect 16224 754277 16248 754290
rect 16292 754277 16316 754290
rect 16360 754277 16384 754290
rect 16428 754277 16452 754290
rect 16496 754277 16520 754290
rect 16564 754277 16588 754290
rect 16632 754277 16656 754290
rect 17290 754277 17314 754290
rect 17358 754277 17382 754290
rect 17426 754277 17450 754290
rect 17494 754277 17518 754290
rect 17562 754277 17586 754290
rect 17630 754277 17654 754290
rect 17698 754277 17722 754290
rect 17766 754277 17790 754290
rect 17834 754277 17858 754290
rect 17902 754277 17926 754290
rect 17970 754277 17994 754290
rect 18038 754277 18062 754290
rect 18106 754277 18130 754290
rect 18174 754277 18198 754290
rect 21413 754217 22813 754345
rect 23685 754217 25085 754345
rect 21413 754054 22813 754182
rect 23685 754054 25085 754182
rect 25936 754132 26936 754182
rect 27274 754033 27358 754036
rect 13899 753998 14059 754002
rect 7389 753887 8389 753943
rect 8990 753887 9990 753943
rect 15678 753932 16678 753988
rect 17278 753932 18278 753988
rect 7389 753815 8389 753871
rect 8990 753815 9990 753871
rect 15678 753860 16678 753916
rect 17278 753860 18278 753916
rect 21413 753891 22813 754019
rect 23685 753891 25085 754019
rect 25936 753976 26936 754032
rect 27158 753983 27358 754033
rect 13899 753852 14059 753856
rect 25936 753820 26936 753876
rect 27158 753807 27358 753935
rect 21413 753741 22813 753784
rect 23685 753741 25085 753784
rect 25936 753664 26936 753720
rect 7389 753513 8389 753585
rect 8990 753513 9990 753585
rect 15678 753558 16678 753630
rect 17278 753558 18278 753630
rect 21413 753605 22813 753648
rect 23685 753605 25085 753648
rect 27158 753631 27358 753687
rect 15748 753547 15782 753558
rect 15816 753547 15850 753558
rect 15884 753547 15918 753558
rect 15952 753547 15986 753558
rect 16020 753547 16054 753558
rect 16088 753547 16122 753558
rect 16156 753547 16190 753558
rect 16224 753547 16258 753558
rect 16292 753547 16326 753558
rect 16360 753547 16394 753558
rect 16428 753547 16462 753558
rect 16496 753547 16530 753558
rect 16564 753547 16598 753558
rect 16632 753547 16666 753558
rect 17290 753547 17324 753558
rect 17358 753547 17392 753558
rect 17426 753547 17460 753558
rect 17494 753547 17528 753558
rect 17562 753547 17596 753558
rect 17630 753547 17664 753558
rect 17698 753547 17732 753558
rect 17766 753547 17800 753558
rect 17834 753547 17868 753558
rect 17902 753547 17936 753558
rect 17970 753547 18004 753558
rect 18038 753547 18072 753558
rect 18106 753547 18140 753558
rect 18174 753547 18208 753558
rect 15748 753537 15806 753547
rect 15816 753537 15874 753547
rect 15884 753537 15942 753547
rect 15952 753537 16010 753547
rect 16020 753537 16078 753547
rect 16088 753537 16146 753547
rect 16156 753537 16214 753547
rect 16224 753537 16282 753547
rect 16292 753537 16350 753547
rect 16360 753537 16418 753547
rect 16428 753537 16486 753547
rect 16496 753537 16554 753547
rect 16564 753537 16622 753547
rect 16632 753537 16690 753547
rect 17290 753537 17348 753547
rect 17358 753537 17416 753547
rect 17426 753537 17484 753547
rect 17494 753537 17552 753547
rect 17562 753537 17620 753547
rect 17630 753537 17688 753547
rect 17698 753537 17756 753547
rect 17766 753537 17824 753547
rect 17834 753537 17892 753547
rect 17902 753537 17960 753547
rect 17970 753537 18028 753547
rect 18038 753537 18096 753547
rect 18106 753537 18164 753547
rect 18174 753537 18232 753547
rect 15724 753513 16690 753537
rect 17266 753513 18232 753537
rect 15748 753498 15772 753513
rect 15816 753498 15840 753513
rect 15884 753498 15908 753513
rect 15952 753498 15976 753513
rect 16020 753498 16044 753513
rect 16088 753498 16112 753513
rect 16156 753498 16180 753513
rect 16224 753498 16248 753513
rect 16292 753498 16316 753513
rect 16360 753498 16384 753513
rect 16428 753498 16452 753513
rect 16496 753498 16520 753513
rect 16564 753498 16588 753513
rect 16632 753498 16656 753513
rect 17290 753498 17314 753513
rect 17358 753498 17382 753513
rect 17426 753498 17450 753513
rect 17494 753498 17518 753513
rect 17562 753498 17586 753513
rect 17630 753498 17654 753513
rect 17698 753498 17722 753513
rect 17766 753498 17790 753513
rect 17834 753498 17858 753513
rect 17902 753498 17926 753513
rect 17970 753498 17994 753513
rect 18038 753498 18062 753513
rect 18106 753498 18130 753513
rect 18174 753498 18198 753513
rect 15678 753343 16678 753498
rect 7389 753253 8389 753313
rect 8990 753253 9990 753313
rect 15678 753309 16690 753343
rect 17278 753333 18278 753498
rect 21413 753442 22813 753570
rect 23685 753442 25085 753570
rect 25936 753514 26936 753564
rect 26393 753511 26477 753514
rect 26726 753511 26810 753514
rect 27158 753455 27358 753583
rect 17266 753309 18278 753333
rect 15678 753298 16678 753309
rect 17278 753298 18278 753309
rect 15748 753285 15772 753298
rect 15816 753285 15840 753298
rect 15884 753285 15908 753298
rect 15952 753285 15976 753298
rect 16020 753285 16044 753298
rect 16088 753285 16112 753298
rect 16156 753285 16180 753298
rect 16224 753285 16248 753298
rect 16292 753285 16316 753298
rect 16360 753285 16384 753298
rect 16428 753285 16452 753298
rect 16496 753285 16520 753298
rect 16564 753285 16588 753298
rect 16632 753285 16656 753298
rect 17290 753285 17314 753298
rect 17358 753285 17382 753298
rect 17426 753285 17450 753298
rect 17494 753285 17518 753298
rect 17562 753285 17586 753298
rect 17630 753285 17654 753298
rect 17698 753285 17722 753298
rect 17766 753285 17790 753298
rect 17834 753285 17858 753298
rect 17902 753285 17926 753298
rect 17970 753285 17994 753298
rect 18038 753285 18062 753298
rect 18106 753285 18130 753298
rect 18174 753285 18198 753298
rect 21413 753279 22813 753407
rect 23685 753279 25085 753407
rect 27158 753279 27358 753335
rect 21413 753116 22813 753244
rect 23685 753116 25085 753244
rect 27158 753103 27358 753231
rect 26393 753100 26477 753103
rect 26726 753100 26810 753103
rect 12543 753069 12881 753085
rect 12559 752967 12865 753069
rect 7389 752895 8389 752951
rect 8990 752895 9990 752951
rect 15678 752940 16678 752996
rect 17278 752940 18278 752996
rect 21413 752953 22813 753081
rect 23685 752953 25085 753081
rect 25936 753050 26936 753100
rect 27622 753095 27672 754095
rect 27772 753095 27828 754095
rect 27928 753095 27984 754095
rect 28084 753095 28140 754095
rect 28240 753095 28296 754095
rect 28396 753637 28446 754095
rect 28396 753553 28449 753637
rect 28396 753305 28446 753553
rect 29778 753320 29802 753344
rect 28396 753221 28449 753305
rect 29802 753296 29826 753309
rect 29880 753299 29914 753333
rect 29778 753261 29802 753285
rect 29890 753275 29914 753299
rect 28396 753095 28446 753221
rect 7389 752823 8389 752879
rect 8990 752823 9990 752879
rect 15678 752868 16678 752924
rect 17278 752868 18278 752924
rect 21413 752790 22813 752918
rect 23685 752790 25085 752918
rect 25936 752894 26936 752950
rect 27158 752927 27358 752983
rect 13899 752656 14059 752660
rect 7389 752521 8389 752593
rect 8990 752521 9990 752593
rect 15678 752566 16678 752638
rect 17278 752566 18278 752638
rect 21413 752627 22813 752755
rect 23685 752627 25085 752755
rect 25936 752738 26936 752794
rect 27158 752751 27358 752879
rect 27912 752757 27962 752873
rect 27909 752673 27962 752757
rect 28082 752673 28210 752873
rect 28258 752673 28314 752873
rect 28434 752673 28562 752873
rect 28610 752673 28660 752873
rect 27917 752669 27951 752673
rect 29880 752672 29914 752706
rect 25936 752582 26936 752638
rect 27158 752581 27358 752631
rect 27274 752578 27358 752581
rect 15748 752555 15782 752566
rect 15816 752555 15850 752566
rect 15884 752555 15918 752566
rect 15952 752555 15986 752566
rect 16020 752555 16054 752566
rect 16088 752555 16122 752566
rect 16156 752555 16190 752566
rect 16224 752555 16258 752566
rect 16292 752555 16326 752566
rect 16360 752555 16394 752566
rect 16428 752555 16462 752566
rect 16496 752555 16530 752566
rect 16564 752555 16598 752566
rect 16632 752555 16666 752566
rect 17290 752555 17324 752566
rect 17358 752555 17392 752566
rect 17426 752555 17460 752566
rect 17494 752555 17528 752566
rect 17562 752555 17596 752566
rect 17630 752555 17664 752566
rect 17698 752555 17732 752566
rect 17766 752555 17800 752566
rect 17834 752555 17868 752566
rect 17902 752555 17936 752566
rect 17970 752555 18004 752566
rect 18038 752555 18072 752566
rect 18106 752555 18140 752566
rect 18174 752555 18208 752566
rect 15748 752545 15806 752555
rect 15816 752545 15874 752555
rect 15884 752545 15942 752555
rect 15952 752545 16010 752555
rect 16020 752545 16078 752555
rect 16088 752545 16146 752555
rect 16156 752545 16214 752555
rect 16224 752545 16282 752555
rect 16292 752545 16350 752555
rect 16360 752545 16418 752555
rect 16428 752545 16486 752555
rect 16496 752545 16554 752555
rect 16564 752545 16622 752555
rect 16632 752545 16690 752555
rect 17290 752545 17348 752555
rect 17358 752545 17416 752555
rect 17426 752545 17484 752555
rect 17494 752545 17552 752555
rect 17562 752545 17620 752555
rect 17630 752545 17688 752555
rect 17698 752545 17756 752555
rect 17766 752545 17824 752555
rect 17834 752545 17892 752555
rect 17902 752545 17960 752555
rect 17970 752545 18028 752555
rect 18038 752545 18096 752555
rect 18106 752545 18164 752555
rect 18174 752545 18232 752555
rect 15724 752521 16690 752545
rect 17266 752521 18232 752545
rect 13901 752510 14061 752514
rect 15748 752506 15772 752521
rect 15816 752506 15840 752521
rect 15884 752506 15908 752521
rect 15952 752506 15976 752521
rect 16020 752506 16044 752521
rect 16088 752506 16112 752521
rect 16156 752506 16180 752521
rect 16224 752506 16248 752521
rect 16292 752506 16316 752521
rect 16360 752506 16384 752521
rect 16428 752506 16452 752521
rect 16496 752506 16520 752521
rect 16564 752506 16588 752521
rect 16632 752506 16656 752521
rect 17290 752506 17314 752521
rect 17358 752506 17382 752521
rect 17426 752506 17450 752521
rect 17494 752506 17518 752521
rect 17562 752506 17586 752521
rect 17630 752506 17654 752521
rect 17698 752506 17722 752521
rect 17766 752506 17790 752521
rect 17834 752506 17858 752521
rect 17902 752506 17926 752521
rect 17970 752506 17994 752521
rect 18038 752506 18062 752521
rect 18106 752506 18130 752521
rect 18174 752506 18198 752521
rect 15678 752351 16678 752506
rect 7389 752261 8389 752321
rect 8990 752261 9990 752321
rect 15678 752317 16690 752351
rect 17278 752341 18278 752506
rect 21413 752470 22813 752520
rect 23685 752470 25085 752520
rect 25936 752432 26936 752482
rect 21349 752390 21373 752414
rect 21407 752390 21431 752414
rect 25067 752390 25091 752414
rect 25125 752390 25149 752414
rect 21383 752356 21397 752390
rect 25101 752356 25115 752390
rect 17266 752317 18278 752341
rect 21349 752332 21373 752356
rect 21407 752332 21431 752356
rect 25067 752332 25091 752356
rect 25125 752332 25149 752356
rect 27917 752325 27951 752329
rect 15678 752306 16678 752317
rect 17278 752306 18278 752317
rect 15748 752293 15772 752306
rect 15816 752293 15840 752306
rect 15884 752293 15908 752306
rect 15952 752293 15976 752306
rect 16020 752293 16044 752306
rect 16088 752293 16112 752306
rect 16156 752293 16180 752306
rect 16224 752293 16248 752306
rect 16292 752293 16316 752306
rect 16360 752293 16384 752306
rect 16428 752293 16452 752306
rect 16496 752293 16520 752306
rect 16564 752293 16588 752306
rect 16632 752293 16656 752306
rect 17290 752293 17314 752306
rect 17358 752293 17382 752306
rect 17426 752293 17450 752306
rect 17494 752293 17518 752306
rect 17562 752293 17586 752306
rect 17630 752293 17654 752306
rect 17698 752293 17722 752306
rect 17766 752293 17790 752306
rect 17834 752293 17858 752306
rect 17902 752293 17926 752306
rect 17970 752293 17994 752306
rect 18038 752293 18062 752306
rect 18106 752293 18130 752306
rect 18174 752293 18198 752306
rect 27909 752241 27962 752325
rect 21634 752101 24864 752203
rect 27912 752125 27962 752241
rect 28082 752125 28210 752325
rect 28258 752125 28314 752325
rect 28434 752125 28562 752325
rect 28610 752125 28660 752325
rect 21186 752047 21210 752071
rect 25288 752047 25312 752071
rect 21162 752023 21186 752037
rect 25312 752023 25336 752037
rect 7389 751903 8389 751959
rect 8990 751903 9990 751959
rect 15678 751948 16678 752004
rect 17278 751948 18278 752004
rect 21072 751989 21084 752013
rect 21186 751989 21210 752013
rect 25288 751989 25312 752013
rect 25414 751989 25426 752013
rect 21385 751944 21403 751948
rect 7389 751831 8389 751887
rect 8990 751831 9990 751887
rect 15678 751876 16678 751932
rect 17278 751876 18278 751932
rect 20250 751914 20316 751930
rect 21377 751914 21403 751944
rect 21385 751904 21403 751914
rect 21383 751880 21403 751904
rect 21407 751880 21415 751914
rect 25113 751904 25121 751944
rect 25101 751880 25121 751904
rect 25125 751880 25143 751948
rect 21383 751846 21419 751880
rect 25101 751846 25147 751880
rect 21383 751812 21403 751846
rect 21407 751812 21415 751846
rect 21383 751778 21419 751812
rect 21481 751784 22881 751834
rect 23617 751784 25017 751834
rect 25101 751812 25121 751846
rect 25125 751812 25143 751846
rect 25101 751778 25147 751812
rect 21383 751744 21403 751778
rect 21407 751744 21415 751778
rect 21383 751710 21419 751744
rect 21383 751676 21403 751710
rect 21407 751676 21415 751710
rect 7389 751529 8389 751601
rect 8990 751529 9990 751601
rect 15678 751574 16678 751646
rect 17278 751574 18278 751646
rect 21383 751642 21419 751676
rect 21383 751608 21403 751642
rect 21407 751608 21415 751642
rect 21481 751621 22881 751749
rect 23617 751621 25017 751749
rect 25101 751744 25121 751778
rect 25125 751744 25143 751778
rect 25101 751710 25147 751744
rect 25101 751676 25121 751710
rect 25125 751676 25143 751710
rect 25101 751642 25147 751676
rect 25101 751608 25121 751642
rect 25125 751608 25143 751642
rect 21383 751574 21419 751608
rect 15748 751563 15782 751574
rect 15816 751563 15850 751574
rect 15884 751563 15918 751574
rect 15952 751563 15986 751574
rect 16020 751563 16054 751574
rect 16088 751563 16122 751574
rect 16156 751563 16190 751574
rect 16224 751563 16258 751574
rect 16292 751563 16326 751574
rect 16360 751563 16394 751574
rect 16428 751563 16462 751574
rect 16496 751563 16530 751574
rect 16564 751563 16598 751574
rect 16632 751563 16666 751574
rect 17290 751563 17324 751574
rect 17358 751563 17392 751574
rect 17426 751563 17460 751574
rect 17494 751563 17528 751574
rect 17562 751563 17596 751574
rect 17630 751563 17664 751574
rect 17698 751563 17732 751574
rect 17766 751563 17800 751574
rect 17834 751563 17868 751574
rect 17902 751563 17936 751574
rect 17970 751563 18004 751574
rect 18038 751563 18072 751574
rect 18106 751563 18140 751574
rect 18174 751563 18208 751574
rect 15748 751553 15806 751563
rect 15816 751553 15874 751563
rect 15884 751553 15942 751563
rect 15952 751553 16010 751563
rect 16020 751553 16078 751563
rect 16088 751553 16146 751563
rect 16156 751553 16214 751563
rect 16224 751553 16282 751563
rect 16292 751553 16350 751563
rect 16360 751553 16418 751563
rect 16428 751553 16486 751563
rect 16496 751553 16554 751563
rect 16564 751553 16622 751563
rect 16632 751553 16690 751563
rect 17290 751553 17348 751563
rect 17358 751553 17416 751563
rect 17426 751553 17484 751563
rect 17494 751553 17552 751563
rect 17562 751553 17620 751563
rect 17630 751553 17688 751563
rect 17698 751553 17756 751563
rect 17766 751553 17824 751563
rect 17834 751553 17892 751563
rect 17902 751553 17960 751563
rect 17970 751553 18028 751563
rect 18038 751553 18096 751563
rect 18106 751553 18164 751563
rect 18174 751553 18232 751563
rect 15724 751529 16690 751553
rect 17266 751529 18232 751553
rect 21383 751540 21403 751574
rect 21407 751540 21415 751574
rect 15748 751514 15772 751529
rect 15816 751514 15840 751529
rect 15884 751514 15908 751529
rect 15952 751514 15976 751529
rect 16020 751514 16044 751529
rect 16088 751514 16112 751529
rect 16156 751514 16180 751529
rect 16224 751514 16248 751529
rect 16292 751514 16316 751529
rect 16360 751514 16384 751529
rect 16428 751514 16452 751529
rect 16496 751514 16520 751529
rect 16564 751514 16588 751529
rect 16632 751514 16656 751529
rect 17290 751514 17314 751529
rect 17358 751514 17382 751529
rect 17426 751514 17450 751529
rect 17494 751514 17518 751529
rect 17562 751514 17586 751529
rect 17630 751514 17654 751529
rect 17698 751514 17722 751529
rect 17766 751514 17790 751529
rect 17834 751514 17858 751529
rect 17902 751514 17926 751529
rect 17970 751514 17994 751529
rect 18038 751514 18062 751529
rect 18106 751514 18130 751529
rect 18174 751514 18198 751529
rect 5937 751318 6089 751386
rect 15678 751359 16678 751514
rect 6005 751315 6089 751318
rect 5967 751305 6059 751315
rect 6005 751275 6021 751305
rect 1288 749503 1338 750503
rect 1438 749503 1566 750503
rect 1594 749503 1644 750503
rect 5995 749493 6021 751275
rect 7389 751269 8389 751329
rect 8990 751269 9990 751329
rect 15678 751325 16690 751359
rect 17278 751349 18278 751514
rect 17266 751325 18278 751349
rect 15678 751314 16678 751325
rect 17278 751314 18278 751325
rect 21383 751506 21419 751540
rect 21383 751472 21403 751506
rect 21407 751472 21415 751506
rect 21383 751438 21419 751472
rect 21481 751458 22881 751586
rect 23617 751458 25017 751586
rect 25101 751574 25147 751608
rect 25101 751540 25121 751574
rect 25125 751540 25143 751574
rect 25101 751506 25147 751540
rect 25101 751472 25121 751506
rect 25125 751472 25143 751506
rect 25101 751438 25147 751472
rect 21383 751404 21403 751438
rect 21407 751404 21415 751438
rect 21383 751370 21419 751404
rect 21383 751336 21403 751370
rect 21407 751336 21415 751370
rect 15748 751301 15772 751314
rect 15816 751301 15840 751314
rect 15884 751301 15908 751314
rect 15952 751301 15976 751314
rect 16020 751301 16044 751314
rect 16088 751301 16112 751314
rect 16156 751301 16180 751314
rect 16224 751301 16248 751314
rect 16292 751301 16316 751314
rect 16360 751301 16384 751314
rect 16428 751301 16452 751314
rect 16496 751301 16520 751314
rect 16564 751301 16588 751314
rect 16632 751301 16656 751314
rect 17290 751301 17314 751314
rect 17358 751301 17382 751314
rect 17426 751301 17450 751314
rect 17494 751301 17518 751314
rect 17562 751301 17586 751314
rect 17630 751301 17654 751314
rect 17698 751301 17722 751314
rect 17766 751301 17790 751314
rect 17834 751301 17858 751314
rect 17902 751301 17926 751314
rect 17970 751301 17994 751314
rect 18038 751301 18062 751314
rect 18106 751301 18130 751314
rect 18174 751301 18198 751314
rect 21383 751302 21419 751336
rect 21383 751268 21403 751302
rect 21407 751268 21415 751302
rect 21481 751295 22881 751423
rect 23617 751295 25017 751423
rect 25101 751404 25121 751438
rect 25125 751404 25143 751438
rect 25101 751370 25147 751404
rect 25101 751336 25121 751370
rect 25125 751336 25143 751370
rect 25101 751302 25147 751336
rect 25101 751268 25121 751302
rect 25125 751268 25143 751302
rect 21383 751234 21419 751268
rect 21383 751200 21403 751234
rect 21407 751200 21415 751234
rect 21383 751166 21419 751200
rect 21383 751132 21403 751166
rect 21407 751132 21415 751166
rect 21481 751132 22881 751260
rect 23617 751132 25017 751260
rect 25101 751234 25147 751268
rect 25101 751200 25121 751234
rect 25125 751200 25143 751234
rect 25101 751166 25147 751200
rect 25101 751132 25121 751166
rect 25125 751132 25143 751166
rect 21383 751098 21419 751132
rect 25101 751098 25147 751132
rect 21383 751064 21403 751098
rect 21407 751064 21415 751098
rect 21383 751030 21419 751064
rect 7389 750911 8389 750967
rect 8990 750911 9990 750967
rect 15678 750956 16678 751012
rect 17278 750956 18278 751012
rect 21383 750996 21403 751030
rect 21407 750996 21415 751030
rect 21383 750962 21419 750996
rect 21481 750969 22881 751097
rect 23617 750969 25017 751097
rect 25101 751064 25121 751098
rect 25125 751064 25143 751098
rect 25101 751030 25147 751064
rect 25101 750996 25121 751030
rect 25125 750996 25143 751030
rect 25101 750962 25147 750996
rect 26478 750985 26648 751291
rect 7389 750839 8389 750895
rect 8990 750839 9990 750895
rect 15678 750884 16678 750940
rect 17278 750884 18278 750940
rect 21383 750928 21403 750962
rect 21407 750928 21415 750962
rect 21383 750894 21419 750928
rect 21383 750860 21403 750894
rect 21407 750860 21415 750894
rect 21383 750826 21419 750860
rect 21383 750792 21403 750826
rect 21407 750792 21415 750826
rect 21481 750806 22881 750934
rect 23617 750806 25017 750934
rect 25101 750928 25121 750962
rect 25125 750928 25143 750962
rect 25101 750894 25147 750928
rect 27622 750903 27672 751903
rect 27772 750903 27828 751903
rect 27928 750903 27984 751903
rect 28084 750903 28140 751903
rect 28240 750903 28296 751903
rect 28396 751777 28446 751903
rect 28396 751693 28449 751777
rect 28396 751445 28446 751693
rect 30015 751523 30027 757246
rect 32596 757239 33596 757367
rect 35255 757345 36255 757401
rect 30135 757062 30735 757112
rect 31049 757042 32049 757092
rect 32596 757083 33596 757211
rect 35255 757169 36255 757297
rect 35255 756993 36255 757121
rect 30135 756886 30735 756942
rect 31049 756886 32049 756942
rect 32596 756927 33596 756983
rect 37998 756979 38148 756991
rect 38317 756979 38467 756991
rect 30135 756716 30735 756766
rect 31049 756736 32049 756786
rect 32596 756777 33596 756827
rect 35255 756823 36255 756873
rect 37998 756866 38598 756916
rect 35255 756754 36255 756766
rect 37998 756690 38598 756746
rect 30135 756600 30735 756650
rect 31049 756600 32049 756650
rect 32596 756575 33196 756625
rect 35255 756621 36255 756671
rect 30135 756424 30735 756480
rect 31049 756444 32049 756500
rect 30135 756248 30735 756376
rect 31049 756288 32049 756344
rect 30135 756072 30735 756200
rect 31049 756132 32049 756188
rect 32596 756141 33196 756191
rect 30135 755896 30735 756024
rect 31049 755982 32049 756032
rect 31049 755866 32049 755916
rect 30135 755726 30735 755776
rect 31049 755710 32049 755838
rect 30135 755610 30735 755660
rect 30135 755434 30735 755562
rect 31049 755554 32049 755682
rect 31049 755398 32049 755526
rect 34152 755490 34202 756478
rect 34322 755490 34372 756478
rect 34492 756465 35092 756515
rect 35255 756445 36255 756573
rect 37998 756520 38598 756570
rect 36785 756496 36797 756500
rect 36785 756485 36800 756496
rect 36970 756485 36985 756500
rect 34492 756289 35092 756345
rect 35255 756269 36255 756325
rect 36785 756305 36985 756485
rect 36785 756294 36800 756305
rect 36785 756290 36797 756294
rect 36970 756290 36985 756305
rect 37083 756485 37098 756500
rect 37083 756305 37120 756485
rect 37083 756290 37098 756305
rect 36785 756260 36797 756264
rect 36785 756249 36800 756260
rect 36970 756249 36985 756264
rect 34492 756119 35092 756169
rect 35255 756099 36255 756149
rect 36785 756069 36985 756249
rect 696597 756200 696600 756320
rect 37993 756094 38593 756144
rect 36785 756058 36800 756069
rect 36785 756054 36797 756058
rect 36970 756054 36985 756069
rect 692376 755983 692396 756017
rect 692463 755993 692532 756017
rect 696191 755993 696239 756017
rect 692487 755983 692532 755993
rect 696204 755983 696239 755993
rect 696340 755983 696360 756017
rect 34491 755849 35091 755899
rect 35255 755883 35855 755933
rect 37993 755924 38593 755974
rect 692487 755915 692502 755939
rect 696200 755915 696215 755939
rect 692454 755891 692478 755915
rect 696224 755891 696248 755915
rect 686755 755800 687355 755850
rect 34491 755673 35091 755729
rect 35255 755707 35855 755763
rect 36785 755748 37385 755798
rect 38920 755761 38946 755787
rect 692487 755748 692505 755752
rect 692479 755718 692505 755748
rect 692487 755698 692505 755718
rect 34491 755503 35091 755553
rect 35255 755531 35855 755659
rect 36785 755572 37385 755628
rect 686755 755624 687355 755680
rect 692485 755674 692505 755698
rect 692509 755674 692517 755718
rect 696215 755698 696223 755748
rect 696203 755674 696223 755698
rect 696227 755674 696245 755752
rect 692485 755640 692521 755674
rect 696203 755640 696249 755674
rect 34019 755418 34029 755490
rect 34152 755478 34372 755490
rect 34091 755415 34101 755418
rect 30135 755258 30735 755314
rect 31049 755242 32049 755370
rect 34091 755365 35091 755415
rect 35255 755361 35855 755411
rect 36785 755396 37385 755452
rect 686755 755448 687355 755504
rect 686755 755278 687355 755328
rect 30135 755082 30735 755210
rect 31049 755086 32049 755214
rect 34091 755195 35091 755245
rect 36785 755226 37385 755276
rect 34091 755192 34101 755195
rect 34202 755192 34302 755195
rect 35255 755159 35855 755209
rect 30135 754912 30735 754962
rect 31049 754930 32049 754986
rect 30135 754796 30735 754846
rect 31049 754774 32049 754902
rect 32481 754898 33081 754948
rect 30135 754620 30735 754748
rect 31049 754618 32049 754746
rect 32481 754742 33081 754870
rect 30135 754444 30735 754572
rect 31049 754462 32049 754590
rect 32481 754586 33081 754714
rect 34152 754532 34202 755132
rect 34302 754532 34352 755132
rect 34491 755066 35091 755116
rect 35255 755003 35855 755131
rect 36785 755094 37385 755144
rect 685547 755102 686147 755152
rect 687155 755007 687170 755022
rect 687343 755018 687355 755022
rect 687340 755007 687355 755018
rect 34491 754890 35091 754946
rect 36785 754918 37385 754974
rect 685547 754932 686147 754982
rect 35255 754847 35855 754903
rect 687155 754827 687355 755007
rect 34491 754720 35091 754770
rect 35255 754691 35855 754819
rect 687155 754812 687170 754827
rect 687340 754816 687355 754827
rect 687343 754812 687355 754816
rect 36785 754742 37385 754798
rect 687042 754771 687057 754786
rect 35255 754541 35855 754591
rect 36785 754572 37385 754622
rect 687020 754591 687057 754771
rect 687155 754771 687170 754786
rect 687343 754782 687355 754786
rect 687340 754771 687355 754782
rect 687155 754591 687355 754771
rect 688210 754630 688260 755630
rect 688360 754740 688488 755630
rect 688516 754740 688644 755630
rect 688672 754740 688800 755630
rect 688828 754740 688956 755630
rect 688984 754740 689112 755630
rect 689140 754740 689268 755630
rect 689296 754740 689424 755630
rect 689452 754740 689580 755630
rect 689608 754740 689736 755630
rect 689764 754740 689892 755630
rect 689920 754740 690048 755630
rect 690076 754740 690204 755630
rect 690232 754740 690360 755630
rect 690388 754630 690438 755630
rect 692485 755606 692505 755640
rect 692509 755606 692517 755640
rect 696203 755606 696223 755640
rect 696227 755606 696245 755640
rect 691275 755523 691875 755573
rect 692485 755572 692521 755606
rect 696203 755572 696249 755606
rect 692485 755538 692505 755572
rect 692509 755538 692517 755572
rect 692485 755504 692521 755538
rect 692583 755528 693983 755571
rect 694719 755528 696119 755571
rect 696203 755538 696223 755572
rect 696227 755538 696245 755572
rect 696203 755504 696249 755538
rect 692485 755470 692505 755504
rect 692509 755470 692517 755504
rect 692485 755436 692521 755470
rect 691275 755373 691875 755423
rect 692485 755402 692505 755436
rect 692509 755402 692517 755436
rect 692485 755368 692521 755402
rect 692485 755334 692505 755368
rect 692509 755334 692517 755368
rect 692583 755365 693983 755493
rect 694719 755365 696119 755493
rect 696203 755470 696223 755504
rect 696227 755470 696245 755504
rect 696203 755436 696249 755470
rect 707624 755441 707658 755475
rect 707695 755441 707729 755475
rect 707769 755441 707803 755475
rect 707840 755441 707874 755475
rect 707914 755441 707948 755475
rect 707985 755441 708019 755475
rect 708059 755441 708093 755475
rect 708130 755441 708164 755475
rect 708204 755441 708238 755475
rect 708275 755441 708309 755475
rect 708369 755441 708403 755475
rect 708446 755441 708480 755475
rect 708520 755441 708554 755465
rect 708588 755441 708610 755465
rect 709211 755441 709234 755465
rect 709270 755441 709304 755475
rect 709364 755441 709398 755475
rect 709435 755441 709469 755475
rect 709509 755441 709543 755475
rect 709580 755441 709614 755475
rect 709654 755441 709688 755475
rect 709725 755441 709759 755475
rect 709799 755441 709833 755475
rect 709870 755441 709904 755475
rect 709944 755441 709978 755475
rect 710015 755441 710049 755475
rect 710089 755441 710123 755475
rect 710160 755441 710194 755475
rect 696203 755402 696223 755436
rect 696227 755402 696245 755436
rect 707610 755431 707624 755441
rect 707658 755431 707695 755441
rect 707729 755431 707769 755441
rect 707803 755431 707840 755441
rect 707874 755431 707914 755441
rect 707948 755431 707985 755441
rect 708019 755431 708059 755441
rect 708093 755431 708130 755441
rect 708164 755431 708204 755441
rect 708238 755431 708275 755441
rect 708309 755431 708369 755441
rect 708403 755431 708446 755441
rect 708480 755431 708520 755441
rect 708554 755431 708588 755441
rect 708610 755431 708634 755441
rect 709211 755431 709270 755441
rect 709304 755431 709364 755441
rect 709398 755431 709435 755441
rect 709469 755431 709509 755441
rect 709543 755431 709580 755441
rect 709614 755431 709654 755441
rect 709688 755431 709725 755441
rect 709759 755431 709799 755441
rect 709833 755431 709870 755441
rect 709904 755431 709944 755441
rect 709978 755431 710015 755441
rect 710049 755431 710089 755441
rect 710123 755431 710160 755441
rect 710194 755431 710211 755441
rect 696203 755368 696249 755402
rect 696203 755334 696223 755368
rect 696227 755334 696245 755368
rect 707610 755337 708610 755431
rect 709211 755337 710211 755431
rect 691275 755251 691875 755301
rect 692485 755300 692521 755334
rect 692485 755266 692505 755300
rect 692509 755266 692517 755300
rect 692485 755232 692521 755266
rect 692485 755198 692505 755232
rect 692509 755198 692517 755232
rect 692583 755202 693983 755330
rect 694719 755202 696119 755330
rect 696203 755300 696249 755334
rect 711579 755317 712463 755331
rect 711579 755307 711619 755317
rect 696203 755266 696223 755300
rect 696227 755266 696245 755300
rect 701730 755290 701747 755292
rect 696203 755232 696249 755266
rect 696203 755198 696223 755232
rect 696227 755198 696245 755232
rect 701692 755220 701722 755254
rect 701730 755220 701760 755290
rect 707610 755241 708610 755301
rect 709211 755241 710211 755301
rect 692485 755164 692521 755198
rect 691275 755101 691875 755151
rect 692485 755130 692505 755164
rect 692509 755130 692517 755164
rect 692485 755096 692521 755130
rect 692485 755062 692505 755096
rect 692509 755062 692517 755096
rect 692485 755028 692521 755062
rect 692583 755039 693983 755167
rect 694719 755039 696119 755167
rect 696203 755164 696249 755198
rect 696203 755130 696223 755164
rect 696227 755130 696245 755164
rect 696203 755096 696249 755130
rect 696203 755062 696223 755096
rect 696227 755062 696245 755096
rect 699322 755064 700322 755097
rect 700922 755064 701922 755097
rect 696203 755028 696249 755062
rect 707610 755044 708610 755048
rect 709211 755044 710211 755048
rect 691275 754975 691875 755025
rect 692485 754994 692505 755028
rect 692509 754994 692517 755028
rect 692485 754960 692521 754994
rect 692485 754926 692505 754960
rect 692509 754926 692517 754960
rect 692485 754892 692521 754926
rect 691275 754825 691875 754875
rect 692485 754858 692505 754892
rect 692509 754858 692517 754892
rect 692583 754876 693983 755004
rect 694719 754876 696119 755004
rect 696203 754994 696223 755028
rect 696227 754994 696245 755028
rect 707574 754994 708646 755030
rect 696203 754960 696249 754994
rect 696203 754926 696223 754960
rect 696227 754926 696245 754960
rect 707574 754953 707610 754994
rect 708610 754953 708646 754994
rect 696203 754892 696249 754926
rect 697284 754894 697350 754910
rect 707574 754897 708646 754953
rect 696203 754858 696223 754892
rect 696227 754858 696245 754892
rect 699322 754877 700322 754894
rect 700922 754877 701922 754894
rect 707574 754881 707610 754897
rect 708610 754881 708646 754897
rect 692485 754824 692521 754858
rect 692485 754790 692505 754824
rect 692509 754790 692517 754824
rect 692485 754756 692521 754790
rect 691275 754703 691875 754753
rect 692485 754740 692505 754756
rect 692509 754740 692517 754756
rect 692583 754740 693983 754841
rect 694719 754740 696119 754841
rect 696203 754824 696249 754858
rect 707574 754825 708646 754881
rect 696203 754790 696223 754824
rect 696227 754790 696245 754824
rect 696203 754756 696249 754790
rect 696203 754740 696223 754756
rect 696227 754740 696245 754756
rect 699322 754740 700322 754811
rect 700922 754740 701922 754811
rect 707574 754788 707610 754825
rect 708610 754788 708646 754825
rect 707574 754748 708646 754788
rect 709175 754994 710247 755030
rect 709175 754953 709211 754994
rect 710211 754953 710247 754994
rect 709175 754897 710247 754953
rect 709175 754881 709211 754897
rect 710211 754881 710247 754897
rect 709175 754825 710247 754881
rect 709175 754788 709211 754825
rect 710211 754788 710247 754825
rect 709175 754748 710247 754788
rect 685542 754506 686142 754556
rect 691275 754553 691875 754603
rect 32481 754436 33081 754486
rect 30135 754268 30735 754396
rect 31049 754306 32049 754434
rect 34491 754379 35091 754429
rect 37993 754396 38593 754446
rect 32481 754306 33081 754356
rect 33261 754287 33861 754323
rect 30135 754092 30735 754220
rect 31049 754150 32049 754278
rect 32481 754150 33081 754278
rect 34491 754203 35091 754331
rect 35255 754287 35855 754337
rect 685542 754330 686142 754386
rect 36785 754312 36797 754316
rect 36785 754301 36800 754312
rect 36970 754301 36985 754316
rect 35255 754131 35855 754259
rect 36785 754121 36985 754301
rect 37993 754226 38593 754276
rect 692583 754237 693983 754280
rect 694719 754237 696119 754280
rect 699322 754278 700322 754418
rect 700922 754278 701922 754418
rect 685542 754160 686142 754210
rect 36785 754110 36800 754121
rect 36785 754106 36797 754110
rect 36970 754106 36985 754121
rect 30135 753916 30735 754044
rect 31049 753994 32049 754050
rect 32481 753994 33081 754050
rect 34491 754027 35091 754083
rect 31049 753818 32049 753946
rect 32481 753838 33081 753966
rect 33261 753907 33861 753963
rect 34491 753851 35091 753979
rect 35255 753975 35855 754103
rect 692583 754101 693983 754144
rect 694719 754101 696119 754144
rect 36785 754076 36797 754080
rect 36785 754065 36800 754076
rect 36970 754065 36985 754080
rect 36785 753885 36985 754065
rect 35255 753819 35855 753875
rect 36785 753874 36800 753885
rect 36785 753870 36797 753874
rect 36970 753870 36985 753885
rect 37083 754065 37098 754080
rect 37083 753885 37120 754065
rect 37083 753870 37098 753885
rect 37998 753800 38598 753850
rect 30135 753740 30735 753796
rect 30135 753564 30735 753692
rect 31049 753642 32049 753770
rect 32481 753688 33081 753738
rect 33261 753723 33861 753773
rect 34491 753681 35091 753731
rect 35255 753669 35855 753719
rect 37998 753624 38598 753680
rect 680215 753678 680815 753728
rect 30135 753388 30735 753516
rect 31049 753466 32049 753594
rect 32481 753558 33081 753608
rect 30135 753212 30735 753340
rect 31049 753290 32049 753418
rect 32481 753402 33081 753458
rect 37998 753454 38598 753504
rect 680215 753502 680815 753558
rect 685551 753516 686551 753566
rect 689154 753480 689204 753897
rect 689304 753480 689360 753897
rect 689460 753480 689516 753897
rect 689616 753480 689672 753897
rect 689772 753480 689828 753897
rect 689928 753480 689978 753897
rect 699322 753860 700322 753916
rect 700922 753860 701922 753916
rect 707610 753905 708610 753961
rect 709211 753905 710211 753961
rect 699322 753788 700322 753844
rect 700922 753788 701922 753844
rect 707610 753833 708610 753889
rect 709211 753833 710211 753889
rect 711579 753525 711605 755307
rect 715956 754297 716006 755297
rect 716106 754740 716234 755297
rect 716262 754297 716312 755297
rect 711579 753480 711595 753495
rect 712409 753480 712431 753485
rect 713640 753480 713641 753785
rect 713750 753772 714750 753822
rect 713750 753562 714750 753612
rect 713750 753480 714750 753496
rect 37998 753451 38220 753454
rect 38245 753451 38539 753454
rect 32481 753252 33081 753302
rect 34427 753259 35027 753309
rect 30135 753036 30735 753164
rect 31049 753114 32049 753242
rect 33672 753183 34272 753233
rect 34427 753083 35027 753211
rect 30135 752860 30735 752988
rect 31049 752938 32049 753066
rect 33672 753007 34272 753063
rect 31049 752762 32049 752890
rect 33672 752831 34272 752959
rect 34427 752907 35027 753035
rect 30135 752684 30735 752740
rect 34427 752731 35027 752859
rect 37998 752825 38148 752837
rect 38317 752825 38467 752837
rect 37998 752712 38598 752762
rect 33672 752655 34272 752711
rect 30135 752508 30735 752636
rect 31049 752592 32049 752642
rect 34427 752555 35027 752683
rect 37998 752536 38598 752592
rect 31049 752476 32049 752526
rect 33672 752479 34272 752535
rect 30135 752332 30735 752388
rect 31049 752320 32049 752448
rect 34427 752379 35027 752435
rect 37998 752366 38598 752416
rect 33672 752303 34272 752359
rect 36785 752342 36797 752346
rect 36785 752331 36800 752342
rect 36970 752331 36985 752346
rect 30135 752156 30735 752284
rect 31049 752164 32049 752292
rect 30135 751980 30735 752036
rect 31049 752008 32049 752136
rect 33672 752127 34272 752255
rect 34427 752203 35027 752331
rect 36785 752151 36985 752331
rect 36785 752140 36800 752151
rect 36785 752136 36797 752140
rect 36970 752136 36985 752151
rect 37083 752331 37098 752346
rect 37083 752151 37120 752331
rect 37083 752136 37098 752151
rect 36785 752106 36797 752110
rect 36785 752095 36800 752106
rect 36970 752095 36985 752110
rect 34427 752033 35027 752083
rect 33672 751957 34272 752007
rect 30135 751804 30735 751932
rect 36785 751915 36985 752095
rect 37993 751940 38593 751990
rect 31049 751852 32049 751908
rect 36785 751904 36800 751915
rect 36785 751900 36797 751904
rect 36970 751900 36985 751915
rect 31049 751696 32049 751824
rect 37993 751770 38593 751820
rect 30135 751634 30735 751684
rect 31049 751540 32049 751668
rect 36785 751594 37385 751644
rect 28396 751361 28449 751445
rect 31049 751384 32049 751512
rect 36785 751418 37385 751474
rect 28396 750903 28446 751361
rect 31049 751234 32049 751284
rect 36785 751242 37385 751298
rect 36785 751072 37385 751122
rect 37939 751039 37963 751063
rect 38085 751039 38109 751063
rect 29925 751003 29931 751032
rect 30271 751003 30305 751027
rect 30342 751003 30376 751027
rect 30413 751003 30447 751027
rect 30484 751003 30518 751027
rect 30555 751003 30589 751027
rect 30626 751003 30660 751027
rect 30697 751003 30731 751027
rect 37963 751015 37987 751038
rect 38061 751015 38085 751038
rect 29931 750962 29939 750986
rect 29955 750962 29961 751003
rect 29891 750938 29915 750962
rect 25101 750860 25121 750894
rect 25125 750860 25143 750894
rect 37759 750867 37783 750891
rect 25101 750826 25147 750860
rect 37792 750843 37807 750867
rect 25101 750792 25121 750826
rect 25125 750792 25143 750826
rect 21383 750758 21419 750792
rect 25101 750758 25147 750792
rect 21383 750724 21403 750758
rect 21407 750724 21415 750758
rect 25101 750724 25121 750758
rect 25125 750724 25143 750758
rect 21383 750690 21419 750724
rect 21383 750656 21403 750690
rect 21407 750656 21415 750690
rect 21481 750656 22881 750699
rect 22892 750675 22920 750703
rect 23617 750656 25017 750699
rect 25101 750690 25147 750724
rect 31458 750703 31608 750715
rect 31777 750703 31927 750715
rect 25101 750656 25121 750690
rect 25125 750656 25143 750690
rect 7389 750628 8389 750632
rect 8990 750628 9990 750632
rect 7353 750578 8425 750614
rect 7353 750537 7389 750578
rect 8389 750537 8425 750578
rect 7353 750501 8425 750537
rect 8954 750578 10026 750614
rect 15678 750582 16678 750654
rect 17278 750582 18278 750654
rect 21383 750622 21419 750656
rect 25101 750622 25147 750656
rect 21383 750588 21403 750622
rect 21407 750588 21415 750622
rect 25101 750588 25121 750622
rect 25125 750588 25143 750622
rect 8954 750537 8990 750578
rect 9990 750537 10026 750578
rect 15748 750571 15782 750582
rect 15816 750571 15850 750582
rect 15884 750571 15918 750582
rect 15952 750571 15986 750582
rect 16020 750571 16054 750582
rect 16088 750571 16122 750582
rect 16156 750571 16190 750582
rect 16224 750571 16258 750582
rect 16292 750571 16326 750582
rect 16360 750571 16394 750582
rect 16428 750571 16462 750582
rect 16496 750571 16530 750582
rect 16564 750571 16598 750582
rect 16632 750571 16666 750582
rect 17290 750571 17324 750582
rect 17358 750571 17392 750582
rect 17426 750571 17460 750582
rect 17494 750571 17528 750582
rect 17562 750571 17596 750582
rect 17630 750571 17664 750582
rect 17698 750571 17732 750582
rect 17766 750571 17800 750582
rect 17834 750571 17868 750582
rect 17902 750571 17936 750582
rect 17970 750571 18004 750582
rect 18038 750571 18072 750582
rect 18106 750571 18140 750582
rect 18174 750571 18208 750582
rect 15748 750561 15806 750571
rect 15816 750561 15874 750571
rect 15884 750561 15942 750571
rect 15952 750561 16010 750571
rect 16020 750561 16078 750571
rect 16088 750561 16146 750571
rect 16156 750561 16214 750571
rect 16224 750561 16282 750571
rect 16292 750561 16350 750571
rect 16360 750561 16418 750571
rect 16428 750561 16486 750571
rect 16496 750561 16554 750571
rect 16564 750561 16622 750571
rect 16632 750561 16690 750571
rect 17290 750561 17348 750571
rect 17358 750561 17416 750571
rect 17426 750561 17484 750571
rect 17494 750561 17552 750571
rect 17562 750561 17620 750571
rect 17630 750561 17688 750571
rect 17698 750561 17756 750571
rect 17766 750561 17824 750571
rect 17834 750561 17892 750571
rect 17902 750561 17960 750571
rect 17970 750561 18028 750571
rect 18038 750561 18096 750571
rect 18106 750561 18164 750571
rect 18174 750561 18232 750571
rect 15724 750537 16690 750561
rect 17266 750537 18232 750561
rect 21383 750554 21419 750588
rect 8954 750501 10026 750537
rect 15748 750522 15772 750537
rect 15816 750522 15840 750537
rect 15884 750522 15908 750537
rect 15952 750522 15976 750537
rect 16020 750522 16044 750537
rect 16088 750522 16112 750537
rect 16156 750522 16180 750537
rect 16224 750522 16248 750537
rect 16292 750522 16316 750537
rect 16360 750522 16384 750537
rect 16428 750522 16452 750537
rect 16496 750522 16520 750537
rect 16564 750522 16588 750537
rect 16632 750522 16656 750537
rect 17290 750522 17314 750537
rect 17358 750522 17382 750537
rect 17426 750522 17450 750537
rect 17494 750522 17518 750537
rect 17562 750522 17586 750537
rect 17630 750522 17654 750537
rect 17698 750522 17722 750537
rect 17766 750522 17790 750537
rect 17834 750522 17858 750537
rect 17902 750522 17926 750537
rect 17970 750522 17994 750537
rect 18038 750522 18062 750537
rect 18106 750522 18130 750537
rect 18174 750522 18198 750537
rect 15678 750367 16678 750522
rect 7389 750277 8389 750337
rect 8990 750277 9990 750337
rect 15678 750333 16690 750367
rect 17278 750357 18278 750522
rect 17266 750333 18278 750357
rect 15678 750322 16678 750333
rect 17278 750322 18278 750333
rect 21383 750520 21403 750554
rect 21407 750520 21415 750554
rect 21481 750520 22881 750563
rect 23617 750520 25017 750563
rect 25101 750554 25147 750588
rect 25414 750573 25438 750607
rect 31458 750590 32058 750640
rect 25101 750520 25121 750554
rect 25125 750520 25143 750554
rect 21383 750486 21419 750520
rect 25101 750486 25147 750520
rect 21383 750452 21403 750486
rect 21407 750452 21415 750486
rect 21383 750418 21419 750452
rect 21383 750384 21403 750418
rect 21407 750384 21415 750418
rect 21383 750350 21419 750384
rect 21481 750357 22881 750485
rect 23617 750357 25017 750485
rect 25101 750452 25121 750486
rect 25125 750452 25143 750486
rect 37792 750470 37807 750494
rect 25101 750418 25147 750452
rect 25101 750384 25121 750418
rect 25125 750384 25143 750418
rect 31458 750414 32058 750470
rect 37759 750446 37783 750470
rect 25101 750350 25147 750384
rect 15748 750309 15772 750322
rect 15816 750309 15840 750322
rect 15884 750309 15908 750322
rect 15952 750309 15976 750322
rect 16020 750309 16044 750322
rect 16088 750309 16112 750322
rect 16156 750309 16180 750322
rect 16224 750309 16248 750322
rect 16292 750309 16316 750322
rect 16360 750309 16384 750322
rect 16428 750309 16452 750322
rect 16496 750309 16520 750322
rect 16564 750309 16588 750322
rect 16632 750309 16656 750322
rect 17290 750309 17314 750322
rect 17358 750309 17382 750322
rect 17426 750309 17450 750322
rect 17494 750309 17518 750322
rect 17562 750309 17586 750322
rect 17630 750309 17654 750322
rect 17698 750309 17722 750322
rect 17766 750309 17790 750322
rect 17834 750309 17858 750322
rect 17902 750309 17926 750322
rect 17970 750309 17994 750322
rect 18038 750309 18062 750322
rect 18106 750309 18130 750322
rect 18174 750309 18198 750322
rect 21383 750316 21403 750350
rect 21407 750316 21415 750350
rect 21383 750282 21419 750316
rect 21383 750248 21403 750282
rect 21407 750248 21415 750282
rect 21383 750214 21419 750248
rect 21383 750180 21403 750214
rect 21407 750180 21415 750214
rect 21481 750194 22881 750322
rect 23617 750194 25017 750322
rect 25101 750316 25121 750350
rect 25125 750316 25143 750350
rect 25101 750282 25147 750316
rect 25101 750248 25121 750282
rect 25125 750248 25143 750282
rect 25101 750214 25147 750248
rect 25101 750180 25121 750214
rect 25125 750180 25143 750214
rect 25725 750197 26325 750247
rect 31458 750244 32058 750294
rect 30245 750220 30257 750224
rect 30245 750209 30260 750220
rect 30430 750209 30445 750224
rect 21383 750146 21419 750180
rect 7389 750066 8389 750070
rect 8990 750066 9990 750070
rect 15678 750061 16678 750133
rect 17278 750061 18278 750133
rect 21383 750112 21403 750146
rect 21407 750112 21415 750146
rect 21383 750078 21419 750112
rect 7353 750016 8425 750052
rect 7353 749975 7389 750016
rect 8389 749975 8425 750016
rect 7353 749919 8425 749975
rect 7353 749903 7389 749919
rect 8389 749903 8425 749919
rect 7353 749847 8425 749903
rect 7353 749810 7389 749847
rect 8389 749810 8425 749847
rect 7353 749770 8425 749810
rect 8954 750016 10026 750052
rect 8954 749975 8990 750016
rect 9990 749975 10026 750016
rect 8954 749919 10026 749975
rect 21383 750044 21403 750078
rect 21407 750044 21415 750078
rect 21383 750010 21419 750044
rect 21481 750031 22881 750159
rect 23617 750031 25017 750159
rect 25101 750146 25147 750180
rect 25101 750112 25121 750146
rect 25125 750112 25143 750146
rect 25101 750078 25147 750112
rect 25101 750044 25121 750078
rect 25125 750044 25143 750078
rect 25725 750047 26325 750097
rect 25101 750010 25147 750044
rect 21383 749976 21403 750010
rect 21407 749976 21415 750010
rect 21383 749942 21419 749976
rect 8954 749903 8990 749919
rect 9990 749903 10026 749919
rect 15678 749906 16678 749923
rect 17278 749906 18278 749923
rect 21383 749908 21403 749942
rect 21407 749908 21415 749942
rect 8954 749847 10026 749903
rect 20250 749890 20316 749906
rect 8954 749810 8990 749847
rect 9990 749810 10026 749847
rect 8954 749770 10026 749810
rect 21383 749874 21419 749908
rect 21383 749840 21403 749874
rect 21407 749840 21415 749874
rect 21481 749868 22881 749996
rect 23617 749868 25017 749996
rect 25101 749976 25121 750010
rect 25125 749976 25143 750010
rect 25101 749942 25147 749976
rect 25101 749908 25121 749942
rect 25125 749908 25143 749942
rect 25725 749925 26325 749975
rect 25101 749874 25147 749908
rect 25101 749840 25121 749874
rect 25125 749840 25143 749874
rect 21383 749806 21419 749840
rect 21383 749772 21403 749806
rect 21407 749772 21415 749806
rect 21383 749738 21419 749772
rect 15678 749703 16678 749736
rect 17278 749703 18278 749736
rect 21383 749704 21403 749738
rect 21407 749704 21415 749738
rect 21481 749705 22881 749833
rect 23617 749705 25017 749833
rect 25101 749806 25147 749840
rect 25101 749772 25121 749806
rect 25125 749772 25143 749806
rect 25725 749775 26325 749825
rect 25101 749738 25147 749772
rect 25101 749704 25121 749738
rect 25125 749704 25143 749738
rect 21383 749670 21419 749704
rect 25101 749670 25147 749704
rect 21383 749636 21403 749670
rect 21407 749636 21415 749670
rect 7389 749559 8389 749631
rect 8990 749559 9990 749631
rect 21383 749602 21419 749636
rect 15840 749510 15870 749580
rect 15878 749546 15908 749580
rect 21383 749568 21403 749602
rect 21407 749568 21415 749602
rect 15853 749508 15870 749510
rect 21383 749534 21419 749568
rect 21481 749542 22881 749670
rect 23617 749542 25017 749670
rect 25101 749636 25121 749670
rect 25125 749636 25143 749670
rect 25725 749649 26325 749699
rect 25101 749602 25147 749636
rect 25101 749568 25121 749602
rect 25125 749568 25143 749602
rect 25101 749534 25147 749568
rect 5981 749483 6021 749493
rect 5137 749469 6021 749483
rect 21383 749500 21403 749534
rect 21407 749500 21415 749534
rect 21383 749466 21419 749500
rect 7389 749369 8389 749463
rect 7389 749359 8413 749369
rect 8990 749359 9990 749463
rect 21383 749432 21403 749466
rect 21407 749432 21415 749466
rect 21383 749398 21419 749432
rect 21383 749364 21403 749398
rect 21407 749364 21415 749398
rect 21481 749379 22881 749507
rect 23617 749379 25017 749507
rect 25101 749500 25121 749534
rect 25125 749500 25143 749534
rect 25101 749466 25147 749500
rect 25725 749499 26325 749549
rect 25101 749432 25121 749466
rect 25125 749432 25143 749466
rect 25101 749398 25147 749432
rect 25101 749364 25121 749398
rect 25125 749364 25143 749398
rect 25725 749377 26325 749427
rect 21383 749330 21419 749364
rect 25101 749330 25147 749364
rect 21383 749296 21403 749330
rect 21407 749296 21415 749330
rect 25101 749296 25121 749330
rect 25125 749296 25143 749330
rect 21383 749262 21419 749296
rect 21383 749228 21403 749262
rect 21407 749228 21415 749262
rect 21481 749229 22881 749272
rect 23617 749229 25017 749272
rect 25101 749262 25147 749296
rect 25101 749228 25121 749262
rect 25125 749228 25143 749262
rect 21383 749194 21419 749228
rect 25101 749194 25147 749228
rect 25725 749227 26325 749277
rect 21383 749160 21403 749194
rect 21407 749160 21415 749194
rect 25101 749160 25121 749194
rect 25125 749160 25143 749194
rect 27162 749170 27212 750170
rect 27312 749170 27440 750170
rect 27468 749170 27596 750170
rect 27624 749170 27752 750170
rect 27780 749170 27908 750170
rect 27936 749170 28064 750170
rect 28092 749170 28220 750170
rect 28248 749170 28376 750170
rect 28404 749170 28532 750170
rect 28560 749170 28688 750170
rect 28716 749170 28844 750170
rect 28872 749170 29000 750170
rect 29028 749170 29156 750170
rect 29184 749170 29312 750170
rect 29340 749170 29390 750170
rect 30245 750029 30445 750209
rect 30245 750018 30260 750029
rect 30245 750014 30257 750018
rect 30430 750014 30445 750029
rect 30543 750209 30558 750224
rect 30543 750029 30580 750209
rect 30543 750014 30558 750029
rect 30245 749984 30257 749988
rect 30245 749973 30260 749984
rect 30430 749973 30445 749988
rect 30245 749793 30445 749973
rect 31453 749818 32053 749868
rect 30245 749782 30260 749793
rect 30245 749778 30257 749782
rect 30430 749778 30445 749793
rect 31453 749648 32053 749698
rect 30245 749472 30845 749522
rect 30245 749296 30845 749352
rect 21383 749126 21419 749160
rect 25101 749126 25147 749160
rect 21383 749102 21403 749126
rect 21385 749048 21403 749102
rect 21407 749082 21415 749126
rect 25101 749102 25121 749126
rect 25113 749082 25121 749102
rect 25125 749048 25143 749126
rect 30245 749120 30845 749176
rect 30245 748950 30845 749000
rect 21000 748800 21003 748920
rect 21352 748885 21376 748909
rect 25122 748885 25146 748909
rect 21385 748861 21400 748885
rect 25098 748861 25113 748885
rect 21274 748783 21294 748851
rect 21410 748817 21430 748851
rect 25068 748817 25088 748851
rect 25204 748817 25224 748851
rect 21385 748807 21430 748817
rect 25102 748807 25137 748817
rect 21361 748783 21430 748807
rect 25089 748783 25137 748807
rect 25238 748783 25258 748817
rect 680480 742427 680517 742520
rect 680615 742427 680815 742520
rect 685793 742483 685993 742520
rect 686053 742483 686253 742520
rect 686607 742440 687607 742490
rect 692427 742392 693027 742448
rect 679007 742216 679607 742266
rect 680615 742191 680815 742371
rect 686829 742301 687429 742351
rect 684004 742243 685004 742293
rect 695201 742282 695251 742520
rect 696287 742282 696337 742520
rect 682890 742161 683490 742211
rect 684004 742127 685004 742177
rect 686829 742125 687429 742181
rect 679007 742046 679607 742096
rect 684004 741971 685004 742027
rect 686829 741955 687429 742005
rect 680215 741870 680815 741920
rect 681713 741881 682313 741931
rect 682921 741899 683521 741949
rect 692427 741930 693027 741980
rect 684004 741821 685004 741871
rect 680215 741694 680815 741750
rect 681713 741705 682313 741761
rect 682921 741743 683521 741799
rect 685537 741749 686137 741799
rect 697088 741749 697138 742520
rect 697706 741749 697756 742520
rect 699322 742374 700322 742514
rect 700922 742374 701922 742514
rect 707610 742098 708610 742099
rect 699322 741956 700322 742012
rect 700922 741956 701922 742012
rect 707610 742001 708610 742057
rect 709211 742001 710211 742057
rect 707610 741959 708610 741960
rect 699322 741884 700322 741940
rect 700922 741884 701922 741940
rect 709211 741936 710211 741960
rect 682921 741593 683521 741643
rect 684070 741599 684670 741649
rect 685537 741593 686137 741649
rect 699322 741623 700322 741673
rect 700922 741623 701922 741673
rect 680215 741518 680815 741574
rect 707610 741523 708610 741617
rect 709211 741523 710211 741591
rect 707610 741513 707624 741523
rect 707658 741513 707695 741523
rect 707729 741513 707769 741523
rect 707803 741513 707840 741523
rect 707874 741513 707914 741523
rect 707948 741513 707985 741523
rect 708019 741513 708059 741523
rect 708093 741513 708130 741523
rect 708164 741513 708204 741523
rect 708238 741513 708275 741523
rect 708309 741513 708369 741523
rect 708403 741513 708446 741523
rect 708480 741513 708522 741523
rect 708556 741513 708604 741523
rect 709219 741513 709270 741523
rect 709304 741513 709364 741523
rect 709398 741513 709435 741523
rect 709469 741513 709509 741523
rect 709543 741513 709580 741523
rect 709614 741513 709654 741523
rect 709688 741513 709725 741523
rect 709759 741513 709799 741523
rect 709833 741513 709870 741523
rect 709904 741513 709944 741523
rect 709978 741513 710015 741523
rect 710049 741513 710089 741523
rect 710123 741513 710160 741523
rect 710194 741513 710211 741523
rect 684070 741443 684670 741499
rect 685537 741443 686137 741493
rect 692428 741442 693028 741492
rect 680215 741348 680815 741398
rect 681713 741359 682313 741409
rect 684070 741293 684670 741343
rect 692428 741292 693028 741342
rect 705107 741336 705173 741352
rect 711579 741301 711595 742520
rect 711892 741697 711942 742520
rect 712062 741697 712112 742520
rect 716071 742357 716074 742358
rect 714645 742323 714752 742357
rect 716071 742356 716072 742357
rect 716073 742356 716074 742357
rect 716071 742355 716074 742356
rect 716208 742357 716211 742358
rect 716208 742356 716209 742357
rect 716210 742356 716211 742357
rect 716208 742355 716211 742356
rect 714964 742247 715998 742329
rect 716284 742247 717318 742329
rect 714175 741398 714225 741998
rect 714425 741398 714475 741998
rect 680215 741232 680815 741282
rect 698017 741232 698053 741260
rect 692428 741162 693028 741212
rect 698030 741198 698077 741232
rect 698017 741164 698053 741198
rect 680215 741056 680815 741112
rect 692428 741006 693028 741134
rect 698030 741130 698077 741164
rect 698017 741096 698053 741130
rect 698030 741062 698077 741096
rect 698017 740983 698053 741062
rect 698084 740983 698120 741260
rect 714781 741191 714863 742226
rect 715134 741955 715828 742037
rect 714686 741123 714863 741191
rect 714645 741089 714863 741123
rect 680215 740880 680815 740936
rect 686719 740893 686739 740917
rect 686743 740893 686753 740917
rect 686719 740859 686757 740893
rect 686719 740822 686739 740859
rect 686743 740822 686753 740859
rect 692428 740850 693028 740978
rect 698017 740947 698210 740983
rect 698084 740935 698210 740947
rect 702756 740959 703645 740983
rect 702756 740935 702853 740959
rect 698084 740828 702853 740935
rect 686719 740788 686757 740822
rect 680215 740704 680815 740760
rect 686719 740751 686739 740788
rect 686743 740751 686753 740788
rect 686719 740741 686757 740751
rect 686699 740717 686767 740741
rect 686719 740704 686739 740717
rect 686743 740704 686753 740717
rect 686719 740695 686753 740704
rect 686719 740693 686743 740695
rect 692428 740694 693028 740750
rect 686685 740656 686709 740680
rect 686743 740656 686767 740680
rect 678799 740503 679399 740553
rect 680215 740534 680815 740584
rect 692428 740538 693028 740666
rect 680593 740531 680815 740534
rect 682009 740501 682069 740516
rect 682024 740465 682054 740501
rect 683708 740387 684308 740437
rect 678799 740327 679399 740383
rect 692428 740382 693028 740510
rect 714781 740308 714863 741089
rect 715063 740609 715145 741915
rect 715289 740777 715339 741719
rect 715633 740777 715683 741719
rect 715382 740672 715422 740756
rect 715542 740672 715582 740756
rect 715342 740632 715382 740672
rect 715582 740632 715622 740672
rect 715815 740609 715897 741915
rect 715134 740387 715828 740469
rect 716100 740308 716182 742226
rect 716454 741955 717148 742037
rect 716385 740609 716467 741915
rect 716599 740777 716649 741719
rect 716943 740777 716993 741719
rect 716700 740672 716740 740756
rect 716860 740672 716900 740756
rect 716660 740632 716700 740672
rect 716900 740632 716940 740672
rect 717137 740609 717219 741915
rect 716454 740387 717148 740469
rect 717419 740308 717501 742226
rect 683708 740237 684308 740287
rect 692428 740232 693028 740282
rect 678799 740157 679399 740207
rect 684565 740160 684790 740168
rect 696597 740000 696600 740120
rect 714964 740095 715998 740177
rect 716284 740095 717318 740177
rect 21000 713000 21003 713120
rect 282 712623 1316 712705
rect 1602 712623 2636 712705
rect 32810 712662 33035 712670
rect 38201 712593 38801 712643
rect 24572 712518 25172 712568
rect 33292 712513 33892 712563
rect 99 710574 181 712492
rect 452 712331 1146 712413
rect 381 710885 463 712191
rect 660 712128 700 712168
rect 900 712128 940 712168
rect 700 712044 740 712128
rect 860 712044 900 712128
rect 607 711081 657 712023
rect 951 711081 1001 712023
rect 1133 710885 1215 712191
rect 452 710763 1146 710845
rect 1418 710574 1500 712492
rect 1772 712331 2466 712413
rect 1703 710885 1785 712191
rect 1978 712128 2018 712168
rect 2218 712128 2258 712168
rect 2018 712044 2058 712128
rect 2178 712044 2218 712128
rect 1917 711081 1967 712023
rect 2261 711081 2311 712023
rect 2455 710885 2537 712191
rect 2737 711779 2819 712492
rect 24572 712362 25172 712490
rect 38201 712417 38801 712473
rect 33292 712363 33892 712413
rect 24572 712206 25172 712334
rect 35546 712299 35576 712335
rect 36785 712329 36935 712341
rect 35531 712284 35591 712299
rect 36785 712216 37385 712266
rect 38201 712247 38801 712297
rect 30833 712120 30857 712144
rect 30891 712120 30915 712144
rect 24572 712050 25172 712106
rect 30857 712105 30881 712107
rect 30857 712096 30887 712105
rect 30867 712083 30887 712096
rect 30891 712083 30907 712120
rect 30833 712059 30857 712083
rect 30867 712049 30911 712083
rect 14747 711865 19516 711972
rect 24572 711894 25172 712022
rect 30867 712012 30887 712049
rect 30891 712012 30907 712049
rect 36785 712040 37385 712096
rect 30867 711978 30911 712012
rect 30867 711941 30887 711978
rect 30891 711941 30907 711978
rect 30867 711907 30911 711941
rect 30867 711883 30887 711907
rect 30891 711883 30907 711907
rect 14747 711841 14844 711865
rect 13955 711817 14844 711841
rect 19390 711853 19516 711865
rect 19390 711841 19583 711853
rect 19390 711817 19605 711841
rect 19639 711817 19673 711841
rect 19707 711817 19741 711841
rect 19775 711817 19809 711841
rect 19843 711817 19877 711841
rect 19911 711817 19945 711841
rect 19979 711817 20013 711841
rect 20047 711817 20081 711841
rect 20115 711817 20149 711841
rect 20183 711817 20217 711841
rect 20251 711817 20285 711841
rect 20319 711817 20353 711841
rect 20387 711817 20421 711841
rect 20455 711817 20489 711841
rect 20523 711817 20557 711841
rect 20591 711817 20625 711841
rect 20659 711817 20693 711841
rect 2737 711711 2914 711779
rect 1772 710763 2466 710845
rect 2737 710574 2819 711711
rect 2848 711677 2955 711711
rect 19480 711540 19516 711817
rect 19547 711540 19583 711817
rect 24572 711738 25172 711866
rect 36785 711864 37385 711920
rect 36785 711688 37385 711744
rect 20809 711650 20833 711684
rect 20809 711582 20833 711616
rect 24572 711588 25172 711638
rect 20809 711540 20833 711548
rect 36785 711518 37385 711568
rect 3125 710802 3175 711402
rect 3375 710802 3425 711402
rect 282 710471 1316 710553
rect 1602 710471 2636 710553
rect 1389 710444 1392 710445
rect 1389 710443 1390 710444
rect 1391 710443 1392 710444
rect 1389 710442 1392 710443
rect 1526 710444 1529 710445
rect 1526 710443 1527 710444
rect 1528 710443 1529 710444
rect 2848 710443 2955 710477
rect 1526 710442 1529 710443
rect 5488 710280 5538 711103
rect 5658 710280 5708 711103
rect 6005 710280 6021 711499
rect 12427 711448 12493 711464
rect 24572 711458 25172 711508
rect 32930 711457 33530 711507
rect 35287 711391 35887 711441
rect 36785 711402 37385 711452
rect 24572 711308 25172 711358
rect 31463 711307 32063 711357
rect 32930 711301 33530 711357
rect 7389 711277 7406 711287
rect 7440 711277 7477 711287
rect 7511 711277 7551 711287
rect 7585 711277 7622 711287
rect 7656 711277 7696 711287
rect 7730 711277 7767 711287
rect 7801 711277 7841 711287
rect 7875 711277 7912 711287
rect 7946 711277 7986 711287
rect 8020 711277 8057 711287
rect 8091 711277 8131 711287
rect 8165 711277 8202 711287
rect 8236 711277 8296 711287
rect 8330 711277 8381 711287
rect 8996 711277 9044 711287
rect 9078 711277 9120 711287
rect 9154 711277 9197 711287
rect 9231 711277 9291 711287
rect 9325 711277 9362 711287
rect 9396 711277 9436 711287
rect 9470 711277 9507 711287
rect 9541 711277 9581 711287
rect 9615 711277 9652 711287
rect 9686 711277 9726 711287
rect 9760 711277 9797 711287
rect 9831 711277 9871 711287
rect 9905 711277 9942 711287
rect 9976 711277 9990 711287
rect 7389 711209 8389 711277
rect 8990 711183 9990 711277
rect 36785 711226 37385 711282
rect 15678 711127 16678 711177
rect 17278 711127 18278 711177
rect 31463 711151 32063 711207
rect 32930 711151 33530 711201
rect 34079 711157 34679 711207
rect 7389 710840 8389 710864
rect 15678 710860 16678 710916
rect 17278 710860 18278 710916
rect 8990 710840 9990 710841
rect 7389 710743 8389 710799
rect 8990 710743 9990 710799
rect 15678 710788 16678 710844
rect 17278 710788 18278 710844
rect 8990 710701 9990 710702
rect 15678 710286 16678 710426
rect 17278 710286 18278 710426
rect 19844 710280 19894 711051
rect 20462 710280 20512 711051
rect 31463 711001 32063 711051
rect 34079 711001 34679 711057
rect 35287 711039 35887 711095
rect 36785 711050 37385 711106
rect 32596 710929 33596 710979
rect 24573 710820 25173 710870
rect 34079 710851 34679 710901
rect 35287 710869 35887 710919
rect 36785 710880 37385 710930
rect 30171 710795 30771 710845
rect 32596 710773 33596 710829
rect 37993 710704 38593 710754
rect 30171 710619 30771 710675
rect 32596 710623 33596 710673
rect 34110 710589 34710 710639
rect 21263 710280 21313 710518
rect 22349 710280 22399 710518
rect 32596 710507 33596 710557
rect 30171 710449 30771 710499
rect 36785 710429 36985 710609
rect 37993 710534 38593 710584
rect 24573 710352 25173 710408
rect 29993 710310 30993 710360
rect 31347 710280 31547 710317
rect 31607 710280 31807 710317
rect 36785 710280 36985 710373
rect 37083 710280 37120 710373
rect 696597 708200 696600 708320
rect 692376 707983 692396 708017
rect 692463 707993 692532 708017
rect 696191 707993 696239 708017
rect 692487 707983 692532 707993
rect 696204 707983 696239 707993
rect 696340 707983 696360 708017
rect 692487 707915 692502 707939
rect 696200 707915 696215 707939
rect 692454 707891 692478 707915
rect 696224 707891 696248 707915
rect 686755 707800 687355 707850
rect 692487 707748 692505 707752
rect 692479 707718 692505 707748
rect 692487 707698 692505 707718
rect 686755 707624 687355 707680
rect 692485 707674 692505 707698
rect 692509 707674 692517 707718
rect 696215 707698 696223 707748
rect 696203 707674 696223 707698
rect 696227 707674 696245 707752
rect 692485 707640 692521 707674
rect 696203 707640 696249 707674
rect 686755 707448 687355 707504
rect 686755 707278 687355 707328
rect 685547 707102 686147 707152
rect 687155 707007 687170 707022
rect 687343 707018 687355 707022
rect 687340 707007 687355 707018
rect 685547 706932 686147 706982
rect 687155 706827 687355 707007
rect 687155 706812 687170 706827
rect 687340 706816 687355 706827
rect 687343 706812 687355 706816
rect 687042 706771 687057 706786
rect 687020 706591 687057 706771
rect 687155 706771 687170 706786
rect 687343 706782 687355 706786
rect 687340 706771 687355 706782
rect 687155 706591 687355 706771
rect 688210 706630 688260 707630
rect 688360 706740 688488 707630
rect 688516 706740 688644 707630
rect 688672 706740 688800 707630
rect 688828 706740 688956 707630
rect 688984 706740 689112 707630
rect 689140 706740 689268 707630
rect 689296 706740 689424 707630
rect 689452 706740 689580 707630
rect 689608 706740 689736 707630
rect 689764 706740 689892 707630
rect 689920 706740 690048 707630
rect 690076 706740 690204 707630
rect 690232 706740 690360 707630
rect 690388 706630 690438 707630
rect 692485 707606 692505 707640
rect 692509 707606 692517 707640
rect 696203 707606 696223 707640
rect 696227 707606 696245 707640
rect 691275 707523 691875 707573
rect 692485 707572 692521 707606
rect 696203 707572 696249 707606
rect 692485 707538 692505 707572
rect 692509 707538 692517 707572
rect 692485 707504 692521 707538
rect 692583 707528 693983 707571
rect 694719 707528 696119 707571
rect 696203 707538 696223 707572
rect 696227 707538 696245 707572
rect 696203 707504 696249 707538
rect 692485 707470 692505 707504
rect 692509 707470 692517 707504
rect 692485 707436 692521 707470
rect 691275 707373 691875 707423
rect 692485 707402 692505 707436
rect 692509 707402 692517 707436
rect 692485 707368 692521 707402
rect 692485 707334 692505 707368
rect 692509 707334 692517 707368
rect 692583 707365 693983 707493
rect 694719 707365 696119 707493
rect 696203 707470 696223 707504
rect 696227 707470 696245 707504
rect 696203 707436 696249 707470
rect 707624 707441 707658 707475
rect 707695 707441 707729 707475
rect 707769 707441 707803 707475
rect 707840 707441 707874 707475
rect 707914 707441 707948 707475
rect 707985 707441 708019 707475
rect 708059 707441 708093 707475
rect 708130 707441 708164 707475
rect 708204 707441 708238 707475
rect 708275 707441 708309 707475
rect 708369 707441 708403 707475
rect 708446 707441 708480 707475
rect 708520 707441 708554 707465
rect 708588 707441 708610 707465
rect 709211 707441 709234 707465
rect 709270 707441 709304 707475
rect 709364 707441 709398 707475
rect 709435 707441 709469 707475
rect 709509 707441 709543 707475
rect 709580 707441 709614 707475
rect 709654 707441 709688 707475
rect 709725 707441 709759 707475
rect 709799 707441 709833 707475
rect 709870 707441 709904 707475
rect 709944 707441 709978 707475
rect 710015 707441 710049 707475
rect 710089 707441 710123 707475
rect 710160 707441 710194 707475
rect 696203 707402 696223 707436
rect 696227 707402 696245 707436
rect 707610 707431 707624 707441
rect 707658 707431 707695 707441
rect 707729 707431 707769 707441
rect 707803 707431 707840 707441
rect 707874 707431 707914 707441
rect 707948 707431 707985 707441
rect 708019 707431 708059 707441
rect 708093 707431 708130 707441
rect 708164 707431 708204 707441
rect 708238 707431 708275 707441
rect 708309 707431 708369 707441
rect 708403 707431 708446 707441
rect 708480 707431 708520 707441
rect 708554 707431 708588 707441
rect 708610 707431 708634 707441
rect 709211 707431 709270 707441
rect 709304 707431 709364 707441
rect 709398 707431 709435 707441
rect 709469 707431 709509 707441
rect 709543 707431 709580 707441
rect 709614 707431 709654 707441
rect 709688 707431 709725 707441
rect 709759 707431 709799 707441
rect 709833 707431 709870 707441
rect 709904 707431 709944 707441
rect 709978 707431 710015 707441
rect 710049 707431 710089 707441
rect 710123 707431 710160 707441
rect 710194 707431 710211 707441
rect 696203 707368 696249 707402
rect 696203 707334 696223 707368
rect 696227 707334 696245 707368
rect 707610 707337 708610 707431
rect 709211 707337 710211 707431
rect 691275 707251 691875 707301
rect 692485 707300 692521 707334
rect 692485 707266 692505 707300
rect 692509 707266 692517 707300
rect 692485 707232 692521 707266
rect 692485 707198 692505 707232
rect 692509 707198 692517 707232
rect 692583 707202 693983 707330
rect 694719 707202 696119 707330
rect 696203 707300 696249 707334
rect 711579 707317 712463 707331
rect 711579 707307 711619 707317
rect 696203 707266 696223 707300
rect 696227 707266 696245 707300
rect 701730 707290 701747 707292
rect 696203 707232 696249 707266
rect 696203 707198 696223 707232
rect 696227 707198 696245 707232
rect 701692 707220 701722 707254
rect 701730 707220 701760 707290
rect 707610 707241 708610 707301
rect 709211 707241 710211 707301
rect 692485 707164 692521 707198
rect 691275 707101 691875 707151
rect 692485 707130 692505 707164
rect 692509 707130 692517 707164
rect 692485 707096 692521 707130
rect 692485 707062 692505 707096
rect 692509 707062 692517 707096
rect 692485 707028 692521 707062
rect 692583 707039 693983 707167
rect 694719 707039 696119 707167
rect 696203 707164 696249 707198
rect 696203 707130 696223 707164
rect 696227 707130 696245 707164
rect 696203 707096 696249 707130
rect 696203 707062 696223 707096
rect 696227 707062 696245 707096
rect 699322 707064 700322 707097
rect 700922 707064 701922 707097
rect 696203 707028 696249 707062
rect 707610 707044 708610 707048
rect 709211 707044 710211 707048
rect 691275 706975 691875 707025
rect 692485 706994 692505 707028
rect 692509 706994 692517 707028
rect 692485 706960 692521 706994
rect 692485 706926 692505 706960
rect 692509 706926 692517 706960
rect 692485 706892 692521 706926
rect 691275 706825 691875 706875
rect 692485 706858 692505 706892
rect 692509 706858 692517 706892
rect 692583 706876 693983 707004
rect 694719 706876 696119 707004
rect 696203 706994 696223 707028
rect 696227 706994 696245 707028
rect 707574 706994 708646 707030
rect 696203 706960 696249 706994
rect 696203 706926 696223 706960
rect 696227 706926 696245 706960
rect 707574 706953 707610 706994
rect 708610 706953 708646 706994
rect 696203 706892 696249 706926
rect 697284 706894 697350 706910
rect 707574 706897 708646 706953
rect 696203 706858 696223 706892
rect 696227 706858 696245 706892
rect 699322 706877 700322 706894
rect 700922 706877 701922 706894
rect 707574 706881 707610 706897
rect 708610 706881 708646 706897
rect 692485 706824 692521 706858
rect 692485 706790 692505 706824
rect 692509 706790 692517 706824
rect 692485 706756 692521 706790
rect 691275 706703 691875 706753
rect 692485 706740 692505 706756
rect 692509 706740 692517 706756
rect 692583 706740 693983 706841
rect 694719 706740 696119 706841
rect 696203 706824 696249 706858
rect 707574 706825 708646 706881
rect 696203 706790 696223 706824
rect 696227 706790 696245 706824
rect 696203 706756 696249 706790
rect 696203 706740 696223 706756
rect 696227 706740 696245 706756
rect 699322 706740 700322 706811
rect 700922 706740 701922 706811
rect 707574 706788 707610 706825
rect 708610 706788 708646 706825
rect 707574 706748 708646 706788
rect 709175 706994 710247 707030
rect 709175 706953 709211 706994
rect 710211 706953 710247 706994
rect 709175 706897 710247 706953
rect 709175 706881 709211 706897
rect 710211 706881 710247 706897
rect 709175 706825 710247 706881
rect 709175 706788 709211 706825
rect 710211 706788 710247 706825
rect 709175 706748 710247 706788
rect 685542 706506 686142 706556
rect 691275 706553 691875 706603
rect 685542 706330 686142 706386
rect 692583 706237 693983 706280
rect 694719 706237 696119 706280
rect 699322 706278 700322 706418
rect 700922 706278 701922 706418
rect 685542 706160 686142 706210
rect 692583 706101 693983 706144
rect 694719 706101 696119 706144
rect 680215 705678 680815 705728
rect 680215 705502 680815 705558
rect 685551 705516 686551 705566
rect 689154 705480 689204 705897
rect 689304 705480 689360 705897
rect 689460 705480 689516 705897
rect 689616 705480 689672 705897
rect 689772 705480 689828 705897
rect 689928 705480 689978 705897
rect 699322 705860 700322 705916
rect 700922 705860 701922 705916
rect 707610 705905 708610 705961
rect 709211 705905 710211 705961
rect 699322 705788 700322 705844
rect 700922 705788 701922 705844
rect 707610 705833 708610 705889
rect 709211 705833 710211 705889
rect 711579 705525 711605 707307
rect 715956 706297 716006 707297
rect 716106 706740 716234 707297
rect 716262 706297 716312 707297
rect 711579 705480 711595 705495
rect 712409 705480 712431 705485
rect 713640 705480 713641 705785
rect 713750 705772 714750 705822
rect 713750 705562 714750 705612
rect 713750 705480 714750 705496
rect 2850 699304 3850 699320
rect 2850 699188 3850 699238
rect 2850 698978 3850 699028
rect 3959 699015 3960 699320
rect 5169 699315 5191 699320
rect 6005 699305 6021 699320
rect 1288 697503 1338 698503
rect 1438 697503 1566 698060
rect 1594 697503 1644 698503
rect 5995 697493 6021 699275
rect 7389 698911 8389 698967
rect 8990 698911 9990 698967
rect 15678 698956 16678 699012
rect 17278 698956 18278 699012
rect 7389 698839 8389 698895
rect 8990 698839 9990 698895
rect 15678 698884 16678 698940
rect 17278 698884 18278 698940
rect 27622 698903 27672 699320
rect 27772 698903 27828 699320
rect 27928 698903 27984 699320
rect 28084 698903 28140 699320
rect 28240 698903 28296 699320
rect 28396 698903 28446 699320
rect 31049 699234 32049 699284
rect 36785 699242 37385 699298
rect 36785 699072 37385 699122
rect 21481 698656 22881 698699
rect 23617 698656 25017 698699
rect 31458 698590 32058 698640
rect 15678 698382 16678 698522
rect 17278 698382 18278 698522
rect 21481 698520 22881 698563
rect 23617 698520 25017 698563
rect 31458 698414 32058 698470
rect 25725 698197 26325 698247
rect 31458 698244 32058 698294
rect 7353 698016 8425 698052
rect 7353 697975 7389 698016
rect 8389 697975 8425 698016
rect 7353 697919 8425 697975
rect 7353 697903 7389 697919
rect 8389 697903 8425 697919
rect 7353 697847 8425 697903
rect 7353 697810 7389 697847
rect 8389 697810 8425 697847
rect 7353 697770 8425 697810
rect 8954 698016 10026 698052
rect 8954 697975 8990 698016
rect 9990 697975 10026 698016
rect 8954 697919 10026 697975
rect 21383 698044 21403 698060
rect 21407 698044 21415 698060
rect 21383 698010 21419 698044
rect 21481 698031 22881 698060
rect 23617 698031 25017 698060
rect 25101 698044 25121 698060
rect 25125 698044 25143 698060
rect 25725 698047 26325 698097
rect 25101 698010 25147 698044
rect 21383 697976 21403 698010
rect 21407 697976 21415 698010
rect 21383 697942 21419 697976
rect 8954 697903 8990 697919
rect 9990 697903 10026 697919
rect 15678 697906 16678 697923
rect 17278 697906 18278 697923
rect 21383 697908 21403 697942
rect 21407 697908 21415 697942
rect 8954 697847 10026 697903
rect 20250 697890 20316 697906
rect 8954 697810 8990 697847
rect 9990 697810 10026 697847
rect 8954 697770 10026 697810
rect 21383 697874 21419 697908
rect 21383 697840 21403 697874
rect 21407 697840 21415 697874
rect 21481 697868 22881 697996
rect 23617 697868 25017 697996
rect 25101 697976 25121 698010
rect 25125 697976 25143 698010
rect 25101 697942 25147 697976
rect 25101 697908 25121 697942
rect 25125 697908 25143 697942
rect 25725 697925 26325 697975
rect 25101 697874 25147 697908
rect 25101 697840 25121 697874
rect 25125 697840 25143 697874
rect 21383 697806 21419 697840
rect 21383 697772 21403 697806
rect 21407 697772 21415 697806
rect 21383 697738 21419 697772
rect 15678 697703 16678 697736
rect 17278 697703 18278 697736
rect 21383 697704 21403 697738
rect 21407 697704 21415 697738
rect 21481 697705 22881 697833
rect 23617 697705 25017 697833
rect 25101 697806 25147 697840
rect 25101 697772 25121 697806
rect 25125 697772 25143 697806
rect 25725 697775 26325 697825
rect 25101 697738 25147 697772
rect 25101 697704 25121 697738
rect 25125 697704 25143 697738
rect 21383 697670 21419 697704
rect 25101 697670 25147 697704
rect 21383 697636 21403 697670
rect 21407 697636 21415 697670
rect 7389 697559 8389 697631
rect 8990 697559 9990 697631
rect 21383 697602 21419 697636
rect 15840 697510 15870 697580
rect 15878 697546 15908 697580
rect 21383 697568 21403 697602
rect 21407 697568 21415 697602
rect 15853 697508 15870 697510
rect 21383 697534 21419 697568
rect 21481 697542 22881 697670
rect 23617 697542 25017 697670
rect 25101 697636 25121 697670
rect 25125 697636 25143 697670
rect 25725 697649 26325 697699
rect 25101 697602 25147 697636
rect 25101 697568 25121 697602
rect 25125 697568 25143 697602
rect 25101 697534 25147 697568
rect 5981 697483 6021 697493
rect 5137 697469 6021 697483
rect 21383 697500 21403 697534
rect 21407 697500 21415 697534
rect 21383 697466 21419 697500
rect 7389 697369 8389 697463
rect 7389 697359 8413 697369
rect 8990 697359 9990 697463
rect 21383 697432 21403 697466
rect 21407 697432 21415 697466
rect 21383 697398 21419 697432
rect 21383 697364 21403 697398
rect 21407 697364 21415 697398
rect 21481 697379 22881 697507
rect 23617 697379 25017 697507
rect 25101 697500 25121 697534
rect 25125 697500 25143 697534
rect 25101 697466 25147 697500
rect 25725 697499 26325 697549
rect 25101 697432 25121 697466
rect 25125 697432 25143 697466
rect 25101 697398 25147 697432
rect 25101 697364 25121 697398
rect 25125 697364 25143 697398
rect 25725 697377 26325 697427
rect 21383 697330 21419 697364
rect 25101 697330 25147 697364
rect 21383 697296 21403 697330
rect 21407 697296 21415 697330
rect 25101 697296 25121 697330
rect 25125 697296 25143 697330
rect 21383 697262 21419 697296
rect 21383 697228 21403 697262
rect 21407 697228 21415 697262
rect 21481 697229 22881 697272
rect 23617 697229 25017 697272
rect 25101 697262 25147 697296
rect 25101 697228 25121 697262
rect 25125 697228 25143 697262
rect 21383 697194 21419 697228
rect 25101 697194 25147 697228
rect 25725 697227 26325 697277
rect 21383 697160 21403 697194
rect 21407 697160 21415 697194
rect 25101 697160 25121 697194
rect 25125 697160 25143 697194
rect 27162 697170 27212 698170
rect 27312 697170 27440 698060
rect 27468 697170 27596 698060
rect 27624 697170 27752 698060
rect 27780 697170 27908 698060
rect 27936 697170 28064 698060
rect 28092 697170 28220 698060
rect 28248 697170 28376 698060
rect 28404 697170 28532 698060
rect 28560 697170 28688 698060
rect 28716 697170 28844 698060
rect 28872 697170 29000 698060
rect 29028 697170 29156 698060
rect 29184 697170 29312 698060
rect 29340 697170 29390 698170
rect 30245 698029 30445 698209
rect 30245 698018 30260 698029
rect 30245 698014 30257 698018
rect 30430 698014 30445 698029
rect 30543 698029 30580 698209
rect 30543 698014 30558 698029
rect 30245 697984 30257 697988
rect 30245 697973 30260 697984
rect 30430 697973 30445 697988
rect 30245 697793 30445 697973
rect 31453 697818 32053 697868
rect 30245 697782 30260 697793
rect 30245 697778 30257 697782
rect 30430 697778 30445 697793
rect 31453 697648 32053 697698
rect 30245 697472 30845 697522
rect 30245 697296 30845 697352
rect 21383 697126 21419 697160
rect 25101 697126 25147 697160
rect 21383 697102 21403 697126
rect 21385 697048 21403 697102
rect 21407 697082 21415 697126
rect 25101 697102 25121 697126
rect 25113 697082 25121 697102
rect 25125 697048 25143 697126
rect 30245 697120 30845 697176
rect 30245 696950 30845 697000
rect 21000 696800 21003 696920
rect 21352 696885 21376 696909
rect 25122 696885 25146 696909
rect 21385 696861 21400 696885
rect 25098 696861 25113 696885
rect 21274 696783 21294 696851
rect 21410 696817 21430 696851
rect 25068 696817 25088 696851
rect 25204 696817 25224 696851
rect 21385 696807 21430 696817
rect 25102 696807 25137 696817
rect 21361 696783 21430 696807
rect 25089 696783 25137 696807
rect 25238 696783 25258 696817
rect 680480 694427 680517 694520
rect 680615 694427 680815 694520
rect 685793 694483 685993 694520
rect 686053 694483 686253 694520
rect 686607 694440 687607 694490
rect 692427 694392 693027 694448
rect 679007 694216 679607 694266
rect 680615 694191 680815 694371
rect 686829 694301 687429 694351
rect 684004 694243 685004 694293
rect 695201 694282 695251 694520
rect 696287 694282 696337 694520
rect 682890 694161 683490 694211
rect 684004 694127 685004 694177
rect 686829 694125 687429 694181
rect 679007 694046 679607 694096
rect 684004 693971 685004 694027
rect 686829 693955 687429 694005
rect 680215 693870 680815 693920
rect 681713 693881 682313 693931
rect 682921 693899 683521 693949
rect 692427 693930 693027 693980
rect 684004 693821 685004 693871
rect 680215 693694 680815 693750
rect 681713 693705 682313 693761
rect 682921 693743 683521 693799
rect 685537 693749 686137 693799
rect 697088 693749 697138 694520
rect 697706 693749 697756 694520
rect 699322 694374 700322 694514
rect 700922 694374 701922 694514
rect 707610 694098 708610 694099
rect 699322 693956 700322 694012
rect 700922 693956 701922 694012
rect 707610 694001 708610 694057
rect 709211 694001 710211 694057
rect 707610 693959 708610 693960
rect 699322 693884 700322 693940
rect 700922 693884 701922 693940
rect 709211 693936 710211 693960
rect 682921 693593 683521 693643
rect 684070 693599 684670 693649
rect 685537 693593 686137 693649
rect 699322 693623 700322 693673
rect 700922 693623 701922 693673
rect 680215 693518 680815 693574
rect 707610 693523 708610 693617
rect 709211 693523 710211 693591
rect 707610 693513 707624 693523
rect 707658 693513 707695 693523
rect 707729 693513 707769 693523
rect 707803 693513 707840 693523
rect 707874 693513 707914 693523
rect 707948 693513 707985 693523
rect 708019 693513 708059 693523
rect 708093 693513 708130 693523
rect 708164 693513 708204 693523
rect 708238 693513 708275 693523
rect 708309 693513 708369 693523
rect 708403 693513 708446 693523
rect 708480 693513 708522 693523
rect 708556 693513 708604 693523
rect 709219 693513 709270 693523
rect 709304 693513 709364 693523
rect 709398 693513 709435 693523
rect 709469 693513 709509 693523
rect 709543 693513 709580 693523
rect 709614 693513 709654 693523
rect 709688 693513 709725 693523
rect 709759 693513 709799 693523
rect 709833 693513 709870 693523
rect 709904 693513 709944 693523
rect 709978 693513 710015 693523
rect 710049 693513 710089 693523
rect 710123 693513 710160 693523
rect 710194 693513 710211 693523
rect 684070 693443 684670 693499
rect 685537 693443 686137 693493
rect 692428 693442 693028 693492
rect 680215 693348 680815 693398
rect 681713 693359 682313 693409
rect 684070 693293 684670 693343
rect 692428 693292 693028 693342
rect 705107 693336 705173 693352
rect 711579 693301 711595 694520
rect 711892 693697 711942 694520
rect 712062 693697 712112 694520
rect 716071 694357 716074 694358
rect 714645 694323 714752 694357
rect 716071 694356 716072 694357
rect 716073 694356 716074 694357
rect 716071 694355 716074 694356
rect 716208 694357 716211 694358
rect 716208 694356 716209 694357
rect 716210 694356 716211 694357
rect 716208 694355 716211 694356
rect 714964 694247 715998 694329
rect 716284 694247 717318 694329
rect 714175 693398 714225 693998
rect 714425 693398 714475 693998
rect 680215 693232 680815 693282
rect 698017 693232 698053 693260
rect 692428 693162 693028 693212
rect 698030 693198 698077 693232
rect 698017 693164 698053 693198
rect 680215 693056 680815 693112
rect 692428 693006 693028 693134
rect 698030 693130 698077 693164
rect 698017 693096 698053 693130
rect 698030 693062 698077 693096
rect 698017 692983 698053 693062
rect 698084 692983 698120 693260
rect 714781 693191 714863 694226
rect 715134 693955 715828 694037
rect 714686 693123 714863 693191
rect 714645 693089 714863 693123
rect 680215 692880 680815 692936
rect 686719 692893 686739 692917
rect 686743 692893 686753 692917
rect 686719 692859 686757 692893
rect 686719 692822 686739 692859
rect 686743 692822 686753 692859
rect 692428 692850 693028 692978
rect 698017 692947 698210 692983
rect 698084 692935 698210 692947
rect 702756 692959 703645 692983
rect 702756 692935 702853 692959
rect 698084 692828 702853 692935
rect 686719 692788 686757 692822
rect 680215 692704 680815 692760
rect 686719 692751 686739 692788
rect 686743 692751 686753 692788
rect 686719 692741 686757 692751
rect 686699 692717 686767 692741
rect 686719 692704 686739 692717
rect 686743 692704 686753 692717
rect 686719 692695 686753 692704
rect 686719 692693 686743 692695
rect 692428 692694 693028 692750
rect 686685 692656 686709 692680
rect 686743 692656 686767 692680
rect 678799 692503 679399 692553
rect 680215 692534 680815 692584
rect 692428 692538 693028 692666
rect 680593 692531 680815 692534
rect 682009 692501 682069 692516
rect 682024 692465 682054 692501
rect 683708 692387 684308 692437
rect 678799 692327 679399 692383
rect 692428 692382 693028 692510
rect 714781 692308 714863 693089
rect 715063 692609 715145 693915
rect 715289 692777 715339 693719
rect 715633 692777 715683 693719
rect 715382 692672 715422 692756
rect 715542 692672 715582 692756
rect 715342 692632 715382 692672
rect 715582 692632 715622 692672
rect 715815 692609 715897 693915
rect 715134 692387 715828 692469
rect 716100 692308 716182 694226
rect 716454 693955 717148 694037
rect 716385 692609 716467 693915
rect 716599 692777 716649 693719
rect 716943 692777 716993 693719
rect 716700 692672 716740 692756
rect 716860 692672 716900 692756
rect 716660 692632 716700 692672
rect 716900 692632 716940 692672
rect 717137 692609 717219 693915
rect 716454 692387 717148 692469
rect 717419 692308 717501 694226
rect 683708 692237 684308 692287
rect 692428 692232 693028 692282
rect 678799 692157 679399 692207
rect 684565 692160 684790 692168
rect 696597 692000 696600 692120
rect 714964 692095 715998 692177
rect 716284 692095 717318 692177
rect 21000 665000 21003 665120
rect 282 664623 1316 664705
rect 1602 664623 2636 664705
rect 32810 664662 33035 664670
rect 38201 664593 38801 664643
rect 24572 664518 25172 664568
rect 33292 664513 33892 664563
rect 99 662574 181 664492
rect 452 664331 1146 664413
rect 381 662885 463 664191
rect 660 664128 700 664168
rect 900 664128 940 664168
rect 700 664044 740 664128
rect 860 664044 900 664128
rect 607 663081 657 664023
rect 700 663048 740 663132
rect 860 663048 900 663132
rect 951 663081 1001 664023
rect 660 663008 700 663048
rect 900 663008 940 663048
rect 1133 662885 1215 664191
rect 452 662763 1146 662845
rect 1418 662574 1500 664492
rect 1772 664331 2466 664413
rect 1703 662885 1785 664191
rect 1978 664128 2018 664168
rect 2218 664128 2258 664168
rect 2018 664044 2058 664128
rect 2178 664044 2218 664128
rect 1917 663081 1967 664023
rect 2018 663048 2058 663132
rect 2178 663048 2218 663132
rect 2261 663081 2311 664023
rect 1978 663008 2018 663048
rect 2218 663008 2258 663048
rect 2455 662885 2537 664191
rect 2737 663779 2819 664492
rect 24572 664362 25172 664490
rect 38201 664417 38801 664473
rect 33292 664363 33892 664413
rect 24572 664206 25172 664334
rect 35546 664299 35576 664335
rect 36785 664329 36935 664341
rect 35531 664284 35591 664299
rect 36785 664216 37385 664266
rect 38201 664247 38801 664297
rect 30833 664120 30857 664144
rect 30891 664120 30915 664144
rect 24572 664050 25172 664106
rect 30857 664105 30881 664107
rect 30857 664096 30887 664105
rect 30867 664083 30887 664096
rect 30891 664083 30907 664120
rect 30833 664059 30857 664083
rect 30867 664049 30911 664083
rect 14747 663865 19516 663972
rect 24572 663894 25172 664022
rect 30867 664012 30887 664049
rect 30891 664012 30907 664049
rect 36785 664040 37385 664096
rect 30867 663978 30911 664012
rect 30867 663941 30887 663978
rect 30891 663941 30907 663978
rect 30867 663907 30911 663941
rect 30867 663883 30887 663907
rect 30891 663883 30907 663907
rect 14747 663841 14844 663865
rect 13955 663817 14844 663841
rect 19390 663853 19516 663865
rect 19390 663841 19583 663853
rect 19390 663817 19605 663841
rect 19639 663817 19673 663841
rect 19707 663817 19741 663841
rect 19775 663817 19809 663841
rect 19843 663817 19877 663841
rect 19911 663817 19945 663841
rect 19979 663817 20013 663841
rect 20047 663817 20081 663841
rect 20115 663817 20149 663841
rect 20183 663817 20217 663841
rect 20251 663817 20285 663841
rect 20319 663817 20353 663841
rect 20387 663817 20421 663841
rect 20455 663817 20489 663841
rect 20523 663817 20557 663841
rect 20591 663817 20625 663841
rect 20659 663817 20693 663841
rect 2737 663711 2914 663779
rect 1772 662763 2466 662845
rect 2737 662574 2819 663711
rect 2848 663677 2955 663711
rect 6005 663498 6021 663499
rect 3125 662802 3175 663402
rect 3375 662802 3425 663402
rect 5967 663363 6059 663498
rect 12427 663448 12493 663464
rect 282 662471 1316 662553
rect 1602 662471 2636 662553
rect 2806 662477 2914 662545
rect 1389 662444 1392 662445
rect 1389 662443 1390 662444
rect 1391 662443 1392 662444
rect 1389 662442 1392 662443
rect 1526 662444 1529 662445
rect 1526 662443 1527 662444
rect 1528 662443 1529 662444
rect 2848 662443 2955 662477
rect 1526 662442 1529 662443
rect 5488 662103 5538 663103
rect 5658 662103 5708 663103
rect 183 661602 1183 661652
rect 2850 661632 3850 661682
rect 183 661446 1183 661574
rect 2850 661416 3850 661544
rect 183 661296 1183 661346
rect 183 661180 1183 661230
rect 2850 661200 3850 661328
rect 183 660964 1183 661020
rect 2850 660984 3850 661112
rect 5488 660993 5538 661993
rect 5658 660993 5708 661993
rect 183 660748 1183 660804
rect 2850 660768 3850 660896
rect 183 660592 1183 660720
rect 2850 660552 3850 660608
rect 183 660442 1183 660492
rect 2850 660336 3850 660392
rect 183 660276 1183 660326
rect 2850 660120 3850 660248
rect 183 660060 1183 660116
rect 183 659904 1183 660032
rect 2850 659904 3850 660032
rect 5488 659872 5538 660872
rect 5658 659872 5708 660872
rect 183 659748 1183 659804
rect 183 659592 1183 659720
rect 2850 659688 3850 659816
rect 183 659436 1183 659492
rect 2850 659472 3850 659600
rect 183 659286 1183 659336
rect 2850 659256 3850 659312
rect 583 659170 1183 659220
rect 583 659020 1183 659070
rect 2850 659040 3850 659168
rect 183 658904 1183 658954
rect 2850 658824 3850 658952
rect 183 658748 1183 658804
rect 5488 658751 5538 659751
rect 5658 658751 5708 659751
rect 183 658598 1183 658648
rect 2850 658608 3850 658736
rect 5971 658489 6059 663363
rect 7406 663287 7440 663321
rect 7477 663287 7511 663321
rect 7551 663287 7585 663321
rect 7622 663287 7656 663321
rect 7696 663287 7730 663321
rect 7767 663287 7801 663321
rect 7841 663287 7875 663321
rect 7912 663287 7946 663321
rect 7986 663287 8020 663321
rect 8057 663287 8091 663321
rect 8131 663287 8165 663321
rect 8202 663287 8236 663321
rect 8296 663287 8330 663321
rect 8381 663311 8423 663321
rect 8381 663287 8389 663311
rect 8415 663287 8423 663311
rect 8956 663311 8996 663321
rect 8956 663287 8962 663311
rect 8990 663287 8996 663311
rect 9044 663287 9078 663321
rect 9120 663287 9154 663321
rect 9197 663287 9231 663321
rect 9291 663287 9325 663321
rect 9362 663287 9396 663321
rect 9436 663287 9470 663321
rect 9507 663287 9541 663321
rect 9581 663287 9615 663321
rect 9652 663287 9686 663321
rect 9726 663287 9760 663321
rect 9797 663287 9831 663321
rect 9871 663287 9905 663321
rect 9942 663287 9976 663321
rect 7389 663277 7406 663287
rect 7440 663277 7477 663287
rect 7511 663277 7551 663287
rect 7585 663277 7622 663287
rect 7656 663277 7696 663287
rect 7730 663277 7767 663287
rect 7801 663277 7841 663287
rect 7875 663277 7912 663287
rect 7946 663277 7986 663287
rect 8020 663277 8057 663287
rect 8091 663277 8131 663287
rect 8165 663277 8202 663287
rect 8236 663277 8296 663287
rect 8330 663277 8381 663287
rect 8389 663277 8423 663287
rect 8990 663277 9044 663287
rect 9078 663277 9120 663287
rect 9154 663277 9197 663287
rect 9231 663277 9291 663287
rect 9325 663277 9362 663287
rect 9396 663277 9436 663287
rect 9470 663277 9507 663287
rect 9541 663277 9581 663287
rect 9615 663277 9652 663287
rect 9686 663277 9726 663287
rect 9760 663277 9797 663287
rect 9831 663277 9871 663287
rect 9905 663277 9942 663287
rect 9976 663277 9990 663287
rect 7389 663209 8389 663277
rect 8990 663183 9990 663277
rect 7389 663087 8389 663147
rect 8990 663087 9990 663147
rect 15678 663127 16678 663177
rect 17278 663127 18278 663177
rect 7353 662864 7389 662876
rect 8389 662864 8425 662876
rect 7353 662840 8425 662864
rect 7353 662799 7389 662840
rect 8389 662799 8425 662840
rect 7353 662743 8425 662799
rect 7353 662706 7389 662743
rect 8389 662706 8425 662743
rect 7353 662666 8425 662706
rect 8954 662841 8990 662876
rect 9990 662841 10026 662876
rect 15678 662860 16678 662916
rect 17278 662860 18278 662916
rect 8954 662840 10026 662841
rect 8954 662799 8990 662840
rect 9990 662799 10026 662840
rect 8954 662743 10026 662799
rect 15678 662788 16678 662844
rect 17278 662788 18278 662844
rect 8954 662706 8990 662743
rect 9990 662706 10026 662743
rect 8954 662701 10026 662706
rect 8954 662666 8990 662701
rect 9990 662666 10026 662701
rect 7389 662441 8389 662513
rect 8990 662441 9990 662513
rect 15678 662486 16678 662558
rect 17278 662486 18278 662558
rect 15748 662475 15782 662486
rect 15816 662475 15850 662486
rect 15884 662475 15918 662486
rect 15952 662475 15986 662486
rect 16020 662475 16054 662486
rect 16088 662475 16122 662486
rect 16156 662475 16190 662486
rect 16224 662475 16258 662486
rect 16292 662475 16326 662486
rect 16360 662475 16394 662486
rect 16428 662475 16462 662486
rect 16496 662475 16530 662486
rect 16564 662475 16598 662486
rect 16632 662475 16666 662486
rect 17290 662475 17324 662486
rect 17358 662475 17392 662486
rect 17426 662475 17460 662486
rect 17494 662475 17528 662486
rect 17562 662475 17596 662486
rect 17630 662475 17664 662486
rect 17698 662475 17732 662486
rect 17766 662475 17800 662486
rect 17834 662475 17868 662486
rect 17902 662475 17936 662486
rect 17970 662475 18004 662486
rect 18038 662475 18072 662486
rect 18106 662475 18140 662486
rect 18174 662475 18208 662486
rect 15748 662465 15806 662475
rect 15816 662465 15874 662475
rect 15884 662465 15942 662475
rect 15952 662465 16010 662475
rect 16020 662465 16078 662475
rect 16088 662465 16146 662475
rect 16156 662465 16214 662475
rect 16224 662465 16282 662475
rect 16292 662465 16350 662475
rect 16360 662465 16418 662475
rect 16428 662465 16486 662475
rect 16496 662465 16554 662475
rect 16564 662465 16622 662475
rect 16632 662465 16690 662475
rect 17290 662465 17348 662475
rect 17358 662465 17416 662475
rect 17426 662465 17484 662475
rect 17494 662465 17552 662475
rect 17562 662465 17620 662475
rect 17630 662465 17688 662475
rect 17698 662465 17756 662475
rect 17766 662465 17824 662475
rect 17834 662465 17892 662475
rect 17902 662465 17960 662475
rect 17970 662465 18028 662475
rect 18038 662465 18096 662475
rect 18106 662465 18164 662475
rect 18174 662465 18232 662475
rect 15724 662441 16690 662465
rect 17266 662441 18232 662465
rect 15748 662426 15772 662441
rect 15816 662426 15840 662441
rect 15884 662426 15908 662441
rect 15952 662426 15976 662441
rect 16020 662426 16044 662441
rect 16088 662426 16112 662441
rect 16156 662426 16180 662441
rect 16224 662426 16248 662441
rect 16292 662426 16316 662441
rect 16360 662426 16384 662441
rect 16428 662426 16452 662441
rect 16496 662426 16520 662441
rect 16564 662426 16588 662441
rect 16632 662426 16656 662441
rect 17290 662426 17314 662441
rect 17358 662426 17382 662441
rect 17426 662426 17450 662441
rect 17494 662426 17518 662441
rect 17562 662426 17586 662441
rect 17630 662426 17654 662441
rect 17698 662426 17722 662441
rect 17766 662426 17790 662441
rect 17834 662426 17858 662441
rect 17902 662426 17926 662441
rect 17970 662426 17994 662441
rect 18038 662426 18062 662441
rect 18106 662426 18130 662441
rect 18174 662426 18198 662441
rect 15678 662271 16678 662426
rect 7389 662181 8389 662241
rect 8990 662181 9990 662241
rect 15678 662237 16690 662271
rect 17278 662261 18278 662426
rect 17266 662237 18278 662261
rect 15678 662226 16678 662237
rect 17278 662226 18278 662237
rect 15748 662213 15772 662226
rect 15816 662213 15840 662226
rect 15884 662213 15908 662226
rect 15952 662213 15976 662226
rect 16020 662213 16044 662226
rect 16088 662213 16112 662226
rect 16156 662213 16180 662226
rect 16224 662213 16248 662226
rect 16292 662213 16316 662226
rect 16360 662213 16384 662226
rect 16428 662213 16452 662226
rect 16496 662213 16520 662226
rect 16564 662213 16588 662226
rect 16632 662213 16656 662226
rect 17290 662213 17314 662226
rect 17358 662213 17382 662226
rect 17426 662213 17450 662226
rect 17494 662213 17518 662226
rect 17562 662213 17586 662226
rect 17630 662213 17654 662226
rect 17698 662213 17722 662226
rect 17766 662213 17790 662226
rect 17834 662213 17858 662226
rect 17902 662213 17926 662226
rect 17970 662213 17994 662226
rect 18038 662213 18062 662226
rect 18106 662213 18130 662226
rect 18174 662213 18198 662226
rect 7389 661823 8389 661879
rect 8990 661823 9990 661879
rect 15678 661868 16678 661924
rect 17278 661868 18278 661924
rect 7389 661751 8389 661807
rect 8990 661751 9990 661807
rect 15678 661796 16678 661852
rect 17278 661796 18278 661852
rect 7389 661449 8389 661521
rect 8990 661449 9990 661521
rect 15678 661494 16678 661566
rect 17278 661494 18278 661566
rect 15748 661483 15782 661494
rect 15816 661483 15850 661494
rect 15884 661483 15918 661494
rect 15952 661483 15986 661494
rect 16020 661483 16054 661494
rect 16088 661483 16122 661494
rect 16156 661483 16190 661494
rect 16224 661483 16258 661494
rect 16292 661483 16326 661494
rect 16360 661483 16394 661494
rect 16428 661483 16462 661494
rect 16496 661483 16530 661494
rect 16564 661483 16598 661494
rect 16632 661483 16666 661494
rect 17290 661483 17324 661494
rect 17358 661483 17392 661494
rect 17426 661483 17460 661494
rect 17494 661483 17528 661494
rect 17562 661483 17596 661494
rect 17630 661483 17664 661494
rect 17698 661483 17732 661494
rect 17766 661483 17800 661494
rect 17834 661483 17868 661494
rect 17902 661483 17936 661494
rect 17970 661483 18004 661494
rect 18038 661483 18072 661494
rect 18106 661483 18140 661494
rect 18174 661483 18208 661494
rect 15748 661473 15806 661483
rect 15816 661473 15874 661483
rect 15884 661473 15942 661483
rect 15952 661473 16010 661483
rect 16020 661473 16078 661483
rect 16088 661473 16146 661483
rect 16156 661473 16214 661483
rect 16224 661473 16282 661483
rect 16292 661473 16350 661483
rect 16360 661473 16418 661483
rect 16428 661473 16486 661483
rect 16496 661473 16554 661483
rect 16564 661473 16622 661483
rect 16632 661473 16690 661483
rect 17290 661473 17348 661483
rect 17358 661473 17416 661483
rect 17426 661473 17484 661483
rect 17494 661473 17552 661483
rect 17562 661473 17620 661483
rect 17630 661473 17688 661483
rect 17698 661473 17756 661483
rect 17766 661473 17824 661483
rect 17834 661473 17892 661483
rect 17902 661473 17960 661483
rect 17970 661473 18028 661483
rect 18038 661473 18096 661483
rect 18106 661473 18164 661483
rect 18174 661473 18232 661483
rect 15724 661449 16690 661473
rect 17266 661449 18232 661473
rect 12427 661424 12493 661440
rect 15748 661434 15772 661449
rect 15816 661434 15840 661449
rect 15884 661434 15908 661449
rect 15952 661434 15976 661449
rect 16020 661434 16044 661449
rect 16088 661434 16112 661449
rect 16156 661434 16180 661449
rect 16224 661434 16248 661449
rect 16292 661434 16316 661449
rect 16360 661434 16384 661449
rect 16428 661434 16452 661449
rect 16496 661434 16520 661449
rect 16564 661434 16588 661449
rect 16632 661434 16656 661449
rect 17290 661434 17314 661449
rect 17358 661434 17382 661449
rect 17426 661434 17450 661449
rect 17494 661434 17518 661449
rect 17562 661434 17586 661449
rect 17630 661434 17654 661449
rect 17698 661434 17722 661449
rect 17766 661434 17790 661449
rect 17834 661434 17858 661449
rect 17902 661434 17926 661449
rect 17970 661434 17994 661449
rect 18038 661434 18062 661449
rect 18106 661434 18130 661449
rect 18174 661434 18198 661449
rect 15678 661279 16678 661434
rect 7389 661189 8389 661249
rect 8990 661189 9990 661249
rect 15678 661245 16690 661279
rect 17278 661269 18278 661434
rect 17266 661245 18278 661269
rect 15678 661234 16678 661245
rect 17278 661234 18278 661245
rect 15748 661221 15772 661234
rect 15816 661221 15840 661234
rect 15884 661221 15908 661234
rect 15952 661221 15976 661234
rect 16020 661221 16044 661234
rect 16088 661221 16112 661234
rect 16156 661221 16180 661234
rect 16224 661221 16248 661234
rect 16292 661221 16316 661234
rect 16360 661221 16384 661234
rect 16428 661221 16452 661234
rect 16496 661221 16520 661234
rect 16564 661221 16588 661234
rect 16632 661221 16656 661234
rect 17290 661221 17314 661234
rect 17358 661221 17382 661234
rect 17426 661221 17450 661234
rect 17494 661221 17518 661234
rect 17562 661221 17586 661234
rect 17630 661221 17654 661234
rect 17698 661221 17722 661234
rect 17766 661221 17790 661234
rect 17834 661221 17858 661234
rect 17902 661221 17926 661234
rect 17970 661221 17994 661234
rect 18038 661221 18062 661234
rect 18106 661221 18130 661234
rect 18174 661221 18198 661234
rect 7389 660831 8389 660887
rect 8990 660831 9990 660887
rect 15678 660876 16678 660932
rect 17278 660876 18278 660932
rect 7389 660759 8389 660815
rect 8990 660759 9990 660815
rect 15678 660804 16678 660860
rect 17278 660804 18278 660860
rect 7389 660457 8389 660529
rect 8990 660457 9990 660529
rect 15678 660502 16678 660574
rect 17278 660502 18278 660574
rect 15748 660491 15782 660502
rect 15816 660491 15850 660502
rect 15884 660491 15918 660502
rect 15952 660491 15986 660502
rect 16020 660491 16054 660502
rect 16088 660491 16122 660502
rect 16156 660491 16190 660502
rect 16224 660491 16258 660502
rect 16292 660491 16326 660502
rect 16360 660491 16394 660502
rect 16428 660491 16462 660502
rect 16496 660491 16530 660502
rect 16564 660491 16598 660502
rect 16632 660491 16666 660502
rect 17290 660491 17324 660502
rect 17358 660491 17392 660502
rect 17426 660491 17460 660502
rect 17494 660491 17528 660502
rect 17562 660491 17596 660502
rect 17630 660491 17664 660502
rect 17698 660491 17732 660502
rect 17766 660491 17800 660502
rect 17834 660491 17868 660502
rect 17902 660491 17936 660502
rect 17970 660491 18004 660502
rect 18038 660491 18072 660502
rect 18106 660491 18140 660502
rect 18174 660491 18208 660502
rect 15748 660481 15806 660491
rect 15816 660481 15874 660491
rect 15884 660481 15942 660491
rect 15952 660481 16010 660491
rect 16020 660481 16078 660491
rect 16088 660481 16146 660491
rect 16156 660481 16214 660491
rect 16224 660481 16282 660491
rect 16292 660481 16350 660491
rect 16360 660481 16418 660491
rect 16428 660481 16486 660491
rect 16496 660481 16554 660491
rect 16564 660481 16622 660491
rect 16632 660481 16690 660491
rect 17290 660481 17348 660491
rect 17358 660481 17416 660491
rect 17426 660481 17484 660491
rect 17494 660481 17552 660491
rect 17562 660481 17620 660491
rect 17630 660481 17688 660491
rect 17698 660481 17756 660491
rect 17766 660481 17824 660491
rect 17834 660481 17892 660491
rect 17902 660481 17960 660491
rect 17970 660481 18028 660491
rect 18038 660481 18096 660491
rect 18106 660481 18164 660491
rect 18174 660481 18232 660491
rect 15724 660457 16690 660481
rect 17266 660457 18232 660481
rect 15748 660442 15772 660457
rect 15816 660442 15840 660457
rect 15884 660442 15908 660457
rect 15952 660442 15976 660457
rect 16020 660442 16044 660457
rect 16088 660442 16112 660457
rect 16156 660442 16180 660457
rect 16224 660442 16248 660457
rect 16292 660442 16316 660457
rect 16360 660442 16384 660457
rect 16428 660442 16452 660457
rect 16496 660442 16520 660457
rect 16564 660442 16588 660457
rect 16632 660442 16656 660457
rect 17290 660442 17314 660457
rect 17358 660442 17382 660457
rect 17426 660442 17450 660457
rect 17494 660442 17518 660457
rect 17562 660442 17586 660457
rect 17630 660442 17654 660457
rect 17698 660442 17722 660457
rect 17766 660442 17790 660457
rect 17834 660442 17858 660457
rect 17902 660442 17926 660457
rect 17970 660442 17994 660457
rect 18038 660442 18062 660457
rect 18106 660442 18130 660457
rect 18174 660442 18198 660457
rect 15678 660287 16678 660442
rect 7389 660197 8389 660257
rect 8990 660197 9990 660257
rect 15678 660253 16690 660287
rect 17278 660277 18278 660442
rect 17266 660253 18278 660277
rect 15678 660242 16678 660253
rect 17278 660242 18278 660253
rect 15748 660229 15772 660242
rect 15816 660229 15840 660242
rect 15884 660229 15908 660242
rect 15952 660229 15976 660242
rect 16020 660229 16044 660242
rect 16088 660229 16112 660242
rect 16156 660229 16180 660242
rect 16224 660229 16248 660242
rect 16292 660229 16316 660242
rect 16360 660229 16384 660242
rect 16428 660229 16452 660242
rect 16496 660229 16520 660242
rect 16564 660229 16588 660242
rect 16632 660229 16656 660242
rect 17290 660229 17314 660242
rect 17358 660229 17382 660242
rect 17426 660229 17450 660242
rect 17494 660229 17518 660242
rect 17562 660229 17586 660242
rect 17630 660229 17654 660242
rect 17698 660229 17722 660242
rect 17766 660229 17790 660242
rect 17834 660229 17858 660242
rect 17902 660229 17926 660242
rect 17970 660229 17994 660242
rect 18038 660229 18062 660242
rect 18106 660229 18130 660242
rect 18174 660229 18198 660242
rect 7389 659839 8389 659895
rect 8990 659839 9990 659895
rect 15678 659884 16678 659940
rect 17278 659884 18278 659940
rect 7389 659767 8389 659823
rect 8990 659767 9990 659823
rect 15678 659812 16678 659868
rect 17278 659812 18278 659868
rect 7389 659465 8389 659537
rect 8990 659465 9990 659537
rect 15678 659510 16678 659582
rect 17278 659510 18278 659582
rect 15748 659499 15782 659510
rect 15816 659499 15850 659510
rect 15884 659499 15918 659510
rect 15952 659499 15986 659510
rect 16020 659499 16054 659510
rect 16088 659499 16122 659510
rect 16156 659499 16190 659510
rect 16224 659499 16258 659510
rect 16292 659499 16326 659510
rect 16360 659499 16394 659510
rect 16428 659499 16462 659510
rect 16496 659499 16530 659510
rect 16564 659499 16598 659510
rect 16632 659499 16666 659510
rect 17290 659499 17324 659510
rect 17358 659499 17392 659510
rect 17426 659499 17460 659510
rect 17494 659499 17528 659510
rect 17562 659499 17596 659510
rect 17630 659499 17664 659510
rect 17698 659499 17732 659510
rect 17766 659499 17800 659510
rect 17834 659499 17868 659510
rect 17902 659499 17936 659510
rect 17970 659499 18004 659510
rect 18038 659499 18072 659510
rect 18106 659499 18140 659510
rect 18174 659499 18208 659510
rect 15748 659489 15806 659499
rect 15816 659489 15874 659499
rect 15884 659489 15942 659499
rect 15952 659489 16010 659499
rect 16020 659489 16078 659499
rect 16088 659489 16146 659499
rect 16156 659489 16214 659499
rect 16224 659489 16282 659499
rect 16292 659489 16350 659499
rect 16360 659489 16418 659499
rect 16428 659489 16486 659499
rect 16496 659489 16554 659499
rect 16564 659489 16622 659499
rect 16632 659489 16690 659499
rect 17290 659489 17348 659499
rect 17358 659489 17416 659499
rect 17426 659489 17484 659499
rect 17494 659489 17552 659499
rect 17562 659489 17620 659499
rect 17630 659489 17688 659499
rect 17698 659489 17756 659499
rect 17766 659489 17824 659499
rect 17834 659489 17892 659499
rect 17902 659489 17960 659499
rect 17970 659489 18028 659499
rect 18038 659489 18096 659499
rect 18106 659489 18164 659499
rect 18174 659489 18232 659499
rect 15724 659465 16690 659489
rect 17266 659465 18232 659489
rect 15748 659450 15772 659465
rect 15816 659450 15840 659465
rect 15884 659450 15908 659465
rect 15952 659450 15976 659465
rect 16020 659450 16044 659465
rect 16088 659450 16112 659465
rect 16156 659450 16180 659465
rect 16224 659450 16248 659465
rect 16292 659450 16316 659465
rect 16360 659450 16384 659465
rect 16428 659450 16452 659465
rect 16496 659450 16520 659465
rect 16564 659450 16588 659465
rect 16632 659450 16656 659465
rect 17290 659450 17314 659465
rect 17358 659450 17382 659465
rect 17426 659450 17450 659465
rect 17494 659450 17518 659465
rect 17562 659450 17586 659465
rect 17630 659450 17654 659465
rect 17698 659450 17722 659465
rect 17766 659450 17790 659465
rect 17834 659450 17858 659465
rect 17902 659450 17926 659465
rect 17970 659450 17994 659465
rect 18038 659450 18062 659465
rect 18106 659450 18130 659465
rect 18174 659450 18198 659465
rect 15678 659295 16678 659450
rect 7389 659205 8389 659265
rect 8990 659205 9990 659265
rect 15678 659261 16690 659295
rect 17278 659285 18278 659450
rect 17266 659261 18278 659285
rect 15678 659250 16678 659261
rect 17278 659250 18278 659261
rect 15748 659237 15772 659250
rect 15816 659237 15840 659250
rect 15884 659237 15908 659250
rect 15952 659237 15976 659250
rect 16020 659237 16044 659250
rect 16088 659237 16112 659250
rect 16156 659237 16180 659250
rect 16224 659237 16248 659250
rect 16292 659237 16316 659250
rect 16360 659237 16384 659250
rect 16428 659237 16452 659250
rect 16496 659237 16520 659250
rect 16564 659237 16588 659250
rect 16632 659237 16656 659250
rect 17290 659237 17314 659250
rect 17358 659237 17382 659250
rect 17426 659237 17450 659250
rect 17494 659237 17518 659250
rect 17562 659237 17586 659250
rect 17630 659237 17654 659250
rect 17698 659237 17722 659250
rect 17766 659237 17790 659250
rect 17834 659237 17858 659250
rect 17902 659237 17926 659250
rect 17970 659237 17994 659250
rect 18038 659237 18062 659250
rect 18106 659237 18130 659250
rect 18174 659237 18198 659250
rect 7389 658847 8389 658903
rect 8990 658847 9990 658903
rect 15678 658892 16678 658948
rect 17278 658892 18278 658948
rect 7389 658775 8389 658831
rect 8990 658775 9990 658831
rect 15678 658820 16678 658876
rect 17278 658820 18278 658876
rect 5967 658455 6059 658489
rect 7389 658473 8389 658545
rect 8990 658473 9990 658545
rect 15678 658518 16678 658590
rect 17278 658518 18278 658590
rect 15748 658507 15782 658518
rect 15816 658507 15850 658518
rect 15884 658507 15918 658518
rect 15952 658507 15986 658518
rect 16020 658507 16054 658518
rect 16088 658507 16122 658518
rect 16156 658507 16190 658518
rect 16224 658507 16258 658518
rect 16292 658507 16326 658518
rect 16360 658507 16394 658518
rect 16428 658507 16462 658518
rect 16496 658507 16530 658518
rect 16564 658507 16598 658518
rect 16632 658507 16666 658518
rect 17290 658507 17324 658518
rect 17358 658507 17392 658518
rect 17426 658507 17460 658518
rect 17494 658507 17528 658518
rect 17562 658507 17596 658518
rect 17630 658507 17664 658518
rect 17698 658507 17732 658518
rect 17766 658507 17800 658518
rect 17834 658507 17868 658518
rect 17902 658507 17936 658518
rect 17970 658507 18004 658518
rect 18038 658507 18072 658518
rect 18106 658507 18140 658518
rect 18174 658507 18208 658518
rect 15748 658497 15806 658507
rect 15816 658497 15874 658507
rect 15884 658497 15942 658507
rect 15952 658497 16010 658507
rect 16020 658497 16078 658507
rect 16088 658497 16146 658507
rect 16156 658497 16214 658507
rect 16224 658497 16282 658507
rect 16292 658497 16350 658507
rect 16360 658497 16418 658507
rect 16428 658497 16486 658507
rect 16496 658497 16554 658507
rect 16564 658497 16622 658507
rect 16632 658497 16690 658507
rect 17290 658497 17348 658507
rect 17358 658497 17416 658507
rect 17426 658497 17484 658507
rect 17494 658497 17552 658507
rect 17562 658497 17620 658507
rect 17630 658497 17688 658507
rect 17698 658497 17756 658507
rect 17766 658497 17824 658507
rect 17834 658497 17892 658507
rect 17902 658497 17960 658507
rect 17970 658497 18028 658507
rect 18038 658497 18096 658507
rect 18106 658497 18164 658507
rect 18174 658497 18232 658507
rect 15724 658473 16690 658497
rect 17266 658473 18232 658497
rect 15748 658458 15772 658473
rect 15816 658458 15840 658473
rect 15884 658458 15908 658473
rect 15952 658458 15976 658473
rect 16020 658458 16044 658473
rect 16088 658458 16112 658473
rect 16156 658458 16180 658473
rect 16224 658458 16248 658473
rect 16292 658458 16316 658473
rect 16360 658458 16384 658473
rect 16428 658458 16452 658473
rect 16496 658458 16520 658473
rect 16564 658458 16588 658473
rect 16632 658458 16656 658473
rect 17290 658458 17314 658473
rect 17358 658458 17382 658473
rect 17426 658458 17450 658473
rect 17494 658458 17518 658473
rect 17562 658458 17586 658473
rect 17630 658458 17654 658473
rect 17698 658458 17722 658473
rect 17766 658458 17790 658473
rect 17834 658458 17858 658473
rect 17902 658458 17926 658473
rect 17970 658458 17994 658473
rect 18038 658458 18062 658473
rect 18106 658458 18130 658473
rect 18174 658458 18198 658473
rect 2850 658398 3850 658448
rect 2850 658282 3850 658332
rect 2850 658072 3850 658122
rect 2850 657956 3850 658006
rect 2850 657746 3850 657796
rect 1153 657660 1187 657718
rect 2850 657630 3850 657680
rect 2850 657420 3850 657470
rect 2850 657417 3107 657420
rect 3250 657304 3850 657354
rect 3250 657048 3850 657104
rect 3250 656892 3850 657020
rect 175 656818 1175 656868
rect 175 656662 1175 656790
rect 3250 656736 3850 656792
rect 175 656506 1175 656634
rect 175 656350 1175 656478
rect 175 656194 1175 656322
rect 175 656044 1175 656094
rect 175 655928 1175 655978
rect 175 655772 1175 655828
rect 175 655622 1175 655672
rect 1578 655609 1628 656609
rect 1728 655609 1856 656609
rect 1884 655609 2012 656609
rect 2040 655609 2090 656609
rect 3250 656580 3850 656708
rect 3250 656430 3850 656480
rect 2850 656314 3850 656364
rect 2850 656158 3850 656214
rect 2850 656008 3850 656058
rect 2850 655880 3850 655930
rect 2850 655724 3850 655852
rect 2850 655568 3850 655696
rect 175 655506 1175 655556
rect 175 655350 1175 655478
rect 2850 655412 3850 655468
rect 2850 655256 3850 655384
rect 175 655194 1175 655250
rect 175 655038 1175 655166
rect 175 654888 1175 654938
rect 175 654772 1175 654822
rect 175 654616 1175 654744
rect 1578 654613 1628 655213
rect 1728 654613 1784 655213
rect 1884 654613 1940 655213
rect 2040 654613 2096 655213
rect 2196 654613 2246 655213
rect 2850 655100 3850 655228
rect 2850 654944 3850 655072
rect 2850 654794 3850 654844
rect 2850 654678 3850 654728
rect 2850 654522 3850 654650
rect 175 654460 1175 654516
rect 175 654304 1175 654432
rect 2850 654366 3850 654494
rect 2850 654210 3850 654338
rect 175 654154 1175 654204
rect 803 654151 1175 654154
rect 2850 654054 3850 654110
rect 2850 653898 3850 654026
rect 2850 653742 3850 653870
rect 2850 653586 3850 653642
rect 2850 653436 3850 653486
rect 3926 653455 3960 653491
rect 3967 653339 3989 653455
rect 1638 651869 1688 652869
rect 1848 651869 1976 652869
rect 2064 651869 2114 652869
rect 2850 652275 3050 652287
rect 2850 652162 3850 652212
rect 2850 651946 3850 652074
rect 2850 651730 3850 651786
rect 2850 651514 3850 651642
rect 2850 651304 3850 651354
rect 2850 651188 3850 651238
rect 2850 650978 3850 651028
rect 3926 651015 3960 653339
rect 5169 651315 5191 658429
rect 5488 657194 5538 658194
rect 5658 657194 5708 658194
rect 5488 656073 5538 657073
rect 5658 656073 5708 657073
rect 5488 654952 5538 655952
rect 5658 654952 5708 655952
rect 5488 653842 5538 654842
rect 5658 653842 5708 654842
rect 5488 652721 5538 653721
rect 5658 652721 5708 653721
rect 5488 651600 5538 652600
rect 5658 651600 5708 652600
rect 5971 651386 6059 658455
rect 15678 658303 16678 658458
rect 7389 658213 8389 658273
rect 8990 658213 9990 658273
rect 15678 658269 16690 658303
rect 17278 658293 18278 658458
rect 17266 658269 18278 658293
rect 15678 658258 16678 658269
rect 17278 658258 18278 658269
rect 15748 658245 15772 658258
rect 15816 658245 15840 658258
rect 15884 658245 15908 658258
rect 15952 658245 15976 658258
rect 16020 658245 16044 658258
rect 16088 658245 16112 658258
rect 16156 658245 16180 658258
rect 16224 658245 16248 658258
rect 16292 658245 16316 658258
rect 16360 658245 16384 658258
rect 16428 658245 16452 658258
rect 16496 658245 16520 658258
rect 16564 658245 16588 658258
rect 16632 658245 16656 658258
rect 17290 658245 17314 658258
rect 17358 658245 17382 658258
rect 17426 658245 17450 658258
rect 17494 658245 17518 658258
rect 17562 658245 17586 658258
rect 17630 658245 17654 658258
rect 17698 658245 17722 658258
rect 17766 658245 17790 658258
rect 17834 658245 17858 658258
rect 17902 658245 17926 658258
rect 17970 658245 17994 658258
rect 18038 658245 18062 658258
rect 18106 658245 18130 658258
rect 18174 658245 18198 658258
rect 7389 657855 8389 657911
rect 8990 657855 9990 657911
rect 15678 657900 16678 657956
rect 17278 657900 18278 657956
rect 7389 657783 8389 657839
rect 8990 657783 9990 657839
rect 15678 657828 16678 657884
rect 17278 657828 18278 657884
rect 7389 657481 8389 657553
rect 8990 657481 9990 657553
rect 15678 657526 16678 657598
rect 17278 657526 18278 657598
rect 15748 657515 15782 657526
rect 15816 657515 15850 657526
rect 15884 657515 15918 657526
rect 15952 657515 15986 657526
rect 16020 657515 16054 657526
rect 16088 657515 16122 657526
rect 16156 657515 16190 657526
rect 16224 657515 16258 657526
rect 16292 657515 16326 657526
rect 16360 657515 16394 657526
rect 16428 657515 16462 657526
rect 16496 657515 16530 657526
rect 16564 657515 16598 657526
rect 16632 657515 16666 657526
rect 17290 657515 17324 657526
rect 17358 657515 17392 657526
rect 17426 657515 17460 657526
rect 17494 657515 17528 657526
rect 17562 657515 17596 657526
rect 17630 657515 17664 657526
rect 17698 657515 17732 657526
rect 17766 657515 17800 657526
rect 17834 657515 17868 657526
rect 17902 657515 17936 657526
rect 17970 657515 18004 657526
rect 18038 657515 18072 657526
rect 18106 657515 18140 657526
rect 18174 657515 18208 657526
rect 15748 657505 15806 657515
rect 15816 657505 15874 657515
rect 15884 657505 15942 657515
rect 15952 657505 16010 657515
rect 16020 657505 16078 657515
rect 16088 657505 16146 657515
rect 16156 657505 16214 657515
rect 16224 657505 16282 657515
rect 16292 657505 16350 657515
rect 16360 657505 16418 657515
rect 16428 657505 16486 657515
rect 16496 657505 16554 657515
rect 16564 657505 16622 657515
rect 16632 657505 16690 657515
rect 17290 657505 17348 657515
rect 17358 657505 17416 657515
rect 17426 657505 17484 657515
rect 17494 657505 17552 657515
rect 17562 657505 17620 657515
rect 17630 657505 17688 657515
rect 17698 657505 17756 657515
rect 17766 657505 17824 657515
rect 17834 657505 17892 657515
rect 17902 657505 17960 657515
rect 17970 657505 18028 657515
rect 18038 657505 18096 657515
rect 18106 657505 18164 657515
rect 18174 657505 18232 657515
rect 15724 657481 16690 657505
rect 17266 657481 18232 657505
rect 15748 657466 15772 657481
rect 15816 657466 15840 657481
rect 15884 657466 15908 657481
rect 15952 657466 15976 657481
rect 16020 657466 16044 657481
rect 16088 657466 16112 657481
rect 16156 657466 16180 657481
rect 16224 657466 16248 657481
rect 16292 657466 16316 657481
rect 16360 657466 16384 657481
rect 16428 657466 16452 657481
rect 16496 657466 16520 657481
rect 16564 657466 16588 657481
rect 16632 657466 16656 657481
rect 17290 657466 17314 657481
rect 17358 657466 17382 657481
rect 17426 657466 17450 657481
rect 17494 657466 17518 657481
rect 17562 657466 17586 657481
rect 17630 657466 17654 657481
rect 17698 657466 17722 657481
rect 17766 657466 17790 657481
rect 17834 657466 17858 657481
rect 17902 657466 17926 657481
rect 17970 657466 17994 657481
rect 18038 657466 18062 657481
rect 18106 657466 18130 657481
rect 18174 657466 18198 657481
rect 15678 657311 16678 657466
rect 7389 657221 8389 657281
rect 8990 657221 9990 657281
rect 15678 657277 16690 657311
rect 17278 657301 18278 657466
rect 17266 657277 18278 657301
rect 15678 657266 16678 657277
rect 17278 657266 18278 657277
rect 15748 657253 15772 657266
rect 15816 657253 15840 657266
rect 15884 657253 15908 657266
rect 15952 657253 15976 657266
rect 16020 657253 16044 657266
rect 16088 657253 16112 657266
rect 16156 657253 16180 657266
rect 16224 657253 16248 657266
rect 16292 657253 16316 657266
rect 16360 657253 16384 657266
rect 16428 657253 16452 657266
rect 16496 657253 16520 657266
rect 16564 657253 16588 657266
rect 16632 657253 16656 657266
rect 17290 657253 17314 657266
rect 17358 657253 17382 657266
rect 17426 657253 17450 657266
rect 17494 657253 17518 657266
rect 17562 657253 17586 657266
rect 17630 657253 17654 657266
rect 17698 657253 17722 657266
rect 17766 657253 17790 657266
rect 17834 657253 17858 657266
rect 17902 657253 17926 657266
rect 17970 657253 17994 657266
rect 18038 657253 18062 657266
rect 18106 657253 18130 657266
rect 18174 657253 18198 657266
rect 7389 656863 8389 656919
rect 8990 656863 9990 656919
rect 15678 656908 16678 656964
rect 17278 656908 18278 656964
rect 7389 656791 8389 656847
rect 8990 656791 9990 656847
rect 15678 656836 16678 656892
rect 17278 656836 18278 656892
rect 19480 656867 19516 663817
rect 19547 656867 19583 663817
rect 24572 663738 25172 663866
rect 36785 663864 37385 663920
rect 36785 663688 37385 663744
rect 20809 663650 20833 663684
rect 20809 663582 20833 663616
rect 24572 663588 25172 663638
rect 20809 663514 20833 663548
rect 36785 663518 37385 663568
rect 20809 663446 20833 663480
rect 24572 663458 25172 663508
rect 32930 663457 33530 663507
rect 20809 663378 20833 663412
rect 35287 663391 35887 663441
rect 36785 663402 37385 663452
rect 20809 663310 20833 663344
rect 24572 663308 25172 663358
rect 31463 663307 32063 663357
rect 32930 663301 33530 663357
rect 20809 663242 20833 663276
rect 35287 663215 35887 663343
rect 36785 663226 37385 663282
rect 20809 663174 20833 663208
rect 31463 663151 32063 663207
rect 32930 663151 33530 663201
rect 34079 663157 34679 663207
rect 20809 663106 20833 663140
rect 19844 662051 19894 663051
rect 19994 662051 20122 663051
rect 20150 662051 20278 663051
rect 20306 662051 20434 663051
rect 20462 662051 20512 663051
rect 20809 663038 20833 663072
rect 20809 662970 20833 663004
rect 20973 663000 21007 663024
rect 21041 663000 21075 663024
rect 21109 663000 21143 663024
rect 21177 663000 21211 663024
rect 21245 663000 21279 663024
rect 21313 663000 21347 663024
rect 21381 663000 21415 663024
rect 21449 663000 21483 663024
rect 21517 663000 21551 663024
rect 21585 663000 21619 663024
rect 21653 663000 21687 663024
rect 21721 663000 21755 663024
rect 21789 663000 21823 663024
rect 21857 663000 21891 663024
rect 21925 663000 21959 663024
rect 21993 663000 22027 663024
rect 22061 663000 22095 663024
rect 22129 663000 22163 663024
rect 22197 663000 22210 663024
rect 31463 663001 32063 663051
rect 34079 663001 34679 663057
rect 35287 663039 35887 663095
rect 36785 663050 37385 663106
rect 20809 662902 20833 662936
rect 32596 662929 33596 662979
rect 20809 662834 20833 662868
rect 24573 662820 25173 662870
rect 34079 662851 34679 662901
rect 35287 662869 35887 662919
rect 36785 662880 37385 662930
rect 35287 662866 35559 662869
rect 35716 662866 35887 662869
rect 20809 662766 20833 662800
rect 30171 662795 30771 662845
rect 20809 662698 20833 662732
rect 24573 662664 25173 662792
rect 32596 662773 33596 662829
rect 37993 662704 38593 662754
rect 19844 660521 19894 661921
rect 19994 660521 20122 661921
rect 20150 660521 20278 661921
rect 20306 660521 20434 661921
rect 20462 660521 20512 661921
rect 20809 660219 20833 660253
rect 19844 658759 19894 660159
rect 19994 658759 20122 660159
rect 20150 658759 20278 660159
rect 20306 658759 20434 660159
rect 20462 658759 20512 660159
rect 20809 660151 20833 660185
rect 20809 660083 20833 660117
rect 20809 660015 20833 660049
rect 20809 659947 20833 659981
rect 20809 659879 20833 659913
rect 20809 659811 20833 659845
rect 20809 659743 20833 659777
rect 20809 659675 20833 659709
rect 20809 659607 20833 659641
rect 20809 659539 20833 659573
rect 21263 659518 21313 662518
rect 21413 659518 21541 662518
rect 21569 659518 21697 662518
rect 21725 659518 21853 662518
rect 21881 659518 22009 662518
rect 22037 659518 22165 662518
rect 22193 659518 22321 662518
rect 22349 659518 22399 662518
rect 24573 662508 25173 662636
rect 30171 662619 30771 662675
rect 32596 662623 33596 662673
rect 34110 662589 34710 662639
rect 36785 662620 36797 662624
rect 36785 662609 36800 662620
rect 36970 662609 36985 662624
rect 26348 662530 26372 662564
rect 32596 662507 33596 662557
rect 26348 662461 26372 662495
rect 30171 662449 30771 662499
rect 24573 662352 25173 662408
rect 24573 662196 25173 662324
rect 29993 662310 30993 662360
rect 32596 662351 33596 662479
rect 34110 662433 34710 662561
rect 36785 662429 36985 662609
rect 37993 662534 38593 662584
rect 36785 662418 36800 662429
rect 36785 662414 36797 662418
rect 36970 662414 36985 662429
rect 31347 662317 31362 662332
rect 31535 662328 31547 662332
rect 31532 662317 31547 662328
rect 24573 662040 25173 662168
rect 26490 662122 26690 662172
rect 29993 662160 30993 662210
rect 31347 662137 31547 662317
rect 31347 662122 31362 662137
rect 31532 662126 31547 662137
rect 31535 662122 31547 662126
rect 31607 662317 31622 662332
rect 31795 662328 31807 662332
rect 31792 662317 31807 662328
rect 31607 662137 31807 662317
rect 32596 662195 33596 662323
rect 34110 662277 34710 662405
rect 36785 662384 36797 662388
rect 36785 662373 36800 662384
rect 36970 662373 36985 662388
rect 31607 662122 31622 662137
rect 31792 662126 31807 662137
rect 31795 662122 31807 662126
rect 31347 662081 31362 662096
rect 31535 662092 31547 662096
rect 31532 662081 31547 662092
rect 22906 661855 23212 662025
rect 23406 661855 23712 662025
rect 26490 661966 26690 662022
rect 29993 662001 30993 662051
rect 24573 661890 25173 661940
rect 31347 661901 31547 662081
rect 26490 661816 26690 661866
rect 29993 661851 30993 661901
rect 31347 661886 31362 661901
rect 31532 661890 31547 661901
rect 31535 661886 31547 661890
rect 31607 662081 31622 662096
rect 31795 662092 31807 662096
rect 31792 662081 31807 662092
rect 31607 661901 31807 662081
rect 32596 662039 33596 662167
rect 34110 662121 34710 662249
rect 36785 662193 36985 662373
rect 36785 662182 36800 662193
rect 36785 662178 36797 662182
rect 36970 662178 36985 662193
rect 37083 662373 37098 662388
rect 37083 662193 37120 662373
rect 37083 662178 37098 662193
rect 37998 662108 38598 662158
rect 34110 661971 34710 662021
rect 31607 661886 31622 661901
rect 31792 661890 31807 661901
rect 31795 661886 31807 661890
rect 32596 661883 33596 661939
rect 37998 661932 38598 661988
rect 34110 661855 34710 661905
rect 24573 661760 25173 661810
rect 27691 661682 28291 661732
rect 30253 661721 30268 661736
rect 30441 661732 30453 661736
rect 30438 661721 30453 661732
rect 24573 661610 25173 661660
rect 27691 661532 28291 661582
rect 30253 661541 30453 661721
rect 30253 661526 30268 661541
rect 30438 661530 30453 661541
rect 30441 661526 30453 661530
rect 30513 661721 30528 661736
rect 30701 661732 30713 661736
rect 30698 661721 30713 661732
rect 30513 661541 30713 661721
rect 30513 661526 30528 661541
rect 30698 661530 30713 661541
rect 30701 661526 30713 661530
rect 30773 661721 30788 661736
rect 30961 661732 30973 661736
rect 30958 661721 30973 661732
rect 30773 661541 30973 661721
rect 30773 661526 30788 661541
rect 30958 661530 30973 661541
rect 30961 661526 30973 661530
rect 31087 661721 31102 661736
rect 31275 661732 31287 661736
rect 31272 661721 31287 661732
rect 31087 661541 31287 661721
rect 31087 661526 31102 661541
rect 31272 661530 31287 661541
rect 31275 661526 31287 661530
rect 31347 661721 31362 661736
rect 31535 661732 31547 661736
rect 31532 661721 31547 661732
rect 31347 661541 31547 661721
rect 31347 661526 31362 661541
rect 31532 661530 31547 661541
rect 31535 661526 31547 661530
rect 31607 661721 31622 661736
rect 31795 661732 31807 661736
rect 31792 661721 31807 661732
rect 31607 661541 31807 661721
rect 31607 661526 31622 661541
rect 31792 661530 31807 661541
rect 31795 661526 31807 661530
rect 31867 661721 31882 661736
rect 32055 661732 32067 661736
rect 32052 661721 32067 661732
rect 32596 661727 33596 661855
rect 31867 661541 32067 661721
rect 34110 661699 34710 661827
rect 37998 661762 38598 661812
rect 37998 661759 38220 661762
rect 38245 661759 38539 661762
rect 32596 661571 33596 661699
rect 34110 661543 34710 661671
rect 31867 661526 31882 661541
rect 32052 661530 32067 661541
rect 32055 661526 32067 661530
rect 22619 661446 22647 661474
rect 24573 661438 25173 661488
rect 26490 661416 26690 661466
rect 27691 661402 28291 661452
rect 32596 661415 33596 661543
rect 34110 661387 34710 661515
rect 24573 661288 25173 661338
rect 26490 661260 26690 661316
rect 27691 661246 28291 661374
rect 30253 661361 30268 661376
rect 30441 661372 30453 661376
rect 30438 661361 30453 661372
rect 30253 661331 30453 661361
rect 30253 661316 30268 661331
rect 30438 661320 30453 661331
rect 30441 661316 30453 661320
rect 30513 661361 30528 661376
rect 30701 661372 30713 661376
rect 30698 661361 30713 661372
rect 30513 661331 30713 661361
rect 30513 661316 30528 661331
rect 30698 661320 30713 661331
rect 30701 661316 30713 661320
rect 30773 661361 30788 661376
rect 31347 661361 31362 661376
rect 31535 661372 31547 661376
rect 31532 661361 31547 661372
rect 30773 661331 30793 661361
rect 31347 661331 31547 661361
rect 30773 661316 30788 661331
rect 31347 661316 31362 661331
rect 31532 661320 31547 661331
rect 31535 661316 31547 661320
rect 31607 661361 31622 661376
rect 31795 661372 31807 661376
rect 31792 661361 31807 661372
rect 31607 661331 31807 661361
rect 31607 661316 31622 661331
rect 31792 661320 31807 661331
rect 31795 661316 31807 661320
rect 31867 661361 31882 661376
rect 31867 661331 31921 661361
rect 31867 661316 31882 661331
rect 30253 661275 30268 661290
rect 30441 661286 30453 661290
rect 30438 661275 30453 661286
rect 30253 661245 30453 661275
rect 30253 661230 30268 661245
rect 30438 661234 30453 661245
rect 30441 661230 30453 661234
rect 30513 661275 30528 661290
rect 30701 661286 30713 661290
rect 30698 661275 30713 661286
rect 30513 661245 30713 661275
rect 30513 661230 30528 661245
rect 30698 661234 30713 661245
rect 30701 661230 30713 661234
rect 30773 661275 30788 661290
rect 31347 661275 31362 661290
rect 31535 661286 31547 661290
rect 31532 661275 31547 661286
rect 30773 661245 30793 661275
rect 31347 661245 31547 661275
rect 30773 661230 30788 661245
rect 31347 661230 31362 661245
rect 31532 661234 31547 661245
rect 31535 661230 31547 661234
rect 31607 661275 31622 661290
rect 31795 661286 31807 661290
rect 31792 661275 31807 661286
rect 31607 661245 31807 661275
rect 31607 661230 31622 661245
rect 31792 661234 31807 661245
rect 31795 661230 31807 661234
rect 31867 661275 31882 661290
rect 31867 661245 31921 661275
rect 32596 661265 33596 661315
rect 31867 661230 31882 661245
rect 34110 661231 34710 661287
rect 22906 661055 23212 661225
rect 23406 661055 23712 661225
rect 24573 661158 25173 661208
rect 24573 661002 25173 661130
rect 26490 661107 26690 661160
rect 27691 661090 28291 661218
rect 31823 661084 32061 661118
rect 31481 661080 32061 661084
rect 31481 661068 31797 661080
rect 32596 661063 33596 661113
rect 34110 661075 34710 661203
rect 37998 661133 38148 661145
rect 38317 661133 38467 661145
rect 24573 660846 25173 660974
rect 27691 660934 28291 660990
rect 32596 660907 33596 661035
rect 34110 660919 34710 661047
rect 37998 661020 38598 661070
rect 27691 660778 28291 660906
rect 25286 660758 25310 660762
rect 32596 660751 33596 660879
rect 34110 660763 34710 660891
rect 37998 660844 38598 660900
rect 24573 660690 25173 660746
rect 25286 660687 25310 660721
rect 24573 660534 25173 660662
rect 25286 660615 25310 660649
rect 27691 660622 28291 660750
rect 32596 660595 33596 660723
rect 35287 660695 35487 660707
rect 37998 660674 38598 660724
rect 34110 660607 34710 660663
rect 36785 660650 36797 660654
rect 36785 660639 36800 660650
rect 36970 660639 36985 660654
rect 35134 660582 35734 660632
rect 25286 660543 25310 660577
rect 22906 660255 23212 660425
rect 23406 660255 23712 660425
rect 24573 660378 25173 660506
rect 25286 660471 25310 660505
rect 27691 660472 28291 660522
rect 32596 660439 33596 660567
rect 34110 660451 34710 660507
rect 35134 660432 35734 660482
rect 36785 660459 36985 660639
rect 36785 660448 36800 660459
rect 36785 660444 36797 660448
rect 36970 660444 36985 660459
rect 37083 660639 37098 660654
rect 37083 660459 37120 660639
rect 37083 660444 37098 660459
rect 36785 660414 36797 660418
rect 32596 660283 33596 660411
rect 36785 660403 36800 660414
rect 36970 660403 36985 660418
rect 34110 660295 34710 660351
rect 35134 660316 35734 660366
rect 24573 660228 25173 660278
rect 32596 660127 33596 660255
rect 34110 660145 34710 660195
rect 35134 660160 35734 660288
rect 32596 659971 33596 660099
rect 34110 660029 34710 660079
rect 35134 660004 35734 660132
rect 31481 659862 31797 659880
rect 34110 659873 34710 660001
rect 31823 659828 32061 659860
rect 32596 659821 33596 659871
rect 35134 659848 35734 659976
rect 36071 659805 36098 660295
rect 36785 660223 36985 660403
rect 37993 660248 38593 660298
rect 36785 660212 36800 660223
rect 36785 660208 36797 660212
rect 36970 660208 36985 660223
rect 696597 660200 696600 660320
rect 37993 660078 38593 660128
rect 692376 659983 692396 660017
rect 692463 659993 692532 660017
rect 696191 659993 696239 660017
rect 692487 659983 692532 659993
rect 696204 659983 696239 659993
rect 696340 659983 696360 660017
rect 36785 659902 37385 659952
rect 692487 659915 692502 659939
rect 696200 659915 696215 659939
rect 692454 659891 692478 659915
rect 696224 659891 696248 659915
rect 686755 659800 687355 659850
rect 34110 659717 34710 659773
rect 30253 659701 30268 659716
rect 30441 659712 30453 659716
rect 30438 659701 30453 659712
rect 30253 659671 30453 659701
rect 30253 659656 30268 659671
rect 30438 659660 30453 659671
rect 30441 659656 30453 659660
rect 30513 659701 30528 659716
rect 30701 659712 30713 659716
rect 30698 659701 30713 659712
rect 30513 659671 30713 659701
rect 30513 659656 30528 659671
rect 30698 659660 30713 659671
rect 30701 659656 30713 659660
rect 30773 659701 30788 659716
rect 31347 659701 31362 659716
rect 31535 659712 31547 659716
rect 31532 659701 31547 659712
rect 30773 659671 30793 659701
rect 31347 659671 31547 659701
rect 30773 659656 30788 659671
rect 31347 659656 31362 659671
rect 31532 659660 31547 659671
rect 31535 659656 31547 659660
rect 31607 659701 31622 659716
rect 31795 659712 31807 659716
rect 31792 659701 31807 659712
rect 31607 659671 31807 659701
rect 31607 659656 31622 659671
rect 31792 659660 31807 659671
rect 31795 659656 31807 659660
rect 31867 659701 31882 659716
rect 31867 659671 31921 659701
rect 35134 659698 35734 659770
rect 36785 659726 37385 659782
rect 692487 659748 692505 659752
rect 692479 659718 692505 659748
rect 692487 659698 692505 659718
rect 31867 659656 31882 659671
rect 30253 659615 30268 659630
rect 30441 659626 30453 659630
rect 30438 659615 30453 659626
rect 30253 659585 30453 659615
rect 30253 659570 30268 659585
rect 30438 659574 30453 659585
rect 30441 659570 30453 659574
rect 30513 659615 30528 659630
rect 30701 659626 30713 659630
rect 30698 659615 30713 659626
rect 30513 659585 30713 659615
rect 30513 659570 30528 659585
rect 30698 659574 30713 659585
rect 30701 659570 30713 659574
rect 30773 659615 30788 659630
rect 31347 659615 31362 659630
rect 31535 659626 31547 659630
rect 31532 659615 31547 659626
rect 30773 659585 30793 659615
rect 31347 659585 31547 659615
rect 30773 659570 30788 659585
rect 31347 659570 31362 659585
rect 31532 659574 31547 659585
rect 31535 659570 31547 659574
rect 31607 659615 31622 659630
rect 31795 659626 31807 659630
rect 31792 659615 31807 659626
rect 31607 659585 31807 659615
rect 31607 659570 31622 659585
rect 31792 659574 31807 659585
rect 31795 659570 31807 659574
rect 31867 659615 31882 659630
rect 32546 659619 33546 659669
rect 31867 659585 31921 659615
rect 31867 659570 31882 659585
rect 20809 659471 20833 659505
rect 32546 659463 33546 659591
rect 34110 659561 34710 659689
rect 35134 659645 36134 659695
rect 686755 659624 687355 659680
rect 692485 659674 692505 659698
rect 692509 659674 692517 659718
rect 696215 659698 696223 659748
rect 696203 659674 696223 659698
rect 696227 659674 696245 659752
rect 692485 659640 692521 659674
rect 696203 659640 696249 659674
rect 35134 659489 36134 659617
rect 36785 659550 37385 659606
rect 20809 659403 20833 659437
rect 30253 659405 30268 659420
rect 30441 659416 30453 659420
rect 30438 659405 30453 659416
rect 20809 659335 20833 659369
rect 20809 659267 20833 659301
rect 20809 659199 20833 659233
rect 30253 659225 30453 659405
rect 30253 659210 30268 659225
rect 30438 659214 30453 659225
rect 30441 659210 30453 659214
rect 30513 659405 30528 659420
rect 30701 659416 30713 659420
rect 30698 659405 30713 659416
rect 30513 659225 30713 659405
rect 30513 659210 30528 659225
rect 30698 659214 30713 659225
rect 30701 659210 30713 659214
rect 30773 659405 30788 659420
rect 30961 659416 30973 659420
rect 30958 659405 30973 659416
rect 30773 659225 30973 659405
rect 30773 659210 30788 659225
rect 30958 659214 30973 659225
rect 30961 659210 30973 659214
rect 31087 659405 31102 659420
rect 31275 659416 31287 659420
rect 31272 659405 31287 659416
rect 31087 659225 31287 659405
rect 31087 659210 31102 659225
rect 31272 659214 31287 659225
rect 31275 659210 31287 659214
rect 31347 659405 31362 659420
rect 31535 659416 31547 659420
rect 31532 659405 31547 659416
rect 31347 659225 31547 659405
rect 31347 659210 31362 659225
rect 31532 659214 31547 659225
rect 31535 659210 31547 659214
rect 31607 659405 31622 659420
rect 31795 659416 31807 659420
rect 31792 659405 31807 659416
rect 31607 659225 31807 659405
rect 31607 659210 31622 659225
rect 31792 659214 31807 659225
rect 31795 659210 31807 659214
rect 31867 659405 31882 659420
rect 32055 659416 32067 659420
rect 32052 659405 32067 659416
rect 31867 659225 32067 659405
rect 32546 659307 33546 659435
rect 34110 659411 34710 659461
rect 686755 659448 687355 659504
rect 35134 659339 36134 659389
rect 36785 659380 37385 659430
rect 31867 659210 31882 659225
rect 32052 659214 32067 659225
rect 32055 659210 32067 659214
rect 20809 659131 20833 659165
rect 32546 659151 33546 659279
rect 36785 659248 37385 659298
rect 686755 659278 687355 659328
rect 35285 659162 35319 659172
rect 35353 659162 35387 659172
rect 35421 659162 35455 659172
rect 35489 659162 35523 659172
rect 35564 659162 35598 659172
rect 35632 659162 35666 659172
rect 35700 659162 35734 659172
rect 35768 659162 35802 659172
rect 35836 659162 35870 659172
rect 35904 659162 35938 659172
rect 35972 659162 36006 659172
rect 36040 659162 36074 659172
rect 36108 659162 36142 659172
rect 36176 659162 36210 659172
rect 35255 659126 36255 659138
rect 20809 659063 20833 659097
rect 20940 659085 20983 659103
rect 20940 659069 20949 659085
rect 20974 659069 20983 659085
rect 25113 659069 25349 659093
rect 25383 659069 25417 659093
rect 20974 659051 21008 659069
rect 20809 658995 20833 659029
rect 20974 659028 21003 659051
rect 21361 659045 21409 659069
rect 20949 659027 20983 659028
rect 21385 658991 21409 659045
rect 25113 658991 25137 659069
rect 29993 659045 30993 659095
rect 31347 659045 31362 659060
rect 31535 659056 31547 659060
rect 31532 659045 31547 659056
rect 21361 658967 21409 658991
rect 25089 658967 25137 658991
rect 20809 658927 20833 658961
rect 20809 658859 20833 658893
rect 20809 658791 20833 658825
rect 20809 658723 20833 658757
rect 20809 658655 20833 658689
rect 21413 658638 22813 658681
rect 23685 658638 25085 658681
rect 19844 657229 19894 658629
rect 19994 657229 20122 658629
rect 20150 657229 20278 658629
rect 20306 657229 20434 658629
rect 20462 657229 20512 658629
rect 20809 658587 20833 658621
rect 20809 658519 20833 658553
rect 20809 658451 20833 658485
rect 21413 658475 22813 658603
rect 23685 658475 25085 658603
rect 20809 658383 20833 658417
rect 20809 658315 20833 658349
rect 21413 658312 22813 658440
rect 23685 658312 25085 658440
rect 20809 658247 20833 658281
rect 20809 658179 20833 658213
rect 21413 658149 22813 658277
rect 23685 658149 25085 658277
rect 20809 658111 20833 658145
rect 20809 658043 20833 658077
rect 20809 657975 20833 658009
rect 21413 657986 22813 658114
rect 23685 657986 25085 658114
rect 20809 657907 20833 657941
rect 20809 657839 20833 657873
rect 21413 657823 22813 657951
rect 23685 657823 25085 657951
rect 20809 657771 20833 657805
rect 20809 657703 20833 657737
rect 21413 657673 22813 657716
rect 23685 657673 25085 657716
rect 20809 657635 20833 657669
rect 20809 657567 20833 657601
rect 21361 657552 21419 657586
rect 25089 657552 25147 657586
rect 20809 657499 20833 657533
rect 20809 657431 20833 657465
rect 20809 657363 20833 657397
rect 21361 657373 21419 657397
rect 25089 657373 25147 657397
rect 21385 657363 21419 657373
rect 25113 657363 25147 657373
rect 20809 657295 20833 657329
rect 21385 657291 21419 657325
rect 25113 657291 25147 657325
rect 20809 657227 20833 657261
rect 21385 657219 21419 657253
rect 25113 657219 25147 657253
rect 20809 657159 20833 657193
rect 21385 657171 21419 657181
rect 25113 657171 25147 657181
rect 21361 657147 21419 657171
rect 25089 657147 25147 657171
rect 20809 657091 20833 657125
rect 20809 657023 20833 657057
rect 20809 656955 20833 656989
rect 21361 656969 21409 656993
rect 25089 656969 25137 656993
rect 20809 656887 20833 656921
rect 21385 656915 21409 656969
rect 25113 656915 25137 656969
rect 21361 656891 21409 656915
rect 25089 656891 25137 656915
rect 19480 656831 19583 656867
rect 21413 656754 22813 656804
rect 23685 656754 25085 656804
rect 7389 656489 8389 656561
rect 8990 656489 9990 656561
rect 15678 656534 16678 656606
rect 17278 656534 18278 656606
rect 21413 656591 22813 656719
rect 23685 656591 25085 656719
rect 15748 656523 15782 656534
rect 15816 656523 15850 656534
rect 15884 656523 15918 656534
rect 15952 656523 15986 656534
rect 16020 656523 16054 656534
rect 16088 656523 16122 656534
rect 16156 656523 16190 656534
rect 16224 656523 16258 656534
rect 16292 656523 16326 656534
rect 16360 656523 16394 656534
rect 16428 656523 16462 656534
rect 16496 656523 16530 656534
rect 16564 656523 16598 656534
rect 16632 656523 16666 656534
rect 17290 656523 17324 656534
rect 17358 656523 17392 656534
rect 17426 656523 17460 656534
rect 17494 656523 17528 656534
rect 17562 656523 17596 656534
rect 17630 656523 17664 656534
rect 17698 656523 17732 656534
rect 17766 656523 17800 656534
rect 17834 656523 17868 656534
rect 17902 656523 17936 656534
rect 17970 656523 18004 656534
rect 18038 656523 18072 656534
rect 18106 656523 18140 656534
rect 18174 656523 18208 656534
rect 15748 656513 15806 656523
rect 15816 656513 15874 656523
rect 15884 656513 15942 656523
rect 15952 656513 16010 656523
rect 16020 656513 16078 656523
rect 16088 656513 16146 656523
rect 16156 656513 16214 656523
rect 16224 656513 16282 656523
rect 16292 656513 16350 656523
rect 16360 656513 16418 656523
rect 16428 656513 16486 656523
rect 16496 656513 16554 656523
rect 16564 656513 16622 656523
rect 16632 656513 16690 656523
rect 17290 656513 17348 656523
rect 17358 656513 17416 656523
rect 17426 656513 17484 656523
rect 17494 656513 17552 656523
rect 17562 656513 17620 656523
rect 17630 656513 17688 656523
rect 17698 656513 17756 656523
rect 17766 656513 17824 656523
rect 17834 656513 17892 656523
rect 17902 656513 17960 656523
rect 17970 656513 18028 656523
rect 18038 656513 18096 656523
rect 18106 656513 18164 656523
rect 18174 656513 18232 656523
rect 15724 656489 16690 656513
rect 17266 656489 18232 656513
rect 15748 656474 15772 656489
rect 15816 656474 15840 656489
rect 15884 656474 15908 656489
rect 15952 656474 15976 656489
rect 16020 656474 16044 656489
rect 16088 656474 16112 656489
rect 16156 656474 16180 656489
rect 16224 656474 16248 656489
rect 16292 656474 16316 656489
rect 16360 656474 16384 656489
rect 16428 656474 16452 656489
rect 16496 656474 16520 656489
rect 16564 656474 16588 656489
rect 16632 656474 16656 656489
rect 17290 656474 17314 656489
rect 17358 656474 17382 656489
rect 17426 656474 17450 656489
rect 17494 656474 17518 656489
rect 17562 656474 17586 656489
rect 17630 656474 17654 656489
rect 17698 656474 17722 656489
rect 17766 656474 17790 656489
rect 17834 656474 17858 656489
rect 17902 656474 17926 656489
rect 17970 656474 17994 656489
rect 18038 656474 18062 656489
rect 18106 656474 18130 656489
rect 18174 656474 18198 656489
rect 15678 656319 16678 656474
rect 7389 656229 8389 656289
rect 8990 656229 9990 656289
rect 15678 656285 16690 656319
rect 17278 656309 18278 656474
rect 21413 656428 22813 656556
rect 23685 656428 25085 656556
rect 17266 656285 18278 656309
rect 15678 656274 16678 656285
rect 17278 656274 18278 656285
rect 15748 656261 15772 656274
rect 15816 656261 15840 656274
rect 15884 656261 15908 656274
rect 15952 656261 15976 656274
rect 16020 656261 16044 656274
rect 16088 656261 16112 656274
rect 16156 656261 16180 656274
rect 16224 656261 16248 656274
rect 16292 656261 16316 656274
rect 16360 656261 16384 656274
rect 16428 656261 16452 656274
rect 16496 656261 16520 656274
rect 16564 656261 16588 656274
rect 16632 656261 16656 656274
rect 17290 656261 17314 656274
rect 17358 656261 17382 656274
rect 17426 656261 17450 656274
rect 17494 656261 17518 656274
rect 17562 656261 17586 656274
rect 17630 656261 17654 656274
rect 17698 656261 17722 656274
rect 17766 656261 17790 656274
rect 17834 656261 17858 656274
rect 17902 656261 17926 656274
rect 17970 656261 17994 656274
rect 18038 656261 18062 656274
rect 18106 656261 18130 656274
rect 18174 656261 18198 656274
rect 21413 656265 22813 656393
rect 23685 656265 25085 656393
rect 21413 656102 22813 656230
rect 23685 656102 25085 656230
rect 7389 655871 8389 655927
rect 8990 655871 9990 655927
rect 15678 655916 16678 655972
rect 17278 655916 18278 655972
rect 21413 655952 22813 655995
rect 23685 655952 25085 655995
rect 7389 655799 8389 655855
rect 8990 655799 9990 655855
rect 15678 655844 16678 655900
rect 17278 655844 18278 655900
rect 21406 655865 21430 655889
rect 25068 655865 25092 655889
rect 21382 655841 21385 655865
rect 25113 655841 25116 655865
rect 21382 655763 21396 655787
rect 25102 655763 25116 655787
rect 21348 655739 21372 655763
rect 21406 655739 21430 655763
rect 25068 655739 25092 655763
rect 25126 655739 25150 655763
rect 25524 655703 25548 659001
rect 29993 658895 30993 658945
rect 31347 658865 31547 659045
rect 31347 658850 31362 658865
rect 31532 658854 31547 658865
rect 31535 658850 31547 658854
rect 31607 659045 31622 659060
rect 31795 659056 31807 659060
rect 31792 659045 31807 659056
rect 31607 658865 31807 659045
rect 32546 658995 33546 659123
rect 36785 659072 37385 659128
rect 685547 659102 686147 659152
rect 35255 659019 36255 659069
rect 687155 659007 687170 659022
rect 687343 659018 687355 659022
rect 687340 659007 687355 659018
rect 31607 658850 31622 658865
rect 31792 658854 31807 658865
rect 31795 658850 31807 658854
rect 32546 658839 33546 658967
rect 35255 658843 36255 658971
rect 36785 658896 37385 658952
rect 685547 658932 686147 658982
rect 687155 658827 687355 659007
rect 31347 658809 31362 658824
rect 31535 658820 31547 658824
rect 31532 658809 31547 658820
rect 29993 658736 30993 658786
rect 29993 658586 30993 658636
rect 31347 658629 31547 658809
rect 31347 658614 31362 658629
rect 31532 658618 31547 658629
rect 31535 658614 31547 658618
rect 31607 658809 31622 658824
rect 31795 658820 31807 658824
rect 31792 658809 31807 658820
rect 687155 658812 687170 658827
rect 687340 658816 687355 658827
rect 687343 658812 687355 658816
rect 31607 658629 31807 658809
rect 32546 658683 33546 658811
rect 35255 658667 36255 658795
rect 36785 658726 37385 658776
rect 687042 658771 687057 658786
rect 31607 658614 31622 658629
rect 31792 658618 31807 658629
rect 31795 658614 31807 658618
rect 32546 658527 33546 658655
rect 37993 658550 38593 658600
rect 687020 658591 687057 658771
rect 687042 658576 687057 658591
rect 687155 658771 687170 658786
rect 687343 658782 687355 658786
rect 687340 658771 687355 658782
rect 687155 658591 687355 658771
rect 688210 658630 688260 659630
rect 688360 658630 688488 659630
rect 688516 658630 688644 659630
rect 688672 658630 688800 659630
rect 688828 658630 688956 659630
rect 688984 658630 689112 659630
rect 689140 658630 689268 659630
rect 689296 658630 689424 659630
rect 689452 658630 689580 659630
rect 689608 658630 689736 659630
rect 689764 658630 689892 659630
rect 689920 658630 690048 659630
rect 690076 658630 690204 659630
rect 690232 658630 690360 659630
rect 690388 658630 690438 659630
rect 692485 659606 692505 659640
rect 692509 659606 692517 659640
rect 696203 659606 696223 659640
rect 696227 659606 696245 659640
rect 691275 659523 691875 659573
rect 692485 659572 692521 659606
rect 696203 659572 696249 659606
rect 692485 659538 692505 659572
rect 692509 659538 692517 659572
rect 692485 659504 692521 659538
rect 692583 659528 693983 659571
rect 694719 659528 696119 659571
rect 696203 659538 696223 659572
rect 696227 659538 696245 659572
rect 696203 659504 696249 659538
rect 692485 659470 692505 659504
rect 692509 659470 692517 659504
rect 692485 659436 692521 659470
rect 691275 659373 691875 659423
rect 692485 659402 692505 659436
rect 692509 659402 692517 659436
rect 692485 659368 692521 659402
rect 692485 659334 692505 659368
rect 692509 659334 692517 659368
rect 692583 659365 693983 659493
rect 694719 659365 696119 659493
rect 696203 659470 696223 659504
rect 696227 659470 696245 659504
rect 696203 659436 696249 659470
rect 707624 659441 707658 659475
rect 707695 659441 707729 659475
rect 707769 659441 707803 659475
rect 707840 659441 707874 659475
rect 707914 659441 707948 659475
rect 707985 659441 708019 659475
rect 708059 659441 708093 659475
rect 708130 659441 708164 659475
rect 708204 659441 708238 659475
rect 708275 659441 708309 659475
rect 708369 659441 708403 659475
rect 708446 659441 708480 659475
rect 708520 659441 708554 659465
rect 708588 659441 708610 659465
rect 709211 659441 709234 659465
rect 709270 659441 709304 659475
rect 709364 659441 709398 659475
rect 709435 659441 709469 659475
rect 709509 659441 709543 659475
rect 709580 659441 709614 659475
rect 709654 659441 709688 659475
rect 709725 659441 709759 659475
rect 709799 659441 709833 659475
rect 709870 659441 709904 659475
rect 709944 659441 709978 659475
rect 710015 659441 710049 659475
rect 710089 659441 710123 659475
rect 710160 659441 710194 659475
rect 696203 659402 696223 659436
rect 696227 659402 696245 659436
rect 707610 659431 707624 659441
rect 707658 659431 707695 659441
rect 707729 659431 707769 659441
rect 707803 659431 707840 659441
rect 707874 659431 707914 659441
rect 707948 659431 707985 659441
rect 708019 659431 708059 659441
rect 708093 659431 708130 659441
rect 708164 659431 708204 659441
rect 708238 659431 708275 659441
rect 708309 659431 708369 659441
rect 708403 659431 708446 659441
rect 708480 659431 708520 659441
rect 708554 659431 708588 659441
rect 708610 659431 708634 659441
rect 709211 659431 709270 659441
rect 709304 659431 709364 659441
rect 709398 659431 709435 659441
rect 709469 659431 709509 659441
rect 709543 659431 709580 659441
rect 709614 659431 709654 659441
rect 709688 659431 709725 659441
rect 709759 659431 709799 659441
rect 709833 659431 709870 659441
rect 709904 659431 709944 659441
rect 709978 659431 710015 659441
rect 710049 659431 710089 659441
rect 710123 659431 710160 659441
rect 710194 659431 710211 659441
rect 696203 659368 696249 659402
rect 696203 659334 696223 659368
rect 696227 659334 696245 659368
rect 707610 659337 708610 659431
rect 709211 659337 710211 659431
rect 691275 659251 691875 659301
rect 692485 659300 692521 659334
rect 692485 659266 692505 659300
rect 692509 659266 692517 659300
rect 692485 659232 692521 659266
rect 692485 659198 692505 659232
rect 692509 659198 692517 659232
rect 692583 659202 693983 659330
rect 694719 659202 696119 659330
rect 696203 659300 696249 659334
rect 711579 659317 712463 659331
rect 711579 659307 711619 659317
rect 696203 659266 696223 659300
rect 696227 659266 696245 659300
rect 701730 659290 701747 659292
rect 696203 659232 696249 659266
rect 696203 659198 696223 659232
rect 696227 659198 696245 659232
rect 701692 659220 701722 659254
rect 701730 659220 701760 659290
rect 707610 659241 708610 659301
rect 709211 659241 710211 659301
rect 692485 659164 692521 659198
rect 691275 659101 691875 659151
rect 692485 659130 692505 659164
rect 692509 659130 692517 659164
rect 692485 659096 692521 659130
rect 692485 659062 692505 659096
rect 692509 659062 692517 659096
rect 692485 659028 692521 659062
rect 692583 659039 693983 659167
rect 694719 659039 696119 659167
rect 696203 659164 696249 659198
rect 696203 659130 696223 659164
rect 696227 659130 696245 659164
rect 696203 659096 696249 659130
rect 696203 659062 696223 659096
rect 696227 659062 696245 659096
rect 699322 659064 700322 659097
rect 700922 659064 701922 659097
rect 696203 659028 696249 659062
rect 707610 659044 708610 659048
rect 709211 659044 710211 659048
rect 691275 658975 691875 659025
rect 692485 658994 692505 659028
rect 692509 658994 692517 659028
rect 692485 658960 692521 658994
rect 692485 658926 692505 658960
rect 692509 658926 692517 658960
rect 692485 658892 692521 658926
rect 691275 658825 691875 658875
rect 692485 658858 692505 658892
rect 692509 658858 692517 658892
rect 692583 658876 693983 659004
rect 694719 658876 696119 659004
rect 696203 658994 696223 659028
rect 696227 658994 696245 659028
rect 707574 658994 708646 659030
rect 696203 658960 696249 658994
rect 696203 658926 696223 658960
rect 696227 658926 696245 658960
rect 707574 658953 707610 658994
rect 708610 658953 708646 658994
rect 696203 658892 696249 658926
rect 697284 658894 697350 658910
rect 707574 658897 708646 658953
rect 696203 658858 696223 658892
rect 696227 658858 696245 658892
rect 699322 658877 700322 658894
rect 700922 658877 701922 658894
rect 707574 658881 707610 658897
rect 708610 658881 708646 658897
rect 692485 658824 692521 658858
rect 692485 658790 692505 658824
rect 692509 658790 692517 658824
rect 692485 658756 692521 658790
rect 691275 658703 691875 658753
rect 692485 658722 692505 658756
rect 692509 658722 692517 658756
rect 692485 658688 692521 658722
rect 692583 658713 693983 658841
rect 694719 658713 696119 658841
rect 696203 658824 696249 658858
rect 707574 658825 708646 658881
rect 696203 658790 696223 658824
rect 696227 658790 696245 658824
rect 696203 658756 696249 658790
rect 696203 658722 696223 658756
rect 696227 658722 696245 658756
rect 699322 658739 700322 658811
rect 700922 658739 701922 658811
rect 707574 658788 707610 658825
rect 708610 658788 708646 658825
rect 707574 658748 708646 658788
rect 709175 658994 710247 659030
rect 709175 658953 709211 658994
rect 710211 658953 710247 658994
rect 709175 658897 710247 658953
rect 709175 658881 709211 658897
rect 710211 658881 710247 658897
rect 709175 658825 710247 658881
rect 709175 658788 709211 658825
rect 710211 658788 710247 658825
rect 709175 658748 710247 658788
rect 696203 658688 696249 658722
rect 692485 658654 692505 658688
rect 692509 658654 692517 658688
rect 692485 658620 692521 658654
rect 687155 658576 687170 658591
rect 687340 658580 687355 658591
rect 687343 658576 687355 658580
rect 28647 658450 28671 658477
rect 30171 658447 30771 658497
rect 35255 658491 36255 658547
rect 685542 658506 686142 658556
rect 691275 658553 691875 658603
rect 692485 658586 692505 658620
rect 692509 658586 692517 658620
rect 692485 658552 692521 658586
rect 692485 658518 692505 658552
rect 692509 658518 692517 658552
rect 692583 658550 693983 658678
rect 694719 658550 696119 658678
rect 696203 658654 696223 658688
rect 696227 658654 696245 658688
rect 696203 658620 696249 658654
rect 696203 658586 696223 658620
rect 696227 658586 696245 658620
rect 696203 658552 696249 658586
rect 696203 658518 696223 658552
rect 696227 658518 696245 658552
rect 692485 658484 692521 658518
rect 36785 658466 36797 658470
rect 36785 658455 36800 658466
rect 36970 658455 36985 658470
rect 28683 658397 28717 658431
rect 32546 658377 33546 658427
rect 28683 658328 28717 658362
rect 28683 658259 28717 658293
rect 30171 658271 30771 658327
rect 35255 658321 36255 658371
rect 36785 658275 36985 658455
rect 692485 658450 692505 658484
rect 692509 658450 692517 658484
rect 37993 658380 38593 658430
rect 692485 658416 692521 658450
rect 679817 658330 679841 658354
rect 685542 658330 686142 658386
rect 692485 658382 692505 658416
rect 692509 658382 692517 658416
rect 692583 658387 693983 658515
rect 694719 658387 696119 658515
rect 696203 658484 696249 658518
rect 696203 658450 696223 658484
rect 696227 658450 696245 658484
rect 699322 658478 700322 658550
rect 700922 658478 701922 658550
rect 707610 658523 708610 658595
rect 709211 658523 710211 658595
rect 699392 658467 699426 658478
rect 699460 658467 699494 658478
rect 699528 658467 699562 658478
rect 699596 658467 699630 658478
rect 699664 658467 699698 658478
rect 699732 658467 699766 658478
rect 699800 658467 699834 658478
rect 699868 658467 699902 658478
rect 699936 658467 699970 658478
rect 700004 658467 700038 658478
rect 700072 658467 700106 658478
rect 700140 658467 700174 658478
rect 700208 658467 700242 658478
rect 700276 658467 700310 658478
rect 700934 658467 700968 658478
rect 701002 658467 701036 658478
rect 701070 658467 701104 658478
rect 701138 658467 701172 658478
rect 701206 658467 701240 658478
rect 701274 658467 701308 658478
rect 701342 658467 701376 658478
rect 701410 658467 701444 658478
rect 701478 658467 701512 658478
rect 701546 658467 701580 658478
rect 701614 658467 701648 658478
rect 701682 658467 701716 658478
rect 701750 658467 701784 658478
rect 701818 658467 701852 658478
rect 699392 658457 699450 658467
rect 699460 658457 699518 658467
rect 699528 658457 699586 658467
rect 699596 658457 699654 658467
rect 699664 658457 699722 658467
rect 699732 658457 699790 658467
rect 699800 658457 699858 658467
rect 699868 658457 699926 658467
rect 699936 658457 699994 658467
rect 700004 658457 700062 658467
rect 700072 658457 700130 658467
rect 700140 658457 700198 658467
rect 700208 658457 700266 658467
rect 700276 658457 700334 658467
rect 700934 658457 700992 658467
rect 701002 658457 701060 658467
rect 701070 658457 701128 658467
rect 701138 658457 701196 658467
rect 701206 658457 701264 658467
rect 701274 658457 701332 658467
rect 701342 658457 701400 658467
rect 701410 658457 701468 658467
rect 701478 658457 701536 658467
rect 701546 658457 701604 658467
rect 701614 658457 701672 658467
rect 701682 658457 701740 658467
rect 701750 658457 701808 658467
rect 701818 658457 701876 658467
rect 696203 658416 696249 658450
rect 699368 658433 700334 658457
rect 700910 658433 701876 658457
rect 699392 658418 699416 658433
rect 699460 658418 699484 658433
rect 699528 658418 699552 658433
rect 699596 658418 699620 658433
rect 699664 658418 699688 658433
rect 699732 658418 699756 658433
rect 699800 658418 699824 658433
rect 699868 658418 699892 658433
rect 699936 658418 699960 658433
rect 700004 658418 700028 658433
rect 700072 658418 700096 658433
rect 700140 658418 700164 658433
rect 700208 658418 700232 658433
rect 700276 658418 700300 658433
rect 700934 658418 700958 658433
rect 701002 658418 701026 658433
rect 701070 658418 701094 658433
rect 701138 658418 701162 658433
rect 701206 658418 701230 658433
rect 701274 658418 701298 658433
rect 701342 658418 701366 658433
rect 701410 658418 701434 658433
rect 701478 658418 701502 658433
rect 701546 658418 701570 658433
rect 701614 658418 701638 658433
rect 701682 658418 701706 658433
rect 701750 658418 701774 658433
rect 701818 658418 701842 658433
rect 696203 658382 696223 658416
rect 696227 658382 696245 658416
rect 692485 658348 692521 658382
rect 696203 658348 696249 658382
rect 679549 658307 679573 658330
rect 679793 658306 679808 658330
rect 692485 658314 692505 658348
rect 692509 658314 692517 658348
rect 696203 658314 696223 658348
rect 696227 658314 696245 658348
rect 36785 658264 36800 658275
rect 36785 658260 36797 658264
rect 36970 658260 36985 658275
rect 692485 658280 692521 658314
rect 696203 658280 696249 658314
rect 679549 658237 679573 658271
rect 692485 658246 692505 658280
rect 692509 658246 692517 658280
rect 36785 658230 36797 658234
rect 28683 658190 28717 658224
rect 32596 658175 33596 658225
rect 35359 658156 35375 658222
rect 36143 658156 36159 658222
rect 36785 658219 36800 658230
rect 36970 658219 36985 658234
rect 28683 658121 28717 658155
rect 30171 658101 30771 658151
rect 28683 658052 28717 658086
rect 32596 658019 33596 658147
rect 28683 657983 28717 658017
rect 33959 657994 33975 658060
rect 36143 657994 36159 658060
rect 36785 658039 36985 658219
rect 36785 658028 36800 658039
rect 36785 658024 36797 658028
rect 36970 658024 36985 658039
rect 37083 658219 37098 658234
rect 37083 658039 37120 658219
rect 692485 658212 692521 658246
rect 692583 658237 693983 658280
rect 694719 658237 696119 658280
rect 696203 658246 696223 658280
rect 696227 658246 696245 658280
rect 699322 658263 700322 658418
rect 696203 658212 696249 658246
rect 699322 658229 700334 658263
rect 700922 658253 701922 658418
rect 700910 658229 701922 658253
rect 699322 658218 700322 658229
rect 700922 658218 701922 658229
rect 707574 658263 708646 658299
rect 707574 658226 707610 658263
rect 708610 658226 708646 658263
rect 679549 658167 679573 658201
rect 685542 658160 686142 658210
rect 685601 658157 685895 658160
rect 685920 658157 686142 658160
rect 692485 658178 692505 658212
rect 692509 658178 692517 658212
rect 696203 658178 696223 658212
rect 696227 658178 696245 658212
rect 699392 658205 699416 658218
rect 699460 658205 699484 658218
rect 699528 658205 699552 658218
rect 699596 658205 699620 658218
rect 699664 658205 699688 658218
rect 699732 658205 699756 658218
rect 699800 658205 699824 658218
rect 699868 658205 699892 658218
rect 699936 658205 699960 658218
rect 700004 658205 700028 658218
rect 700072 658205 700096 658218
rect 700140 658205 700164 658218
rect 700208 658205 700232 658218
rect 700276 658205 700300 658218
rect 700934 658205 700958 658218
rect 701002 658205 701026 658218
rect 701070 658205 701094 658218
rect 701138 658205 701162 658218
rect 701206 658205 701230 658218
rect 701274 658205 701298 658218
rect 701342 658205 701366 658218
rect 701410 658205 701434 658218
rect 701478 658205 701502 658218
rect 701546 658205 701570 658218
rect 701614 658205 701638 658218
rect 701682 658205 701706 658218
rect 701750 658205 701774 658218
rect 701818 658205 701842 658218
rect 707574 658186 708646 658226
rect 709175 658263 710247 658299
rect 709175 658226 709211 658263
rect 710211 658226 710247 658263
rect 709175 658186 710247 658226
rect 692485 658144 692521 658178
rect 696203 658144 696249 658178
rect 679549 658097 679573 658131
rect 692485 658110 692505 658144
rect 692509 658110 692517 658144
rect 692485 658076 692521 658110
rect 692583 658101 693983 658144
rect 694719 658101 696119 658144
rect 696203 658110 696223 658144
rect 696227 658110 696245 658144
rect 696203 658076 696249 658110
rect 37083 658024 37098 658039
rect 679549 658027 679573 658061
rect 692485 658042 692505 658076
rect 692509 658042 692517 658076
rect 692485 658008 692521 658042
rect 28683 657914 28717 657948
rect 31463 657895 32063 657945
rect 28683 657845 28717 657879
rect 32596 657863 33596 657991
rect 37998 657954 38598 658004
rect 679549 657957 679573 657991
rect 692485 657974 692505 658008
rect 692509 657974 692517 658008
rect 679793 657933 679808 657957
rect 692485 657940 692521 657974
rect 679817 657909 679841 657933
rect 692485 657906 692505 657940
rect 692509 657906 692517 657940
rect 692583 657938 693983 658066
rect 694719 657938 696119 658066
rect 696203 658042 696223 658076
rect 696227 658042 696245 658076
rect 696203 658008 696249 658042
rect 696203 657974 696223 658008
rect 696227 657974 696245 658008
rect 696203 657940 696249 657974
rect 696203 657906 696223 657940
rect 696227 657906 696245 657940
rect 28683 657776 28717 657810
rect 28683 657707 28717 657741
rect 31463 657739 32063 657795
rect 32596 657707 33596 657835
rect 33959 657832 33975 657898
rect 36143 657832 36159 657898
rect 687685 657838 687709 657862
rect 37998 657778 38598 657834
rect 687661 657814 687675 657838
rect 687669 657797 687675 657814
rect 679515 657762 679539 657785
rect 679613 657762 679637 657785
rect 679491 657737 679515 657761
rect 679637 657737 679661 657761
rect 28683 657638 28717 657672
rect 28683 657569 28717 657603
rect 31463 657589 32063 657639
rect 32596 657551 33596 657679
rect 35359 657670 35375 657736
rect 36143 657670 36159 657736
rect 680215 657678 680815 657728
rect 37998 657608 38598 657658
rect 37998 657605 38220 657608
rect 38245 657605 38539 657608
rect 28683 657500 28717 657534
rect 28683 657431 28717 657465
rect 28683 657362 28717 657396
rect 32596 657395 33596 657523
rect 35255 657521 36255 657571
rect 680215 657502 680815 657558
rect 685551 657516 686551 657566
rect 28683 657293 28717 657327
rect 28683 657224 28717 657258
rect 30015 657256 30718 657272
rect 30015 657246 30721 657256
rect 28683 657155 28717 657189
rect 28683 657086 28717 657120
rect 28683 657017 28717 657051
rect 28683 656948 28717 656982
rect 28683 656879 28717 656913
rect 28683 656810 28717 656844
rect 28683 656741 28717 656775
rect 28683 656672 28717 656706
rect 28683 656603 28717 656637
rect 28683 656534 28717 656568
rect 28683 656465 28717 656499
rect 28683 656396 28717 656430
rect 28682 656361 28683 656366
rect 28682 656332 28717 656361
rect 28647 656303 28671 656332
rect 28647 656234 28671 656268
rect 28647 656165 28671 656199
rect 28647 656096 28671 656130
rect 28647 656027 28671 656061
rect 28647 655958 28671 655992
rect 28647 655889 28671 655923
rect 28647 655820 28671 655854
rect 28647 655751 28671 655785
rect 28647 655682 28671 655716
rect 29778 655695 29802 655719
rect 29802 655671 29826 655683
rect 29880 655681 29914 655715
rect 25524 655635 25548 655669
rect 7389 655497 8389 655569
rect 8990 655497 9990 655569
rect 15678 655542 16678 655614
rect 17278 655542 18278 655614
rect 28647 655613 28671 655647
rect 29778 655635 29802 655659
rect 21361 655586 21409 655610
rect 25089 655586 25137 655610
rect 15748 655531 15782 655542
rect 15816 655531 15850 655542
rect 15884 655531 15918 655542
rect 15952 655531 15986 655542
rect 16020 655531 16054 655542
rect 16088 655531 16122 655542
rect 16156 655531 16190 655542
rect 16224 655531 16258 655542
rect 16292 655531 16326 655542
rect 16360 655531 16394 655542
rect 16428 655531 16462 655542
rect 16496 655531 16530 655542
rect 16564 655531 16598 655542
rect 16632 655531 16666 655542
rect 17290 655531 17324 655542
rect 17358 655531 17392 655542
rect 17426 655531 17460 655542
rect 17494 655531 17528 655542
rect 17562 655531 17596 655542
rect 17630 655531 17664 655542
rect 17698 655531 17732 655542
rect 17766 655531 17800 655542
rect 17834 655531 17868 655542
rect 17902 655531 17936 655542
rect 17970 655531 18004 655542
rect 18038 655531 18072 655542
rect 18106 655531 18140 655542
rect 18174 655531 18208 655542
rect 21385 655532 21409 655586
rect 25113 655532 25137 655586
rect 28647 655544 28671 655578
rect 15748 655521 15806 655531
rect 15816 655521 15874 655531
rect 15884 655521 15942 655531
rect 15952 655521 16010 655531
rect 16020 655521 16078 655531
rect 16088 655521 16146 655531
rect 16156 655521 16214 655531
rect 16224 655521 16282 655531
rect 16292 655521 16350 655531
rect 16360 655521 16418 655531
rect 16428 655521 16486 655531
rect 16496 655521 16554 655531
rect 16564 655521 16622 655531
rect 16632 655521 16690 655531
rect 17290 655521 17348 655531
rect 17358 655521 17416 655531
rect 17426 655521 17484 655531
rect 17494 655521 17552 655531
rect 17562 655521 17620 655531
rect 17630 655521 17688 655531
rect 17698 655521 17756 655531
rect 17766 655521 17824 655531
rect 17834 655521 17892 655531
rect 17902 655521 17960 655531
rect 17970 655521 18028 655531
rect 18038 655521 18096 655531
rect 18106 655521 18164 655531
rect 18174 655521 18232 655531
rect 15724 655497 16690 655521
rect 17266 655497 18232 655521
rect 21361 655508 21409 655532
rect 25089 655508 25137 655532
rect 15748 655482 15772 655497
rect 15816 655482 15840 655497
rect 15884 655482 15908 655497
rect 15952 655482 15976 655497
rect 16020 655482 16044 655497
rect 16088 655482 16112 655497
rect 16156 655482 16180 655497
rect 16224 655482 16248 655497
rect 16292 655482 16316 655497
rect 16360 655482 16384 655497
rect 16428 655482 16452 655497
rect 16496 655482 16520 655497
rect 16564 655482 16588 655497
rect 16632 655482 16656 655497
rect 17290 655482 17314 655497
rect 17358 655482 17382 655497
rect 17426 655482 17450 655497
rect 17494 655482 17518 655497
rect 17562 655482 17586 655497
rect 17630 655482 17654 655497
rect 17698 655482 17722 655497
rect 17766 655482 17790 655497
rect 17834 655482 17858 655497
rect 17902 655482 17926 655497
rect 17970 655482 17994 655497
rect 18038 655482 18062 655497
rect 18106 655482 18130 655497
rect 18174 655482 18198 655497
rect 7389 655237 8389 655297
rect 8990 655237 9990 655297
rect 12559 655273 12865 655375
rect 15678 655327 16678 655482
rect 15678 655293 16690 655327
rect 17278 655317 18278 655482
rect 28647 655475 28671 655509
rect 28647 655406 28671 655440
rect 28647 655337 28671 655371
rect 17266 655293 18278 655317
rect 15678 655282 16678 655293
rect 17278 655282 18278 655293
rect 12543 655257 12881 655273
rect 15748 655269 15772 655282
rect 15816 655269 15840 655282
rect 15884 655269 15908 655282
rect 15952 655269 15976 655282
rect 16020 655269 16044 655282
rect 16088 655269 16112 655282
rect 16156 655269 16180 655282
rect 16224 655269 16248 655282
rect 16292 655269 16316 655282
rect 16360 655269 16384 655282
rect 16428 655269 16452 655282
rect 16496 655269 16520 655282
rect 16564 655269 16588 655282
rect 16632 655269 16656 655282
rect 17290 655269 17314 655282
rect 17358 655269 17382 655282
rect 17426 655269 17450 655282
rect 17494 655269 17518 655282
rect 17562 655269 17586 655282
rect 17630 655269 17654 655282
rect 17698 655269 17722 655282
rect 17766 655269 17790 655282
rect 17834 655269 17858 655282
rect 17902 655269 17926 655282
rect 17970 655269 17994 655282
rect 18038 655269 18062 655282
rect 18106 655269 18130 655282
rect 18174 655269 18198 655282
rect 19980 655048 20286 655218
rect 7389 654879 8389 654935
rect 8990 654879 9990 654935
rect 15678 654924 16678 654980
rect 17278 654924 18278 654980
rect 7389 654807 8389 654863
rect 8990 654807 9990 654863
rect 15678 654852 16678 654908
rect 17278 654852 18278 654908
rect 20945 654796 25553 655332
rect 28647 655268 28671 655302
rect 28647 655199 28671 655233
rect 28647 655154 28671 655164
rect 21413 654706 22813 654796
rect 23685 654706 25085 654796
rect 7389 654505 8389 654577
rect 8990 654505 9990 654577
rect 15678 654550 16678 654622
rect 17278 654550 18278 654622
rect 15748 654539 15782 654550
rect 15816 654539 15850 654550
rect 15884 654539 15918 654550
rect 15952 654539 15986 654550
rect 16020 654539 16054 654550
rect 16088 654539 16122 654550
rect 16156 654539 16190 654550
rect 16224 654539 16258 654550
rect 16292 654539 16326 654550
rect 16360 654539 16394 654550
rect 16428 654539 16462 654550
rect 16496 654539 16530 654550
rect 16564 654539 16598 654550
rect 16632 654539 16666 654550
rect 17290 654539 17324 654550
rect 17358 654539 17392 654550
rect 17426 654539 17460 654550
rect 17494 654539 17528 654550
rect 17562 654539 17596 654550
rect 17630 654539 17664 654550
rect 17698 654539 17732 654550
rect 17766 654539 17800 654550
rect 17834 654539 17868 654550
rect 17902 654539 17936 654550
rect 17970 654539 18004 654550
rect 18038 654539 18072 654550
rect 18106 654539 18140 654550
rect 18174 654539 18208 654550
rect 21413 654543 22813 654671
rect 23685 654543 25085 654671
rect 15748 654529 15806 654539
rect 15816 654529 15874 654539
rect 15884 654529 15942 654539
rect 15952 654529 16010 654539
rect 16020 654529 16078 654539
rect 16088 654529 16146 654539
rect 16156 654529 16214 654539
rect 16224 654529 16282 654539
rect 16292 654529 16350 654539
rect 16360 654529 16418 654539
rect 16428 654529 16486 654539
rect 16496 654529 16554 654539
rect 16564 654529 16622 654539
rect 16632 654529 16690 654539
rect 17290 654529 17348 654539
rect 17358 654529 17416 654539
rect 17426 654529 17484 654539
rect 17494 654529 17552 654539
rect 17562 654529 17620 654539
rect 17630 654529 17688 654539
rect 17698 654529 17756 654539
rect 17766 654529 17824 654539
rect 17834 654529 17892 654539
rect 17902 654529 17960 654539
rect 17970 654529 18028 654539
rect 18038 654529 18096 654539
rect 18106 654529 18164 654539
rect 18174 654529 18232 654539
rect 15724 654505 16690 654529
rect 17266 654505 18232 654529
rect 15748 654490 15772 654505
rect 15816 654490 15840 654505
rect 15884 654490 15908 654505
rect 15952 654490 15976 654505
rect 16020 654490 16044 654505
rect 16088 654490 16112 654505
rect 16156 654490 16180 654505
rect 16224 654490 16248 654505
rect 16292 654490 16316 654505
rect 16360 654490 16384 654505
rect 16428 654490 16452 654505
rect 16496 654490 16520 654505
rect 16564 654490 16588 654505
rect 16632 654490 16656 654505
rect 17290 654490 17314 654505
rect 17358 654490 17382 654505
rect 17426 654490 17450 654505
rect 17494 654490 17518 654505
rect 17562 654490 17586 654505
rect 17630 654490 17654 654505
rect 17698 654490 17722 654505
rect 17766 654490 17790 654505
rect 17834 654490 17858 654505
rect 17902 654490 17926 654505
rect 17970 654490 17994 654505
rect 18038 654490 18062 654505
rect 18106 654490 18130 654505
rect 18174 654490 18198 654505
rect 15678 654335 16678 654490
rect 7389 654245 8389 654305
rect 8990 654245 9990 654305
rect 15678 654301 16690 654335
rect 17278 654325 18278 654490
rect 21413 654380 22813 654508
rect 23685 654380 25085 654508
rect 17266 654301 18278 654325
rect 15678 654290 16678 654301
rect 17278 654290 18278 654301
rect 15748 654277 15772 654290
rect 15816 654277 15840 654290
rect 15884 654277 15908 654290
rect 15952 654277 15976 654290
rect 16020 654277 16044 654290
rect 16088 654277 16112 654290
rect 16156 654277 16180 654290
rect 16224 654277 16248 654290
rect 16292 654277 16316 654290
rect 16360 654277 16384 654290
rect 16428 654277 16452 654290
rect 16496 654277 16520 654290
rect 16564 654277 16588 654290
rect 16632 654277 16656 654290
rect 17290 654277 17314 654290
rect 17358 654277 17382 654290
rect 17426 654277 17450 654290
rect 17494 654277 17518 654290
rect 17562 654277 17586 654290
rect 17630 654277 17654 654290
rect 17698 654277 17722 654290
rect 17766 654277 17790 654290
rect 17834 654277 17858 654290
rect 17902 654277 17926 654290
rect 17970 654277 17994 654290
rect 18038 654277 18062 654290
rect 18106 654277 18130 654290
rect 18174 654277 18198 654290
rect 21413 654217 22813 654345
rect 23685 654217 25085 654345
rect 21413 654054 22813 654182
rect 23685 654054 25085 654182
rect 25936 654132 26936 654182
rect 27274 654033 27358 654036
rect 13899 653998 14059 654002
rect 7389 653887 8389 653943
rect 8990 653887 9990 653943
rect 15678 653932 16678 653988
rect 17278 653932 18278 653988
rect 7389 653815 8389 653871
rect 8990 653815 9990 653871
rect 15678 653860 16678 653916
rect 17278 653860 18278 653916
rect 21413 653891 22813 654019
rect 23685 653891 25085 654019
rect 25936 653976 26936 654032
rect 27158 653983 27358 654033
rect 13899 653852 14059 653856
rect 25936 653820 26936 653876
rect 27158 653807 27358 653935
rect 21413 653741 22813 653784
rect 23685 653741 25085 653784
rect 25936 653664 26936 653720
rect 7389 653513 8389 653585
rect 8990 653513 9990 653585
rect 15678 653558 16678 653630
rect 17278 653558 18278 653630
rect 21413 653605 22813 653648
rect 23685 653605 25085 653648
rect 27158 653631 27358 653687
rect 15748 653547 15782 653558
rect 15816 653547 15850 653558
rect 15884 653547 15918 653558
rect 15952 653547 15986 653558
rect 16020 653547 16054 653558
rect 16088 653547 16122 653558
rect 16156 653547 16190 653558
rect 16224 653547 16258 653558
rect 16292 653547 16326 653558
rect 16360 653547 16394 653558
rect 16428 653547 16462 653558
rect 16496 653547 16530 653558
rect 16564 653547 16598 653558
rect 16632 653547 16666 653558
rect 17290 653547 17324 653558
rect 17358 653547 17392 653558
rect 17426 653547 17460 653558
rect 17494 653547 17528 653558
rect 17562 653547 17596 653558
rect 17630 653547 17664 653558
rect 17698 653547 17732 653558
rect 17766 653547 17800 653558
rect 17834 653547 17868 653558
rect 17902 653547 17936 653558
rect 17970 653547 18004 653558
rect 18038 653547 18072 653558
rect 18106 653547 18140 653558
rect 18174 653547 18208 653558
rect 15748 653537 15806 653547
rect 15816 653537 15874 653547
rect 15884 653537 15942 653547
rect 15952 653537 16010 653547
rect 16020 653537 16078 653547
rect 16088 653537 16146 653547
rect 16156 653537 16214 653547
rect 16224 653537 16282 653547
rect 16292 653537 16350 653547
rect 16360 653537 16418 653547
rect 16428 653537 16486 653547
rect 16496 653537 16554 653547
rect 16564 653537 16622 653547
rect 16632 653537 16690 653547
rect 17290 653537 17348 653547
rect 17358 653537 17416 653547
rect 17426 653537 17484 653547
rect 17494 653537 17552 653547
rect 17562 653537 17620 653547
rect 17630 653537 17688 653547
rect 17698 653537 17756 653547
rect 17766 653537 17824 653547
rect 17834 653537 17892 653547
rect 17902 653537 17960 653547
rect 17970 653537 18028 653547
rect 18038 653537 18096 653547
rect 18106 653537 18164 653547
rect 18174 653537 18232 653547
rect 15724 653513 16690 653537
rect 17266 653513 18232 653537
rect 15748 653498 15772 653513
rect 15816 653498 15840 653513
rect 15884 653498 15908 653513
rect 15952 653498 15976 653513
rect 16020 653498 16044 653513
rect 16088 653498 16112 653513
rect 16156 653498 16180 653513
rect 16224 653498 16248 653513
rect 16292 653498 16316 653513
rect 16360 653498 16384 653513
rect 16428 653498 16452 653513
rect 16496 653498 16520 653513
rect 16564 653498 16588 653513
rect 16632 653498 16656 653513
rect 17290 653498 17314 653513
rect 17358 653498 17382 653513
rect 17426 653498 17450 653513
rect 17494 653498 17518 653513
rect 17562 653498 17586 653513
rect 17630 653498 17654 653513
rect 17698 653498 17722 653513
rect 17766 653498 17790 653513
rect 17834 653498 17858 653513
rect 17902 653498 17926 653513
rect 17970 653498 17994 653513
rect 18038 653498 18062 653513
rect 18106 653498 18130 653513
rect 18174 653498 18198 653513
rect 15678 653343 16678 653498
rect 7389 653253 8389 653313
rect 8990 653253 9990 653313
rect 15678 653309 16690 653343
rect 17278 653333 18278 653498
rect 21413 653442 22813 653570
rect 23685 653442 25085 653570
rect 25936 653514 26936 653564
rect 26393 653511 26477 653514
rect 26726 653511 26810 653514
rect 27158 653455 27358 653583
rect 17266 653309 18278 653333
rect 15678 653298 16678 653309
rect 17278 653298 18278 653309
rect 15748 653285 15772 653298
rect 15816 653285 15840 653298
rect 15884 653285 15908 653298
rect 15952 653285 15976 653298
rect 16020 653285 16044 653298
rect 16088 653285 16112 653298
rect 16156 653285 16180 653298
rect 16224 653285 16248 653298
rect 16292 653285 16316 653298
rect 16360 653285 16384 653298
rect 16428 653285 16452 653298
rect 16496 653285 16520 653298
rect 16564 653285 16588 653298
rect 16632 653285 16656 653298
rect 17290 653285 17314 653298
rect 17358 653285 17382 653298
rect 17426 653285 17450 653298
rect 17494 653285 17518 653298
rect 17562 653285 17586 653298
rect 17630 653285 17654 653298
rect 17698 653285 17722 653298
rect 17766 653285 17790 653298
rect 17834 653285 17858 653298
rect 17902 653285 17926 653298
rect 17970 653285 17994 653298
rect 18038 653285 18062 653298
rect 18106 653285 18130 653298
rect 18174 653285 18198 653298
rect 21413 653279 22813 653407
rect 23685 653279 25085 653407
rect 27158 653279 27358 653335
rect 21413 653116 22813 653244
rect 23685 653116 25085 653244
rect 27158 653103 27358 653231
rect 26393 653100 26477 653103
rect 26726 653100 26810 653103
rect 12543 653069 12881 653085
rect 12559 652967 12865 653069
rect 7389 652895 8389 652951
rect 8990 652895 9990 652951
rect 15678 652940 16678 652996
rect 17278 652940 18278 652996
rect 21413 652953 22813 653081
rect 23685 652953 25085 653081
rect 25936 653050 26936 653100
rect 27622 653095 27672 654095
rect 27772 653095 27828 654095
rect 27928 653095 27984 654095
rect 28084 653095 28140 654095
rect 28240 653095 28296 654095
rect 28396 653637 28446 654095
rect 28396 653553 28449 653637
rect 28396 653305 28446 653553
rect 29778 653320 29802 653344
rect 28396 653221 28449 653305
rect 29802 653296 29826 653309
rect 29880 653299 29914 653333
rect 29778 653261 29802 653285
rect 29890 653275 29914 653299
rect 28396 653095 28446 653221
rect 7389 652823 8389 652879
rect 8990 652823 9990 652879
rect 15678 652868 16678 652924
rect 17278 652868 18278 652924
rect 21413 652790 22813 652918
rect 23685 652790 25085 652918
rect 25936 652894 26936 652950
rect 27158 652927 27358 652983
rect 13899 652656 14059 652660
rect 7389 652521 8389 652593
rect 8990 652521 9990 652593
rect 15678 652566 16678 652638
rect 17278 652566 18278 652638
rect 21413 652627 22813 652755
rect 23685 652627 25085 652755
rect 25936 652738 26936 652794
rect 27158 652751 27358 652879
rect 27912 652757 27962 652873
rect 27909 652673 27962 652757
rect 28082 652673 28210 652873
rect 28258 652673 28314 652873
rect 28434 652673 28562 652873
rect 28610 652673 28660 652873
rect 27917 652669 27951 652673
rect 29880 652672 29914 652706
rect 25936 652582 26936 652638
rect 27158 652581 27358 652631
rect 27274 652578 27358 652581
rect 15748 652555 15782 652566
rect 15816 652555 15850 652566
rect 15884 652555 15918 652566
rect 15952 652555 15986 652566
rect 16020 652555 16054 652566
rect 16088 652555 16122 652566
rect 16156 652555 16190 652566
rect 16224 652555 16258 652566
rect 16292 652555 16326 652566
rect 16360 652555 16394 652566
rect 16428 652555 16462 652566
rect 16496 652555 16530 652566
rect 16564 652555 16598 652566
rect 16632 652555 16666 652566
rect 17290 652555 17324 652566
rect 17358 652555 17392 652566
rect 17426 652555 17460 652566
rect 17494 652555 17528 652566
rect 17562 652555 17596 652566
rect 17630 652555 17664 652566
rect 17698 652555 17732 652566
rect 17766 652555 17800 652566
rect 17834 652555 17868 652566
rect 17902 652555 17936 652566
rect 17970 652555 18004 652566
rect 18038 652555 18072 652566
rect 18106 652555 18140 652566
rect 18174 652555 18208 652566
rect 15748 652545 15806 652555
rect 15816 652545 15874 652555
rect 15884 652545 15942 652555
rect 15952 652545 16010 652555
rect 16020 652545 16078 652555
rect 16088 652545 16146 652555
rect 16156 652545 16214 652555
rect 16224 652545 16282 652555
rect 16292 652545 16350 652555
rect 16360 652545 16418 652555
rect 16428 652545 16486 652555
rect 16496 652545 16554 652555
rect 16564 652545 16622 652555
rect 16632 652545 16690 652555
rect 17290 652545 17348 652555
rect 17358 652545 17416 652555
rect 17426 652545 17484 652555
rect 17494 652545 17552 652555
rect 17562 652545 17620 652555
rect 17630 652545 17688 652555
rect 17698 652545 17756 652555
rect 17766 652545 17824 652555
rect 17834 652545 17892 652555
rect 17902 652545 17960 652555
rect 17970 652545 18028 652555
rect 18038 652545 18096 652555
rect 18106 652545 18164 652555
rect 18174 652545 18232 652555
rect 15724 652521 16690 652545
rect 17266 652521 18232 652545
rect 13901 652510 14061 652514
rect 15748 652506 15772 652521
rect 15816 652506 15840 652521
rect 15884 652506 15908 652521
rect 15952 652506 15976 652521
rect 16020 652506 16044 652521
rect 16088 652506 16112 652521
rect 16156 652506 16180 652521
rect 16224 652506 16248 652521
rect 16292 652506 16316 652521
rect 16360 652506 16384 652521
rect 16428 652506 16452 652521
rect 16496 652506 16520 652521
rect 16564 652506 16588 652521
rect 16632 652506 16656 652521
rect 17290 652506 17314 652521
rect 17358 652506 17382 652521
rect 17426 652506 17450 652521
rect 17494 652506 17518 652521
rect 17562 652506 17586 652521
rect 17630 652506 17654 652521
rect 17698 652506 17722 652521
rect 17766 652506 17790 652521
rect 17834 652506 17858 652521
rect 17902 652506 17926 652521
rect 17970 652506 17994 652521
rect 18038 652506 18062 652521
rect 18106 652506 18130 652521
rect 18174 652506 18198 652521
rect 15678 652351 16678 652506
rect 7389 652261 8389 652321
rect 8990 652261 9990 652321
rect 15678 652317 16690 652351
rect 17278 652341 18278 652506
rect 21413 652470 22813 652520
rect 23685 652470 25085 652520
rect 25936 652432 26936 652482
rect 21349 652390 21373 652414
rect 21407 652390 21431 652414
rect 25067 652390 25091 652414
rect 25125 652390 25149 652414
rect 21383 652356 21397 652390
rect 25101 652356 25115 652390
rect 17266 652317 18278 652341
rect 21349 652332 21373 652356
rect 21407 652332 21431 652356
rect 25067 652332 25091 652356
rect 25125 652332 25149 652356
rect 27917 652325 27951 652329
rect 15678 652306 16678 652317
rect 17278 652306 18278 652317
rect 15748 652293 15772 652306
rect 15816 652293 15840 652306
rect 15884 652293 15908 652306
rect 15952 652293 15976 652306
rect 16020 652293 16044 652306
rect 16088 652293 16112 652306
rect 16156 652293 16180 652306
rect 16224 652293 16248 652306
rect 16292 652293 16316 652306
rect 16360 652293 16384 652306
rect 16428 652293 16452 652306
rect 16496 652293 16520 652306
rect 16564 652293 16588 652306
rect 16632 652293 16656 652306
rect 17290 652293 17314 652306
rect 17358 652293 17382 652306
rect 17426 652293 17450 652306
rect 17494 652293 17518 652306
rect 17562 652293 17586 652306
rect 17630 652293 17654 652306
rect 17698 652293 17722 652306
rect 17766 652293 17790 652306
rect 17834 652293 17858 652306
rect 17902 652293 17926 652306
rect 17970 652293 17994 652306
rect 18038 652293 18062 652306
rect 18106 652293 18130 652306
rect 18174 652293 18198 652306
rect 27909 652241 27962 652325
rect 21634 652101 24864 652203
rect 27912 652125 27962 652241
rect 28082 652125 28210 652325
rect 28258 652125 28314 652325
rect 28434 652125 28562 652325
rect 28610 652125 28660 652325
rect 21186 652047 21210 652071
rect 25288 652047 25312 652071
rect 21162 652023 21186 652037
rect 25312 652023 25336 652037
rect 7389 651903 8389 651959
rect 8990 651903 9990 651959
rect 15678 651948 16678 652004
rect 17278 651948 18278 652004
rect 21072 651989 21084 652013
rect 21186 651989 21210 652013
rect 25288 651989 25312 652013
rect 25414 651989 25426 652013
rect 21385 651944 21403 651948
rect 7389 651831 8389 651887
rect 8990 651831 9990 651887
rect 15678 651876 16678 651932
rect 17278 651876 18278 651932
rect 20250 651914 20316 651930
rect 21377 651914 21403 651944
rect 21385 651904 21403 651914
rect 21383 651880 21403 651904
rect 21407 651880 21415 651914
rect 25113 651904 25121 651944
rect 25101 651880 25121 651904
rect 25125 651880 25143 651948
rect 21383 651846 21419 651880
rect 25101 651846 25147 651880
rect 21383 651812 21403 651846
rect 21407 651812 21415 651846
rect 21383 651778 21419 651812
rect 21481 651784 22881 651834
rect 23617 651784 25017 651834
rect 25101 651812 25121 651846
rect 25125 651812 25143 651846
rect 25101 651778 25147 651812
rect 21383 651744 21403 651778
rect 21407 651744 21415 651778
rect 21383 651710 21419 651744
rect 21383 651676 21403 651710
rect 21407 651676 21415 651710
rect 7389 651529 8389 651601
rect 8990 651529 9990 651601
rect 15678 651574 16678 651646
rect 17278 651574 18278 651646
rect 21383 651642 21419 651676
rect 21383 651608 21403 651642
rect 21407 651608 21415 651642
rect 21481 651621 22881 651749
rect 23617 651621 25017 651749
rect 25101 651744 25121 651778
rect 25125 651744 25143 651778
rect 25101 651710 25147 651744
rect 25101 651676 25121 651710
rect 25125 651676 25143 651710
rect 25101 651642 25147 651676
rect 25101 651608 25121 651642
rect 25125 651608 25143 651642
rect 21383 651574 21419 651608
rect 15748 651563 15782 651574
rect 15816 651563 15850 651574
rect 15884 651563 15918 651574
rect 15952 651563 15986 651574
rect 16020 651563 16054 651574
rect 16088 651563 16122 651574
rect 16156 651563 16190 651574
rect 16224 651563 16258 651574
rect 16292 651563 16326 651574
rect 16360 651563 16394 651574
rect 16428 651563 16462 651574
rect 16496 651563 16530 651574
rect 16564 651563 16598 651574
rect 16632 651563 16666 651574
rect 17290 651563 17324 651574
rect 17358 651563 17392 651574
rect 17426 651563 17460 651574
rect 17494 651563 17528 651574
rect 17562 651563 17596 651574
rect 17630 651563 17664 651574
rect 17698 651563 17732 651574
rect 17766 651563 17800 651574
rect 17834 651563 17868 651574
rect 17902 651563 17936 651574
rect 17970 651563 18004 651574
rect 18038 651563 18072 651574
rect 18106 651563 18140 651574
rect 18174 651563 18208 651574
rect 15748 651553 15806 651563
rect 15816 651553 15874 651563
rect 15884 651553 15942 651563
rect 15952 651553 16010 651563
rect 16020 651553 16078 651563
rect 16088 651553 16146 651563
rect 16156 651553 16214 651563
rect 16224 651553 16282 651563
rect 16292 651553 16350 651563
rect 16360 651553 16418 651563
rect 16428 651553 16486 651563
rect 16496 651553 16554 651563
rect 16564 651553 16622 651563
rect 16632 651553 16690 651563
rect 17290 651553 17348 651563
rect 17358 651553 17416 651563
rect 17426 651553 17484 651563
rect 17494 651553 17552 651563
rect 17562 651553 17620 651563
rect 17630 651553 17688 651563
rect 17698 651553 17756 651563
rect 17766 651553 17824 651563
rect 17834 651553 17892 651563
rect 17902 651553 17960 651563
rect 17970 651553 18028 651563
rect 18038 651553 18096 651563
rect 18106 651553 18164 651563
rect 18174 651553 18232 651563
rect 15724 651529 16690 651553
rect 17266 651529 18232 651553
rect 21383 651540 21403 651574
rect 21407 651540 21415 651574
rect 15748 651514 15772 651529
rect 15816 651514 15840 651529
rect 15884 651514 15908 651529
rect 15952 651514 15976 651529
rect 16020 651514 16044 651529
rect 16088 651514 16112 651529
rect 16156 651514 16180 651529
rect 16224 651514 16248 651529
rect 16292 651514 16316 651529
rect 16360 651514 16384 651529
rect 16428 651514 16452 651529
rect 16496 651514 16520 651529
rect 16564 651514 16588 651529
rect 16632 651514 16656 651529
rect 17290 651514 17314 651529
rect 17358 651514 17382 651529
rect 17426 651514 17450 651529
rect 17494 651514 17518 651529
rect 17562 651514 17586 651529
rect 17630 651514 17654 651529
rect 17698 651514 17722 651529
rect 17766 651514 17790 651529
rect 17834 651514 17858 651529
rect 17902 651514 17926 651529
rect 17970 651514 17994 651529
rect 18038 651514 18062 651529
rect 18106 651514 18130 651529
rect 18174 651514 18198 651529
rect 5937 651318 6089 651386
rect 15678 651359 16678 651514
rect 6005 651315 6089 651318
rect 5967 651305 6059 651315
rect 6005 651275 6021 651305
rect 1288 649503 1338 650503
rect 1438 649503 1566 650503
rect 1594 649503 1644 650503
rect 5995 649493 6021 651275
rect 7389 651269 8389 651329
rect 8990 651269 9990 651329
rect 15678 651325 16690 651359
rect 17278 651349 18278 651514
rect 17266 651325 18278 651349
rect 15678 651314 16678 651325
rect 17278 651314 18278 651325
rect 21383 651506 21419 651540
rect 21383 651472 21403 651506
rect 21407 651472 21415 651506
rect 21383 651438 21419 651472
rect 21481 651458 22881 651586
rect 23617 651458 25017 651586
rect 25101 651574 25147 651608
rect 25101 651540 25121 651574
rect 25125 651540 25143 651574
rect 25101 651506 25147 651540
rect 25101 651472 25121 651506
rect 25125 651472 25143 651506
rect 25101 651438 25147 651472
rect 21383 651404 21403 651438
rect 21407 651404 21415 651438
rect 21383 651370 21419 651404
rect 21383 651336 21403 651370
rect 21407 651336 21415 651370
rect 15748 651301 15772 651314
rect 15816 651301 15840 651314
rect 15884 651301 15908 651314
rect 15952 651301 15976 651314
rect 16020 651301 16044 651314
rect 16088 651301 16112 651314
rect 16156 651301 16180 651314
rect 16224 651301 16248 651314
rect 16292 651301 16316 651314
rect 16360 651301 16384 651314
rect 16428 651301 16452 651314
rect 16496 651301 16520 651314
rect 16564 651301 16588 651314
rect 16632 651301 16656 651314
rect 17290 651301 17314 651314
rect 17358 651301 17382 651314
rect 17426 651301 17450 651314
rect 17494 651301 17518 651314
rect 17562 651301 17586 651314
rect 17630 651301 17654 651314
rect 17698 651301 17722 651314
rect 17766 651301 17790 651314
rect 17834 651301 17858 651314
rect 17902 651301 17926 651314
rect 17970 651301 17994 651314
rect 18038 651301 18062 651314
rect 18106 651301 18130 651314
rect 18174 651301 18198 651314
rect 21383 651302 21419 651336
rect 21383 651268 21403 651302
rect 21407 651268 21415 651302
rect 21481 651295 22881 651423
rect 23617 651295 25017 651423
rect 25101 651404 25121 651438
rect 25125 651404 25143 651438
rect 25101 651370 25147 651404
rect 25101 651336 25121 651370
rect 25125 651336 25143 651370
rect 25101 651302 25147 651336
rect 25101 651268 25121 651302
rect 25125 651268 25143 651302
rect 21383 651234 21419 651268
rect 21383 651200 21403 651234
rect 21407 651200 21415 651234
rect 21383 651166 21419 651200
rect 21383 651132 21403 651166
rect 21407 651132 21415 651166
rect 21481 651132 22881 651260
rect 23617 651132 25017 651260
rect 25101 651234 25147 651268
rect 25101 651200 25121 651234
rect 25125 651200 25143 651234
rect 25101 651166 25147 651200
rect 25101 651132 25121 651166
rect 25125 651132 25143 651166
rect 21383 651098 21419 651132
rect 25101 651098 25147 651132
rect 21383 651064 21403 651098
rect 21407 651064 21415 651098
rect 21383 651030 21419 651064
rect 7389 650911 8389 650967
rect 8990 650911 9990 650967
rect 15678 650956 16678 651012
rect 17278 650956 18278 651012
rect 21383 650996 21403 651030
rect 21407 650996 21415 651030
rect 21383 650962 21419 650996
rect 21481 650969 22881 651097
rect 23617 650969 25017 651097
rect 25101 651064 25121 651098
rect 25125 651064 25143 651098
rect 25101 651030 25147 651064
rect 25101 650996 25121 651030
rect 25125 650996 25143 651030
rect 25101 650962 25147 650996
rect 26478 650985 26648 651291
rect 7389 650839 8389 650895
rect 8990 650839 9990 650895
rect 15678 650884 16678 650940
rect 17278 650884 18278 650940
rect 21383 650928 21403 650962
rect 21407 650928 21415 650962
rect 21383 650894 21419 650928
rect 21383 650860 21403 650894
rect 21407 650860 21415 650894
rect 21383 650826 21419 650860
rect 21383 650792 21403 650826
rect 21407 650792 21415 650826
rect 21481 650806 22881 650934
rect 23617 650806 25017 650934
rect 25101 650928 25121 650962
rect 25125 650928 25143 650962
rect 25101 650894 25147 650928
rect 27622 650903 27672 651903
rect 27772 650903 27828 651903
rect 27928 650903 27984 651903
rect 28084 650903 28140 651903
rect 28240 650903 28296 651903
rect 28396 651777 28446 651903
rect 28396 651693 28449 651777
rect 28396 651445 28446 651693
rect 30015 651523 30027 657246
rect 32596 657239 33596 657367
rect 35255 657345 36255 657401
rect 680215 657326 680815 657382
rect 685551 657360 686551 657488
rect 689154 657439 689204 657897
rect 689151 657355 689204 657439
rect 30135 657062 30735 657112
rect 31049 657042 32049 657092
rect 32596 657083 33596 657211
rect 35255 657169 36255 657297
rect 680215 657156 680815 657206
rect 685551 657204 686551 657332
rect 35255 656993 36255 657121
rect 685551 657048 686551 657176
rect 686865 657116 687465 657166
rect 30135 656886 30735 656942
rect 31049 656886 32049 656942
rect 32596 656927 33596 656983
rect 37998 656979 38148 656991
rect 38317 656979 38467 656991
rect 679007 656980 679607 657030
rect 30135 656716 30735 656766
rect 31049 656736 32049 656786
rect 32596 656777 33596 656827
rect 35255 656823 36255 656873
rect 37998 656866 38598 656916
rect 680615 656885 680630 656900
rect 680803 656896 680815 656900
rect 680800 656885 680815 656896
rect 685551 656892 686551 656948
rect 686865 656940 687465 657068
rect 679007 656810 679607 656860
rect 35255 656754 36255 656766
rect 37998 656690 38598 656746
rect 680615 656705 680815 656885
rect 683328 656793 683928 656843
rect 682573 656717 683173 656767
rect 680615 656690 680630 656705
rect 680800 656694 680815 656705
rect 680803 656690 680815 656694
rect 30135 656600 30735 656650
rect 31049 656600 32049 656650
rect 32596 656575 33196 656625
rect 35255 656621 36255 656671
rect 680502 656649 680517 656664
rect 30135 656424 30735 656480
rect 31049 656444 32049 656500
rect 30135 656248 30735 656376
rect 31049 656288 32049 656344
rect 30135 656072 30735 656200
rect 31049 656132 32049 656188
rect 32596 656141 33196 656191
rect 30135 655896 30735 656024
rect 31049 655982 32049 656032
rect 31049 655866 32049 655916
rect 30135 655726 30735 655776
rect 31049 655710 32049 655838
rect 30135 655610 30735 655660
rect 30135 655434 30735 655562
rect 31049 655554 32049 655682
rect 31049 655398 32049 655526
rect 34152 655490 34202 656478
rect 34322 655490 34372 656478
rect 34492 656465 35092 656515
rect 35255 656445 36255 656573
rect 37998 656520 38598 656570
rect 36785 656496 36797 656500
rect 36785 656485 36800 656496
rect 36970 656485 36985 656500
rect 34492 656289 35092 656345
rect 35255 656269 36255 656325
rect 36785 656305 36985 656485
rect 36785 656294 36800 656305
rect 36785 656290 36797 656294
rect 36970 656290 36985 656305
rect 37083 656485 37098 656500
rect 37083 656305 37120 656485
rect 680480 656469 680517 656649
rect 680502 656454 680517 656469
rect 680615 656649 680630 656664
rect 680803 656660 680815 656664
rect 680800 656649 680815 656660
rect 680615 656469 680815 656649
rect 682573 656541 683173 656669
rect 683328 656617 683928 656745
rect 685551 656736 686551 656864
rect 686865 656764 687465 656820
rect 685551 656580 686551 656708
rect 686865 656588 687465 656716
rect 680615 656454 680630 656469
rect 680800 656458 680815 656469
rect 680803 656454 680815 656458
rect 683328 656441 683928 656497
rect 679002 656384 679602 656434
rect 685551 656424 686551 656552
rect 682573 656365 683173 656421
rect 686865 656412 687465 656468
rect 37083 656290 37098 656305
rect 36785 656260 36797 656264
rect 36785 656249 36800 656260
rect 36970 656249 36985 656264
rect 34492 656119 35092 656169
rect 35255 656099 36255 656149
rect 36785 656069 36985 656249
rect 679002 656208 679602 656264
rect 682573 656189 683173 656317
rect 683328 656265 683928 656321
rect 685551 656274 686551 656324
rect 686865 656236 687465 656364
rect 685551 656158 686551 656208
rect 37993 656094 38593 656144
rect 678680 656123 678704 656157
rect 36785 656058 36800 656069
rect 36785 656054 36797 656058
rect 36970 656054 36985 656069
rect 678680 656055 678704 656089
rect 679002 656038 679602 656088
rect 679061 656035 679355 656038
rect 679380 656035 679602 656038
rect 678680 655987 678704 656021
rect 682573 656013 683173 656141
rect 683328 656089 683928 656145
rect 34491 655849 35091 655899
rect 35255 655883 35855 655933
rect 37993 655924 38593 655974
rect 678680 655919 678704 655953
rect 678680 655851 678704 655885
rect 682573 655837 683173 655965
rect 683328 655913 683928 656041
rect 685551 655982 686551 656110
rect 686865 656060 687465 656116
rect 34491 655673 35091 655729
rect 35255 655707 35855 655763
rect 36785 655748 37385 655798
rect 38920 655761 38946 655787
rect 678680 655783 678704 655817
rect 685551 655806 686551 655934
rect 686865 655884 687465 656012
rect 678680 655715 678704 655749
rect 34491 655503 35091 655553
rect 35255 655531 35855 655659
rect 678680 655647 678704 655681
rect 682573 655661 683173 655789
rect 683328 655737 683928 655793
rect 685551 655630 686551 655758
rect 686865 655708 687465 655836
rect 36785 655572 37385 655628
rect 678680 655579 678704 655613
rect 683328 655567 683928 655617
rect 678680 655511 678704 655545
rect 682573 655491 683173 655541
rect 684519 655498 685119 655548
rect 34019 655418 34029 655490
rect 34152 655478 34372 655490
rect 34091 655415 34101 655418
rect 30135 655258 30735 655314
rect 31049 655242 32049 655370
rect 34091 655365 35091 655415
rect 35255 655361 35855 655411
rect 36785 655396 37385 655452
rect 678680 655443 678704 655477
rect 685551 655454 686551 655582
rect 686865 655532 687465 655660
rect 679133 655409 679283 655421
rect 679452 655409 679602 655421
rect 678680 655375 678704 655409
rect 678680 655307 678704 655341
rect 679002 655296 679602 655346
rect 684519 655342 685119 655398
rect 685551 655278 686551 655406
rect 686865 655356 687465 655484
rect 30135 655082 30735 655210
rect 31049 655086 32049 655214
rect 34091 655195 35091 655245
rect 36785 655226 37385 655276
rect 678680 655239 678704 655273
rect 34091 655192 34101 655195
rect 34202 655192 34302 655195
rect 35255 655159 35855 655209
rect 678680 655171 678704 655205
rect 684519 655192 685119 655242
rect 30135 654912 30735 654962
rect 31049 654930 32049 654986
rect 30135 654796 30735 654846
rect 31049 654774 32049 654902
rect 32481 654898 33081 654948
rect 30135 654620 30735 654748
rect 31049 654618 32049 654746
rect 32481 654742 33081 654870
rect 30135 654444 30735 654572
rect 31049 654462 32049 654590
rect 32481 654586 33081 654714
rect 34152 654532 34202 655132
rect 34302 654532 34352 655132
rect 34491 655066 35091 655116
rect 35255 655003 35855 655131
rect 36785 655094 37385 655144
rect 678680 655103 678704 655137
rect 679002 655120 679602 655176
rect 681745 655081 682345 655131
rect 682509 655069 683109 655119
rect 678680 655035 678704 655069
rect 683739 655027 684339 655077
rect 684519 655062 685119 655112
rect 685551 655102 686551 655230
rect 686865 655180 687465 655308
rect 34491 654890 35091 654946
rect 36785 654918 37385 654974
rect 678680 654967 678704 655001
rect 679002 654950 679602 655000
rect 35255 654847 35855 654903
rect 678680 654899 678704 654933
rect 680502 654915 680517 654930
rect 678680 654831 678704 654865
rect 34491 654720 35091 654770
rect 35255 654691 35855 654819
rect 36785 654742 37385 654798
rect 678680 654763 678704 654797
rect 680480 654735 680517 654915
rect 678680 654695 678704 654729
rect 680502 654720 680517 654735
rect 680615 654915 680630 654930
rect 680803 654926 680815 654930
rect 680800 654915 680815 654926
rect 681745 654925 682345 654981
rect 680615 654735 680815 654915
rect 681745 654769 682345 654897
rect 682509 654893 683109 655021
rect 684519 654906 685119 655034
rect 685551 654926 686551 655054
rect 686865 655004 687465 655060
rect 683739 654837 684339 654893
rect 686865 654828 687465 654956
rect 680615 654720 680630 654735
rect 680800 654724 680815 654735
rect 680803 654720 680815 654724
rect 680615 654679 680630 654694
rect 680803 654690 680815 654694
rect 680800 654679 680815 654690
rect 678680 654627 678704 654661
rect 35255 654541 35855 654591
rect 36785 654572 37385 654622
rect 678680 654559 678704 654593
rect 678680 654491 678704 654525
rect 679007 654524 679607 654574
rect 680615 654499 680815 654679
rect 681745 654613 682345 654741
rect 682509 654717 683109 654773
rect 684519 654750 685119 654806
rect 685551 654750 686551 654806
rect 682509 654541 683109 654669
rect 684519 654594 685119 654722
rect 685551 654594 686551 654722
rect 686865 654652 687465 654780
rect 32481 654436 33081 654486
rect 680615 654484 680630 654499
rect 680800 654488 680815 654499
rect 680803 654484 680815 654488
rect 681745 654463 682345 654513
rect 683739 654477 684339 654513
rect 30135 654268 30735 654396
rect 31049 654306 32049 654434
rect 34491 654379 35091 654429
rect 37993 654396 38593 654446
rect 678680 654423 678704 654457
rect 684519 654444 685119 654494
rect 685551 654438 686551 654566
rect 686865 654476 687465 654604
rect 32481 654306 33081 654356
rect 678680 654355 678704 654389
rect 679007 654354 679607 654404
rect 682509 654371 683109 654421
rect 33261 654287 33861 654323
rect 30135 654092 30735 654220
rect 31049 654150 32049 654278
rect 32481 654150 33081 654278
rect 34491 654203 35091 654331
rect 35255 654287 35855 654337
rect 36785 654312 36797 654316
rect 36785 654301 36800 654312
rect 36970 654301 36985 654316
rect 35255 654131 35855 654259
rect 36785 654121 36985 654301
rect 678680 654287 678704 654321
rect 684519 654314 685119 654364
rect 37993 654226 38593 654276
rect 678680 654219 678704 654253
rect 678680 654151 678704 654185
rect 680215 654178 680815 654228
rect 681745 654209 682345 654259
rect 36785 654110 36800 654121
rect 36785 654106 36797 654110
rect 36970 654106 36985 654121
rect 30135 653916 30735 654044
rect 31049 653994 32049 654050
rect 32481 653994 33081 654050
rect 34491 654027 35091 654083
rect 31049 653818 32049 653946
rect 32481 653838 33081 653966
rect 33261 653907 33861 653963
rect 34491 653851 35091 653979
rect 35255 653975 35855 654103
rect 678680 654083 678704 654117
rect 36785 654076 36797 654080
rect 36785 654065 36800 654076
rect 36970 654065 36985 654080
rect 36785 653885 36985 654065
rect 35255 653819 35855 653875
rect 36785 653874 36800 653885
rect 36785 653870 36797 653874
rect 36970 653870 36985 653885
rect 37083 654065 37098 654080
rect 37083 653885 37120 654065
rect 678680 654015 678704 654049
rect 680215 654002 680815 654058
rect 681745 654053 682345 654181
rect 682509 654030 683109 654080
rect 678680 653947 678704 653981
rect 37083 653870 37098 653885
rect 678680 653879 678704 653913
rect 681745 653897 682345 653953
rect 37998 653800 38598 653850
rect 678680 653811 678704 653845
rect 680215 653826 680815 653882
rect 30135 653740 30735 653796
rect 30135 653564 30735 653692
rect 31049 653642 32049 653770
rect 32481 653688 33081 653738
rect 33261 653723 33861 653773
rect 678680 653743 678704 653777
rect 681745 653741 682345 653869
rect 682509 653854 683109 653910
rect 34491 653681 35091 653731
rect 35255 653669 35855 653719
rect 37998 653624 38598 653680
rect 678680 653675 678704 653709
rect 680215 653656 680815 653706
rect 682509 653684 683109 653734
rect 683248 653680 683298 654268
rect 683398 653680 683448 654268
rect 684519 654158 685119 654286
rect 685551 654282 686551 654410
rect 686865 654300 687465 654428
rect 684519 654002 685119 654130
rect 685551 654126 686551 654254
rect 686865 654124 687465 654252
rect 685551 653970 686551 654098
rect 686865 653954 687465 654004
rect 684519 653852 685119 653902
rect 685551 653814 686551 653870
rect 686865 653838 687465 653888
rect 683248 653668 683448 653680
rect 685551 653658 686551 653786
rect 686865 653662 687465 653790
rect 30135 653388 30735 653516
rect 31049 653466 32049 653594
rect 32481 653558 33081 653608
rect 678680 653607 678704 653641
rect 681745 653591 682345 653641
rect 683571 653605 683581 653646
rect 678680 653539 678704 653573
rect 680215 653524 680815 653574
rect 682509 653555 683509 653605
rect 30135 653212 30735 653340
rect 31049 653290 32049 653418
rect 32481 653402 33081 653458
rect 37998 653454 38598 653504
rect 678680 653471 678704 653505
rect 685551 653502 686551 653630
rect 686865 653486 687465 653542
rect 37998 653451 38220 653454
rect 38245 653451 38539 653454
rect 678680 653403 678704 653437
rect 678680 653335 678704 653369
rect 680215 653348 680815 653404
rect 681745 653389 682345 653439
rect 682509 653385 683509 653435
rect 683278 653382 683398 653385
rect 683571 653382 683581 653385
rect 685551 653346 686551 653474
rect 32481 653252 33081 653302
rect 34427 653259 35027 653309
rect 678680 653267 678704 653301
rect 30135 653036 30735 653164
rect 31049 653114 32049 653242
rect 33672 653183 34272 653233
rect 34427 653083 35027 653211
rect 678680 653199 678704 653233
rect 680215 653172 680815 653228
rect 681745 653213 682345 653341
rect 682509 653247 683109 653297
rect 678680 653131 678704 653165
rect 30135 652860 30735 652988
rect 31049 652938 32049 653066
rect 678680 653063 678704 653097
rect 33672 653007 34272 653063
rect 31049 652762 32049 652890
rect 33672 652831 34272 652959
rect 34427 652907 35027 653035
rect 678654 653013 678680 653039
rect 680215 653002 680815 653052
rect 681745 653037 682345 653093
rect 682509 653071 683109 653127
rect 678680 652929 678704 652963
rect 678680 652861 678704 652895
rect 30135 652684 30735 652740
rect 34427 652731 35027 652859
rect 37998 652825 38148 652837
rect 38317 652825 38467 652837
rect 678680 652793 678704 652827
rect 679007 652826 679607 652876
rect 681745 652867 682345 652917
rect 682509 652901 683109 652951
rect 37998 652712 38598 652762
rect 678680 652725 678704 652759
rect 680615 652731 680630 652746
rect 680803 652742 680815 652746
rect 680800 652731 680815 652742
rect 33672 652655 34272 652711
rect 30135 652508 30735 652636
rect 31049 652592 32049 652642
rect 34427 652555 35027 652683
rect 678680 652657 678704 652691
rect 679007 652656 679607 652706
rect 37998 652536 38598 652592
rect 678680 652589 678704 652623
rect 31049 652476 32049 652526
rect 33672 652479 34272 652535
rect 678680 652521 678704 652555
rect 680615 652551 680815 652731
rect 681345 652651 682345 652701
rect 682508 652631 683108 652681
rect 680615 652536 680630 652551
rect 680800 652540 680815 652551
rect 680803 652536 680815 652540
rect 680502 652495 680517 652510
rect 678680 652453 678704 652487
rect 30135 652332 30735 652388
rect 31049 652320 32049 652448
rect 34427 652379 35027 652435
rect 37998 652366 38598 652416
rect 678680 652385 678704 652419
rect 33672 652303 34272 652359
rect 36785 652342 36797 652346
rect 36785 652331 36800 652342
rect 36970 652331 36985 652346
rect 30135 652156 30735 652284
rect 31049 652164 32049 652292
rect 30135 651980 30735 652036
rect 31049 652008 32049 652136
rect 33672 652127 34272 652255
rect 34427 652203 35027 652331
rect 36785 652151 36985 652331
rect 36785 652140 36800 652151
rect 36785 652136 36797 652140
rect 36970 652136 36985 652151
rect 37083 652331 37098 652346
rect 37083 652151 37120 652331
rect 678680 652317 678704 652351
rect 680480 652315 680517 652495
rect 680502 652300 680517 652315
rect 680615 652495 680630 652510
rect 680803 652506 680815 652510
rect 680800 652495 680815 652506
rect 680615 652315 680815 652495
rect 681345 652475 682345 652531
rect 682508 652455 683108 652511
rect 680615 652300 680630 652315
rect 680800 652304 680815 652315
rect 680803 652300 680815 652304
rect 681345 652299 682345 652427
rect 682508 652285 683108 652335
rect 683228 652322 683278 653322
rect 683398 652322 683448 653322
rect 685551 653190 686551 653318
rect 686865 653310 687465 653438
rect 685551 653034 686551 653162
rect 686865 653140 687465 653190
rect 686865 653024 687465 653074
rect 685551 652884 686551 652934
rect 686865 652848 687465 652976
rect 685551 652768 686551 652818
rect 686865 652672 687465 652800
rect 684404 652609 685004 652659
rect 685551 652612 686551 652668
rect 685551 652456 686551 652512
rect 686865 652496 687465 652624
rect 685551 652300 686551 652356
rect 686865 652320 687465 652376
rect 678680 652249 678704 652283
rect 679002 652230 679602 652280
rect 678680 652181 678704 652215
rect 37083 652136 37098 652151
rect 678680 652113 678704 652147
rect 681345 652129 682345 652179
rect 684404 652175 685004 652225
rect 685551 652150 686551 652200
rect 686865 652150 687465 652200
rect 36785 652106 36797 652110
rect 36785 652095 36800 652106
rect 36970 652095 36985 652110
rect 34427 652033 35027 652083
rect 33672 651957 34272 652007
rect 30135 651804 30735 651932
rect 36785 651915 36985 652095
rect 678680 652045 678704 652079
rect 679002 652054 679602 652110
rect 681390 652070 681424 652080
rect 681458 652070 681492 652080
rect 681526 652070 681560 652080
rect 681594 652070 681628 652080
rect 681662 652070 681696 652080
rect 681730 652070 681764 652080
rect 681798 652070 681832 652080
rect 681866 652070 681900 652080
rect 681934 652070 681968 652080
rect 682002 652070 682036 652080
rect 682077 652070 682111 652080
rect 682145 652070 682179 652080
rect 682213 652070 682247 652080
rect 682281 652070 682315 652080
rect 681345 652034 682345 652046
rect 37993 651940 38593 651990
rect 678680 651977 678704 652011
rect 31049 651852 32049 651908
rect 36785 651904 36800 651915
rect 36785 651900 36797 651904
rect 36970 651900 36985 651915
rect 678680 651909 678704 651943
rect 679002 651884 679602 651934
rect 681345 651927 682345 651977
rect 684004 651973 685004 652023
rect 685551 652014 686551 652064
rect 686865 652034 687465 652084
rect 679061 651881 679355 651884
rect 679380 651881 679602 651884
rect 678680 651841 678704 651875
rect 31049 651696 32049 651824
rect 37993 651770 38593 651820
rect 678680 651773 678704 651807
rect 681345 651751 682345 651879
rect 684004 651817 685004 651873
rect 685551 651858 686551 651914
rect 686865 651858 687465 651914
rect 686686 651812 686714 651840
rect 678680 651705 678704 651739
rect 30135 651634 30735 651684
rect 31049 651540 32049 651668
rect 36785 651594 37385 651644
rect 678680 651637 678704 651671
rect 678680 651569 678704 651603
rect 681345 651575 682345 651703
rect 684004 651661 685004 651789
rect 685551 651708 686551 651758
rect 686865 651688 687465 651738
rect 28396 651361 28449 651445
rect 31049 651384 32049 651512
rect 678680 651501 678704 651535
rect 684004 651505 685004 651633
rect 687573 651554 687585 657277
rect 689154 657107 689204 657355
rect 689151 657023 689204 657107
rect 689154 656897 689204 657023
rect 689304 656897 689360 657897
rect 689460 656897 689516 657897
rect 689616 656897 689672 657897
rect 689772 656897 689828 657897
rect 689928 656897 689978 657897
rect 692485 657872 692521 657906
rect 692485 657838 692505 657872
rect 692509 657838 692517 657872
rect 690952 657509 691122 657815
rect 692485 657804 692521 657838
rect 692485 657770 692505 657804
rect 692509 657770 692517 657804
rect 692583 657775 693983 657903
rect 694719 657775 696119 657903
rect 696203 657872 696249 657906
rect 696203 657838 696223 657872
rect 696227 657838 696245 657872
rect 699322 657860 700322 657916
rect 700922 657860 701922 657916
rect 707610 657905 708610 657961
rect 709211 657905 710211 657961
rect 696203 657804 696249 657838
rect 696203 657770 696223 657804
rect 696227 657770 696245 657804
rect 699322 657788 700322 657844
rect 700922 657788 701922 657844
rect 707610 657833 708610 657889
rect 709211 657833 710211 657889
rect 692485 657736 692521 657770
rect 692485 657702 692505 657736
rect 692509 657702 692517 657736
rect 692485 657668 692521 657702
rect 692485 657634 692505 657668
rect 692509 657634 692517 657668
rect 692485 657600 692521 657634
rect 692583 657612 693983 657740
rect 694719 657612 696119 657740
rect 696203 657736 696249 657770
rect 696203 657702 696223 657736
rect 696227 657702 696245 657736
rect 696203 657668 696249 657702
rect 696203 657634 696223 657668
rect 696227 657634 696245 657668
rect 696203 657600 696249 657634
rect 692485 657566 692505 657600
rect 692509 657566 692517 657600
rect 692485 657532 692521 657566
rect 692485 657498 692505 657532
rect 692509 657498 692517 657532
rect 692485 657464 692521 657498
rect 692485 657430 692505 657464
rect 692509 657430 692517 657464
rect 692583 657449 693983 657577
rect 694719 657449 696119 657577
rect 696203 657566 696223 657600
rect 696227 657566 696245 657600
rect 696203 657532 696249 657566
rect 696203 657498 696223 657532
rect 696227 657498 696245 657532
rect 696203 657464 696249 657498
rect 699322 657486 700322 657558
rect 700922 657486 701922 657558
rect 707610 657531 708610 657603
rect 709211 657531 710211 657603
rect 711579 657553 711605 659307
rect 715956 658297 716006 659297
rect 716106 658297 716234 659297
rect 716262 658297 716312 659297
rect 699392 657475 699426 657486
rect 699460 657475 699494 657486
rect 699528 657475 699562 657486
rect 699596 657475 699630 657486
rect 699664 657475 699698 657486
rect 699732 657475 699766 657486
rect 699800 657475 699834 657486
rect 699868 657475 699902 657486
rect 699936 657475 699970 657486
rect 700004 657475 700038 657486
rect 700072 657475 700106 657486
rect 700140 657475 700174 657486
rect 700208 657475 700242 657486
rect 700276 657475 700310 657486
rect 700934 657475 700968 657486
rect 701002 657475 701036 657486
rect 701070 657475 701104 657486
rect 701138 657475 701172 657486
rect 701206 657475 701240 657486
rect 701274 657475 701308 657486
rect 701342 657475 701376 657486
rect 701410 657475 701444 657486
rect 701478 657475 701512 657486
rect 701546 657475 701580 657486
rect 701614 657475 701648 657486
rect 701682 657475 701716 657486
rect 701750 657475 701784 657486
rect 701818 657475 701852 657486
rect 711511 657485 711663 657553
rect 712447 657501 712557 657511
rect 711579 657482 711663 657485
rect 699392 657465 699450 657475
rect 699460 657465 699518 657475
rect 699528 657465 699586 657475
rect 699596 657465 699654 657475
rect 699664 657465 699722 657475
rect 699732 657465 699790 657475
rect 699800 657465 699858 657475
rect 699868 657465 699926 657475
rect 699936 657465 699994 657475
rect 700004 657465 700062 657475
rect 700072 657465 700130 657475
rect 700140 657465 700198 657475
rect 700208 657465 700266 657475
rect 700276 657465 700334 657475
rect 700934 657465 700992 657475
rect 701002 657465 701060 657475
rect 701070 657465 701128 657475
rect 701138 657465 701196 657475
rect 701206 657465 701264 657475
rect 701274 657465 701332 657475
rect 701342 657465 701400 657475
rect 701410 657465 701468 657475
rect 701478 657465 701536 657475
rect 701546 657465 701604 657475
rect 701614 657465 701672 657475
rect 701682 657465 701740 657475
rect 701750 657465 701808 657475
rect 701818 657465 701876 657475
rect 696203 657430 696223 657464
rect 696227 657430 696245 657464
rect 699368 657441 700334 657465
rect 700910 657441 701876 657465
rect 711541 657461 711633 657482
rect 692485 657396 692521 657430
rect 692485 657362 692505 657396
rect 692509 657362 692517 657396
rect 692485 657328 692521 657362
rect 692485 657294 692505 657328
rect 692509 657294 692517 657328
rect 692485 657260 692521 657294
rect 692583 657286 693983 657414
rect 694719 657286 696119 657414
rect 696203 657396 696249 657430
rect 699392 657426 699416 657441
rect 699460 657426 699484 657441
rect 699528 657426 699552 657441
rect 699596 657426 699620 657441
rect 699664 657426 699688 657441
rect 699732 657426 699756 657441
rect 699800 657426 699824 657441
rect 699868 657426 699892 657441
rect 699936 657426 699960 657441
rect 700004 657426 700028 657441
rect 700072 657426 700096 657441
rect 700140 657426 700164 657441
rect 700208 657426 700232 657441
rect 700276 657426 700300 657441
rect 700934 657426 700958 657441
rect 701002 657426 701026 657441
rect 701070 657426 701094 657441
rect 701138 657426 701162 657441
rect 701206 657426 701230 657441
rect 701274 657426 701298 657441
rect 701342 657426 701366 657441
rect 701410 657426 701434 657441
rect 701478 657426 701502 657441
rect 701546 657426 701570 657441
rect 701614 657426 701638 657441
rect 701682 657426 701706 657441
rect 701750 657426 701774 657441
rect 701818 657426 701842 657441
rect 696203 657362 696223 657396
rect 696227 657362 696245 657396
rect 696203 657328 696249 657362
rect 696203 657294 696223 657328
rect 696227 657294 696245 657328
rect 696203 657260 696249 657294
rect 699322 657271 700322 657426
rect 692485 657226 692505 657260
rect 692509 657226 692517 657260
rect 692485 657192 692521 657226
rect 692485 657158 692505 657192
rect 692509 657158 692517 657192
rect 692485 657124 692521 657158
rect 692485 657090 692505 657124
rect 692509 657090 692517 657124
rect 692583 657123 693983 657251
rect 694719 657123 696119 657251
rect 696203 657226 696223 657260
rect 696227 657226 696245 657260
rect 699322 657237 700334 657271
rect 700922 657261 701922 657426
rect 707610 657271 708610 657331
rect 709211 657271 710211 657331
rect 700910 657237 701922 657261
rect 699322 657226 700322 657237
rect 700922 657226 701922 657237
rect 696203 657192 696249 657226
rect 699392 657213 699416 657226
rect 699460 657213 699484 657226
rect 699528 657213 699552 657226
rect 699596 657213 699620 657226
rect 699664 657213 699688 657226
rect 699732 657213 699756 657226
rect 699800 657213 699824 657226
rect 699868 657213 699892 657226
rect 699936 657213 699960 657226
rect 700004 657213 700028 657226
rect 700072 657213 700096 657226
rect 700140 657213 700164 657226
rect 700208 657213 700232 657226
rect 700276 657213 700300 657226
rect 700934 657213 700958 657226
rect 701002 657213 701026 657226
rect 701070 657213 701094 657226
rect 701138 657213 701162 657226
rect 701206 657213 701230 657226
rect 701274 657213 701298 657226
rect 701342 657213 701366 657226
rect 701410 657213 701434 657226
rect 701478 657213 701502 657226
rect 701546 657213 701570 657226
rect 701614 657213 701638 657226
rect 701682 657213 701706 657226
rect 701750 657213 701774 657226
rect 701818 657213 701842 657226
rect 696203 657158 696223 657192
rect 696227 657158 696245 657192
rect 696203 657124 696249 657158
rect 696203 657090 696223 657124
rect 696227 657090 696245 657124
rect 692485 657056 692521 657090
rect 696203 657056 696249 657090
rect 692485 657022 692505 657056
rect 692509 657022 692517 657056
rect 696203 657022 696223 657056
rect 696227 657022 696245 657056
rect 692485 656988 692521 657022
rect 692485 656954 692505 656988
rect 692509 656954 692517 656988
rect 692583 656966 693983 657016
rect 694719 656966 696119 657016
rect 696203 656988 696249 657022
rect 696203 656954 696223 656988
rect 696227 656954 696245 656988
rect 692485 656920 692521 656954
rect 696203 656920 696249 656954
rect 692485 656896 692505 656920
rect 692487 656852 692505 656896
rect 692509 656886 692517 656920
rect 696203 656896 696223 656920
rect 696215 656886 696223 656896
rect 696227 656852 696245 656920
rect 697284 656870 697350 656886
rect 699322 656868 700322 656924
rect 700922 656868 701922 656924
rect 707610 656913 708610 656969
rect 709211 656913 710211 656969
rect 692174 656787 692186 656811
rect 692288 656787 692312 656811
rect 696390 656787 696414 656811
rect 696516 656787 696528 656811
rect 699322 656796 700322 656852
rect 700922 656796 701922 656852
rect 707610 656841 708610 656897
rect 709211 656841 710211 656897
rect 692264 656763 692288 656777
rect 696414 656763 696438 656777
rect 692288 656729 692312 656753
rect 696390 656729 696414 656753
rect 688940 656475 688990 656675
rect 689110 656475 689238 656675
rect 689286 656475 689342 656675
rect 689462 656475 689590 656675
rect 689638 656559 689688 656675
rect 692736 656597 695966 656699
rect 689638 656475 689691 656559
rect 699322 656494 700322 656566
rect 700922 656494 701922 656566
rect 707610 656539 708610 656611
rect 709211 656539 710211 656611
rect 699392 656483 699426 656494
rect 699460 656483 699494 656494
rect 699528 656483 699562 656494
rect 699596 656483 699630 656494
rect 699664 656483 699698 656494
rect 699732 656483 699766 656494
rect 699800 656483 699834 656494
rect 699868 656483 699902 656494
rect 699936 656483 699970 656494
rect 700004 656483 700038 656494
rect 700072 656483 700106 656494
rect 700140 656483 700174 656494
rect 700208 656483 700242 656494
rect 700276 656483 700310 656494
rect 700934 656483 700968 656494
rect 701002 656483 701036 656494
rect 701070 656483 701104 656494
rect 701138 656483 701172 656494
rect 701206 656483 701240 656494
rect 701274 656483 701308 656494
rect 701342 656483 701376 656494
rect 701410 656483 701444 656494
rect 701478 656483 701512 656494
rect 701546 656483 701580 656494
rect 701614 656483 701648 656494
rect 701682 656483 701716 656494
rect 701750 656483 701784 656494
rect 701818 656483 701852 656494
rect 689649 656471 689683 656475
rect 699392 656473 699450 656483
rect 699460 656473 699518 656483
rect 699528 656473 699586 656483
rect 699596 656473 699654 656483
rect 699664 656473 699722 656483
rect 699732 656473 699790 656483
rect 699800 656473 699858 656483
rect 699868 656473 699926 656483
rect 699936 656473 699994 656483
rect 700004 656473 700062 656483
rect 700072 656473 700130 656483
rect 700140 656473 700198 656483
rect 700208 656473 700266 656483
rect 700276 656473 700334 656483
rect 700934 656473 700992 656483
rect 701002 656473 701060 656483
rect 701070 656473 701128 656483
rect 701138 656473 701196 656483
rect 701206 656473 701264 656483
rect 701274 656473 701332 656483
rect 701342 656473 701400 656483
rect 701410 656473 701468 656483
rect 701478 656473 701536 656483
rect 701546 656473 701604 656483
rect 701614 656473 701672 656483
rect 701682 656473 701740 656483
rect 701750 656473 701808 656483
rect 701818 656473 701876 656483
rect 692451 656444 692475 656468
rect 692509 656444 692533 656468
rect 696169 656444 696193 656468
rect 696227 656444 696251 656468
rect 699368 656449 700334 656473
rect 700910 656449 701876 656473
rect 692485 656410 692499 656444
rect 696203 656410 696217 656444
rect 699392 656434 699416 656449
rect 699460 656434 699484 656449
rect 699528 656434 699552 656449
rect 699596 656434 699620 656449
rect 699664 656434 699688 656449
rect 699732 656434 699756 656449
rect 699800 656434 699824 656449
rect 699868 656434 699892 656449
rect 699936 656434 699960 656449
rect 700004 656434 700028 656449
rect 700072 656434 700096 656449
rect 700140 656434 700164 656449
rect 700208 656434 700232 656449
rect 700276 656434 700300 656449
rect 700934 656434 700958 656449
rect 701002 656434 701026 656449
rect 701070 656434 701094 656449
rect 701138 656434 701162 656449
rect 701206 656434 701230 656449
rect 701274 656434 701298 656449
rect 701342 656434 701366 656449
rect 701410 656434 701434 656449
rect 701478 656434 701502 656449
rect 701546 656434 701570 656449
rect 701614 656434 701638 656449
rect 701682 656434 701706 656449
rect 701750 656434 701774 656449
rect 701818 656434 701842 656449
rect 692451 656386 692475 656410
rect 692509 656386 692533 656410
rect 696169 656386 696193 656410
rect 696227 656386 696251 656410
rect 690664 656318 691664 656368
rect 692515 656280 693915 656330
rect 694787 656280 696187 656330
rect 699322 656279 700322 656434
rect 699322 656245 700334 656279
rect 700922 656269 701922 656434
rect 703539 656286 703699 656290
rect 707610 656279 708610 656339
rect 709211 656279 710211 656339
rect 700910 656245 701922 656269
rect 690242 656219 690326 656222
rect 690242 656214 690442 656219
rect 690238 656180 690442 656214
rect 690242 656169 690442 656180
rect 690664 656162 691664 656218
rect 687686 656128 687720 656162
rect 687686 656104 687710 656128
rect 689649 656127 689683 656131
rect 688940 655927 688990 656127
rect 689110 655927 689238 656127
rect 689286 655927 689342 656127
rect 689462 655927 689590 656127
rect 689638 656043 689691 656127
rect 689638 655927 689688 656043
rect 690242 655993 690442 656121
rect 692515 656117 693915 656245
rect 694787 656117 696187 656245
rect 699322 656234 700322 656245
rect 700922 656234 701922 656245
rect 699392 656221 699416 656234
rect 699460 656221 699484 656234
rect 699528 656221 699552 656234
rect 699596 656221 699620 656234
rect 699664 656221 699688 656234
rect 699732 656221 699756 656234
rect 699800 656221 699824 656234
rect 699868 656221 699892 656234
rect 699936 656221 699960 656234
rect 700004 656221 700028 656234
rect 700072 656221 700096 656234
rect 700140 656221 700164 656234
rect 700208 656221 700232 656234
rect 700276 656221 700300 656234
rect 700934 656221 700958 656234
rect 701002 656221 701026 656234
rect 701070 656221 701094 656234
rect 701138 656221 701162 656234
rect 701206 656221 701230 656234
rect 701274 656221 701298 656234
rect 701342 656221 701366 656234
rect 701410 656221 701434 656234
rect 701478 656221 701502 656234
rect 701546 656221 701570 656234
rect 701614 656221 701638 656234
rect 701682 656221 701706 656234
rect 701750 656221 701774 656234
rect 701818 656221 701842 656234
rect 703541 656140 703701 656144
rect 690664 656006 691664 656062
rect 692515 655954 693915 656082
rect 694787 655954 696187 656082
rect 690242 655817 690442 655873
rect 690664 655850 691664 655906
rect 692515 655791 693915 655919
rect 694787 655791 696187 655919
rect 699322 655876 700322 655932
rect 700922 655876 701922 655932
rect 707610 655921 708610 655977
rect 709211 655921 710211 655977
rect 699322 655804 700322 655860
rect 700922 655804 701922 655860
rect 707610 655849 708610 655905
rect 709211 655849 710211 655905
rect 689154 655579 689204 655705
rect 687686 655501 687720 655535
rect 687798 655515 687822 655539
rect 687774 655491 687798 655504
rect 689151 655495 689204 655579
rect 687798 655456 687822 655480
rect 689154 655247 689204 655495
rect 689151 655163 689204 655247
rect 689154 654705 689204 655163
rect 689304 654705 689360 655705
rect 689460 654705 689516 655705
rect 689616 654705 689672 655705
rect 689772 654705 689828 655705
rect 689928 654705 689978 655705
rect 690242 655641 690442 655769
rect 690664 655700 691664 655750
rect 690790 655697 690874 655700
rect 691123 655697 691207 655700
rect 692515 655628 693915 655756
rect 694787 655628 696187 655756
rect 704735 655731 705041 655833
rect 704719 655715 705057 655731
rect 690242 655465 690442 655521
rect 692515 655465 693915 655593
rect 694787 655465 696187 655593
rect 699322 655502 700322 655574
rect 700922 655502 701922 655574
rect 707610 655547 708610 655619
rect 709211 655547 710211 655619
rect 699392 655491 699426 655502
rect 699460 655491 699494 655502
rect 699528 655491 699562 655502
rect 699596 655491 699630 655502
rect 699664 655491 699698 655502
rect 699732 655491 699766 655502
rect 699800 655491 699834 655502
rect 699868 655491 699902 655502
rect 699936 655491 699970 655502
rect 700004 655491 700038 655502
rect 700072 655491 700106 655502
rect 700140 655491 700174 655502
rect 700208 655491 700242 655502
rect 700276 655491 700310 655502
rect 700934 655491 700968 655502
rect 701002 655491 701036 655502
rect 701070 655491 701104 655502
rect 701138 655491 701172 655502
rect 701206 655491 701240 655502
rect 701274 655491 701308 655502
rect 701342 655491 701376 655502
rect 701410 655491 701444 655502
rect 701478 655491 701512 655502
rect 701546 655491 701580 655502
rect 701614 655491 701648 655502
rect 701682 655491 701716 655502
rect 701750 655491 701784 655502
rect 701818 655491 701852 655502
rect 699392 655481 699450 655491
rect 699460 655481 699518 655491
rect 699528 655481 699586 655491
rect 699596 655481 699654 655491
rect 699664 655481 699722 655491
rect 699732 655481 699790 655491
rect 699800 655481 699858 655491
rect 699868 655481 699926 655491
rect 699936 655481 699994 655491
rect 700004 655481 700062 655491
rect 700072 655481 700130 655491
rect 700140 655481 700198 655491
rect 700208 655481 700266 655491
rect 700276 655481 700334 655491
rect 700934 655481 700992 655491
rect 701002 655481 701060 655491
rect 701070 655481 701128 655491
rect 701138 655481 701196 655491
rect 701206 655481 701264 655491
rect 701274 655481 701332 655491
rect 701342 655481 701400 655491
rect 701410 655481 701468 655491
rect 701478 655481 701536 655491
rect 701546 655481 701604 655491
rect 701614 655481 701672 655491
rect 701682 655481 701740 655491
rect 701750 655481 701808 655491
rect 701818 655481 701876 655491
rect 699368 655457 700334 655481
rect 700910 655457 701876 655481
rect 699392 655442 699416 655457
rect 699460 655442 699484 655457
rect 699528 655442 699552 655457
rect 699596 655442 699620 655457
rect 699664 655442 699688 655457
rect 699732 655442 699756 655457
rect 699800 655442 699824 655457
rect 699868 655442 699892 655457
rect 699936 655442 699960 655457
rect 700004 655442 700028 655457
rect 700072 655442 700096 655457
rect 700140 655442 700164 655457
rect 700208 655442 700232 655457
rect 700276 655442 700300 655457
rect 700934 655442 700958 655457
rect 701002 655442 701026 655457
rect 701070 655442 701094 655457
rect 701138 655442 701162 655457
rect 701206 655442 701230 655457
rect 701274 655442 701298 655457
rect 701342 655442 701366 655457
rect 701410 655442 701434 655457
rect 701478 655442 701502 655457
rect 701546 655442 701570 655457
rect 701614 655442 701638 655457
rect 701682 655442 701706 655457
rect 701750 655442 701774 655457
rect 701818 655442 701842 655457
rect 690242 655289 690442 655417
rect 692515 655302 693915 655430
rect 694787 655302 696187 655430
rect 690790 655286 690874 655289
rect 691123 655286 691207 655289
rect 699322 655287 700322 655442
rect 690664 655236 691664 655286
rect 699322 655253 700334 655287
rect 700922 655277 701922 655442
rect 707610 655287 708610 655347
rect 709211 655287 710211 655347
rect 700910 655253 701922 655277
rect 699322 655242 700322 655253
rect 700922 655242 701922 655253
rect 699392 655229 699416 655242
rect 699460 655229 699484 655242
rect 699528 655229 699552 655242
rect 699596 655229 699620 655242
rect 699664 655229 699688 655242
rect 699732 655229 699756 655242
rect 699800 655229 699824 655242
rect 699868 655229 699892 655242
rect 699936 655229 699960 655242
rect 700004 655229 700028 655242
rect 700072 655229 700096 655242
rect 700140 655229 700164 655242
rect 700208 655229 700232 655242
rect 700276 655229 700300 655242
rect 700934 655229 700958 655242
rect 701002 655229 701026 655242
rect 701070 655229 701094 655242
rect 701138 655229 701162 655242
rect 701206 655229 701230 655242
rect 701274 655229 701298 655242
rect 701342 655229 701366 655242
rect 701410 655229 701434 655242
rect 701478 655229 701502 655242
rect 701546 655229 701570 655242
rect 701614 655229 701638 655242
rect 701682 655229 701706 655242
rect 701750 655229 701774 655242
rect 701818 655229 701842 655242
rect 690242 655113 690442 655169
rect 692515 655152 693915 655195
rect 694787 655152 696187 655195
rect 690664 655080 691664 655136
rect 690242 654937 690442 655065
rect 692515 655016 693915 655059
rect 694787 655016 696187 655059
rect 690664 654924 691664 654980
rect 692515 654853 693915 654981
rect 694787 654853 696187 654981
rect 703541 654944 703701 654948
rect 699322 654884 700322 654940
rect 700922 654884 701922 654940
rect 707610 654929 708610 654985
rect 709211 654929 710211 654985
rect 690242 654806 690442 654817
rect 690238 654772 690442 654806
rect 690242 654767 690442 654772
rect 690664 654768 691664 654824
rect 690242 654764 690326 654767
rect 692515 654690 693915 654818
rect 694787 654690 696187 654818
rect 699322 654812 700322 654868
rect 700922 654812 701922 654868
rect 707610 654857 708610 654913
rect 709211 654857 710211 654913
rect 703541 654798 703701 654802
rect 690664 654618 691664 654668
rect 692515 654527 693915 654655
rect 694787 654527 696187 654655
rect 699322 654510 700322 654582
rect 700922 654510 701922 654582
rect 707610 654555 708610 654627
rect 709211 654555 710211 654627
rect 699392 654499 699426 654510
rect 699460 654499 699494 654510
rect 699528 654499 699562 654510
rect 699596 654499 699630 654510
rect 699664 654499 699698 654510
rect 699732 654499 699766 654510
rect 699800 654499 699834 654510
rect 699868 654499 699902 654510
rect 699936 654499 699970 654510
rect 700004 654499 700038 654510
rect 700072 654499 700106 654510
rect 700140 654499 700174 654510
rect 700208 654499 700242 654510
rect 700276 654499 700310 654510
rect 700934 654499 700968 654510
rect 701002 654499 701036 654510
rect 701070 654499 701104 654510
rect 701138 654499 701172 654510
rect 701206 654499 701240 654510
rect 701274 654499 701308 654510
rect 701342 654499 701376 654510
rect 701410 654499 701444 654510
rect 701478 654499 701512 654510
rect 701546 654499 701580 654510
rect 701614 654499 701648 654510
rect 701682 654499 701716 654510
rect 701750 654499 701784 654510
rect 701818 654499 701852 654510
rect 692515 654364 693915 654492
rect 694787 654364 696187 654492
rect 699392 654489 699450 654499
rect 699460 654489 699518 654499
rect 699528 654489 699586 654499
rect 699596 654489 699654 654499
rect 699664 654489 699722 654499
rect 699732 654489 699790 654499
rect 699800 654489 699858 654499
rect 699868 654489 699926 654499
rect 699936 654489 699994 654499
rect 700004 654489 700062 654499
rect 700072 654489 700130 654499
rect 700140 654489 700198 654499
rect 700208 654489 700266 654499
rect 700276 654489 700334 654499
rect 700934 654489 700992 654499
rect 701002 654489 701060 654499
rect 701070 654489 701128 654499
rect 701138 654489 701196 654499
rect 701206 654489 701264 654499
rect 701274 654489 701332 654499
rect 701342 654489 701400 654499
rect 701410 654489 701468 654499
rect 701478 654489 701536 654499
rect 701546 654489 701604 654499
rect 701614 654489 701672 654499
rect 701682 654489 701740 654499
rect 701750 654489 701808 654499
rect 701818 654489 701876 654499
rect 699368 654465 700334 654489
rect 700910 654465 701876 654489
rect 699392 654450 699416 654465
rect 699460 654450 699484 654465
rect 699528 654450 699552 654465
rect 699596 654450 699620 654465
rect 699664 654450 699688 654465
rect 699732 654450 699756 654465
rect 699800 654450 699824 654465
rect 699868 654450 699892 654465
rect 699936 654450 699960 654465
rect 700004 654450 700028 654465
rect 700072 654450 700096 654465
rect 700140 654450 700164 654465
rect 700208 654450 700232 654465
rect 700276 654450 700300 654465
rect 700934 654450 700958 654465
rect 701002 654450 701026 654465
rect 701070 654450 701094 654465
rect 701138 654450 701162 654465
rect 701206 654450 701230 654465
rect 701274 654450 701298 654465
rect 701342 654450 701366 654465
rect 701410 654450 701434 654465
rect 701478 654450 701502 654465
rect 701546 654450 701570 654465
rect 701614 654450 701638 654465
rect 701682 654450 701706 654465
rect 701750 654450 701774 654465
rect 701818 654450 701842 654465
rect 692515 654201 693915 654329
rect 694787 654201 696187 654329
rect 699322 654295 700322 654450
rect 699322 654261 700334 654295
rect 700922 654285 701922 654450
rect 707610 654295 708610 654355
rect 709211 654295 710211 654355
rect 700910 654261 701922 654285
rect 699322 654250 700322 654261
rect 700922 654250 701922 654261
rect 699392 654237 699416 654250
rect 699460 654237 699484 654250
rect 699528 654237 699552 654250
rect 699596 654237 699620 654250
rect 699664 654237 699688 654250
rect 699732 654237 699756 654250
rect 699800 654237 699824 654250
rect 699868 654237 699892 654250
rect 699936 654237 699960 654250
rect 700004 654237 700028 654250
rect 700072 654237 700096 654250
rect 700140 654237 700164 654250
rect 700208 654237 700232 654250
rect 700276 654237 700300 654250
rect 700934 654237 700958 654250
rect 701002 654237 701026 654250
rect 701070 654237 701094 654250
rect 701138 654237 701162 654250
rect 701206 654237 701230 654250
rect 701274 654237 701298 654250
rect 701342 654237 701366 654250
rect 701410 654237 701434 654250
rect 701478 654237 701502 654250
rect 701546 654237 701570 654250
rect 701614 654237 701638 654250
rect 701682 654237 701706 654250
rect 701750 654237 701774 654250
rect 701818 654237 701842 654250
rect 692515 654038 693915 654166
rect 694787 654038 696187 654166
rect 692047 653468 696655 654004
rect 699322 653892 700322 653948
rect 700922 653892 701922 653948
rect 707610 653937 708610 653993
rect 709211 653937 710211 653993
rect 699322 653820 700322 653876
rect 700922 653820 701922 653876
rect 707610 653865 708610 653921
rect 709211 653865 710211 653921
rect 697314 653582 697620 653752
rect 699322 653518 700322 653590
rect 700922 653518 701922 653590
rect 707610 653563 708610 653635
rect 709211 653563 710211 653635
rect 704719 653527 705057 653543
rect 699392 653507 699426 653518
rect 699460 653507 699494 653518
rect 699528 653507 699562 653518
rect 699596 653507 699630 653518
rect 699664 653507 699698 653518
rect 699732 653507 699766 653518
rect 699800 653507 699834 653518
rect 699868 653507 699902 653518
rect 699936 653507 699970 653518
rect 700004 653507 700038 653518
rect 700072 653507 700106 653518
rect 700140 653507 700174 653518
rect 700208 653507 700242 653518
rect 700276 653507 700310 653518
rect 700934 653507 700968 653518
rect 701002 653507 701036 653518
rect 701070 653507 701104 653518
rect 701138 653507 701172 653518
rect 701206 653507 701240 653518
rect 701274 653507 701308 653518
rect 701342 653507 701376 653518
rect 701410 653507 701444 653518
rect 701478 653507 701512 653518
rect 701546 653507 701580 653518
rect 701614 653507 701648 653518
rect 701682 653507 701716 653518
rect 701750 653507 701784 653518
rect 701818 653507 701852 653518
rect 699392 653497 699450 653507
rect 699460 653497 699518 653507
rect 699528 653497 699586 653507
rect 699596 653497 699654 653507
rect 699664 653497 699722 653507
rect 699732 653497 699790 653507
rect 699800 653497 699858 653507
rect 699868 653497 699926 653507
rect 699936 653497 699994 653507
rect 700004 653497 700062 653507
rect 700072 653497 700130 653507
rect 700140 653497 700198 653507
rect 700208 653497 700266 653507
rect 700276 653497 700334 653507
rect 700934 653497 700992 653507
rect 701002 653497 701060 653507
rect 701070 653497 701128 653507
rect 701138 653497 701196 653507
rect 701206 653497 701264 653507
rect 701274 653497 701332 653507
rect 701342 653497 701400 653507
rect 701410 653497 701468 653507
rect 701478 653497 701536 653507
rect 701546 653497 701604 653507
rect 701614 653497 701672 653507
rect 701682 653497 701740 653507
rect 701750 653497 701808 653507
rect 701818 653497 701876 653507
rect 699368 653473 700334 653497
rect 700910 653473 701876 653497
rect 699392 653458 699416 653473
rect 699460 653458 699484 653473
rect 699528 653458 699552 653473
rect 699596 653458 699620 653473
rect 699664 653458 699688 653473
rect 699732 653458 699756 653473
rect 699800 653458 699824 653473
rect 699868 653458 699892 653473
rect 699936 653458 699960 653473
rect 700004 653458 700028 653473
rect 700072 653458 700096 653473
rect 700140 653458 700164 653473
rect 700208 653458 700232 653473
rect 700276 653458 700300 653473
rect 700934 653458 700958 653473
rect 701002 653458 701026 653473
rect 701070 653458 701094 653473
rect 701138 653458 701162 653473
rect 701206 653458 701230 653473
rect 701274 653458 701298 653473
rect 701342 653458 701366 653473
rect 701410 653458 701434 653473
rect 701478 653458 701502 653473
rect 701546 653458 701570 653473
rect 701614 653458 701638 653473
rect 701682 653458 701706 653473
rect 701750 653458 701774 653473
rect 701818 653458 701842 653473
rect 699322 653303 700322 653458
rect 692463 653268 692511 653292
rect 696191 653268 696239 653292
rect 692487 653214 692511 653268
rect 696215 653214 696239 653268
rect 699322 653269 700334 653303
rect 700922 653293 701922 653458
rect 704735 653425 705041 653527
rect 707610 653303 708610 653363
rect 709211 653303 710211 653363
rect 700910 653269 701922 653293
rect 699322 653258 700322 653269
rect 700922 653258 701922 653269
rect 699392 653245 699416 653258
rect 699460 653245 699484 653258
rect 699528 653245 699552 653258
rect 699596 653245 699620 653258
rect 699664 653245 699688 653258
rect 699732 653245 699756 653258
rect 699800 653245 699824 653258
rect 699868 653245 699892 653258
rect 699936 653245 699960 653258
rect 700004 653245 700028 653258
rect 700072 653245 700096 653258
rect 700140 653245 700164 653258
rect 700208 653245 700232 653258
rect 700276 653245 700300 653258
rect 700934 653245 700958 653258
rect 701002 653245 701026 653258
rect 701070 653245 701094 653258
rect 701138 653245 701162 653258
rect 701206 653245 701230 653258
rect 701274 653245 701298 653258
rect 701342 653245 701366 653258
rect 701410 653245 701434 653258
rect 701478 653245 701502 653258
rect 701546 653245 701570 653258
rect 701614 653245 701638 653258
rect 701682 653245 701706 653258
rect 701750 653245 701774 653258
rect 701818 653245 701842 653258
rect 692463 653190 692511 653214
rect 696191 653190 696239 653214
rect 687686 653119 687720 653153
rect 687798 653141 687822 653165
rect 687686 653095 687710 653119
rect 687774 653117 687798 653129
rect 687798 653081 687822 653105
rect 692450 653037 692474 653061
rect 692508 653037 692532 653061
rect 696170 653037 696194 653061
rect 696228 653037 696252 653061
rect 692484 653013 692498 653037
rect 696204 653013 696218 653037
rect 692484 652935 692487 652959
rect 696215 652935 696218 652959
rect 692508 652911 692532 652935
rect 696170 652911 696194 652935
rect 699322 652900 700322 652956
rect 700922 652900 701922 652956
rect 707610 652945 708610 653001
rect 709211 652945 710211 653001
rect 692515 652805 693915 652848
rect 694787 652805 696187 652848
rect 699322 652828 700322 652884
rect 700922 652828 701922 652884
rect 707610 652873 708610 652929
rect 709211 652873 710211 652929
rect 692515 652642 693915 652770
rect 694787 652642 696187 652770
rect 688883 652473 688918 652502
rect 692515 652479 693915 652607
rect 694787 652479 696187 652607
rect 699322 652526 700322 652598
rect 700922 652526 701922 652598
rect 707610 652571 708610 652643
rect 709211 652571 710211 652643
rect 699392 652515 699426 652526
rect 699460 652515 699494 652526
rect 699528 652515 699562 652526
rect 699596 652515 699630 652526
rect 699664 652515 699698 652526
rect 699732 652515 699766 652526
rect 699800 652515 699834 652526
rect 699868 652515 699902 652526
rect 699936 652515 699970 652526
rect 700004 652515 700038 652526
rect 700072 652515 700106 652526
rect 700140 652515 700174 652526
rect 700208 652515 700242 652526
rect 700276 652515 700310 652526
rect 700934 652515 700968 652526
rect 701002 652515 701036 652526
rect 701070 652515 701104 652526
rect 701138 652515 701172 652526
rect 701206 652515 701240 652526
rect 701274 652515 701308 652526
rect 701342 652515 701376 652526
rect 701410 652515 701444 652526
rect 701478 652515 701512 652526
rect 701546 652515 701580 652526
rect 701614 652515 701648 652526
rect 701682 652515 701716 652526
rect 701750 652515 701784 652526
rect 701818 652515 701852 652526
rect 699392 652505 699450 652515
rect 699460 652505 699518 652515
rect 699528 652505 699586 652515
rect 699596 652505 699654 652515
rect 699664 652505 699722 652515
rect 699732 652505 699790 652515
rect 699800 652505 699858 652515
rect 699868 652505 699926 652515
rect 699936 652505 699994 652515
rect 700004 652505 700062 652515
rect 700072 652505 700130 652515
rect 700140 652505 700198 652515
rect 700208 652505 700266 652515
rect 700276 652505 700334 652515
rect 700934 652505 700992 652515
rect 701002 652505 701060 652515
rect 701070 652505 701128 652515
rect 701138 652505 701196 652515
rect 701206 652505 701264 652515
rect 701274 652505 701332 652515
rect 701342 652505 701400 652515
rect 701410 652505 701468 652515
rect 701478 652505 701536 652515
rect 701546 652505 701604 652515
rect 701614 652505 701672 652515
rect 701682 652505 701740 652515
rect 701750 652505 701808 652515
rect 701818 652505 701876 652515
rect 699368 652481 700334 652505
rect 700910 652481 701876 652505
rect 688883 652468 688884 652473
rect 688917 652468 688918 652473
rect 688917 652439 688951 652468
rect 699392 652466 699416 652481
rect 699460 652466 699484 652481
rect 699528 652466 699552 652481
rect 699596 652466 699620 652481
rect 699664 652466 699688 652481
rect 699732 652466 699756 652481
rect 699800 652466 699824 652481
rect 699868 652466 699892 652481
rect 699936 652466 699960 652481
rect 700004 652466 700028 652481
rect 700072 652466 700096 652481
rect 700140 652466 700164 652481
rect 700208 652466 700232 652481
rect 700276 652466 700300 652481
rect 700934 652466 700958 652481
rect 701002 652466 701026 652481
rect 701070 652466 701094 652481
rect 701138 652466 701162 652481
rect 701206 652466 701230 652481
rect 701274 652466 701298 652481
rect 701342 652466 701366 652481
rect 701410 652466 701434 652481
rect 701478 652466 701502 652481
rect 701546 652466 701570 652481
rect 701614 652466 701638 652481
rect 701682 652466 701706 652481
rect 701750 652466 701774 652481
rect 701818 652466 701842 652481
rect 688917 652370 688951 652404
rect 688917 652301 688951 652335
rect 692515 652316 693915 652444
rect 694787 652316 696187 652444
rect 699322 652311 700322 652466
rect 688917 652232 688951 652266
rect 688917 652163 688951 652197
rect 692515 652153 693915 652281
rect 694787 652153 696187 652281
rect 699322 652277 700334 652311
rect 700922 652301 701922 652466
rect 707610 652311 708610 652371
rect 709211 652311 710211 652371
rect 700910 652277 701922 652301
rect 699322 652266 700322 652277
rect 700922 652266 701922 652277
rect 699392 652253 699416 652266
rect 699460 652253 699484 652266
rect 699528 652253 699552 652266
rect 699596 652253 699620 652266
rect 699664 652253 699688 652266
rect 699732 652253 699756 652266
rect 699800 652253 699824 652266
rect 699868 652253 699892 652266
rect 699936 652253 699960 652266
rect 700004 652253 700028 652266
rect 700072 652253 700096 652266
rect 700140 652253 700164 652266
rect 700208 652253 700232 652266
rect 700276 652253 700300 652266
rect 700934 652253 700958 652266
rect 701002 652253 701026 652266
rect 701070 652253 701094 652266
rect 701138 652253 701162 652266
rect 701206 652253 701230 652266
rect 701274 652253 701298 652266
rect 701342 652253 701366 652266
rect 701410 652253 701434 652266
rect 701478 652253 701502 652266
rect 701546 652253 701570 652266
rect 701614 652253 701638 652266
rect 701682 652253 701706 652266
rect 701750 652253 701774 652266
rect 701818 652253 701842 652266
rect 688917 652094 688951 652128
rect 688917 652025 688951 652059
rect 692515 651996 693915 652046
rect 694787 651996 696187 652046
rect 688917 651956 688951 651990
rect 698017 651933 698120 651969
rect 688917 651887 688951 651921
rect 692463 651885 692511 651909
rect 696191 651885 696239 651909
rect 688917 651818 688951 651852
rect 692487 651831 692511 651885
rect 696215 651831 696239 651885
rect 698017 651858 698053 651933
rect 692463 651807 692511 651831
rect 696191 651807 696239 651831
rect 698030 651824 698077 651858
rect 698017 651790 698053 651824
rect 688917 651749 688951 651783
rect 698030 651756 698077 651790
rect 698017 651722 698053 651756
rect 688917 651680 688951 651714
rect 698030 651688 698077 651722
rect 698017 651654 698053 651688
rect 688917 651611 688951 651645
rect 692463 651629 692521 651653
rect 696191 651629 696249 651653
rect 692487 651619 692521 651629
rect 696215 651619 696249 651629
rect 698030 651620 698077 651654
rect 698017 651586 698053 651620
rect 686879 651544 687585 651554
rect 686882 651528 687585 651544
rect 688917 651542 688951 651576
rect 692487 651547 692521 651581
rect 696215 651547 696249 651581
rect 36785 651418 37385 651474
rect 678680 651433 678704 651467
rect 681345 651399 682345 651455
rect 678680 651365 678704 651399
rect 28396 650903 28446 651361
rect 684004 651349 685004 651477
rect 688917 651473 688951 651507
rect 692487 651475 692521 651509
rect 696215 651475 696249 651509
rect 688917 651404 688951 651438
rect 692487 651427 692521 651437
rect 696215 651427 696249 651437
rect 692463 651403 692521 651427
rect 696191 651403 696249 651427
rect 688917 651335 688951 651369
rect 31049 651234 32049 651284
rect 36785 651242 37385 651298
rect 678680 651297 678704 651331
rect 678680 651229 678704 651263
rect 679133 651255 679283 651267
rect 679452 651255 679602 651267
rect 681345 651229 682345 651279
rect 678680 651161 678704 651195
rect 684004 651193 685004 651321
rect 688917 651266 688951 651300
rect 679002 651142 679602 651192
rect 36785 651072 37385 651122
rect 678680 651093 678704 651127
rect 681441 651064 681457 651130
rect 682225 651064 682241 651130
rect 37939 651039 37963 651063
rect 38085 651039 38109 651063
rect 29925 651003 29931 651032
rect 30271 651003 30305 651027
rect 30342 651003 30376 651027
rect 30413 651003 30447 651027
rect 30484 651003 30518 651027
rect 30555 651003 30589 651027
rect 30626 651003 30660 651027
rect 30697 651003 30731 651027
rect 37963 651015 37987 651038
rect 38061 651015 38085 651038
rect 678680 651025 678704 651059
rect 684004 651037 685004 651165
rect 685537 651161 686137 651211
rect 688917 651197 688951 651231
rect 692463 651214 692521 651248
rect 696191 651214 696249 651248
rect 688917 651128 688951 651162
rect 29931 650962 29939 650986
rect 29955 650962 29961 651003
rect 29891 650938 29915 650962
rect 678680 650957 678704 650991
rect 679002 650966 679602 651022
rect 25101 650860 25121 650894
rect 25125 650860 25143 650894
rect 37759 650867 37783 650891
rect 678680 650889 678704 650923
rect 681441 650902 681457 650968
rect 683625 650902 683641 650968
rect 684004 650881 685004 651009
rect 685537 651005 686137 651061
rect 688917 651059 688951 651093
rect 692515 651084 693915 651127
rect 694787 651084 696187 651127
rect 688917 650990 688951 651024
rect 688917 650921 688951 650955
rect 692515 650921 693915 651049
rect 694787 650921 696187 651049
rect 25101 650826 25147 650860
rect 37792 650843 37807 650867
rect 685537 650855 686137 650905
rect 25101 650792 25121 650826
rect 25125 650792 25143 650826
rect 678680 650821 678704 650855
rect 679002 650796 679602 650846
rect 21383 650758 21419 650792
rect 25101 650758 25147 650792
rect 21383 650724 21403 650758
rect 21407 650724 21415 650758
rect 25101 650724 25121 650758
rect 25125 650724 25143 650758
rect 678680 650753 678704 650787
rect 680502 650761 680517 650776
rect 21383 650690 21419 650724
rect 21383 650656 21403 650690
rect 21407 650656 21415 650690
rect 21481 650656 22881 650699
rect 22892 650675 22920 650703
rect 23617 650656 25017 650699
rect 25101 650690 25147 650724
rect 31458 650703 31608 650715
rect 31777 650703 31927 650715
rect 25101 650656 25121 650690
rect 25125 650656 25143 650690
rect 678680 650685 678704 650719
rect 7389 650628 8389 650632
rect 8990 650628 9990 650632
rect 7353 650578 8425 650614
rect 7353 650537 7389 650578
rect 8389 650537 8425 650578
rect 7353 650501 8425 650537
rect 8954 650578 10026 650614
rect 15678 650582 16678 650654
rect 17278 650582 18278 650654
rect 21383 650622 21419 650656
rect 25101 650622 25147 650656
rect 21383 650588 21403 650622
rect 21407 650588 21415 650622
rect 25101 650588 25121 650622
rect 25125 650588 25143 650622
rect 8954 650537 8990 650578
rect 9990 650537 10026 650578
rect 15748 650571 15782 650582
rect 15816 650571 15850 650582
rect 15884 650571 15918 650582
rect 15952 650571 15986 650582
rect 16020 650571 16054 650582
rect 16088 650571 16122 650582
rect 16156 650571 16190 650582
rect 16224 650571 16258 650582
rect 16292 650571 16326 650582
rect 16360 650571 16394 650582
rect 16428 650571 16462 650582
rect 16496 650571 16530 650582
rect 16564 650571 16598 650582
rect 16632 650571 16666 650582
rect 17290 650571 17324 650582
rect 17358 650571 17392 650582
rect 17426 650571 17460 650582
rect 17494 650571 17528 650582
rect 17562 650571 17596 650582
rect 17630 650571 17664 650582
rect 17698 650571 17732 650582
rect 17766 650571 17800 650582
rect 17834 650571 17868 650582
rect 17902 650571 17936 650582
rect 17970 650571 18004 650582
rect 18038 650571 18072 650582
rect 18106 650571 18140 650582
rect 18174 650571 18208 650582
rect 15748 650561 15806 650571
rect 15816 650561 15874 650571
rect 15884 650561 15942 650571
rect 15952 650561 16010 650571
rect 16020 650561 16078 650571
rect 16088 650561 16146 650571
rect 16156 650561 16214 650571
rect 16224 650561 16282 650571
rect 16292 650561 16350 650571
rect 16360 650561 16418 650571
rect 16428 650561 16486 650571
rect 16496 650561 16554 650571
rect 16564 650561 16622 650571
rect 16632 650561 16690 650571
rect 17290 650561 17348 650571
rect 17358 650561 17416 650571
rect 17426 650561 17484 650571
rect 17494 650561 17552 650571
rect 17562 650561 17620 650571
rect 17630 650561 17688 650571
rect 17698 650561 17756 650571
rect 17766 650561 17824 650571
rect 17834 650561 17892 650571
rect 17902 650561 17960 650571
rect 17970 650561 18028 650571
rect 18038 650561 18096 650571
rect 18106 650561 18164 650571
rect 18174 650561 18232 650571
rect 15724 650537 16690 650561
rect 17266 650537 18232 650561
rect 21383 650554 21419 650588
rect 8954 650501 10026 650537
rect 15748 650522 15772 650537
rect 15816 650522 15840 650537
rect 15884 650522 15908 650537
rect 15952 650522 15976 650537
rect 16020 650522 16044 650537
rect 16088 650522 16112 650537
rect 16156 650522 16180 650537
rect 16224 650522 16248 650537
rect 16292 650522 16316 650537
rect 16360 650522 16384 650537
rect 16428 650522 16452 650537
rect 16496 650522 16520 650537
rect 16564 650522 16588 650537
rect 16632 650522 16656 650537
rect 17290 650522 17314 650537
rect 17358 650522 17382 650537
rect 17426 650522 17450 650537
rect 17494 650522 17518 650537
rect 17562 650522 17586 650537
rect 17630 650522 17654 650537
rect 17698 650522 17722 650537
rect 17766 650522 17790 650537
rect 17834 650522 17858 650537
rect 17902 650522 17926 650537
rect 17970 650522 17994 650537
rect 18038 650522 18062 650537
rect 18106 650522 18130 650537
rect 18174 650522 18198 650537
rect 15678 650367 16678 650522
rect 7389 650277 8389 650337
rect 8990 650277 9990 650337
rect 15678 650333 16690 650367
rect 17278 650357 18278 650522
rect 17266 650333 18278 650357
rect 15678 650322 16678 650333
rect 17278 650322 18278 650333
rect 21383 650520 21403 650554
rect 21407 650520 21415 650554
rect 21481 650520 22881 650563
rect 23617 650520 25017 650563
rect 25101 650554 25147 650588
rect 25414 650573 25438 650607
rect 31458 650590 32058 650640
rect 678680 650617 678704 650651
rect 25101 650520 25121 650554
rect 25125 650520 25143 650554
rect 678680 650549 678704 650583
rect 680480 650581 680517 650761
rect 680502 650566 680517 650581
rect 680615 650761 680630 650776
rect 680803 650772 680815 650776
rect 680800 650761 680815 650772
rect 680615 650581 680815 650761
rect 681441 650740 681457 650806
rect 683625 650740 683641 650806
rect 684004 650725 685004 650853
rect 688917 650852 688951 650886
rect 688917 650783 688951 650817
rect 692515 650758 693915 650886
rect 694787 650758 696187 650886
rect 688917 650714 688951 650748
rect 686829 650649 687429 650699
rect 688917 650645 688951 650679
rect 680615 650566 680630 650581
rect 680800 650570 680815 650581
rect 681441 650578 681457 650644
rect 682225 650578 682241 650644
rect 684004 650575 685004 650625
rect 688917 650576 688951 650610
rect 692515 650595 693915 650723
rect 694787 650595 696187 650723
rect 680803 650566 680815 650570
rect 680615 650525 680630 650540
rect 680803 650536 680815 650540
rect 680800 650525 680815 650536
rect 21383 650486 21419 650520
rect 25101 650486 25147 650520
rect 21383 650452 21403 650486
rect 21407 650452 21415 650486
rect 21383 650418 21419 650452
rect 21383 650384 21403 650418
rect 21407 650384 21415 650418
rect 21383 650350 21419 650384
rect 21481 650357 22881 650485
rect 23617 650357 25017 650485
rect 25101 650452 25121 650486
rect 25125 650452 25143 650486
rect 37792 650470 37807 650494
rect 678680 650481 678704 650515
rect 25101 650418 25147 650452
rect 25101 650384 25121 650418
rect 25125 650384 25143 650418
rect 31458 650414 32058 650470
rect 37759 650446 37783 650470
rect 678680 650413 678704 650447
rect 25101 650350 25147 650384
rect 15748 650309 15772 650322
rect 15816 650309 15840 650322
rect 15884 650309 15908 650322
rect 15952 650309 15976 650322
rect 16020 650309 16044 650322
rect 16088 650309 16112 650322
rect 16156 650309 16180 650322
rect 16224 650309 16248 650322
rect 16292 650309 16316 650322
rect 16360 650309 16384 650322
rect 16428 650309 16452 650322
rect 16496 650309 16520 650322
rect 16564 650309 16588 650322
rect 16632 650309 16656 650322
rect 17290 650309 17314 650322
rect 17358 650309 17382 650322
rect 17426 650309 17450 650322
rect 17494 650309 17518 650322
rect 17562 650309 17586 650322
rect 17630 650309 17654 650322
rect 17698 650309 17722 650322
rect 17766 650309 17790 650322
rect 17834 650309 17858 650322
rect 17902 650309 17926 650322
rect 17970 650309 17994 650322
rect 18038 650309 18062 650322
rect 18106 650309 18130 650322
rect 18174 650309 18198 650322
rect 21383 650316 21403 650350
rect 21407 650316 21415 650350
rect 21383 650282 21419 650316
rect 21383 650248 21403 650282
rect 21407 650248 21415 650282
rect 21383 650214 21419 650248
rect 21383 650180 21403 650214
rect 21407 650180 21415 650214
rect 21481 650194 22881 650322
rect 23617 650194 25017 650322
rect 25101 650316 25121 650350
rect 25125 650316 25143 650350
rect 678680 650345 678704 650379
rect 679007 650370 679607 650420
rect 680615 650345 680815 650525
rect 681345 650429 682345 650479
rect 686829 650473 687429 650529
rect 688917 650507 688951 650541
rect 688917 650438 688951 650472
rect 692515 650432 693915 650560
rect 694787 650432 696187 650560
rect 684054 650373 685054 650423
rect 688917 650393 688951 650403
rect 688893 650369 688951 650393
rect 680615 650330 680630 650345
rect 680800 650334 680815 650345
rect 680803 650330 680815 650334
rect 25101 650282 25147 650316
rect 25101 650248 25121 650282
rect 25125 650248 25143 650282
rect 25101 650214 25147 650248
rect 25101 650180 25121 650214
rect 25125 650180 25143 650214
rect 25725 650197 26325 650247
rect 31458 650244 32058 650294
rect 678680 650277 678704 650311
rect 681345 650253 682345 650309
rect 30245 650220 30257 650224
rect 30245 650209 30260 650220
rect 30430 650209 30445 650224
rect 21383 650146 21419 650180
rect 7389 650066 8389 650070
rect 8990 650066 9990 650070
rect 15678 650061 16678 650133
rect 17278 650061 18278 650133
rect 21383 650112 21403 650146
rect 21407 650112 21415 650146
rect 21383 650078 21419 650112
rect 7353 650016 8425 650052
rect 7353 649975 7389 650016
rect 8389 649975 8425 650016
rect 7353 649919 8425 649975
rect 7353 649903 7389 649919
rect 8389 649903 8425 649919
rect 7353 649847 8425 649903
rect 7353 649810 7389 649847
rect 8389 649810 8425 649847
rect 7353 649770 8425 649810
rect 8954 650016 10026 650052
rect 8954 649975 8990 650016
rect 9990 649975 10026 650016
rect 8954 649919 10026 649975
rect 21383 650044 21403 650078
rect 21407 650044 21415 650078
rect 21383 650010 21419 650044
rect 21481 650031 22881 650159
rect 23617 650031 25017 650159
rect 25101 650146 25147 650180
rect 25101 650112 25121 650146
rect 25125 650112 25143 650146
rect 25101 650078 25147 650112
rect 25101 650044 25121 650078
rect 25125 650044 25143 650078
rect 25725 650047 26325 650097
rect 25101 650010 25147 650044
rect 21383 649976 21403 650010
rect 21407 649976 21415 650010
rect 21383 649942 21419 649976
rect 8954 649903 8990 649919
rect 9990 649903 10026 649919
rect 15678 649906 16678 649923
rect 17278 649906 18278 649923
rect 21383 649908 21403 649942
rect 21407 649908 21415 649942
rect 8954 649847 10026 649903
rect 20250 649890 20316 649906
rect 8954 649810 8990 649847
rect 9990 649810 10026 649847
rect 8954 649770 10026 649810
rect 21383 649874 21419 649908
rect 21383 649840 21403 649874
rect 21407 649840 21415 649874
rect 21481 649868 22881 649996
rect 23617 649868 25017 649996
rect 25101 649976 25121 650010
rect 25125 649976 25143 650010
rect 25101 649942 25147 649976
rect 25101 649908 25121 649942
rect 25125 649908 25143 649942
rect 25725 649925 26325 649975
rect 25101 649874 25147 649908
rect 25101 649840 25121 649874
rect 25125 649840 25143 649874
rect 21383 649806 21419 649840
rect 21383 649772 21403 649806
rect 21407 649772 21415 649806
rect 21383 649738 21419 649772
rect 15678 649703 16678 649736
rect 17278 649703 18278 649736
rect 21383 649704 21403 649738
rect 21407 649704 21415 649738
rect 21481 649705 22881 649833
rect 23617 649705 25017 649833
rect 25101 649806 25147 649840
rect 25101 649772 25121 649806
rect 25125 649772 25143 649806
rect 25725 649775 26325 649825
rect 25101 649738 25147 649772
rect 25101 649704 25121 649738
rect 25125 649704 25143 649738
rect 21383 649670 21419 649704
rect 25101 649670 25147 649704
rect 21383 649636 21403 649670
rect 21407 649636 21415 649670
rect 7389 649559 8389 649631
rect 8990 649559 9990 649631
rect 21383 649602 21419 649636
rect 15840 649510 15870 649580
rect 15878 649546 15908 649580
rect 21383 649568 21403 649602
rect 21407 649568 21415 649602
rect 15853 649508 15870 649510
rect 21383 649534 21419 649568
rect 21481 649542 22881 649670
rect 23617 649542 25017 649670
rect 25101 649636 25121 649670
rect 25125 649636 25143 649670
rect 25725 649649 26325 649699
rect 25101 649602 25147 649636
rect 25101 649568 25121 649602
rect 25125 649568 25143 649602
rect 25101 649534 25147 649568
rect 5981 649483 6021 649493
rect 5137 649469 6021 649483
rect 21383 649500 21403 649534
rect 21407 649500 21415 649534
rect 21383 649466 21419 649500
rect 7389 649369 8389 649463
rect 7389 649359 8413 649369
rect 8990 649359 9990 649463
rect 21383 649432 21403 649466
rect 21407 649432 21415 649466
rect 21383 649398 21419 649432
rect 21383 649364 21403 649398
rect 21407 649364 21415 649398
rect 21481 649379 22881 649507
rect 23617 649379 25017 649507
rect 25101 649500 25121 649534
rect 25125 649500 25143 649534
rect 25101 649466 25147 649500
rect 25725 649499 26325 649549
rect 25101 649432 25121 649466
rect 25125 649432 25143 649466
rect 25101 649398 25147 649432
rect 25101 649364 25121 649398
rect 25125 649364 25143 649398
rect 25725 649377 26325 649427
rect 21383 649330 21419 649364
rect 25101 649330 25147 649364
rect 21383 649296 21403 649330
rect 21407 649296 21415 649330
rect 25101 649296 25121 649330
rect 25125 649296 25143 649330
rect 21383 649262 21419 649296
rect 21383 649228 21403 649262
rect 21407 649228 21415 649262
rect 21481 649229 22881 649272
rect 23617 649229 25017 649272
rect 25101 649262 25147 649296
rect 25101 649228 25121 649262
rect 25125 649228 25143 649262
rect 21383 649194 21419 649228
rect 25101 649194 25147 649228
rect 25725 649227 26325 649277
rect 21383 649160 21403 649194
rect 21407 649160 21415 649194
rect 25101 649160 25121 649194
rect 25125 649160 25143 649194
rect 27162 649170 27212 650170
rect 27312 649170 27440 650170
rect 27468 649170 27596 650170
rect 27624 649170 27752 650170
rect 27780 649170 27908 650170
rect 27936 649170 28064 650170
rect 28092 649170 28220 650170
rect 28248 649170 28376 650170
rect 28404 649170 28532 650170
rect 28560 649170 28688 650170
rect 28716 649170 28844 650170
rect 28872 649170 29000 650170
rect 29028 649170 29156 650170
rect 29184 649170 29312 650170
rect 29340 649170 29390 650170
rect 30245 650029 30445 650209
rect 30245 650018 30260 650029
rect 30245 650014 30257 650018
rect 30430 650014 30445 650029
rect 30543 650209 30558 650224
rect 678680 650209 678704 650243
rect 30543 650029 30580 650209
rect 679007 650200 679607 650250
rect 684054 650217 685054 650345
rect 686829 650303 687429 650353
rect 692515 650269 693915 650397
rect 694787 650269 696187 650397
rect 678680 650141 678704 650175
rect 678680 650073 678704 650107
rect 681345 650077 682345 650205
rect 30543 650014 30558 650029
rect 678680 650005 678704 650039
rect 680215 650024 680815 650074
rect 684054 650061 685054 650189
rect 685793 650182 685805 650186
rect 685793 650171 685808 650182
rect 685978 650171 685993 650186
rect 30245 649984 30257 649988
rect 30245 649973 30260 649984
rect 30430 649973 30445 649988
rect 30245 649793 30445 649973
rect 678680 649937 678704 649971
rect 678680 649869 678704 649903
rect 31453 649818 32053 649868
rect 680215 649848 680815 649904
rect 681345 649901 682345 650029
rect 684054 649905 685054 650033
rect 685793 649991 685993 650171
rect 685793 649980 685808 649991
rect 685793 649976 685805 649980
rect 685978 649976 685993 649991
rect 686053 650182 686065 650186
rect 686053 650171 686068 650182
rect 686238 650171 686253 650186
rect 686053 649991 686253 650171
rect 686607 650164 687607 650214
rect 697088 650171 697138 651571
rect 697238 650171 697366 651571
rect 697394 650171 697522 651571
rect 697550 650171 697678 651571
rect 697706 650171 697756 651571
rect 698030 651552 698077 651586
rect 698017 651518 698053 651552
rect 698030 651484 698077 651518
rect 698017 651450 698053 651484
rect 698030 651416 698077 651450
rect 698017 651382 698053 651416
rect 698030 651348 698077 651382
rect 698017 651314 698053 651348
rect 698030 651280 698077 651314
rect 698017 651246 698053 651280
rect 698030 651212 698077 651246
rect 698017 651178 698053 651212
rect 698030 651144 698077 651178
rect 698017 651110 698053 651144
rect 698030 651076 698077 651110
rect 698017 651042 698053 651076
rect 698030 651008 698077 651042
rect 698017 650974 698053 651008
rect 698030 650940 698077 650974
rect 698017 650906 698053 650940
rect 698030 650872 698077 650906
rect 698017 650838 698053 650872
rect 698030 650804 698077 650838
rect 698017 650770 698053 650804
rect 698030 650736 698077 650770
rect 698017 650702 698053 650736
rect 698030 650668 698077 650702
rect 698017 650634 698053 650668
rect 698030 650600 698077 650634
rect 698017 650566 698053 650600
rect 698030 650532 698077 650566
rect 698017 650498 698053 650532
rect 698030 650464 698077 650498
rect 698017 650430 698053 650464
rect 698030 650396 698077 650430
rect 698017 650362 698053 650396
rect 698030 650328 698077 650362
rect 698017 650294 698053 650328
rect 698030 650260 698077 650294
rect 698017 650226 698053 650260
rect 698030 650192 698077 650226
rect 692515 650119 693915 650162
rect 694787 650119 696187 650162
rect 698017 650158 698053 650192
rect 698030 650124 698077 650158
rect 698017 650090 698053 650124
rect 686607 650014 687607 650064
rect 698030 650056 698077 650090
rect 686053 649980 686068 649991
rect 686053 649976 686065 649980
rect 686238 649976 686253 649991
rect 685793 649946 685805 649950
rect 685793 649935 685808 649946
rect 685978 649935 685993 649950
rect 678680 649801 678704 649835
rect 30245 649782 30260 649793
rect 30245 649778 30257 649782
rect 30430 649778 30445 649793
rect 678680 649733 678704 649767
rect 681345 649731 682345 649781
rect 684054 649749 685054 649877
rect 685793 649755 685993 649935
rect 685793 649744 685808 649755
rect 685793 649740 685805 649744
rect 685978 649740 685993 649755
rect 686053 649946 686065 649950
rect 686053 649935 686068 649946
rect 686238 649935 686253 649950
rect 686053 649755 686253 649935
rect 686607 649855 687607 649905
rect 692463 649809 692511 649833
rect 696191 649809 696239 649833
rect 686053 649744 686068 649755
rect 686053 649740 686065 649744
rect 686238 649740 686253 649755
rect 31453 649648 32053 649698
rect 678680 649665 678704 649699
rect 680215 649672 680815 649728
rect 681345 649662 682345 649674
rect 678680 649597 678704 649631
rect 684054 649593 685054 649721
rect 686607 649705 687607 649755
rect 692487 649731 692511 649809
rect 696215 649755 696239 649809
rect 696191 649731 696239 649755
rect 696617 649772 696651 649773
rect 696617 649749 696626 649772
rect 696617 649731 696675 649749
rect 696651 649715 696675 649731
rect 696651 649647 696675 649681
rect 685533 649586 685545 649590
rect 685533 649575 685548 649586
rect 685718 649575 685733 649590
rect 678680 649529 678704 649563
rect 30245 649472 30845 649522
rect 680215 649502 680815 649552
rect 678680 649461 678704 649495
rect 678680 649393 678704 649427
rect 680215 649370 680815 649420
rect 681466 649411 682466 649461
rect 684054 649437 685054 649565
rect 30245 649296 30845 649352
rect 678680 649325 678704 649359
rect 678680 649257 678704 649291
rect 681466 649255 682466 649383
rect 682890 649339 683490 649389
rect 678680 649189 678704 649223
rect 680215 649194 680815 649250
rect 682890 649183 683490 649311
rect 684054 649281 685054 649409
rect 685533 649395 685733 649575
rect 685533 649384 685548 649395
rect 685533 649380 685545 649384
rect 685718 649380 685733 649395
rect 685793 649586 685805 649590
rect 685793 649575 685808 649586
rect 685978 649575 685993 649590
rect 685793 649395 685993 649575
rect 685793 649384 685808 649395
rect 685793 649380 685805 649384
rect 685978 649380 685993 649395
rect 686053 649586 686065 649590
rect 686053 649575 686068 649586
rect 686238 649575 686253 649590
rect 686053 649395 686253 649575
rect 686053 649384 686068 649395
rect 686053 649380 686065 649384
rect 686238 649380 686253 649395
rect 686313 649586 686325 649590
rect 686313 649575 686328 649586
rect 686498 649575 686513 649590
rect 686313 649395 686513 649575
rect 686313 649384 686328 649395
rect 686313 649380 686325 649384
rect 686498 649380 686513 649395
rect 686627 649586 686639 649590
rect 686627 649575 686642 649586
rect 686812 649575 686827 649590
rect 686627 649395 686827 649575
rect 686627 649384 686642 649395
rect 686627 649380 686639 649384
rect 686812 649380 686827 649395
rect 686887 649586 686899 649590
rect 686887 649575 686902 649586
rect 687072 649575 687087 649590
rect 686887 649395 687087 649575
rect 686887 649384 686902 649395
rect 686887 649380 686899 649384
rect 687072 649380 687087 649395
rect 687147 649586 687159 649590
rect 687147 649575 687162 649586
rect 687332 649575 687347 649590
rect 696651 649579 696675 649613
rect 687147 649395 687347 649575
rect 696651 649511 696675 649545
rect 696651 649443 696675 649477
rect 687147 649384 687162 649395
rect 687147 649380 687159 649384
rect 687332 649380 687347 649395
rect 696651 649375 696675 649409
rect 696651 649307 696675 649341
rect 685718 649215 685733 649230
rect 685679 649185 685733 649215
rect 21383 649126 21419 649160
rect 25101 649126 25147 649160
rect 21383 649102 21403 649126
rect 21385 649048 21403 649102
rect 21407 649082 21415 649126
rect 25101 649102 25121 649126
rect 25113 649082 25121 649102
rect 25125 649048 25143 649126
rect 30245 649120 30845 649176
rect 678680 649121 678704 649155
rect 681466 649105 682466 649155
rect 684054 649131 685054 649181
rect 685718 649170 685733 649185
rect 685793 649226 685805 649230
rect 685793 649215 685808 649226
rect 685978 649215 685993 649230
rect 685793 649185 685993 649215
rect 685793 649174 685808 649185
rect 685793 649170 685805 649174
rect 685978 649170 685993 649185
rect 686053 649226 686065 649230
rect 686053 649215 686068 649226
rect 686238 649215 686253 649230
rect 686812 649215 686827 649230
rect 686053 649185 686253 649215
rect 686807 649185 686827 649215
rect 686053 649174 686068 649185
rect 686053 649170 686065 649174
rect 686238 649170 686253 649185
rect 686812 649170 686827 649185
rect 686887 649226 686899 649230
rect 686887 649215 686902 649226
rect 687072 649215 687087 649230
rect 686887 649185 687087 649215
rect 686887 649174 686902 649185
rect 686887 649170 686899 649174
rect 687072 649170 687087 649185
rect 687147 649226 687159 649230
rect 687147 649215 687162 649226
rect 687332 649215 687347 649230
rect 687147 649185 687347 649215
rect 687147 649174 687162 649185
rect 687147 649170 687159 649174
rect 687332 649170 687347 649185
rect 685718 649129 685733 649144
rect 681794 649102 682466 649105
rect 685679 649099 685733 649129
rect 678680 649053 678704 649087
rect 685718 649084 685733 649099
rect 685793 649140 685805 649144
rect 685793 649129 685808 649140
rect 685978 649129 685993 649144
rect 685793 649099 685993 649129
rect 685793 649088 685808 649099
rect 685793 649084 685805 649088
rect 685978 649084 685993 649099
rect 686053 649140 686065 649144
rect 686053 649129 686068 649140
rect 686238 649129 686253 649144
rect 686812 649129 686827 649144
rect 686053 649099 686253 649129
rect 686807 649099 686827 649129
rect 686053 649088 686068 649099
rect 686053 649084 686065 649088
rect 686238 649084 686253 649099
rect 686812 649084 686827 649099
rect 686887 649140 686899 649144
rect 686887 649129 686902 649140
rect 687072 649129 687087 649144
rect 686887 649099 687087 649129
rect 686887 649088 686902 649099
rect 686887 649084 686899 649088
rect 687072 649084 687087 649099
rect 687147 649140 687159 649144
rect 687147 649129 687162 649140
rect 687332 649129 687347 649144
rect 687147 649099 687347 649129
rect 687147 649088 687162 649099
rect 687147 649084 687159 649088
rect 687332 649084 687347 649099
rect 30245 648950 30845 649000
rect 678680 648985 678704 649019
rect 680215 649018 680815 649074
rect 682890 649027 683490 649083
rect 21000 648800 21003 648920
rect 678680 648917 678704 648951
rect 21352 648885 21376 648909
rect 25122 648885 25146 648909
rect 21385 648861 21400 648885
rect 25098 648861 25113 648885
rect 21274 648783 21294 648851
rect 21410 648817 21430 648851
rect 25068 648817 25088 648851
rect 25204 648817 25224 648851
rect 678680 648849 678704 648883
rect 680215 648848 680815 648898
rect 21385 648807 21430 648817
rect 25102 648807 25137 648817
rect 21361 648783 21430 648807
rect 25089 648783 25137 648807
rect 25238 648783 25258 648817
rect 678680 648781 678704 648815
rect 678680 648713 678704 648747
rect 678680 648645 678704 648679
rect 679007 648672 679607 648722
rect 678680 648577 678704 648611
rect 680615 648577 680630 648592
rect 680803 648588 680815 648592
rect 680800 648577 680815 648588
rect 678680 648509 678704 648543
rect 679007 648502 679607 648552
rect 678680 648441 678704 648475
rect 678680 648373 678704 648407
rect 680615 648397 680815 648577
rect 681502 648505 681529 648995
rect 681866 648896 682466 649024
rect 682890 648871 683490 648999
rect 684004 648929 685004 648979
rect 685539 648940 685777 648972
rect 685803 648920 686119 648938
rect 681866 648740 682466 648868
rect 684004 648773 685004 648901
rect 682890 648721 683490 648771
rect 681866 648584 682466 648712
rect 682890 648605 683490 648655
rect 684004 648617 685004 648745
rect 681866 648434 682466 648484
rect 682890 648449 683490 648505
rect 684004 648461 685004 648589
rect 692427 648522 693027 648572
rect 680615 648382 680630 648397
rect 680800 648386 680815 648397
rect 680803 648382 680815 648386
rect 680502 648341 680517 648356
rect 678680 648305 678704 648339
rect 678680 648237 678704 648271
rect 678680 648169 678704 648203
rect 680480 648161 680517 648341
rect 680502 648146 680517 648161
rect 680615 648341 680630 648356
rect 680803 648352 680815 648356
rect 680800 648341 680815 648352
rect 680615 648161 680815 648341
rect 681866 648318 682466 648368
rect 682890 648293 683490 648349
rect 684004 648305 685004 648433
rect 692427 648366 693027 648494
rect 693888 648375 694194 648545
rect 694388 648375 694694 648545
rect 689309 648278 689909 648328
rect 681866 648168 682466 648218
rect 682041 648165 682385 648168
rect 680615 648146 680630 648161
rect 680800 648150 680815 648161
rect 680803 648146 680815 648150
rect 682890 648137 683490 648193
rect 684004 648149 685004 648277
rect 678680 648101 678704 648135
rect 679002 648076 679602 648126
rect 689309 648122 689909 648250
rect 692427 648210 693027 648338
rect 678680 648033 678704 648067
rect 678680 647965 678704 647999
rect 682890 647981 683490 648109
rect 684004 647993 685004 648121
rect 689309 647966 689909 648094
rect 692427 648054 693027 648110
rect 678680 647897 678704 647931
rect 679002 647900 679602 647956
rect 678680 647829 678704 647863
rect 682890 647825 683490 647953
rect 684004 647837 685004 647965
rect 692427 647898 693027 648026
rect 689309 647810 689909 647866
rect 678680 647761 678704 647795
rect 679002 647730 679602 647780
rect 679061 647727 679355 647730
rect 679380 647727 679602 647730
rect 678680 647693 678704 647727
rect 682890 647669 683490 647797
rect 684004 647687 685004 647737
rect 685803 647720 686119 647732
rect 685539 647716 686119 647720
rect 685513 647682 685537 647716
rect 685539 647682 685777 647716
rect 678680 647625 678704 647659
rect 689309 647654 689909 647782
rect 690910 647754 691110 647765
rect 692427 647742 693027 647870
rect 690910 647640 691110 647690
rect 678680 647557 678704 647591
rect 678680 647489 678704 647523
rect 682890 647513 683490 647569
rect 685718 647555 685733 647570
rect 684004 647485 685004 647535
rect 685679 647525 685733 647555
rect 685718 647510 685733 647525
rect 685793 647566 685805 647570
rect 685793 647555 685808 647566
rect 685978 647555 685993 647570
rect 685793 647525 685993 647555
rect 685793 647514 685808 647525
rect 685793 647510 685805 647514
rect 685978 647510 685993 647525
rect 686053 647566 686065 647570
rect 686053 647555 686068 647566
rect 686238 647555 686253 647570
rect 686812 647555 686827 647570
rect 686053 647525 686253 647555
rect 686807 647525 686827 647555
rect 686053 647514 686068 647525
rect 686053 647510 686065 647514
rect 686238 647510 686253 647525
rect 686812 647510 686827 647525
rect 686887 647566 686899 647570
rect 686887 647555 686902 647566
rect 687072 647555 687087 647570
rect 686887 647525 687087 647555
rect 686887 647514 686902 647525
rect 686887 647510 686899 647514
rect 687072 647510 687087 647525
rect 687147 647566 687159 647570
rect 687147 647555 687162 647566
rect 687332 647555 687347 647570
rect 687147 647525 687347 647555
rect 687147 647514 687162 647525
rect 687147 647510 687159 647514
rect 687332 647510 687347 647525
rect 689309 647498 689909 647626
rect 692427 647592 693027 647642
rect 693888 647575 694194 647745
rect 694388 647575 694694 647745
rect 678680 647421 678704 647455
rect 678680 647353 678704 647387
rect 682890 647357 683490 647485
rect 690910 647484 691110 647540
rect 685718 647469 685733 647484
rect 684004 647329 685004 647457
rect 685679 647439 685733 647469
rect 685718 647424 685733 647439
rect 685793 647480 685805 647484
rect 685793 647469 685808 647480
rect 685978 647469 685993 647484
rect 685793 647439 685993 647469
rect 685793 647428 685808 647439
rect 685793 647424 685805 647428
rect 685978 647424 685993 647439
rect 686053 647480 686065 647484
rect 686053 647469 686068 647480
rect 686238 647469 686253 647484
rect 686812 647469 686827 647484
rect 686053 647439 686253 647469
rect 686807 647439 686827 647469
rect 686053 647428 686068 647439
rect 686053 647424 686065 647428
rect 686238 647424 686253 647439
rect 686812 647424 686827 647439
rect 686887 647480 686899 647484
rect 686887 647469 686902 647480
rect 687072 647469 687087 647484
rect 686887 647439 687087 647469
rect 686887 647428 686902 647439
rect 686887 647424 686899 647428
rect 687072 647424 687087 647439
rect 687147 647480 687159 647484
rect 687147 647469 687162 647480
rect 687332 647469 687347 647484
rect 687147 647439 687347 647469
rect 692427 647462 693027 647512
rect 687147 647428 687162 647439
rect 687147 647424 687159 647428
rect 687332 647424 687347 647439
rect 689309 647348 689909 647398
rect 690910 647334 691110 647384
rect 678680 647285 678704 647319
rect 678680 647217 678704 647251
rect 682890 647201 683490 647329
rect 692427 647312 693027 647362
rect 678680 647149 678704 647183
rect 684004 647173 685004 647301
rect 685533 647270 685545 647274
rect 685533 647259 685548 647270
rect 685718 647259 685733 647274
rect 678680 647081 678704 647115
rect 679133 647101 679283 647113
rect 679452 647101 679602 647113
rect 678680 647013 678704 647047
rect 682890 647045 683490 647173
rect 679002 646988 679602 647038
rect 684004 647017 685004 647145
rect 685533 647079 685733 647259
rect 685533 647068 685548 647079
rect 685533 647064 685545 647068
rect 685718 647064 685733 647079
rect 685793 647270 685805 647274
rect 685793 647259 685808 647270
rect 685978 647259 685993 647274
rect 685793 647079 685993 647259
rect 685793 647068 685808 647079
rect 685793 647064 685805 647068
rect 685978 647064 685993 647079
rect 686053 647270 686065 647274
rect 686053 647259 686068 647270
rect 686238 647259 686253 647274
rect 686053 647079 686253 647259
rect 686053 647068 686068 647079
rect 686053 647064 686065 647068
rect 686238 647064 686253 647079
rect 686313 647270 686325 647274
rect 686313 647259 686328 647270
rect 686498 647259 686513 647274
rect 686313 647079 686513 647259
rect 686313 647068 686328 647079
rect 686313 647064 686325 647068
rect 686498 647064 686513 647079
rect 686627 647270 686639 647274
rect 686627 647259 686642 647270
rect 686812 647259 686827 647274
rect 686627 647079 686827 647259
rect 686627 647068 686642 647079
rect 686627 647064 686639 647068
rect 686812 647064 686827 647079
rect 686887 647270 686899 647274
rect 686887 647259 686902 647270
rect 687072 647259 687087 647274
rect 686887 647079 687087 647259
rect 686887 647068 686902 647079
rect 686887 647064 686899 647068
rect 687072 647064 687087 647079
rect 687147 647270 687159 647274
rect 687147 647259 687162 647270
rect 687332 647259 687347 647274
rect 687147 647079 687347 647259
rect 689309 647218 689909 647268
rect 692427 647140 693027 647190
rect 687147 647068 687162 647079
rect 687147 647064 687159 647068
rect 687332 647064 687347 647079
rect 689309 647068 689909 647118
rect 692427 646990 693027 647040
rect 678680 646945 678704 646979
rect 678680 646877 678704 646911
rect 682890 646895 683490 646945
rect 678680 646809 678704 646843
rect 679002 646812 679602 646868
rect 684004 646861 685004 646917
rect 685793 646910 685805 646914
rect 685793 646899 685808 646910
rect 685978 646899 685993 646914
rect 682890 646779 683490 646829
rect 678680 646741 678704 646775
rect 678680 646673 678704 646707
rect 679002 646642 679602 646692
rect 678680 646605 678704 646639
rect 682890 646623 683490 646751
rect 684004 646705 685004 646833
rect 685793 646719 685993 646899
rect 685793 646708 685808 646719
rect 685793 646704 685805 646708
rect 685978 646704 685993 646719
rect 686053 646910 686065 646914
rect 686053 646899 686068 646910
rect 686238 646899 686253 646914
rect 686607 646899 687607 646949
rect 690910 646934 691110 646984
rect 686053 646719 686253 646899
rect 692427 646860 693027 646910
rect 686607 646749 687607 646799
rect 690910 646778 691110 646834
rect 686053 646708 686068 646719
rect 686053 646704 686065 646708
rect 686238 646704 686253 646719
rect 692427 646704 693027 646832
rect 693888 646775 694194 646945
rect 694388 646775 694694 646945
rect 680502 646607 680517 646622
rect 678680 646537 678704 646571
rect 678680 646469 678704 646503
rect 678680 646401 678704 646435
rect 680480 646427 680517 646607
rect 680502 646412 680517 646427
rect 680615 646607 680630 646622
rect 680803 646618 680815 646622
rect 680800 646607 680815 646618
rect 680615 646427 680815 646607
rect 682890 646467 683490 646595
rect 684004 646549 685004 646677
rect 685793 646674 685805 646678
rect 685793 646663 685808 646674
rect 685978 646663 685993 646678
rect 680615 646412 680630 646427
rect 680800 646416 680815 646427
rect 680803 646412 680815 646416
rect 680615 646371 680630 646386
rect 680803 646382 680815 646386
rect 680800 646371 680815 646382
rect 678680 646333 678704 646367
rect 678680 646265 678704 646299
rect 678680 646197 678704 646231
rect 679007 646216 679607 646266
rect 680615 646191 680815 646371
rect 682890 646311 683490 646439
rect 684004 646393 685004 646521
rect 685793 646483 685993 646663
rect 685793 646472 685808 646483
rect 685793 646468 685805 646472
rect 685978 646468 685993 646483
rect 686053 646674 686065 646678
rect 686053 646663 686068 646674
rect 686238 646663 686253 646678
rect 686053 646483 686253 646663
rect 686607 646590 687607 646640
rect 690910 646628 691110 646678
rect 692427 646548 693027 646676
rect 686053 646472 686068 646483
rect 686053 646468 686065 646472
rect 686238 646468 686253 646483
rect 686607 646440 687607 646490
rect 692427 646392 693027 646448
rect 686829 646301 687429 646351
rect 684004 646243 685004 646293
rect 692427 646236 693027 646364
rect 695201 646282 695251 649282
rect 695351 646282 695479 649282
rect 695507 646282 695635 649282
rect 695663 646282 695791 649282
rect 695819 646282 695947 649282
rect 695975 646282 696103 649282
rect 696131 646282 696259 649282
rect 696287 646282 696337 649282
rect 696651 649239 696675 649273
rect 696651 649171 696675 649205
rect 696651 649103 696675 649137
rect 696651 649035 696675 649069
rect 696651 648967 696675 649001
rect 696651 648899 696675 648933
rect 696651 648831 696675 648865
rect 696651 648763 696675 648797
rect 696651 648695 696675 648729
rect 696651 648627 696675 648661
rect 697088 648641 697138 650041
rect 697238 648641 697366 650041
rect 697394 648641 697522 650041
rect 697550 648641 697678 650041
rect 697706 648641 697756 650041
rect 698017 650022 698053 650056
rect 698030 649988 698077 650022
rect 698017 649954 698053 649988
rect 698030 649920 698077 649954
rect 698017 649886 698053 649920
rect 698030 649852 698077 649886
rect 698017 649818 698053 649852
rect 698030 649784 698077 649818
rect 698017 649750 698053 649784
rect 698030 649716 698077 649750
rect 698017 649682 698053 649716
rect 698030 649648 698077 649682
rect 698017 649614 698053 649648
rect 698030 649580 698077 649614
rect 698017 649546 698053 649580
rect 698030 649512 698077 649546
rect 698017 649478 698053 649512
rect 698030 649444 698077 649478
rect 698017 649410 698053 649444
rect 698030 649376 698077 649410
rect 698017 649342 698053 649376
rect 698030 649308 698077 649342
rect 698017 649274 698053 649308
rect 698030 649240 698077 649274
rect 698017 649206 698053 649240
rect 698030 649172 698077 649206
rect 698017 649138 698053 649172
rect 698030 649104 698077 649138
rect 698017 649070 698053 649104
rect 698030 649036 698077 649070
rect 698017 649002 698053 649036
rect 698030 648968 698077 649002
rect 698017 648934 698053 648968
rect 698030 648900 698077 648934
rect 698017 648866 698053 648900
rect 698030 648832 698077 648866
rect 698017 648798 698053 648832
rect 698030 648764 698077 648798
rect 698017 648730 698053 648764
rect 698030 648696 698077 648730
rect 698017 648662 698053 648696
rect 698030 648628 698077 648662
rect 698017 648594 698053 648628
rect 696651 648559 696675 648593
rect 698030 648560 698077 648594
rect 698017 648526 698053 648560
rect 696651 648491 696675 648525
rect 698030 648492 698077 648526
rect 696651 648423 696675 648457
rect 698017 648428 698053 648492
rect 698030 648394 698077 648428
rect 696651 648355 696675 648389
rect 698017 648360 698053 648394
rect 698030 648326 698077 648360
rect 696651 648287 696675 648321
rect 698017 648292 698053 648326
rect 696651 648219 696675 648253
rect 696651 648151 696675 648185
rect 696651 648083 696675 648117
rect 696651 648015 696675 648049
rect 696651 647947 696675 647981
rect 696651 647879 696675 647913
rect 696651 647811 696675 647845
rect 696651 647743 696675 647777
rect 696651 647675 696675 647709
rect 696651 647607 696675 647641
rect 696651 647539 696675 647573
rect 696651 647471 696675 647505
rect 696651 647403 696675 647437
rect 696651 647335 696675 647369
rect 696651 647267 696675 647301
rect 696651 647199 696675 647233
rect 696651 647131 696675 647165
rect 696651 647063 696675 647097
rect 696651 646995 696675 647029
rect 696651 646927 696675 646961
rect 696651 646859 696675 646893
rect 697088 646879 697138 648279
rect 697238 646879 697366 648279
rect 697394 646879 697522 648279
rect 697550 646879 697678 648279
rect 697706 646879 697756 648279
rect 698030 648258 698077 648292
rect 698017 648224 698053 648258
rect 698030 648190 698077 648224
rect 698017 648156 698053 648190
rect 698030 648122 698077 648156
rect 698017 648088 698053 648122
rect 698030 648054 698077 648088
rect 698017 648020 698053 648054
rect 698030 647986 698077 648020
rect 698017 647952 698053 647986
rect 698030 647918 698077 647952
rect 698017 647884 698053 647918
rect 698030 647850 698077 647884
rect 698017 647816 698053 647850
rect 698030 647782 698077 647816
rect 698017 647748 698053 647782
rect 698030 647714 698077 647748
rect 698017 647680 698053 647714
rect 698030 647646 698077 647680
rect 698017 647612 698053 647646
rect 698030 647578 698077 647612
rect 698017 647544 698053 647578
rect 698030 647510 698077 647544
rect 698017 647476 698053 647510
rect 698030 647442 698077 647476
rect 698017 647408 698053 647442
rect 698030 647374 698077 647408
rect 698017 647340 698053 647374
rect 698030 647306 698077 647340
rect 698017 647272 698053 647306
rect 698030 647238 698077 647272
rect 698017 647204 698053 647238
rect 698030 647170 698077 647204
rect 698017 647136 698053 647170
rect 698030 647102 698077 647136
rect 698017 647068 698053 647102
rect 698030 647034 698077 647068
rect 698017 647000 698053 647034
rect 698030 646966 698077 647000
rect 698017 646932 698053 646966
rect 698030 646898 698077 646932
rect 698017 646864 698053 646898
rect 698030 646830 698077 646864
rect 696651 646791 696675 646825
rect 698017 646796 698053 646830
rect 698030 646762 698077 646796
rect 696651 646723 696675 646757
rect 696651 646655 696675 646689
rect 696651 646587 696675 646621
rect 696651 646519 696675 646553
rect 696651 646451 696675 646485
rect 696651 646383 696675 646417
rect 696651 646315 696675 646349
rect 696651 646247 696675 646281
rect 680615 646176 680630 646191
rect 680800 646180 680815 646191
rect 680803 646176 680815 646180
rect 678680 646129 678704 646163
rect 682890 646161 683490 646211
rect 684004 646127 685004 646177
rect 686829 646125 687429 646181
rect 678680 646061 678704 646095
rect 679007 646046 679607 646096
rect 692427 646080 693027 646208
rect 696651 646179 696675 646213
rect 696651 646111 696675 646145
rect 696651 646043 696675 646077
rect 678680 645993 678704 646027
rect 681664 646002 681812 646006
rect 681641 645994 681812 646002
rect 682113 645994 682313 646006
rect 684004 645971 685004 646027
rect 678680 645925 678704 645959
rect 686829 645955 687429 646005
rect 678680 645857 678704 645891
rect 680215 645870 680815 645920
rect 681713 645881 682313 645931
rect 682921 645899 683521 645949
rect 692427 645930 693027 645980
rect 696651 645975 696675 646009
rect 696651 645907 696675 645941
rect 678680 645789 678704 645823
rect 684004 645821 685004 645871
rect 678680 645721 678704 645755
rect 680215 645694 680815 645750
rect 681713 645705 682313 645761
rect 682921 645743 683521 645799
rect 685537 645749 686137 645799
rect 697088 645749 697138 646749
rect 697238 645749 697366 646749
rect 697394 645749 697522 646749
rect 697550 645749 697678 646749
rect 697706 645749 697756 646749
rect 698017 646728 698053 646762
rect 698030 646694 698077 646728
rect 698017 646660 698053 646694
rect 698030 646626 698077 646660
rect 698017 646592 698053 646626
rect 698030 646558 698077 646592
rect 698017 646524 698053 646558
rect 698030 646490 698077 646524
rect 698017 646456 698053 646490
rect 698030 646422 698077 646456
rect 698017 646388 698053 646422
rect 698030 646354 698077 646388
rect 698017 646320 698053 646354
rect 698030 646286 698077 646320
rect 698017 646252 698053 646286
rect 698030 646218 698077 646252
rect 698017 646184 698053 646218
rect 698030 646150 698077 646184
rect 698017 646116 698053 646150
rect 698030 646082 698077 646116
rect 698017 646048 698053 646082
rect 698030 646014 698077 646048
rect 698017 645980 698053 646014
rect 698030 645946 698077 645980
rect 698017 645912 698053 645946
rect 698030 645878 698077 645912
rect 698017 645844 698053 645878
rect 698030 645810 698077 645844
rect 698017 645776 698053 645810
rect 698030 645742 698077 645776
rect 698017 645708 698053 645742
rect 678680 645653 678704 645687
rect 698030 645674 698077 645708
rect 678680 645585 678704 645619
rect 680215 645518 680815 645574
rect 681713 645529 682313 645657
rect 682921 645593 683521 645643
rect 684070 645599 684670 645649
rect 685537 645593 686137 645649
rect 698017 645640 698053 645674
rect 698030 645606 698077 645640
rect 698017 645572 698053 645606
rect 698030 645538 698077 645572
rect 698017 645504 698053 645538
rect 684070 645443 684670 645499
rect 685537 645443 686137 645493
rect 692428 645442 693028 645492
rect 698030 645470 698077 645504
rect 698017 645436 698053 645470
rect 680215 645348 680815 645398
rect 681713 645359 682313 645409
rect 698030 645402 698077 645436
rect 698017 645368 698053 645402
rect 684070 645293 684670 645343
rect 692428 645292 693028 645342
rect 698030 645334 698077 645368
rect 698017 645300 698053 645334
rect 680215 645232 680815 645282
rect 698030 645266 698077 645300
rect 698017 645232 698053 645266
rect 692428 645162 693028 645212
rect 698030 645198 698077 645232
rect 698017 645164 698053 645198
rect 680215 645056 680815 645112
rect 692428 645006 693028 645134
rect 698030 645130 698077 645164
rect 698017 645096 698053 645130
rect 698030 645062 698077 645096
rect 698017 644983 698053 645062
rect 698084 644983 698120 651933
rect 699322 651908 700322 651964
rect 700922 651908 701922 651964
rect 707610 651953 708610 652009
rect 709211 651953 710211 652009
rect 699322 651836 700322 651892
rect 700922 651836 701922 651892
rect 707610 651881 708610 651937
rect 709211 651881 710211 651937
rect 699322 651534 700322 651606
rect 700922 651534 701922 651606
rect 707610 651579 708610 651651
rect 709211 651579 710211 651651
rect 699392 651523 699426 651534
rect 699460 651523 699494 651534
rect 699528 651523 699562 651534
rect 699596 651523 699630 651534
rect 699664 651523 699698 651534
rect 699732 651523 699766 651534
rect 699800 651523 699834 651534
rect 699868 651523 699902 651534
rect 699936 651523 699970 651534
rect 700004 651523 700038 651534
rect 700072 651523 700106 651534
rect 700140 651523 700174 651534
rect 700208 651523 700242 651534
rect 700276 651523 700310 651534
rect 700934 651523 700968 651534
rect 701002 651523 701036 651534
rect 701070 651523 701104 651534
rect 701138 651523 701172 651534
rect 701206 651523 701240 651534
rect 701274 651523 701308 651534
rect 701342 651523 701376 651534
rect 701410 651523 701444 651534
rect 701478 651523 701512 651534
rect 701546 651523 701580 651534
rect 701614 651523 701648 651534
rect 701682 651523 701716 651534
rect 701750 651523 701784 651534
rect 701818 651523 701852 651534
rect 699392 651513 699450 651523
rect 699460 651513 699518 651523
rect 699528 651513 699586 651523
rect 699596 651513 699654 651523
rect 699664 651513 699722 651523
rect 699732 651513 699790 651523
rect 699800 651513 699858 651523
rect 699868 651513 699926 651523
rect 699936 651513 699994 651523
rect 700004 651513 700062 651523
rect 700072 651513 700130 651523
rect 700140 651513 700198 651523
rect 700208 651513 700266 651523
rect 700276 651513 700334 651523
rect 700934 651513 700992 651523
rect 701002 651513 701060 651523
rect 701070 651513 701128 651523
rect 701138 651513 701196 651523
rect 701206 651513 701264 651523
rect 701274 651513 701332 651523
rect 701342 651513 701400 651523
rect 701410 651513 701468 651523
rect 701478 651513 701536 651523
rect 701546 651513 701604 651523
rect 701614 651513 701672 651523
rect 701682 651513 701740 651523
rect 701750 651513 701808 651523
rect 701818 651513 701876 651523
rect 699368 651489 700334 651513
rect 700910 651489 701876 651513
rect 699392 651474 699416 651489
rect 699460 651474 699484 651489
rect 699528 651474 699552 651489
rect 699596 651474 699620 651489
rect 699664 651474 699688 651489
rect 699732 651474 699756 651489
rect 699800 651474 699824 651489
rect 699868 651474 699892 651489
rect 699936 651474 699960 651489
rect 700004 651474 700028 651489
rect 700072 651474 700096 651489
rect 700140 651474 700164 651489
rect 700208 651474 700232 651489
rect 700276 651474 700300 651489
rect 700934 651474 700958 651489
rect 701002 651474 701026 651489
rect 701070 651474 701094 651489
rect 701138 651474 701162 651489
rect 701206 651474 701230 651489
rect 701274 651474 701298 651489
rect 701342 651474 701366 651489
rect 701410 651474 701434 651489
rect 701478 651474 701502 651489
rect 701546 651474 701570 651489
rect 701614 651474 701638 651489
rect 701682 651474 701706 651489
rect 701750 651474 701774 651489
rect 701818 651474 701842 651489
rect 699322 651319 700322 651474
rect 699322 651285 700334 651319
rect 700922 651309 701922 651474
rect 707610 651319 708610 651379
rect 709211 651319 710211 651379
rect 700910 651285 701922 651309
rect 699322 651274 700322 651285
rect 700922 651274 701922 651285
rect 699392 651261 699416 651274
rect 699460 651261 699484 651274
rect 699528 651261 699552 651274
rect 699596 651261 699620 651274
rect 699664 651261 699688 651274
rect 699732 651261 699756 651274
rect 699800 651261 699824 651274
rect 699868 651261 699892 651274
rect 699936 651261 699960 651274
rect 700004 651261 700028 651274
rect 700072 651261 700096 651274
rect 700140 651261 700164 651274
rect 700208 651261 700232 651274
rect 700276 651261 700300 651274
rect 700934 651261 700958 651274
rect 701002 651261 701026 651274
rect 701070 651261 701094 651274
rect 701138 651261 701162 651274
rect 701206 651261 701230 651274
rect 701274 651261 701298 651274
rect 701342 651261 701366 651274
rect 701410 651261 701434 651274
rect 701478 651261 701502 651274
rect 701546 651261 701570 651274
rect 701614 651261 701638 651274
rect 701682 651261 701706 651274
rect 701750 651261 701774 651274
rect 701818 651261 701842 651274
rect 699322 650916 700322 650972
rect 700922 650916 701922 650972
rect 707610 650961 708610 651017
rect 709211 650961 710211 651017
rect 699322 650844 700322 650900
rect 700922 650844 701922 650900
rect 707610 650889 708610 650945
rect 709211 650889 710211 650945
rect 699322 650542 700322 650614
rect 700922 650542 701922 650614
rect 707610 650587 708610 650659
rect 709211 650587 710211 650659
rect 699392 650531 699426 650542
rect 699460 650531 699494 650542
rect 699528 650531 699562 650542
rect 699596 650531 699630 650542
rect 699664 650531 699698 650542
rect 699732 650531 699766 650542
rect 699800 650531 699834 650542
rect 699868 650531 699902 650542
rect 699936 650531 699970 650542
rect 700004 650531 700038 650542
rect 700072 650531 700106 650542
rect 700140 650531 700174 650542
rect 700208 650531 700242 650542
rect 700276 650531 700310 650542
rect 700934 650531 700968 650542
rect 701002 650531 701036 650542
rect 701070 650531 701104 650542
rect 701138 650531 701172 650542
rect 701206 650531 701240 650542
rect 701274 650531 701308 650542
rect 701342 650531 701376 650542
rect 701410 650531 701444 650542
rect 701478 650531 701512 650542
rect 701546 650531 701580 650542
rect 701614 650531 701648 650542
rect 701682 650531 701716 650542
rect 701750 650531 701784 650542
rect 701818 650531 701852 650542
rect 699392 650521 699450 650531
rect 699460 650521 699518 650531
rect 699528 650521 699586 650531
rect 699596 650521 699654 650531
rect 699664 650521 699722 650531
rect 699732 650521 699790 650531
rect 699800 650521 699858 650531
rect 699868 650521 699926 650531
rect 699936 650521 699994 650531
rect 700004 650521 700062 650531
rect 700072 650521 700130 650531
rect 700140 650521 700198 650531
rect 700208 650521 700266 650531
rect 700276 650521 700334 650531
rect 700934 650521 700992 650531
rect 701002 650521 701060 650531
rect 701070 650521 701128 650531
rect 701138 650521 701196 650531
rect 701206 650521 701264 650531
rect 701274 650521 701332 650531
rect 701342 650521 701400 650531
rect 701410 650521 701468 650531
rect 701478 650521 701536 650531
rect 701546 650521 701604 650531
rect 701614 650521 701672 650531
rect 701682 650521 701740 650531
rect 701750 650521 701808 650531
rect 701818 650521 701876 650531
rect 699368 650497 700334 650521
rect 700910 650497 701876 650521
rect 699392 650482 699416 650497
rect 699460 650482 699484 650497
rect 699528 650482 699552 650497
rect 699596 650482 699620 650497
rect 699664 650482 699688 650497
rect 699732 650482 699756 650497
rect 699800 650482 699824 650497
rect 699868 650482 699892 650497
rect 699936 650482 699960 650497
rect 700004 650482 700028 650497
rect 700072 650482 700096 650497
rect 700140 650482 700164 650497
rect 700208 650482 700232 650497
rect 700276 650482 700300 650497
rect 700934 650482 700958 650497
rect 701002 650482 701026 650497
rect 701070 650482 701094 650497
rect 701138 650482 701162 650497
rect 701206 650482 701230 650497
rect 701274 650482 701298 650497
rect 701342 650482 701366 650497
rect 701410 650482 701434 650497
rect 701478 650482 701502 650497
rect 701546 650482 701570 650497
rect 701614 650482 701638 650497
rect 701682 650482 701706 650497
rect 701750 650482 701774 650497
rect 701818 650482 701842 650497
rect 699322 650327 700322 650482
rect 699322 650293 700334 650327
rect 700922 650317 701922 650482
rect 707610 650327 708610 650387
rect 709211 650327 710211 650387
rect 711541 650345 711629 657461
rect 711892 656200 711942 657200
rect 712062 656200 712112 657200
rect 711892 655079 711942 656079
rect 712062 655079 712112 656079
rect 711892 653958 711942 654958
rect 712062 653958 712112 654958
rect 711892 652848 711942 653848
rect 712062 652848 712112 653848
rect 711892 651727 711942 652727
rect 712062 651727 712112 652727
rect 711892 650606 711942 651606
rect 712062 650606 712112 651606
rect 712409 650371 712431 657485
rect 712469 657459 712487 657501
rect 712499 657459 712505 657467
rect 712499 657455 712511 657459
rect 712539 657455 712557 657501
rect 713640 655461 713674 657785
rect 713750 657772 714750 657822
rect 717367 657820 717413 657853
rect 717367 657819 717379 657820
rect 717401 657819 717413 657820
rect 717401 657809 717600 657819
rect 717401 657786 717413 657809
rect 713750 657562 714750 657612
rect 713750 657446 714750 657496
rect 713750 657230 714750 657358
rect 713750 657014 714750 657070
rect 713750 656798 714750 656926
rect 713750 656588 714750 656638
rect 714478 656585 714750 656588
rect 715486 655931 715536 656931
rect 715696 655931 715824 656931
rect 715912 655931 715962 656931
rect 713641 655345 713663 655461
rect 713640 655309 713674 655345
rect 713750 655314 714750 655364
rect 713750 655158 714750 655214
rect 713750 655002 714750 655130
rect 713750 654846 714750 654974
rect 713750 654690 714750 654746
rect 716425 654709 716725 654721
rect 713750 654534 714750 654662
rect 716425 654596 717425 654646
rect 713750 654378 714750 654506
rect 716425 654440 717425 654568
rect 713750 654222 714750 654350
rect 716425 654284 717425 654340
rect 713750 654072 714750 654122
rect 713750 653956 714750 654006
rect 713750 653800 714750 653928
rect 713750 653644 714750 653772
rect 713750 653488 714750 653616
rect 715354 653587 715404 654187
rect 715504 653587 715560 654187
rect 715660 653587 715716 654187
rect 715816 653587 715872 654187
rect 715972 653587 716022 654187
rect 716425 654128 717425 654256
rect 716425 653978 717425 654028
rect 716425 653862 717425 653912
rect 716425 653706 717425 653834
rect 716425 653550 717425 653606
rect 716425 653394 717425 653522
rect 713750 653332 714750 653388
rect 713750 653176 714750 653304
rect 716425 653244 717425 653294
rect 713750 653020 714750 653148
rect 713750 652870 714750 652920
rect 713750 652742 714750 652792
rect 713750 652586 714750 652642
rect 713750 652436 714750 652486
rect 713750 652320 714350 652370
rect 713750 652164 714350 652292
rect 715510 652191 715560 653191
rect 715660 652191 715788 653191
rect 715816 652191 715944 653191
rect 715972 652191 716022 653191
rect 716425 653128 717425 653178
rect 716425 652972 717425 653028
rect 716425 652822 717425 652872
rect 716425 652706 717425 652756
rect 716425 652550 717425 652678
rect 716425 652394 717425 652522
rect 716425 652238 717425 652366
rect 716425 652082 717425 652210
rect 713750 652008 714350 652064
rect 713750 651852 714350 651980
rect 716425 651932 717425 651982
rect 713750 651696 714350 651752
rect 713750 651446 714350 651496
rect 714565 651443 714765 651455
rect 713750 651330 714750 651380
rect 713750 651120 714750 651170
rect 716413 651092 716447 651150
rect 713750 651004 714750 651054
rect 713750 650794 714750 650844
rect 713750 650678 714750 650728
rect 713750 650468 714750 650518
rect 713750 650352 714750 650402
rect 700910 650293 701922 650317
rect 699322 650282 700322 650293
rect 700922 650282 701922 650293
rect 711541 650311 711633 650345
rect 699392 650269 699416 650282
rect 699460 650269 699484 650282
rect 699528 650269 699552 650282
rect 699596 650269 699620 650282
rect 699664 650269 699688 650282
rect 699732 650269 699756 650282
rect 699800 650269 699824 650282
rect 699868 650269 699892 650282
rect 699936 650269 699960 650282
rect 700004 650269 700028 650282
rect 700072 650269 700096 650282
rect 700140 650269 700164 650282
rect 700208 650269 700232 650282
rect 700276 650269 700300 650282
rect 700934 650269 700958 650282
rect 701002 650269 701026 650282
rect 701070 650269 701094 650282
rect 701138 650269 701162 650282
rect 701206 650269 701230 650282
rect 701274 650269 701298 650282
rect 701342 650269 701366 650282
rect 701410 650269 701434 650282
rect 701478 650269 701502 650282
rect 701546 650269 701570 650282
rect 701614 650269 701638 650282
rect 701682 650269 701706 650282
rect 701750 650269 701774 650282
rect 701818 650269 701842 650282
rect 699322 649924 700322 649980
rect 700922 649924 701922 649980
rect 707610 649969 708610 650025
rect 709211 649969 710211 650025
rect 699322 649852 700322 649908
rect 700922 649852 701922 649908
rect 707610 649897 708610 649953
rect 709211 649897 710211 649953
rect 699322 649550 700322 649622
rect 700922 649550 701922 649622
rect 707610 649595 708610 649667
rect 709211 649595 710211 649667
rect 699392 649539 699426 649550
rect 699460 649539 699494 649550
rect 699528 649539 699562 649550
rect 699596 649539 699630 649550
rect 699664 649539 699698 649550
rect 699732 649539 699766 649550
rect 699800 649539 699834 649550
rect 699868 649539 699902 649550
rect 699936 649539 699970 649550
rect 700004 649539 700038 649550
rect 700072 649539 700106 649550
rect 700140 649539 700174 649550
rect 700208 649539 700242 649550
rect 700276 649539 700310 649550
rect 700934 649539 700968 649550
rect 701002 649539 701036 649550
rect 701070 649539 701104 649550
rect 701138 649539 701172 649550
rect 701206 649539 701240 649550
rect 701274 649539 701308 649550
rect 701342 649539 701376 649550
rect 701410 649539 701444 649550
rect 701478 649539 701512 649550
rect 701546 649539 701580 649550
rect 701614 649539 701648 649550
rect 701682 649539 701716 649550
rect 701750 649539 701784 649550
rect 701818 649539 701852 649550
rect 699392 649529 699450 649539
rect 699460 649529 699518 649539
rect 699528 649529 699586 649539
rect 699596 649529 699654 649539
rect 699664 649529 699722 649539
rect 699732 649529 699790 649539
rect 699800 649529 699858 649539
rect 699868 649529 699926 649539
rect 699936 649529 699994 649539
rect 700004 649529 700062 649539
rect 700072 649529 700130 649539
rect 700140 649529 700198 649539
rect 700208 649529 700266 649539
rect 700276 649529 700334 649539
rect 700934 649529 700992 649539
rect 701002 649529 701060 649539
rect 701070 649529 701128 649539
rect 701138 649529 701196 649539
rect 701206 649529 701264 649539
rect 701274 649529 701332 649539
rect 701342 649529 701400 649539
rect 701410 649529 701468 649539
rect 701478 649529 701536 649539
rect 701546 649529 701604 649539
rect 701614 649529 701672 649539
rect 701682 649529 701740 649539
rect 701750 649529 701808 649539
rect 701818 649529 701876 649539
rect 699368 649505 700334 649529
rect 700910 649505 701876 649529
rect 699392 649490 699416 649505
rect 699460 649490 699484 649505
rect 699528 649490 699552 649505
rect 699596 649490 699620 649505
rect 699664 649490 699688 649505
rect 699732 649490 699756 649505
rect 699800 649490 699824 649505
rect 699868 649490 699892 649505
rect 699936 649490 699960 649505
rect 700004 649490 700028 649505
rect 700072 649490 700096 649505
rect 700140 649490 700164 649505
rect 700208 649490 700232 649505
rect 700276 649490 700300 649505
rect 700934 649490 700958 649505
rect 701002 649490 701026 649505
rect 701070 649490 701094 649505
rect 701138 649490 701162 649505
rect 701206 649490 701230 649505
rect 701274 649490 701298 649505
rect 701342 649490 701366 649505
rect 701410 649490 701434 649505
rect 701478 649490 701502 649505
rect 701546 649490 701570 649505
rect 701614 649490 701638 649505
rect 701682 649490 701706 649505
rect 701750 649490 701774 649505
rect 701818 649490 701842 649505
rect 699322 649335 700322 649490
rect 699322 649301 700334 649335
rect 700922 649325 701922 649490
rect 707610 649335 708610 649395
rect 709211 649335 710211 649395
rect 700910 649301 701922 649325
rect 699322 649290 700322 649301
rect 700922 649290 701922 649301
rect 699392 649277 699416 649290
rect 699460 649277 699484 649290
rect 699528 649277 699552 649290
rect 699596 649277 699620 649290
rect 699664 649277 699688 649290
rect 699732 649277 699756 649290
rect 699800 649277 699824 649290
rect 699868 649277 699892 649290
rect 699936 649277 699960 649290
rect 700004 649277 700028 649290
rect 700072 649277 700096 649290
rect 700140 649277 700164 649290
rect 700208 649277 700232 649290
rect 700276 649277 700300 649290
rect 700934 649277 700958 649290
rect 701002 649277 701026 649290
rect 701070 649277 701094 649290
rect 701138 649277 701162 649290
rect 701206 649277 701230 649290
rect 701274 649277 701298 649290
rect 701342 649277 701366 649290
rect 701410 649277 701434 649290
rect 701478 649277 701502 649290
rect 701546 649277 701570 649290
rect 701614 649277 701638 649290
rect 701682 649277 701706 649290
rect 701750 649277 701774 649290
rect 701818 649277 701842 649290
rect 699322 648932 700322 648988
rect 700922 648932 701922 648988
rect 707610 648977 708610 649033
rect 709211 648977 710211 649033
rect 699322 648860 700322 648916
rect 700922 648860 701922 648916
rect 707610 648905 708610 648961
rect 709211 648905 710211 648961
rect 699322 648558 700322 648630
rect 700922 648558 701922 648630
rect 707610 648603 708610 648675
rect 709211 648603 710211 648675
rect 699392 648547 699426 648558
rect 699460 648547 699494 648558
rect 699528 648547 699562 648558
rect 699596 648547 699630 648558
rect 699664 648547 699698 648558
rect 699732 648547 699766 648558
rect 699800 648547 699834 648558
rect 699868 648547 699902 648558
rect 699936 648547 699970 648558
rect 700004 648547 700038 648558
rect 700072 648547 700106 648558
rect 700140 648547 700174 648558
rect 700208 648547 700242 648558
rect 700276 648547 700310 648558
rect 700934 648547 700968 648558
rect 701002 648547 701036 648558
rect 701070 648547 701104 648558
rect 701138 648547 701172 648558
rect 701206 648547 701240 648558
rect 701274 648547 701308 648558
rect 701342 648547 701376 648558
rect 701410 648547 701444 648558
rect 701478 648547 701512 648558
rect 701546 648547 701580 648558
rect 701614 648547 701648 648558
rect 701682 648547 701716 648558
rect 701750 648547 701784 648558
rect 701818 648547 701852 648558
rect 699392 648537 699450 648547
rect 699460 648537 699518 648547
rect 699528 648537 699586 648547
rect 699596 648537 699654 648547
rect 699664 648537 699722 648547
rect 699732 648537 699790 648547
rect 699800 648537 699858 648547
rect 699868 648537 699926 648547
rect 699936 648537 699994 648547
rect 700004 648537 700062 648547
rect 700072 648537 700130 648547
rect 700140 648537 700198 648547
rect 700208 648537 700266 648547
rect 700276 648537 700334 648547
rect 700934 648537 700992 648547
rect 701002 648537 701060 648547
rect 701070 648537 701128 648547
rect 701138 648537 701196 648547
rect 701206 648537 701264 648547
rect 701274 648537 701332 648547
rect 701342 648537 701400 648547
rect 701410 648537 701468 648547
rect 701478 648537 701536 648547
rect 701546 648537 701604 648547
rect 701614 648537 701672 648547
rect 701682 648537 701740 648547
rect 701750 648537 701808 648547
rect 701818 648537 701876 648547
rect 699368 648513 700334 648537
rect 700910 648513 701876 648537
rect 699392 648498 699416 648513
rect 699460 648498 699484 648513
rect 699528 648498 699552 648513
rect 699596 648498 699620 648513
rect 699664 648498 699688 648513
rect 699732 648498 699756 648513
rect 699800 648498 699824 648513
rect 699868 648498 699892 648513
rect 699936 648498 699960 648513
rect 700004 648498 700028 648513
rect 700072 648498 700096 648513
rect 700140 648498 700164 648513
rect 700208 648498 700232 648513
rect 700276 648498 700300 648513
rect 700934 648498 700958 648513
rect 701002 648498 701026 648513
rect 701070 648498 701094 648513
rect 701138 648498 701162 648513
rect 701206 648498 701230 648513
rect 701274 648498 701298 648513
rect 701342 648498 701366 648513
rect 701410 648498 701434 648513
rect 701478 648498 701502 648513
rect 701546 648498 701570 648513
rect 701614 648498 701638 648513
rect 701682 648498 701706 648513
rect 701750 648498 701774 648513
rect 701818 648498 701842 648513
rect 699322 648343 700322 648498
rect 699322 648309 700334 648343
rect 700922 648333 701922 648498
rect 707610 648343 708610 648403
rect 709211 648343 710211 648403
rect 700910 648309 701922 648333
rect 699322 648298 700322 648309
rect 700922 648298 701922 648309
rect 699392 648285 699416 648298
rect 699460 648285 699484 648298
rect 699528 648285 699552 648298
rect 699596 648285 699620 648298
rect 699664 648285 699688 648298
rect 699732 648285 699756 648298
rect 699800 648285 699824 648298
rect 699868 648285 699892 648298
rect 699936 648285 699960 648298
rect 700004 648285 700028 648298
rect 700072 648285 700096 648298
rect 700140 648285 700164 648298
rect 700208 648285 700232 648298
rect 700276 648285 700300 648298
rect 700934 648285 700958 648298
rect 701002 648285 701026 648298
rect 701070 648285 701094 648298
rect 701138 648285 701162 648298
rect 701206 648285 701230 648298
rect 701274 648285 701298 648298
rect 701342 648285 701366 648298
rect 701410 648285 701434 648298
rect 701478 648285 701502 648298
rect 701546 648285 701570 648298
rect 701614 648285 701638 648298
rect 701682 648285 701706 648298
rect 701750 648285 701774 648298
rect 701818 648285 701842 648298
rect 699322 647940 700322 647996
rect 700922 647940 701922 647996
rect 707610 647985 708610 648041
rect 709211 647985 710211 648041
rect 699322 647868 700322 647924
rect 700922 647868 701922 647924
rect 707610 647913 708610 647969
rect 709211 647913 710211 647969
rect 699322 647566 700322 647638
rect 700922 647566 701922 647638
rect 707610 647611 708610 647683
rect 709211 647611 710211 647683
rect 699392 647555 699426 647566
rect 699460 647555 699494 647566
rect 699528 647555 699562 647566
rect 699596 647555 699630 647566
rect 699664 647555 699698 647566
rect 699732 647555 699766 647566
rect 699800 647555 699834 647566
rect 699868 647555 699902 647566
rect 699936 647555 699970 647566
rect 700004 647555 700038 647566
rect 700072 647555 700106 647566
rect 700140 647555 700174 647566
rect 700208 647555 700242 647566
rect 700276 647555 700310 647566
rect 700934 647555 700968 647566
rect 701002 647555 701036 647566
rect 701070 647555 701104 647566
rect 701138 647555 701172 647566
rect 701206 647555 701240 647566
rect 701274 647555 701308 647566
rect 701342 647555 701376 647566
rect 701410 647555 701444 647566
rect 701478 647555 701512 647566
rect 701546 647555 701580 647566
rect 701614 647555 701648 647566
rect 701682 647555 701716 647566
rect 701750 647555 701784 647566
rect 701818 647555 701852 647566
rect 699392 647545 699450 647555
rect 699460 647545 699518 647555
rect 699528 647545 699586 647555
rect 699596 647545 699654 647555
rect 699664 647545 699722 647555
rect 699732 647545 699790 647555
rect 699800 647545 699858 647555
rect 699868 647545 699926 647555
rect 699936 647545 699994 647555
rect 700004 647545 700062 647555
rect 700072 647545 700130 647555
rect 700140 647545 700198 647555
rect 700208 647545 700266 647555
rect 700276 647545 700334 647555
rect 700934 647545 700992 647555
rect 701002 647545 701060 647555
rect 701070 647545 701128 647555
rect 701138 647545 701196 647555
rect 701206 647545 701264 647555
rect 701274 647545 701332 647555
rect 701342 647545 701400 647555
rect 701410 647545 701468 647555
rect 701478 647545 701536 647555
rect 701546 647545 701604 647555
rect 701614 647545 701672 647555
rect 701682 647545 701740 647555
rect 701750 647545 701808 647555
rect 701818 647545 701876 647555
rect 699368 647521 700334 647545
rect 700910 647521 701876 647545
rect 699392 647506 699416 647521
rect 699460 647506 699484 647521
rect 699528 647506 699552 647521
rect 699596 647506 699620 647521
rect 699664 647506 699688 647521
rect 699732 647506 699756 647521
rect 699800 647506 699824 647521
rect 699868 647506 699892 647521
rect 699936 647506 699960 647521
rect 700004 647506 700028 647521
rect 700072 647506 700096 647521
rect 700140 647506 700164 647521
rect 700208 647506 700232 647521
rect 700276 647506 700300 647521
rect 700934 647506 700958 647521
rect 701002 647506 701026 647521
rect 701070 647506 701094 647521
rect 701138 647506 701162 647521
rect 701206 647506 701230 647521
rect 701274 647506 701298 647521
rect 701342 647506 701366 647521
rect 701410 647506 701434 647521
rect 701478 647506 701502 647521
rect 701546 647506 701570 647521
rect 701614 647506 701638 647521
rect 701682 647506 701706 647521
rect 701750 647506 701774 647521
rect 701818 647506 701842 647521
rect 699322 647351 700322 647506
rect 699322 647317 700334 647351
rect 700922 647341 701922 647506
rect 705107 647360 705173 647376
rect 707610 647351 708610 647411
rect 709211 647351 710211 647411
rect 700910 647317 701922 647341
rect 699322 647306 700322 647317
rect 700922 647306 701922 647317
rect 699392 647293 699416 647306
rect 699460 647293 699484 647306
rect 699528 647293 699552 647306
rect 699596 647293 699620 647306
rect 699664 647293 699688 647306
rect 699732 647293 699756 647306
rect 699800 647293 699824 647306
rect 699868 647293 699892 647306
rect 699936 647293 699960 647306
rect 700004 647293 700028 647306
rect 700072 647293 700096 647306
rect 700140 647293 700164 647306
rect 700208 647293 700232 647306
rect 700276 647293 700300 647306
rect 700934 647293 700958 647306
rect 701002 647293 701026 647306
rect 701070 647293 701094 647306
rect 701138 647293 701162 647306
rect 701206 647293 701230 647306
rect 701274 647293 701298 647306
rect 701342 647293 701366 647306
rect 701410 647293 701434 647306
rect 701478 647293 701502 647306
rect 701546 647293 701570 647306
rect 701614 647293 701638 647306
rect 701682 647293 701706 647306
rect 701750 647293 701774 647306
rect 701818 647293 701842 647306
rect 699322 646948 700322 647004
rect 700922 646948 701922 647004
rect 707610 646993 708610 647049
rect 709211 646993 710211 647049
rect 699322 646876 700322 646932
rect 700922 646876 701922 646932
rect 707610 646921 708610 646977
rect 709211 646921 710211 646977
rect 699322 646574 700322 646646
rect 700922 646574 701922 646646
rect 707610 646619 708610 646691
rect 709211 646619 710211 646691
rect 699392 646563 699426 646574
rect 699460 646563 699494 646574
rect 699528 646563 699562 646574
rect 699596 646563 699630 646574
rect 699664 646563 699698 646574
rect 699732 646563 699766 646574
rect 699800 646563 699834 646574
rect 699868 646563 699902 646574
rect 699936 646563 699970 646574
rect 700004 646563 700038 646574
rect 700072 646563 700106 646574
rect 700140 646563 700174 646574
rect 700208 646563 700242 646574
rect 700276 646563 700310 646574
rect 700934 646563 700968 646574
rect 701002 646563 701036 646574
rect 701070 646563 701104 646574
rect 701138 646563 701172 646574
rect 701206 646563 701240 646574
rect 701274 646563 701308 646574
rect 701342 646563 701376 646574
rect 701410 646563 701444 646574
rect 701478 646563 701512 646574
rect 701546 646563 701580 646574
rect 701614 646563 701648 646574
rect 701682 646563 701716 646574
rect 701750 646563 701784 646574
rect 701818 646563 701852 646574
rect 699392 646553 699450 646563
rect 699460 646553 699518 646563
rect 699528 646553 699586 646563
rect 699596 646553 699654 646563
rect 699664 646553 699722 646563
rect 699732 646553 699790 646563
rect 699800 646553 699858 646563
rect 699868 646553 699926 646563
rect 699936 646553 699994 646563
rect 700004 646553 700062 646563
rect 700072 646553 700130 646563
rect 700140 646553 700198 646563
rect 700208 646553 700266 646563
rect 700276 646553 700334 646563
rect 700934 646553 700992 646563
rect 701002 646553 701060 646563
rect 701070 646553 701128 646563
rect 701138 646553 701196 646563
rect 701206 646553 701264 646563
rect 701274 646553 701332 646563
rect 701342 646553 701400 646563
rect 701410 646553 701468 646563
rect 701478 646553 701536 646563
rect 701546 646553 701604 646563
rect 701614 646553 701672 646563
rect 701682 646553 701740 646563
rect 701750 646553 701808 646563
rect 701818 646553 701876 646563
rect 699368 646529 700334 646553
rect 700910 646529 701876 646553
rect 699392 646514 699416 646529
rect 699460 646514 699484 646529
rect 699528 646514 699552 646529
rect 699596 646514 699620 646529
rect 699664 646514 699688 646529
rect 699732 646514 699756 646529
rect 699800 646514 699824 646529
rect 699868 646514 699892 646529
rect 699936 646514 699960 646529
rect 700004 646514 700028 646529
rect 700072 646514 700096 646529
rect 700140 646514 700164 646529
rect 700208 646514 700232 646529
rect 700276 646514 700300 646529
rect 700934 646514 700958 646529
rect 701002 646514 701026 646529
rect 701070 646514 701094 646529
rect 701138 646514 701162 646529
rect 701206 646514 701230 646529
rect 701274 646514 701298 646529
rect 701342 646514 701366 646529
rect 701410 646514 701434 646529
rect 701478 646514 701502 646529
rect 701546 646514 701570 646529
rect 701614 646514 701638 646529
rect 701682 646514 701706 646529
rect 701750 646514 701774 646529
rect 701818 646514 701842 646529
rect 699322 646359 700322 646514
rect 699322 646325 700334 646359
rect 700922 646349 701922 646514
rect 707610 646359 708610 646419
rect 709211 646359 710211 646419
rect 700910 646325 701922 646349
rect 699322 646314 700322 646325
rect 700922 646314 701922 646325
rect 699392 646301 699416 646314
rect 699460 646301 699484 646314
rect 699528 646301 699552 646314
rect 699596 646301 699620 646314
rect 699664 646301 699688 646314
rect 699732 646301 699756 646314
rect 699800 646301 699824 646314
rect 699868 646301 699892 646314
rect 699936 646301 699960 646314
rect 700004 646301 700028 646314
rect 700072 646301 700096 646314
rect 700140 646301 700164 646314
rect 700208 646301 700232 646314
rect 700276 646301 700300 646314
rect 700934 646301 700958 646314
rect 701002 646301 701026 646314
rect 701070 646301 701094 646314
rect 701138 646301 701162 646314
rect 701206 646301 701230 646314
rect 701274 646301 701298 646314
rect 701342 646301 701366 646314
rect 701410 646301 701434 646314
rect 701478 646301 701502 646314
rect 701546 646301 701570 646314
rect 701614 646301 701638 646314
rect 701682 646301 701706 646314
rect 701750 646301 701774 646314
rect 701818 646301 701842 646314
rect 709211 646148 710211 646152
rect 707574 646099 707610 646134
rect 708610 646099 708646 646134
rect 707574 646098 708646 646099
rect 707574 646057 707610 646098
rect 708610 646057 708646 646098
rect 699322 645956 700322 646012
rect 700922 645956 701922 646012
rect 707574 646001 708646 646057
rect 707574 645964 707610 646001
rect 708610 645964 708646 646001
rect 707574 645959 708646 645964
rect 699322 645884 700322 645940
rect 700922 645884 701922 645940
rect 707574 645924 707610 645959
rect 708610 645924 708646 645959
rect 709175 646098 710247 646134
rect 709175 646057 709211 646098
rect 710211 646057 710247 646098
rect 709175 646001 710247 646057
rect 709175 645964 709211 646001
rect 710211 645964 710247 646001
rect 709175 645936 710247 645964
rect 709175 645924 709211 645936
rect 710211 645924 710247 645936
rect 707610 645713 708610 645785
rect 709211 645713 710211 645785
rect 699322 645623 700322 645673
rect 700922 645623 701922 645673
rect 707610 645523 708610 645617
rect 707610 645513 708644 645523
rect 709211 645513 710211 645591
rect 711541 645437 711629 650311
rect 713750 650136 714750 650264
rect 716417 650152 717417 650202
rect 711892 649049 711942 650049
rect 712062 649049 712112 650049
rect 713750 649920 714750 650048
rect 716417 649996 717417 650052
rect 716417 649846 717417 649896
rect 713750 649704 714750 649832
rect 716417 649730 717017 649780
rect 716417 649580 717017 649630
rect 713750 649488 714750 649544
rect 716417 649464 717417 649514
rect 713750 649272 714750 649400
rect 716417 649308 717417 649364
rect 713750 649056 714750 649184
rect 716417 649152 717417 649280
rect 716417 648996 717417 649052
rect 711892 647928 711942 648928
rect 712062 647928 712112 648928
rect 713750 648840 714750 648968
rect 716417 648840 717417 648968
rect 713750 648624 714750 648752
rect 716417 648684 717417 648740
rect 716417 648474 717417 648524
rect 713750 648408 714750 648464
rect 716417 648308 717417 648358
rect 713750 648192 714750 648248
rect 716417 648152 717417 648280
rect 713750 647976 714750 648104
rect 716417 647996 717417 648052
rect 711892 646807 711942 647807
rect 712062 646807 712112 647807
rect 713750 647760 714750 647888
rect 716417 647780 717417 647836
rect 713750 647544 714750 647672
rect 716417 647570 717417 647620
rect 713750 647328 714750 647456
rect 716417 647454 717417 647504
rect 716417 647298 717417 647426
rect 713750 647118 714750 647168
rect 716417 647148 717417 647198
rect 711892 645697 711942 646697
rect 712062 645697 712112 646697
rect 714686 646357 714794 646424
rect 714645 646323 714794 646357
rect 716071 646357 716074 646358
rect 716071 646356 716072 646357
rect 716073 646356 716074 646357
rect 716071 646355 716074 646356
rect 716208 646357 716211 646358
rect 716208 646356 716209 646357
rect 716210 646356 716211 646357
rect 716208 646355 716211 646356
rect 714964 646247 715998 646329
rect 716284 646247 717318 646329
rect 705107 645336 705173 645352
rect 711541 645302 711633 645437
rect 714175 645398 714225 645998
rect 714425 645398 714475 645998
rect 711579 645301 711595 645302
rect 714781 645191 714863 646226
rect 715134 645955 715828 646037
rect 714686 645123 714863 645191
rect 714645 645089 714863 645123
rect 680215 644880 680815 644936
rect 686719 644893 686739 644917
rect 686743 644893 686753 644917
rect 686719 644859 686757 644893
rect 686719 644822 686739 644859
rect 686743 644822 686753 644859
rect 692428 644850 693028 644978
rect 698017 644947 698210 644983
rect 698084 644935 698210 644947
rect 702756 644959 703645 644983
rect 702756 644935 702853 644959
rect 698084 644828 702853 644935
rect 686719 644788 686757 644822
rect 680215 644704 680815 644760
rect 686719 644751 686739 644788
rect 686743 644751 686753 644788
rect 686719 644741 686757 644751
rect 686699 644717 686767 644741
rect 686719 644704 686739 644717
rect 686743 644704 686753 644717
rect 686719 644695 686753 644704
rect 686719 644693 686743 644695
rect 692428 644694 693028 644750
rect 686685 644656 686709 644680
rect 686743 644656 686767 644680
rect 678799 644503 679399 644553
rect 680215 644534 680815 644584
rect 692428 644538 693028 644666
rect 680593 644531 680815 644534
rect 682009 644501 682069 644516
rect 682024 644465 682054 644501
rect 683708 644387 684308 644437
rect 678799 644327 679399 644383
rect 692428 644382 693028 644510
rect 714781 644308 714863 645089
rect 715063 644609 715145 645915
rect 715342 645752 715382 645792
rect 715582 645752 715622 645792
rect 715289 644777 715339 645719
rect 715382 645668 715422 645752
rect 715542 645668 715582 645752
rect 715633 644777 715683 645719
rect 715382 644672 715422 644756
rect 715542 644672 715582 644756
rect 715342 644632 715382 644672
rect 715582 644632 715622 644672
rect 715815 644609 715897 645915
rect 715134 644387 715828 644469
rect 716100 644308 716182 646226
rect 716454 645955 717148 646037
rect 716385 644609 716467 645915
rect 716660 645752 716700 645792
rect 716900 645752 716940 645792
rect 716599 644777 716649 645719
rect 716700 645668 716740 645752
rect 716860 645668 716900 645752
rect 716943 644777 716993 645719
rect 716700 644672 716740 644756
rect 716860 644672 716900 644756
rect 716660 644632 716700 644672
rect 716900 644632 716940 644672
rect 717137 644609 717219 645915
rect 716454 644387 717148 644469
rect 717419 644308 717501 646226
rect 683708 644237 684308 644287
rect 692428 644232 693028 644282
rect 678799 644157 679399 644207
rect 684565 644160 684790 644168
rect 696597 644000 696600 644120
rect 714964 644095 715998 644177
rect 716284 644095 717318 644177
rect 21000 617000 21003 617120
rect 282 616623 1316 616705
rect 1602 616623 2636 616705
rect 32810 616662 33035 616670
rect 38201 616593 38801 616643
rect 24572 616518 25172 616568
rect 33292 616513 33892 616563
rect 99 614574 181 616492
rect 452 616331 1146 616413
rect 381 614885 463 616191
rect 660 616128 700 616168
rect 900 616128 940 616168
rect 700 616044 740 616128
rect 860 616044 900 616128
rect 607 615081 657 616023
rect 951 615081 1001 616023
rect 1133 614885 1215 616191
rect 452 614763 1146 614845
rect 1418 614574 1500 616492
rect 1772 616331 2466 616413
rect 1703 614885 1785 616191
rect 1978 616128 2018 616168
rect 2218 616128 2258 616168
rect 2018 616044 2058 616128
rect 2178 616044 2218 616128
rect 1917 615081 1967 616023
rect 2261 615081 2311 616023
rect 2455 614885 2537 616191
rect 2737 615779 2819 616492
rect 24572 616362 25172 616490
rect 38201 616417 38801 616473
rect 33292 616363 33892 616413
rect 24572 616206 25172 616334
rect 35546 616299 35576 616335
rect 36785 616329 36935 616341
rect 35531 616284 35591 616299
rect 36785 616216 37385 616266
rect 38201 616247 38801 616297
rect 30833 616120 30857 616144
rect 30891 616120 30915 616144
rect 24572 616050 25172 616106
rect 30857 616105 30881 616107
rect 30857 616096 30887 616105
rect 30867 616083 30887 616096
rect 30891 616083 30907 616120
rect 30833 616059 30857 616083
rect 30867 616049 30911 616083
rect 14747 615865 19516 615972
rect 24572 615894 25172 616022
rect 30867 616012 30887 616049
rect 30891 616012 30907 616049
rect 36785 616040 37385 616096
rect 30867 615978 30911 616012
rect 30867 615941 30887 615978
rect 30891 615941 30907 615978
rect 30867 615907 30911 615941
rect 30867 615883 30887 615907
rect 30891 615883 30907 615907
rect 14747 615841 14844 615865
rect 13955 615817 14844 615841
rect 19390 615853 19516 615865
rect 19390 615841 19583 615853
rect 19390 615817 19605 615841
rect 19639 615817 19673 615841
rect 19707 615817 19741 615841
rect 19775 615817 19809 615841
rect 19843 615817 19877 615841
rect 19911 615817 19945 615841
rect 19979 615817 20013 615841
rect 20047 615817 20081 615841
rect 20115 615817 20149 615841
rect 20183 615817 20217 615841
rect 20251 615817 20285 615841
rect 20319 615817 20353 615841
rect 20387 615817 20421 615841
rect 20455 615817 20489 615841
rect 20523 615817 20557 615841
rect 20591 615817 20625 615841
rect 20659 615817 20693 615841
rect 2737 615711 2914 615779
rect 1772 614763 2466 614845
rect 2737 614574 2819 615711
rect 2848 615677 2955 615711
rect 19480 615540 19516 615817
rect 19547 615540 19583 615817
rect 24572 615738 25172 615866
rect 36785 615864 37385 615920
rect 36785 615688 37385 615744
rect 20809 615650 20833 615684
rect 20809 615582 20833 615616
rect 24572 615588 25172 615638
rect 20809 615540 20833 615548
rect 36785 615518 37385 615568
rect 3125 614802 3175 615402
rect 3375 614802 3425 615402
rect 282 614471 1316 614553
rect 1602 614471 2636 614553
rect 1389 614444 1392 614445
rect 1389 614443 1390 614444
rect 1391 614443 1392 614444
rect 1389 614442 1392 614443
rect 1526 614444 1529 614445
rect 1526 614443 1527 614444
rect 1528 614443 1529 614444
rect 2848 614443 2955 614477
rect 1526 614442 1529 614443
rect 5488 614280 5538 615103
rect 5658 614280 5708 615103
rect 6005 614280 6021 615499
rect 12427 615448 12493 615464
rect 24572 615458 25172 615508
rect 32930 615457 33530 615507
rect 35287 615391 35887 615441
rect 36785 615402 37385 615452
rect 24572 615308 25172 615358
rect 31463 615307 32063 615357
rect 32930 615301 33530 615357
rect 7389 615277 7406 615287
rect 7440 615277 7477 615287
rect 7511 615277 7551 615287
rect 7585 615277 7622 615287
rect 7656 615277 7696 615287
rect 7730 615277 7767 615287
rect 7801 615277 7841 615287
rect 7875 615277 7912 615287
rect 7946 615277 7986 615287
rect 8020 615277 8057 615287
rect 8091 615277 8131 615287
rect 8165 615277 8202 615287
rect 8236 615277 8296 615287
rect 8330 615277 8381 615287
rect 8996 615277 9044 615287
rect 9078 615277 9120 615287
rect 9154 615277 9197 615287
rect 9231 615277 9291 615287
rect 9325 615277 9362 615287
rect 9396 615277 9436 615287
rect 9470 615277 9507 615287
rect 9541 615277 9581 615287
rect 9615 615277 9652 615287
rect 9686 615277 9726 615287
rect 9760 615277 9797 615287
rect 9831 615277 9871 615287
rect 9905 615277 9942 615287
rect 9976 615277 9990 615287
rect 7389 615209 8389 615277
rect 8990 615183 9990 615277
rect 36785 615226 37385 615282
rect 15678 615127 16678 615177
rect 17278 615127 18278 615177
rect 31463 615151 32063 615207
rect 32930 615151 33530 615201
rect 34079 615157 34679 615207
rect 7389 614840 8389 614864
rect 15678 614860 16678 614916
rect 17278 614860 18278 614916
rect 8990 614840 9990 614841
rect 7389 614743 8389 614799
rect 8990 614743 9990 614799
rect 15678 614788 16678 614844
rect 17278 614788 18278 614844
rect 8990 614701 9990 614702
rect 15678 614286 16678 614426
rect 17278 614286 18278 614426
rect 19844 614280 19894 615051
rect 20462 614280 20512 615051
rect 31463 615001 32063 615051
rect 34079 615001 34679 615057
rect 35287 615039 35887 615095
rect 36785 615050 37385 615106
rect 32596 614929 33596 614979
rect 24573 614820 25173 614870
rect 34079 614851 34679 614901
rect 35287 614869 35887 614919
rect 36785 614880 37385 614930
rect 30171 614795 30771 614845
rect 32596 614773 33596 614829
rect 37993 614704 38593 614754
rect 30171 614619 30771 614675
rect 32596 614623 33596 614673
rect 34110 614589 34710 614639
rect 21263 614280 21313 614518
rect 22349 614280 22399 614518
rect 32596 614507 33596 614557
rect 30171 614449 30771 614499
rect 36785 614429 36985 614609
rect 37993 614534 38593 614584
rect 24573 614352 25173 614408
rect 29993 614310 30993 614360
rect 31347 614280 31547 614317
rect 31607 614280 31807 614317
rect 36785 614280 36985 614373
rect 37083 614280 37120 614373
rect 696597 612200 696600 612320
rect 692376 611983 692396 612017
rect 692463 611993 692532 612017
rect 696191 611993 696239 612017
rect 692487 611983 692532 611993
rect 696204 611983 696239 611993
rect 696340 611983 696360 612017
rect 692487 611915 692502 611939
rect 696200 611915 696215 611939
rect 692454 611891 692478 611915
rect 696224 611891 696248 611915
rect 686755 611800 687355 611850
rect 692487 611748 692505 611752
rect 692479 611718 692505 611748
rect 692487 611698 692505 611718
rect 686755 611624 687355 611680
rect 692485 611674 692505 611698
rect 692509 611674 692517 611718
rect 696215 611698 696223 611748
rect 696203 611674 696223 611698
rect 696227 611674 696245 611752
rect 692485 611640 692521 611674
rect 696203 611640 696249 611674
rect 686755 611448 687355 611504
rect 686755 611278 687355 611328
rect 685547 611102 686147 611152
rect 687155 611007 687170 611022
rect 687343 611018 687355 611022
rect 687340 611007 687355 611018
rect 685547 610932 686147 610982
rect 687155 610827 687355 611007
rect 687155 610812 687170 610827
rect 687340 610816 687355 610827
rect 687343 610812 687355 610816
rect 687042 610771 687057 610786
rect 687020 610591 687057 610771
rect 687155 610771 687170 610786
rect 687343 610782 687355 610786
rect 687340 610771 687355 610782
rect 687155 610591 687355 610771
rect 688210 610630 688260 611630
rect 688360 610740 688488 611630
rect 688516 610740 688644 611630
rect 688672 610740 688800 611630
rect 688828 610740 688956 611630
rect 688984 610740 689112 611630
rect 689140 610740 689268 611630
rect 689296 610740 689424 611630
rect 689452 610740 689580 611630
rect 689608 610740 689736 611630
rect 689764 610740 689892 611630
rect 689920 610740 690048 611630
rect 690076 610740 690204 611630
rect 690232 610740 690360 611630
rect 690388 610630 690438 611630
rect 692485 611606 692505 611640
rect 692509 611606 692517 611640
rect 696203 611606 696223 611640
rect 696227 611606 696245 611640
rect 691275 611523 691875 611573
rect 692485 611572 692521 611606
rect 696203 611572 696249 611606
rect 692485 611538 692505 611572
rect 692509 611538 692517 611572
rect 692485 611504 692521 611538
rect 692583 611528 693983 611571
rect 694719 611528 696119 611571
rect 696203 611538 696223 611572
rect 696227 611538 696245 611572
rect 696203 611504 696249 611538
rect 692485 611470 692505 611504
rect 692509 611470 692517 611504
rect 692485 611436 692521 611470
rect 691275 611373 691875 611423
rect 692485 611402 692505 611436
rect 692509 611402 692517 611436
rect 692485 611368 692521 611402
rect 692485 611334 692505 611368
rect 692509 611334 692517 611368
rect 692583 611365 693983 611493
rect 694719 611365 696119 611493
rect 696203 611470 696223 611504
rect 696227 611470 696245 611504
rect 696203 611436 696249 611470
rect 707624 611441 707658 611475
rect 707695 611441 707729 611475
rect 707769 611441 707803 611475
rect 707840 611441 707874 611475
rect 707914 611441 707948 611475
rect 707985 611441 708019 611475
rect 708059 611441 708093 611475
rect 708130 611441 708164 611475
rect 708204 611441 708238 611475
rect 708275 611441 708309 611475
rect 708369 611441 708403 611475
rect 708446 611441 708480 611475
rect 708520 611441 708554 611465
rect 708588 611441 708610 611465
rect 709211 611441 709234 611465
rect 709270 611441 709304 611475
rect 709364 611441 709398 611475
rect 709435 611441 709469 611475
rect 709509 611441 709543 611475
rect 709580 611441 709614 611475
rect 709654 611441 709688 611475
rect 709725 611441 709759 611475
rect 709799 611441 709833 611475
rect 709870 611441 709904 611475
rect 709944 611441 709978 611475
rect 710015 611441 710049 611475
rect 710089 611441 710123 611475
rect 710160 611441 710194 611475
rect 696203 611402 696223 611436
rect 696227 611402 696245 611436
rect 707610 611431 707624 611441
rect 707658 611431 707695 611441
rect 707729 611431 707769 611441
rect 707803 611431 707840 611441
rect 707874 611431 707914 611441
rect 707948 611431 707985 611441
rect 708019 611431 708059 611441
rect 708093 611431 708130 611441
rect 708164 611431 708204 611441
rect 708238 611431 708275 611441
rect 708309 611431 708369 611441
rect 708403 611431 708446 611441
rect 708480 611431 708520 611441
rect 708554 611431 708588 611441
rect 708610 611431 708634 611441
rect 709211 611431 709270 611441
rect 709304 611431 709364 611441
rect 709398 611431 709435 611441
rect 709469 611431 709509 611441
rect 709543 611431 709580 611441
rect 709614 611431 709654 611441
rect 709688 611431 709725 611441
rect 709759 611431 709799 611441
rect 709833 611431 709870 611441
rect 709904 611431 709944 611441
rect 709978 611431 710015 611441
rect 710049 611431 710089 611441
rect 710123 611431 710160 611441
rect 710194 611431 710211 611441
rect 696203 611368 696249 611402
rect 696203 611334 696223 611368
rect 696227 611334 696245 611368
rect 707610 611337 708610 611431
rect 709211 611337 710211 611431
rect 691275 611251 691875 611301
rect 692485 611300 692521 611334
rect 692485 611266 692505 611300
rect 692509 611266 692517 611300
rect 692485 611232 692521 611266
rect 692485 611198 692505 611232
rect 692509 611198 692517 611232
rect 692583 611202 693983 611330
rect 694719 611202 696119 611330
rect 696203 611300 696249 611334
rect 711579 611317 712463 611331
rect 711579 611307 711619 611317
rect 696203 611266 696223 611300
rect 696227 611266 696245 611300
rect 701730 611290 701747 611292
rect 696203 611232 696249 611266
rect 696203 611198 696223 611232
rect 696227 611198 696245 611232
rect 701692 611220 701722 611254
rect 701730 611220 701760 611290
rect 707610 611241 708610 611301
rect 709211 611241 710211 611301
rect 692485 611164 692521 611198
rect 691275 611101 691875 611151
rect 692485 611130 692505 611164
rect 692509 611130 692517 611164
rect 692485 611096 692521 611130
rect 692485 611062 692505 611096
rect 692509 611062 692517 611096
rect 692485 611028 692521 611062
rect 692583 611039 693983 611167
rect 694719 611039 696119 611167
rect 696203 611164 696249 611198
rect 696203 611130 696223 611164
rect 696227 611130 696245 611164
rect 696203 611096 696249 611130
rect 696203 611062 696223 611096
rect 696227 611062 696245 611096
rect 699322 611064 700322 611097
rect 700922 611064 701922 611097
rect 696203 611028 696249 611062
rect 707610 611044 708610 611048
rect 709211 611044 710211 611048
rect 691275 610975 691875 611025
rect 692485 610994 692505 611028
rect 692509 610994 692517 611028
rect 692485 610960 692521 610994
rect 692485 610926 692505 610960
rect 692509 610926 692517 610960
rect 692485 610892 692521 610926
rect 691275 610825 691875 610875
rect 692485 610858 692505 610892
rect 692509 610858 692517 610892
rect 692583 610876 693983 611004
rect 694719 610876 696119 611004
rect 696203 610994 696223 611028
rect 696227 610994 696245 611028
rect 707574 610994 708646 611030
rect 696203 610960 696249 610994
rect 696203 610926 696223 610960
rect 696227 610926 696245 610960
rect 707574 610953 707610 610994
rect 708610 610953 708646 610994
rect 696203 610892 696249 610926
rect 697284 610894 697350 610910
rect 707574 610897 708646 610953
rect 696203 610858 696223 610892
rect 696227 610858 696245 610892
rect 699322 610877 700322 610894
rect 700922 610877 701922 610894
rect 707574 610881 707610 610897
rect 708610 610881 708646 610897
rect 692485 610824 692521 610858
rect 692485 610790 692505 610824
rect 692509 610790 692517 610824
rect 692485 610756 692521 610790
rect 691275 610703 691875 610753
rect 692485 610740 692505 610756
rect 692509 610740 692517 610756
rect 692583 610740 693983 610841
rect 694719 610740 696119 610841
rect 696203 610824 696249 610858
rect 707574 610825 708646 610881
rect 696203 610790 696223 610824
rect 696227 610790 696245 610824
rect 696203 610756 696249 610790
rect 696203 610740 696223 610756
rect 696227 610740 696245 610756
rect 699322 610740 700322 610811
rect 700922 610740 701922 610811
rect 707574 610788 707610 610825
rect 708610 610788 708646 610825
rect 707574 610748 708646 610788
rect 709175 610994 710247 611030
rect 709175 610953 709211 610994
rect 710211 610953 710247 610994
rect 709175 610897 710247 610953
rect 709175 610881 709211 610897
rect 710211 610881 710247 610897
rect 709175 610825 710247 610881
rect 709175 610788 709211 610825
rect 710211 610788 710247 610825
rect 709175 610748 710247 610788
rect 685542 610506 686142 610556
rect 691275 610553 691875 610603
rect 685542 610330 686142 610386
rect 692583 610237 693983 610280
rect 694719 610237 696119 610280
rect 699322 610278 700322 610418
rect 700922 610278 701922 610418
rect 685542 610160 686142 610210
rect 692583 610101 693983 610144
rect 694719 610101 696119 610144
rect 680215 609678 680815 609728
rect 680215 609502 680815 609558
rect 685551 609516 686551 609566
rect 689154 609480 689204 609897
rect 689304 609480 689360 609897
rect 689460 609480 689516 609897
rect 689616 609480 689672 609897
rect 689772 609480 689828 609897
rect 689928 609480 689978 609897
rect 699322 609860 700322 609916
rect 700922 609860 701922 609916
rect 707610 609905 708610 609961
rect 709211 609905 710211 609961
rect 699322 609788 700322 609844
rect 700922 609788 701922 609844
rect 707610 609833 708610 609889
rect 709211 609833 710211 609889
rect 711579 609525 711605 611307
rect 715956 610297 716006 611297
rect 716106 610740 716234 611297
rect 716262 610297 716312 611297
rect 711579 609480 711595 609495
rect 712409 609480 712431 609485
rect 713640 609480 713641 609785
rect 713750 609772 714750 609822
rect 713750 609562 714750 609612
rect 713750 609480 714750 609496
rect 2850 603304 3850 603320
rect 2850 603188 3850 603238
rect 2850 602978 3850 603028
rect 3959 603015 3960 603320
rect 5169 603315 5191 603320
rect 6005 603305 6021 603320
rect 1288 601503 1338 602503
rect 1438 601503 1566 602060
rect 1594 601503 1644 602503
rect 5995 601493 6021 603275
rect 7389 602911 8389 602967
rect 8990 602911 9990 602967
rect 15678 602956 16678 603012
rect 17278 602956 18278 603012
rect 7389 602839 8389 602895
rect 8990 602839 9990 602895
rect 15678 602884 16678 602940
rect 17278 602884 18278 602940
rect 27622 602903 27672 603320
rect 27772 602903 27828 603320
rect 27928 602903 27984 603320
rect 28084 602903 28140 603320
rect 28240 602903 28296 603320
rect 28396 602903 28446 603320
rect 31049 603234 32049 603284
rect 36785 603242 37385 603298
rect 36785 603072 37385 603122
rect 21481 602656 22881 602699
rect 23617 602656 25017 602699
rect 31458 602590 32058 602640
rect 15678 602382 16678 602522
rect 17278 602382 18278 602522
rect 21481 602520 22881 602563
rect 23617 602520 25017 602563
rect 31458 602414 32058 602470
rect 25725 602197 26325 602247
rect 31458 602244 32058 602294
rect 7353 602016 8425 602052
rect 7353 601975 7389 602016
rect 8389 601975 8425 602016
rect 7353 601919 8425 601975
rect 7353 601903 7389 601919
rect 8389 601903 8425 601919
rect 7353 601847 8425 601903
rect 7353 601810 7389 601847
rect 8389 601810 8425 601847
rect 7353 601770 8425 601810
rect 8954 602016 10026 602052
rect 8954 601975 8990 602016
rect 9990 601975 10026 602016
rect 8954 601919 10026 601975
rect 21383 602044 21403 602060
rect 21407 602044 21415 602060
rect 21383 602010 21419 602044
rect 21481 602031 22881 602060
rect 23617 602031 25017 602060
rect 25101 602044 25121 602060
rect 25125 602044 25143 602060
rect 25725 602047 26325 602097
rect 25101 602010 25147 602044
rect 21383 601976 21403 602010
rect 21407 601976 21415 602010
rect 21383 601942 21419 601976
rect 8954 601903 8990 601919
rect 9990 601903 10026 601919
rect 15678 601906 16678 601923
rect 17278 601906 18278 601923
rect 21383 601908 21403 601942
rect 21407 601908 21415 601942
rect 8954 601847 10026 601903
rect 20250 601890 20316 601906
rect 8954 601810 8990 601847
rect 9990 601810 10026 601847
rect 8954 601770 10026 601810
rect 21383 601874 21419 601908
rect 21383 601840 21403 601874
rect 21407 601840 21415 601874
rect 21481 601868 22881 601996
rect 23617 601868 25017 601996
rect 25101 601976 25121 602010
rect 25125 601976 25143 602010
rect 25101 601942 25147 601976
rect 25101 601908 25121 601942
rect 25125 601908 25143 601942
rect 25725 601925 26325 601975
rect 25101 601874 25147 601908
rect 25101 601840 25121 601874
rect 25125 601840 25143 601874
rect 21383 601806 21419 601840
rect 21383 601772 21403 601806
rect 21407 601772 21415 601806
rect 21383 601738 21419 601772
rect 15678 601703 16678 601736
rect 17278 601703 18278 601736
rect 21383 601704 21403 601738
rect 21407 601704 21415 601738
rect 21481 601705 22881 601833
rect 23617 601705 25017 601833
rect 25101 601806 25147 601840
rect 25101 601772 25121 601806
rect 25125 601772 25143 601806
rect 25725 601775 26325 601825
rect 25101 601738 25147 601772
rect 25101 601704 25121 601738
rect 25125 601704 25143 601738
rect 21383 601670 21419 601704
rect 25101 601670 25147 601704
rect 21383 601636 21403 601670
rect 21407 601636 21415 601670
rect 7389 601559 8389 601631
rect 8990 601559 9990 601631
rect 21383 601602 21419 601636
rect 15840 601510 15870 601580
rect 15878 601546 15908 601580
rect 21383 601568 21403 601602
rect 21407 601568 21415 601602
rect 15853 601508 15870 601510
rect 21383 601534 21419 601568
rect 21481 601542 22881 601670
rect 23617 601542 25017 601670
rect 25101 601636 25121 601670
rect 25125 601636 25143 601670
rect 25725 601649 26325 601699
rect 25101 601602 25147 601636
rect 25101 601568 25121 601602
rect 25125 601568 25143 601602
rect 25101 601534 25147 601568
rect 5981 601483 6021 601493
rect 5137 601469 6021 601483
rect 21383 601500 21403 601534
rect 21407 601500 21415 601534
rect 21383 601466 21419 601500
rect 7389 601369 8389 601463
rect 7389 601359 8413 601369
rect 8990 601359 9990 601463
rect 21383 601432 21403 601466
rect 21407 601432 21415 601466
rect 21383 601398 21419 601432
rect 21383 601364 21403 601398
rect 21407 601364 21415 601398
rect 21481 601379 22881 601507
rect 23617 601379 25017 601507
rect 25101 601500 25121 601534
rect 25125 601500 25143 601534
rect 25101 601466 25147 601500
rect 25725 601499 26325 601549
rect 25101 601432 25121 601466
rect 25125 601432 25143 601466
rect 25101 601398 25147 601432
rect 25101 601364 25121 601398
rect 25125 601364 25143 601398
rect 25725 601377 26325 601427
rect 21383 601330 21419 601364
rect 25101 601330 25147 601364
rect 21383 601296 21403 601330
rect 21407 601296 21415 601330
rect 25101 601296 25121 601330
rect 25125 601296 25143 601330
rect 21383 601262 21419 601296
rect 21383 601228 21403 601262
rect 21407 601228 21415 601262
rect 21481 601229 22881 601272
rect 23617 601229 25017 601272
rect 25101 601262 25147 601296
rect 25101 601228 25121 601262
rect 25125 601228 25143 601262
rect 21383 601194 21419 601228
rect 25101 601194 25147 601228
rect 25725 601227 26325 601277
rect 21383 601160 21403 601194
rect 21407 601160 21415 601194
rect 25101 601160 25121 601194
rect 25125 601160 25143 601194
rect 27162 601170 27212 602170
rect 27312 601170 27440 602060
rect 27468 601170 27596 602060
rect 27624 601170 27752 602060
rect 27780 601170 27908 602060
rect 27936 601170 28064 602060
rect 28092 601170 28220 602060
rect 28248 601170 28376 602060
rect 28404 601170 28532 602060
rect 28560 601170 28688 602060
rect 28716 601170 28844 602060
rect 28872 601170 29000 602060
rect 29028 601170 29156 602060
rect 29184 601170 29312 602060
rect 29340 601170 29390 602170
rect 30245 602029 30445 602209
rect 30245 602018 30260 602029
rect 30245 602014 30257 602018
rect 30430 602014 30445 602029
rect 30543 602029 30580 602209
rect 30543 602014 30558 602029
rect 30245 601984 30257 601988
rect 30245 601973 30260 601984
rect 30430 601973 30445 601988
rect 30245 601793 30445 601973
rect 31453 601818 32053 601868
rect 30245 601782 30260 601793
rect 30245 601778 30257 601782
rect 30430 601778 30445 601793
rect 31453 601648 32053 601698
rect 30245 601472 30845 601522
rect 30245 601296 30845 601352
rect 21383 601126 21419 601160
rect 25101 601126 25147 601160
rect 21383 601102 21403 601126
rect 21385 601048 21403 601102
rect 21407 601082 21415 601126
rect 25101 601102 25121 601126
rect 25113 601082 25121 601102
rect 25125 601048 25143 601126
rect 30245 601120 30845 601176
rect 30245 600950 30845 601000
rect 21000 600800 21003 600920
rect 21352 600885 21376 600909
rect 25122 600885 25146 600909
rect 21385 600861 21400 600885
rect 25098 600861 25113 600885
rect 21274 600783 21294 600851
rect 21410 600817 21430 600851
rect 25068 600817 25088 600851
rect 25204 600817 25224 600851
rect 21385 600807 21430 600817
rect 25102 600807 25137 600817
rect 21361 600783 21430 600807
rect 25089 600783 25137 600807
rect 25238 600783 25258 600817
rect 680480 598427 680517 598520
rect 680615 598427 680815 598520
rect 685793 598483 685993 598520
rect 686053 598483 686253 598520
rect 686607 598440 687607 598490
rect 692427 598392 693027 598448
rect 679007 598216 679607 598266
rect 680615 598191 680815 598371
rect 686829 598301 687429 598351
rect 684004 598243 685004 598293
rect 695201 598282 695251 598520
rect 696287 598282 696337 598520
rect 682890 598161 683490 598211
rect 684004 598127 685004 598177
rect 686829 598125 687429 598181
rect 679007 598046 679607 598096
rect 684004 597971 685004 598027
rect 686829 597955 687429 598005
rect 680215 597870 680815 597920
rect 681713 597881 682313 597931
rect 682921 597899 683521 597949
rect 692427 597930 693027 597980
rect 684004 597821 685004 597871
rect 680215 597694 680815 597750
rect 681713 597705 682313 597761
rect 682921 597743 683521 597799
rect 685537 597749 686137 597799
rect 697088 597749 697138 598520
rect 697706 597749 697756 598520
rect 699322 598374 700322 598514
rect 700922 598374 701922 598514
rect 707610 598098 708610 598099
rect 699322 597956 700322 598012
rect 700922 597956 701922 598012
rect 707610 598001 708610 598057
rect 709211 598001 710211 598057
rect 707610 597959 708610 597960
rect 699322 597884 700322 597940
rect 700922 597884 701922 597940
rect 709211 597936 710211 597960
rect 682921 597593 683521 597643
rect 684070 597599 684670 597649
rect 685537 597593 686137 597649
rect 699322 597623 700322 597673
rect 700922 597623 701922 597673
rect 680215 597518 680815 597574
rect 707610 597523 708610 597617
rect 709211 597523 710211 597591
rect 707610 597513 707624 597523
rect 707658 597513 707695 597523
rect 707729 597513 707769 597523
rect 707803 597513 707840 597523
rect 707874 597513 707914 597523
rect 707948 597513 707985 597523
rect 708019 597513 708059 597523
rect 708093 597513 708130 597523
rect 708164 597513 708204 597523
rect 708238 597513 708275 597523
rect 708309 597513 708369 597523
rect 708403 597513 708446 597523
rect 708480 597513 708522 597523
rect 708556 597513 708604 597523
rect 709219 597513 709270 597523
rect 709304 597513 709364 597523
rect 709398 597513 709435 597523
rect 709469 597513 709509 597523
rect 709543 597513 709580 597523
rect 709614 597513 709654 597523
rect 709688 597513 709725 597523
rect 709759 597513 709799 597523
rect 709833 597513 709870 597523
rect 709904 597513 709944 597523
rect 709978 597513 710015 597523
rect 710049 597513 710089 597523
rect 710123 597513 710160 597523
rect 710194 597513 710211 597523
rect 684070 597443 684670 597499
rect 685537 597443 686137 597493
rect 692428 597442 693028 597492
rect 680215 597348 680815 597398
rect 681713 597359 682313 597409
rect 684070 597293 684670 597343
rect 692428 597292 693028 597342
rect 705107 597336 705173 597352
rect 711579 597301 711595 598520
rect 711892 597697 711942 598520
rect 712062 597697 712112 598520
rect 716071 598357 716074 598358
rect 714645 598323 714752 598357
rect 716071 598356 716072 598357
rect 716073 598356 716074 598357
rect 716071 598355 716074 598356
rect 716208 598357 716211 598358
rect 716208 598356 716209 598357
rect 716210 598356 716211 598357
rect 716208 598355 716211 598356
rect 714964 598247 715998 598329
rect 716284 598247 717318 598329
rect 714175 597398 714225 597998
rect 714425 597398 714475 597998
rect 680215 597232 680815 597282
rect 698017 597232 698053 597260
rect 692428 597162 693028 597212
rect 698030 597198 698077 597232
rect 698017 597164 698053 597198
rect 680215 597056 680815 597112
rect 692428 597006 693028 597134
rect 698030 597130 698077 597164
rect 698017 597096 698053 597130
rect 698030 597062 698077 597096
rect 698017 596983 698053 597062
rect 698084 596983 698120 597260
rect 714781 597191 714863 598226
rect 715134 597955 715828 598037
rect 714686 597123 714863 597191
rect 714645 597089 714863 597123
rect 680215 596880 680815 596936
rect 686719 596893 686739 596917
rect 686743 596893 686753 596917
rect 686719 596859 686757 596893
rect 686719 596822 686739 596859
rect 686743 596822 686753 596859
rect 692428 596850 693028 596978
rect 698017 596947 698210 596983
rect 698084 596935 698210 596947
rect 702756 596959 703645 596983
rect 702756 596935 702853 596959
rect 698084 596828 702853 596935
rect 686719 596788 686757 596822
rect 680215 596704 680815 596760
rect 686719 596751 686739 596788
rect 686743 596751 686753 596788
rect 686719 596741 686757 596751
rect 686699 596717 686767 596741
rect 686719 596704 686739 596717
rect 686743 596704 686753 596717
rect 686719 596695 686753 596704
rect 686719 596693 686743 596695
rect 692428 596694 693028 596750
rect 686685 596656 686709 596680
rect 686743 596656 686767 596680
rect 678799 596503 679399 596553
rect 680215 596534 680815 596584
rect 692428 596538 693028 596666
rect 680593 596531 680815 596534
rect 682009 596501 682069 596516
rect 682024 596465 682054 596501
rect 683708 596387 684308 596437
rect 678799 596327 679399 596383
rect 692428 596382 693028 596510
rect 714781 596308 714863 597089
rect 715063 596609 715145 597915
rect 715289 596777 715339 597719
rect 715633 596777 715683 597719
rect 715382 596672 715422 596756
rect 715542 596672 715582 596756
rect 715342 596632 715382 596672
rect 715582 596632 715622 596672
rect 715815 596609 715897 597915
rect 715134 596387 715828 596469
rect 716100 596308 716182 598226
rect 716454 597955 717148 598037
rect 716385 596609 716467 597915
rect 716599 596777 716649 597719
rect 716943 596777 716993 597719
rect 716700 596672 716740 596756
rect 716860 596672 716900 596756
rect 716660 596632 716700 596672
rect 716900 596632 716940 596672
rect 717137 596609 717219 597915
rect 716454 596387 717148 596469
rect 717419 596308 717501 598226
rect 683708 596237 684308 596287
rect 692428 596232 693028 596282
rect 678799 596157 679399 596207
rect 684565 596160 684790 596168
rect 696597 596000 696600 596120
rect 714964 596095 715998 596177
rect 716284 596095 717318 596177
rect 21000 569000 21003 569120
rect 282 568623 1316 568705
rect 1602 568623 2636 568705
rect 32810 568662 33035 568670
rect 38201 568593 38801 568643
rect 24572 568518 25172 568568
rect 33292 568513 33892 568563
rect 99 566574 181 568492
rect 452 568331 1146 568413
rect 381 566885 463 568191
rect 660 568128 700 568168
rect 900 568128 940 568168
rect 700 568044 740 568128
rect 860 568044 900 568128
rect 607 567081 657 568023
rect 951 567081 1001 568023
rect 1133 566885 1215 568191
rect 452 566763 1146 566845
rect 1418 566574 1500 568492
rect 1772 568331 2466 568413
rect 1703 566885 1785 568191
rect 1978 568128 2018 568168
rect 2218 568128 2258 568168
rect 2018 568044 2058 568128
rect 2178 568044 2218 568128
rect 1917 567081 1967 568023
rect 2261 567081 2311 568023
rect 2455 566885 2537 568191
rect 2737 567779 2819 568492
rect 24572 568362 25172 568490
rect 38201 568417 38801 568473
rect 33292 568363 33892 568413
rect 24572 568206 25172 568334
rect 35546 568299 35576 568335
rect 36785 568329 36935 568341
rect 35531 568284 35591 568299
rect 36785 568216 37385 568266
rect 38201 568247 38801 568297
rect 30833 568120 30857 568144
rect 30891 568120 30915 568144
rect 24572 568050 25172 568106
rect 30857 568105 30881 568107
rect 30857 568096 30887 568105
rect 30867 568083 30887 568096
rect 30891 568083 30907 568120
rect 30833 568059 30857 568083
rect 30867 568049 30911 568083
rect 14747 567865 19516 567972
rect 24572 567894 25172 568022
rect 30867 568012 30887 568049
rect 30891 568012 30907 568049
rect 36785 568040 37385 568096
rect 30867 567978 30911 568012
rect 30867 567941 30887 567978
rect 30891 567941 30907 567978
rect 30867 567907 30911 567941
rect 30867 567883 30887 567907
rect 30891 567883 30907 567907
rect 14747 567841 14844 567865
rect 13955 567817 14844 567841
rect 19390 567853 19516 567865
rect 19390 567841 19583 567853
rect 19390 567817 19605 567841
rect 19639 567817 19673 567841
rect 19707 567817 19741 567841
rect 19775 567817 19809 567841
rect 19843 567817 19877 567841
rect 19911 567817 19945 567841
rect 19979 567817 20013 567841
rect 20047 567817 20081 567841
rect 20115 567817 20149 567841
rect 20183 567817 20217 567841
rect 20251 567817 20285 567841
rect 20319 567817 20353 567841
rect 20387 567817 20421 567841
rect 20455 567817 20489 567841
rect 20523 567817 20557 567841
rect 20591 567817 20625 567841
rect 20659 567817 20693 567841
rect 2737 567711 2914 567779
rect 1772 566763 2466 566845
rect 2737 566574 2819 567711
rect 2848 567677 2955 567711
rect 19480 567540 19516 567817
rect 19547 567540 19583 567817
rect 24572 567738 25172 567866
rect 36785 567864 37385 567920
rect 36785 567688 37385 567744
rect 20809 567650 20833 567684
rect 20809 567582 20833 567616
rect 24572 567588 25172 567638
rect 20809 567540 20833 567548
rect 36785 567518 37385 567568
rect 3125 566802 3175 567402
rect 3375 566802 3425 567402
rect 282 566471 1316 566553
rect 1602 566471 2636 566553
rect 1389 566444 1392 566445
rect 1389 566443 1390 566444
rect 1391 566443 1392 566444
rect 1389 566442 1392 566443
rect 1526 566444 1529 566445
rect 1526 566443 1527 566444
rect 1528 566443 1529 566444
rect 2848 566443 2955 566477
rect 1526 566442 1529 566443
rect 5488 566280 5538 567103
rect 5658 566280 5708 567103
rect 6005 566280 6021 567499
rect 12427 567448 12493 567464
rect 24572 567458 25172 567508
rect 32930 567457 33530 567507
rect 35287 567391 35887 567441
rect 36785 567402 37385 567452
rect 24572 567308 25172 567358
rect 31463 567307 32063 567357
rect 32930 567301 33530 567357
rect 7389 567277 7406 567287
rect 7440 567277 7477 567287
rect 7511 567277 7551 567287
rect 7585 567277 7622 567287
rect 7656 567277 7696 567287
rect 7730 567277 7767 567287
rect 7801 567277 7841 567287
rect 7875 567277 7912 567287
rect 7946 567277 7986 567287
rect 8020 567277 8057 567287
rect 8091 567277 8131 567287
rect 8165 567277 8202 567287
rect 8236 567277 8296 567287
rect 8330 567277 8381 567287
rect 8996 567277 9044 567287
rect 9078 567277 9120 567287
rect 9154 567277 9197 567287
rect 9231 567277 9291 567287
rect 9325 567277 9362 567287
rect 9396 567277 9436 567287
rect 9470 567277 9507 567287
rect 9541 567277 9581 567287
rect 9615 567277 9652 567287
rect 9686 567277 9726 567287
rect 9760 567277 9797 567287
rect 9831 567277 9871 567287
rect 9905 567277 9942 567287
rect 9976 567277 9990 567287
rect 7389 567209 8389 567277
rect 8990 567183 9990 567277
rect 36785 567226 37385 567282
rect 15678 567127 16678 567177
rect 17278 567127 18278 567177
rect 31463 567151 32063 567207
rect 32930 567151 33530 567201
rect 34079 567157 34679 567207
rect 7389 566840 8389 566864
rect 15678 566860 16678 566916
rect 17278 566860 18278 566916
rect 8990 566840 9990 566841
rect 7389 566743 8389 566799
rect 8990 566743 9990 566799
rect 15678 566788 16678 566844
rect 17278 566788 18278 566844
rect 8990 566701 9990 566702
rect 15678 566286 16678 566426
rect 17278 566286 18278 566426
rect 19844 566280 19894 567051
rect 20462 566280 20512 567051
rect 31463 567001 32063 567051
rect 34079 567001 34679 567057
rect 35287 567039 35887 567095
rect 36785 567050 37385 567106
rect 32596 566929 33596 566979
rect 24573 566820 25173 566870
rect 34079 566851 34679 566901
rect 35287 566869 35887 566919
rect 36785 566880 37385 566930
rect 30171 566795 30771 566845
rect 32596 566773 33596 566829
rect 37993 566704 38593 566754
rect 30171 566619 30771 566675
rect 32596 566623 33596 566673
rect 34110 566589 34710 566639
rect 21263 566280 21313 566518
rect 22349 566280 22399 566518
rect 32596 566507 33596 566557
rect 30171 566449 30771 566499
rect 36785 566429 36985 566609
rect 37993 566534 38593 566584
rect 24573 566352 25173 566408
rect 29993 566310 30993 566360
rect 31347 566280 31547 566317
rect 31607 566280 31807 566317
rect 36785 566280 36985 566373
rect 37083 566280 37120 566373
rect 696597 560200 696600 560320
rect 692376 559983 692396 560017
rect 692463 559993 692532 560017
rect 696191 559993 696239 560017
rect 692487 559983 692532 559993
rect 696204 559983 696239 559993
rect 696340 559983 696360 560017
rect 692487 559915 692502 559939
rect 696200 559915 696215 559939
rect 692454 559891 692478 559915
rect 696224 559891 696248 559915
rect 686755 559800 687355 559850
rect 692487 559748 692505 559752
rect 692479 559718 692505 559748
rect 692487 559698 692505 559718
rect 686755 559624 687355 559680
rect 692485 559674 692505 559698
rect 692509 559674 692517 559718
rect 696215 559698 696223 559748
rect 696203 559674 696223 559698
rect 696227 559674 696245 559752
rect 692485 559640 692521 559674
rect 696203 559640 696249 559674
rect 686755 559448 687355 559504
rect 686755 559278 687355 559328
rect 685547 559102 686147 559152
rect 687155 559007 687170 559022
rect 687343 559018 687355 559022
rect 687340 559007 687355 559018
rect 685547 558932 686147 558982
rect 687155 558827 687355 559007
rect 687155 558812 687170 558827
rect 687340 558816 687355 558827
rect 687343 558812 687355 558816
rect 687042 558771 687057 558786
rect 687020 558591 687057 558771
rect 687042 558576 687057 558591
rect 687155 558771 687170 558786
rect 687343 558782 687355 558786
rect 687340 558771 687355 558782
rect 687155 558591 687355 558771
rect 688210 558630 688260 559630
rect 688360 558630 688488 559630
rect 688516 558630 688644 559630
rect 688672 558630 688800 559630
rect 688828 558630 688956 559630
rect 688984 558630 689112 559630
rect 689140 558630 689268 559630
rect 689296 558630 689424 559630
rect 689452 558630 689580 559630
rect 689608 558630 689736 559630
rect 689764 558630 689892 559630
rect 689920 558630 690048 559630
rect 690076 558630 690204 559630
rect 690232 558630 690360 559630
rect 690388 558630 690438 559630
rect 692485 559606 692505 559640
rect 692509 559606 692517 559640
rect 696203 559606 696223 559640
rect 696227 559606 696245 559640
rect 691275 559523 691875 559573
rect 692485 559572 692521 559606
rect 696203 559572 696249 559606
rect 692485 559538 692505 559572
rect 692509 559538 692517 559572
rect 692485 559504 692521 559538
rect 692583 559528 693983 559571
rect 694719 559528 696119 559571
rect 696203 559538 696223 559572
rect 696227 559538 696245 559572
rect 696203 559504 696249 559538
rect 692485 559470 692505 559504
rect 692509 559470 692517 559504
rect 692485 559436 692521 559470
rect 691275 559373 691875 559423
rect 692485 559402 692505 559436
rect 692509 559402 692517 559436
rect 692485 559368 692521 559402
rect 692485 559334 692505 559368
rect 692509 559334 692517 559368
rect 692583 559365 693983 559493
rect 694719 559365 696119 559493
rect 696203 559470 696223 559504
rect 696227 559470 696245 559504
rect 696203 559436 696249 559470
rect 707624 559441 707658 559475
rect 707695 559441 707729 559475
rect 707769 559441 707803 559475
rect 707840 559441 707874 559475
rect 707914 559441 707948 559475
rect 707985 559441 708019 559475
rect 708059 559441 708093 559475
rect 708130 559441 708164 559475
rect 708204 559441 708238 559475
rect 708275 559441 708309 559475
rect 708369 559441 708403 559475
rect 708446 559441 708480 559475
rect 708520 559441 708554 559465
rect 708588 559441 708610 559465
rect 709211 559441 709234 559465
rect 709270 559441 709304 559475
rect 709364 559441 709398 559475
rect 709435 559441 709469 559475
rect 709509 559441 709543 559475
rect 709580 559441 709614 559475
rect 709654 559441 709688 559475
rect 709725 559441 709759 559475
rect 709799 559441 709833 559475
rect 709870 559441 709904 559475
rect 709944 559441 709978 559475
rect 710015 559441 710049 559475
rect 710089 559441 710123 559475
rect 710160 559441 710194 559475
rect 696203 559402 696223 559436
rect 696227 559402 696245 559436
rect 707610 559431 707624 559441
rect 707658 559431 707695 559441
rect 707729 559431 707769 559441
rect 707803 559431 707840 559441
rect 707874 559431 707914 559441
rect 707948 559431 707985 559441
rect 708019 559431 708059 559441
rect 708093 559431 708130 559441
rect 708164 559431 708204 559441
rect 708238 559431 708275 559441
rect 708309 559431 708369 559441
rect 708403 559431 708446 559441
rect 708480 559431 708520 559441
rect 708554 559431 708588 559441
rect 708610 559431 708634 559441
rect 709211 559431 709270 559441
rect 709304 559431 709364 559441
rect 709398 559431 709435 559441
rect 709469 559431 709509 559441
rect 709543 559431 709580 559441
rect 709614 559431 709654 559441
rect 709688 559431 709725 559441
rect 709759 559431 709799 559441
rect 709833 559431 709870 559441
rect 709904 559431 709944 559441
rect 709978 559431 710015 559441
rect 710049 559431 710089 559441
rect 710123 559431 710160 559441
rect 710194 559431 710211 559441
rect 696203 559368 696249 559402
rect 696203 559334 696223 559368
rect 696227 559334 696245 559368
rect 707610 559337 708610 559431
rect 709211 559337 710211 559431
rect 691275 559251 691875 559301
rect 692485 559300 692521 559334
rect 692485 559266 692505 559300
rect 692509 559266 692517 559300
rect 692485 559232 692521 559266
rect 692485 559198 692505 559232
rect 692509 559198 692517 559232
rect 692583 559202 693983 559330
rect 694719 559202 696119 559330
rect 696203 559300 696249 559334
rect 711579 559317 712463 559331
rect 711579 559307 711619 559317
rect 696203 559266 696223 559300
rect 696227 559266 696245 559300
rect 701730 559290 701747 559292
rect 696203 559232 696249 559266
rect 696203 559198 696223 559232
rect 696227 559198 696245 559232
rect 701692 559220 701722 559254
rect 701730 559220 701760 559290
rect 707610 559241 708610 559301
rect 709211 559241 710211 559301
rect 692485 559164 692521 559198
rect 691275 559101 691875 559151
rect 692485 559130 692505 559164
rect 692509 559130 692517 559164
rect 692485 559096 692521 559130
rect 692485 559062 692505 559096
rect 692509 559062 692517 559096
rect 692485 559028 692521 559062
rect 692583 559039 693983 559167
rect 694719 559039 696119 559167
rect 696203 559164 696249 559198
rect 696203 559130 696223 559164
rect 696227 559130 696245 559164
rect 696203 559096 696249 559130
rect 696203 559062 696223 559096
rect 696227 559062 696245 559096
rect 699322 559064 700322 559097
rect 700922 559064 701922 559097
rect 696203 559028 696249 559062
rect 707610 559044 708610 559048
rect 709211 559044 710211 559048
rect 691275 558975 691875 559025
rect 692485 558994 692505 559028
rect 692509 558994 692517 559028
rect 692485 558960 692521 558994
rect 692485 558926 692505 558960
rect 692509 558926 692517 558960
rect 692485 558892 692521 558926
rect 691275 558825 691875 558875
rect 692485 558858 692505 558892
rect 692509 558858 692517 558892
rect 692583 558876 693983 559004
rect 694719 558876 696119 559004
rect 696203 558994 696223 559028
rect 696227 558994 696245 559028
rect 707574 558994 708646 559030
rect 696203 558960 696249 558994
rect 696203 558926 696223 558960
rect 696227 558926 696245 558960
rect 707574 558953 707610 558994
rect 708610 558953 708646 558994
rect 696203 558892 696249 558926
rect 697284 558894 697350 558910
rect 707574 558897 708646 558953
rect 696203 558858 696223 558892
rect 696227 558858 696245 558892
rect 699322 558877 700322 558894
rect 700922 558877 701922 558894
rect 707574 558881 707610 558897
rect 708610 558881 708646 558897
rect 692485 558824 692521 558858
rect 692485 558790 692505 558824
rect 692509 558790 692517 558824
rect 692485 558756 692521 558790
rect 691275 558703 691875 558753
rect 692485 558722 692505 558756
rect 692509 558722 692517 558756
rect 692485 558688 692521 558722
rect 692583 558713 693983 558841
rect 694719 558713 696119 558841
rect 696203 558824 696249 558858
rect 707574 558825 708646 558881
rect 696203 558790 696223 558824
rect 696227 558790 696245 558824
rect 696203 558756 696249 558790
rect 696203 558722 696223 558756
rect 696227 558722 696245 558756
rect 699322 558739 700322 558811
rect 700922 558739 701922 558811
rect 707574 558788 707610 558825
rect 708610 558788 708646 558825
rect 707574 558748 708646 558788
rect 709175 558994 710247 559030
rect 709175 558953 709211 558994
rect 710211 558953 710247 558994
rect 709175 558897 710247 558953
rect 709175 558881 709211 558897
rect 710211 558881 710247 558897
rect 709175 558825 710247 558881
rect 709175 558788 709211 558825
rect 710211 558788 710247 558825
rect 709175 558748 710247 558788
rect 696203 558688 696249 558722
rect 692485 558654 692505 558688
rect 692509 558654 692517 558688
rect 692485 558620 692521 558654
rect 687155 558576 687170 558591
rect 687340 558580 687355 558591
rect 687343 558576 687355 558580
rect 685542 558506 686142 558556
rect 691275 558553 691875 558603
rect 692485 558586 692505 558620
rect 692509 558586 692517 558620
rect 692485 558552 692521 558586
rect 692485 558518 692505 558552
rect 692509 558518 692517 558552
rect 692583 558550 693983 558678
rect 694719 558550 696119 558678
rect 696203 558654 696223 558688
rect 696227 558654 696245 558688
rect 696203 558620 696249 558654
rect 696203 558586 696223 558620
rect 696227 558586 696245 558620
rect 696203 558552 696249 558586
rect 696203 558518 696223 558552
rect 696227 558518 696245 558552
rect 692485 558484 692521 558518
rect 692485 558450 692505 558484
rect 692509 558450 692517 558484
rect 692485 558416 692521 558450
rect 679817 558330 679841 558354
rect 685542 558330 686142 558386
rect 692485 558382 692505 558416
rect 692509 558382 692517 558416
rect 692583 558387 693983 558515
rect 694719 558387 696119 558515
rect 696203 558484 696249 558518
rect 696203 558450 696223 558484
rect 696227 558450 696245 558484
rect 699322 558478 700322 558550
rect 700922 558478 701922 558550
rect 707610 558523 708610 558595
rect 709211 558523 710211 558595
rect 699392 558467 699426 558478
rect 699460 558467 699494 558478
rect 699528 558467 699562 558478
rect 699596 558467 699630 558478
rect 699664 558467 699698 558478
rect 699732 558467 699766 558478
rect 699800 558467 699834 558478
rect 699868 558467 699902 558478
rect 699936 558467 699970 558478
rect 700004 558467 700038 558478
rect 700072 558467 700106 558478
rect 700140 558467 700174 558478
rect 700208 558467 700242 558478
rect 700276 558467 700310 558478
rect 700934 558467 700968 558478
rect 701002 558467 701036 558478
rect 701070 558467 701104 558478
rect 701138 558467 701172 558478
rect 701206 558467 701240 558478
rect 701274 558467 701308 558478
rect 701342 558467 701376 558478
rect 701410 558467 701444 558478
rect 701478 558467 701512 558478
rect 701546 558467 701580 558478
rect 701614 558467 701648 558478
rect 701682 558467 701716 558478
rect 701750 558467 701784 558478
rect 701818 558467 701852 558478
rect 699392 558457 699450 558467
rect 699460 558457 699518 558467
rect 699528 558457 699586 558467
rect 699596 558457 699654 558467
rect 699664 558457 699722 558467
rect 699732 558457 699790 558467
rect 699800 558457 699858 558467
rect 699868 558457 699926 558467
rect 699936 558457 699994 558467
rect 700004 558457 700062 558467
rect 700072 558457 700130 558467
rect 700140 558457 700198 558467
rect 700208 558457 700266 558467
rect 700276 558457 700334 558467
rect 700934 558457 700992 558467
rect 701002 558457 701060 558467
rect 701070 558457 701128 558467
rect 701138 558457 701196 558467
rect 701206 558457 701264 558467
rect 701274 558457 701332 558467
rect 701342 558457 701400 558467
rect 701410 558457 701468 558467
rect 701478 558457 701536 558467
rect 701546 558457 701604 558467
rect 701614 558457 701672 558467
rect 701682 558457 701740 558467
rect 701750 558457 701808 558467
rect 701818 558457 701876 558467
rect 696203 558416 696249 558450
rect 699368 558433 700334 558457
rect 700910 558433 701876 558457
rect 699392 558418 699416 558433
rect 699460 558418 699484 558433
rect 699528 558418 699552 558433
rect 699596 558418 699620 558433
rect 699664 558418 699688 558433
rect 699732 558418 699756 558433
rect 699800 558418 699824 558433
rect 699868 558418 699892 558433
rect 699936 558418 699960 558433
rect 700004 558418 700028 558433
rect 700072 558418 700096 558433
rect 700140 558418 700164 558433
rect 700208 558418 700232 558433
rect 700276 558418 700300 558433
rect 700934 558418 700958 558433
rect 701002 558418 701026 558433
rect 701070 558418 701094 558433
rect 701138 558418 701162 558433
rect 701206 558418 701230 558433
rect 701274 558418 701298 558433
rect 701342 558418 701366 558433
rect 701410 558418 701434 558433
rect 701478 558418 701502 558433
rect 701546 558418 701570 558433
rect 701614 558418 701638 558433
rect 701682 558418 701706 558433
rect 701750 558418 701774 558433
rect 701818 558418 701842 558433
rect 696203 558382 696223 558416
rect 696227 558382 696245 558416
rect 692485 558348 692521 558382
rect 696203 558348 696249 558382
rect 679549 558307 679573 558330
rect 679793 558306 679808 558330
rect 692485 558314 692505 558348
rect 692509 558314 692517 558348
rect 696203 558314 696223 558348
rect 696227 558314 696245 558348
rect 692485 558280 692521 558314
rect 696203 558280 696249 558314
rect 679549 558237 679573 558271
rect 692485 558246 692505 558280
rect 692509 558246 692517 558280
rect 692485 558212 692521 558246
rect 692583 558237 693983 558280
rect 694719 558237 696119 558280
rect 696203 558246 696223 558280
rect 696227 558246 696245 558280
rect 699322 558263 700322 558418
rect 696203 558212 696249 558246
rect 699322 558229 700334 558263
rect 700922 558253 701922 558418
rect 700910 558229 701922 558253
rect 699322 558218 700322 558229
rect 700922 558218 701922 558229
rect 707574 558263 708646 558299
rect 707574 558226 707610 558263
rect 708610 558226 708646 558263
rect 679549 558167 679573 558201
rect 685542 558160 686142 558210
rect 685601 558157 685895 558160
rect 685920 558157 686142 558160
rect 692485 558178 692505 558212
rect 692509 558178 692517 558212
rect 696203 558178 696223 558212
rect 696227 558178 696245 558212
rect 699392 558205 699416 558218
rect 699460 558205 699484 558218
rect 699528 558205 699552 558218
rect 699596 558205 699620 558218
rect 699664 558205 699688 558218
rect 699732 558205 699756 558218
rect 699800 558205 699824 558218
rect 699868 558205 699892 558218
rect 699936 558205 699960 558218
rect 700004 558205 700028 558218
rect 700072 558205 700096 558218
rect 700140 558205 700164 558218
rect 700208 558205 700232 558218
rect 700276 558205 700300 558218
rect 700934 558205 700958 558218
rect 701002 558205 701026 558218
rect 701070 558205 701094 558218
rect 701138 558205 701162 558218
rect 701206 558205 701230 558218
rect 701274 558205 701298 558218
rect 701342 558205 701366 558218
rect 701410 558205 701434 558218
rect 701478 558205 701502 558218
rect 701546 558205 701570 558218
rect 701614 558205 701638 558218
rect 701682 558205 701706 558218
rect 701750 558205 701774 558218
rect 701818 558205 701842 558218
rect 707574 558186 708646 558226
rect 709175 558263 710247 558299
rect 709175 558226 709211 558263
rect 710211 558226 710247 558263
rect 709175 558186 710247 558226
rect 692485 558144 692521 558178
rect 696203 558144 696249 558178
rect 679549 558097 679573 558131
rect 692485 558110 692505 558144
rect 692509 558110 692517 558144
rect 692485 558076 692521 558110
rect 692583 558101 693983 558144
rect 694719 558101 696119 558144
rect 696203 558110 696223 558144
rect 696227 558110 696245 558144
rect 696203 558076 696249 558110
rect 679549 558027 679573 558061
rect 692485 558042 692505 558076
rect 692509 558042 692517 558076
rect 692485 558008 692521 558042
rect 679549 557957 679573 557991
rect 692485 557974 692505 558008
rect 692509 557974 692517 558008
rect 679793 557933 679808 557957
rect 692485 557940 692521 557974
rect 679817 557909 679841 557933
rect 692485 557906 692505 557940
rect 692509 557906 692517 557940
rect 692583 557938 693983 558066
rect 694719 557938 696119 558066
rect 696203 558042 696223 558076
rect 696227 558042 696245 558076
rect 696203 558008 696249 558042
rect 696203 557974 696223 558008
rect 696227 557974 696245 558008
rect 696203 557940 696249 557974
rect 696203 557906 696223 557940
rect 696227 557906 696245 557940
rect 687685 557838 687709 557862
rect 687661 557814 687675 557838
rect 687669 557797 687675 557814
rect 679515 557762 679539 557785
rect 679613 557762 679637 557785
rect 679491 557737 679515 557761
rect 679637 557737 679661 557761
rect 680215 557678 680815 557728
rect 680215 557502 680815 557558
rect 685551 557516 686551 557566
rect 680215 557326 680815 557382
rect 685551 557360 686551 557488
rect 689154 557439 689204 557897
rect 689151 557355 689204 557439
rect 680215 557156 680815 557206
rect 685551 557204 686551 557332
rect 685551 557048 686551 557176
rect 686865 557116 687465 557166
rect 679007 556980 679607 557030
rect 680615 556885 680630 556900
rect 680803 556896 680815 556900
rect 680800 556885 680815 556896
rect 685551 556892 686551 556948
rect 686865 556940 687465 557068
rect 679007 556810 679607 556860
rect 680615 556705 680815 556885
rect 683328 556793 683928 556843
rect 682573 556717 683173 556767
rect 680615 556690 680630 556705
rect 680800 556694 680815 556705
rect 680803 556690 680815 556694
rect 680502 556649 680517 556664
rect 680480 556469 680517 556649
rect 680502 556454 680517 556469
rect 680615 556649 680630 556664
rect 680803 556660 680815 556664
rect 680800 556649 680815 556660
rect 680615 556469 680815 556649
rect 682573 556541 683173 556669
rect 683328 556617 683928 556745
rect 685551 556736 686551 556864
rect 686865 556764 687465 556820
rect 685551 556580 686551 556708
rect 686865 556588 687465 556716
rect 680615 556454 680630 556469
rect 680800 556458 680815 556469
rect 680803 556454 680815 556458
rect 683328 556441 683928 556497
rect 679002 556384 679602 556434
rect 685551 556424 686551 556552
rect 682573 556365 683173 556421
rect 686865 556412 687465 556468
rect 679002 556208 679602 556264
rect 682573 556189 683173 556317
rect 683328 556265 683928 556321
rect 685551 556274 686551 556324
rect 686865 556236 687465 556364
rect 685551 556158 686551 556208
rect 678680 556123 678704 556157
rect 678680 556055 678704 556089
rect 679002 556038 679602 556088
rect 679061 556035 679355 556038
rect 679380 556035 679602 556038
rect 678680 555987 678704 556021
rect 682573 556013 683173 556141
rect 683328 556089 683928 556145
rect 678680 555919 678704 555953
rect 678680 555851 678704 555885
rect 682573 555837 683173 555965
rect 683328 555913 683928 556041
rect 685551 555982 686551 556110
rect 686865 556060 687465 556116
rect 678680 555783 678704 555817
rect 685551 555806 686551 555934
rect 686865 555884 687465 556012
rect 678680 555715 678704 555749
rect 678680 555647 678704 555681
rect 682573 555661 683173 555789
rect 683328 555737 683928 555793
rect 685551 555630 686551 555758
rect 686865 555708 687465 555836
rect 678680 555579 678704 555613
rect 683328 555567 683928 555617
rect 678680 555511 678704 555545
rect 682573 555491 683173 555541
rect 684519 555498 685119 555548
rect 678680 555443 678704 555477
rect 685551 555454 686551 555582
rect 686865 555532 687465 555660
rect 679133 555409 679283 555421
rect 679452 555409 679602 555421
rect 678680 555375 678704 555409
rect 2850 555304 3850 555320
rect 2850 555188 3850 555238
rect 2850 554978 3850 555028
rect 3959 555015 3960 555320
rect 5169 555315 5191 555320
rect 6005 555305 6021 555320
rect 1288 553503 1338 554503
rect 1438 553503 1566 554060
rect 1594 553503 1644 554503
rect 5995 553493 6021 555275
rect 7389 554911 8389 554967
rect 8990 554911 9990 554967
rect 15678 554956 16678 555012
rect 17278 554956 18278 555012
rect 7389 554839 8389 554895
rect 8990 554839 9990 554895
rect 15678 554884 16678 554940
rect 17278 554884 18278 554940
rect 27622 554903 27672 555320
rect 27772 554903 27828 555320
rect 27928 554903 27984 555320
rect 28084 554903 28140 555320
rect 28240 554903 28296 555320
rect 28396 554903 28446 555320
rect 678680 555307 678704 555341
rect 31049 555234 32049 555284
rect 36785 555242 37385 555298
rect 679002 555296 679602 555346
rect 684519 555342 685119 555398
rect 685551 555278 686551 555406
rect 686865 555356 687465 555484
rect 678680 555239 678704 555273
rect 678680 555171 678704 555205
rect 684519 555192 685119 555242
rect 36785 555072 37385 555122
rect 678680 555103 678704 555137
rect 679002 555120 679602 555176
rect 681745 555081 682345 555131
rect 682509 555069 683109 555119
rect 678680 555035 678704 555069
rect 683739 555027 684339 555077
rect 684519 555062 685119 555112
rect 685551 555102 686551 555230
rect 686865 555180 687465 555308
rect 678680 554967 678704 555001
rect 679002 554950 679602 555000
rect 678680 554899 678704 554933
rect 680502 554915 680517 554930
rect 678680 554831 678704 554865
rect 678680 554763 678704 554797
rect 680480 554735 680517 554915
rect 21481 554656 22881 554699
rect 23617 554656 25017 554699
rect 678680 554695 678704 554729
rect 680502 554720 680517 554735
rect 680615 554915 680630 554930
rect 680803 554926 680815 554930
rect 680800 554915 680815 554926
rect 681745 554925 682345 554981
rect 680615 554735 680815 554915
rect 681745 554769 682345 554897
rect 682509 554893 683109 555021
rect 684519 554906 685119 555034
rect 685551 554926 686551 555054
rect 686865 555004 687465 555060
rect 683739 554837 684339 554893
rect 686865 554828 687465 554956
rect 680615 554720 680630 554735
rect 680800 554724 680815 554735
rect 680803 554720 680815 554724
rect 680615 554679 680630 554694
rect 680803 554690 680815 554694
rect 680800 554679 680815 554690
rect 31458 554590 32058 554640
rect 678680 554627 678704 554661
rect 15678 554382 16678 554522
rect 17278 554382 18278 554522
rect 21481 554520 22881 554563
rect 23617 554520 25017 554563
rect 678680 554559 678704 554593
rect 678680 554491 678704 554525
rect 679007 554524 679607 554574
rect 680615 554499 680815 554679
rect 681745 554613 682345 554741
rect 682509 554717 683109 554773
rect 684519 554750 685119 554806
rect 685551 554750 686551 554806
rect 682509 554541 683109 554669
rect 684519 554594 685119 554722
rect 685551 554594 686551 554722
rect 686865 554652 687465 554780
rect 680615 554484 680630 554499
rect 680800 554488 680815 554499
rect 680803 554484 680815 554488
rect 31458 554414 32058 554470
rect 681745 554463 682345 554513
rect 683739 554477 684339 554513
rect 678680 554423 678704 554457
rect 684519 554444 685119 554494
rect 685551 554438 686551 554566
rect 686865 554476 687465 554604
rect 678680 554355 678704 554389
rect 679007 554354 679607 554404
rect 682509 554371 683109 554421
rect 25725 554197 26325 554247
rect 31458 554244 32058 554294
rect 678680 554287 678704 554321
rect 684519 554314 685119 554364
rect 678680 554219 678704 554253
rect 7353 554016 8425 554052
rect 7353 553975 7389 554016
rect 8389 553975 8425 554016
rect 7353 553919 8425 553975
rect 7353 553903 7389 553919
rect 8389 553903 8425 553919
rect 7353 553847 8425 553903
rect 7353 553810 7389 553847
rect 8389 553810 8425 553847
rect 7353 553770 8425 553810
rect 8954 554016 10026 554052
rect 8954 553975 8990 554016
rect 9990 553975 10026 554016
rect 8954 553919 10026 553975
rect 21383 554044 21403 554060
rect 21407 554044 21415 554060
rect 21383 554010 21419 554044
rect 21481 554031 22881 554060
rect 23617 554031 25017 554060
rect 25101 554044 25121 554060
rect 25125 554044 25143 554060
rect 25725 554047 26325 554097
rect 25101 554010 25147 554044
rect 21383 553976 21403 554010
rect 21407 553976 21415 554010
rect 21383 553942 21419 553976
rect 8954 553903 8990 553919
rect 9990 553903 10026 553919
rect 15678 553906 16678 553923
rect 17278 553906 18278 553923
rect 21383 553908 21403 553942
rect 21407 553908 21415 553942
rect 8954 553847 10026 553903
rect 20250 553890 20316 553906
rect 8954 553810 8990 553847
rect 9990 553810 10026 553847
rect 8954 553770 10026 553810
rect 21383 553874 21419 553908
rect 21383 553840 21403 553874
rect 21407 553840 21415 553874
rect 21481 553868 22881 553996
rect 23617 553868 25017 553996
rect 25101 553976 25121 554010
rect 25125 553976 25143 554010
rect 25101 553942 25147 553976
rect 25101 553908 25121 553942
rect 25125 553908 25143 553942
rect 25725 553925 26325 553975
rect 25101 553874 25147 553908
rect 25101 553840 25121 553874
rect 25125 553840 25143 553874
rect 21383 553806 21419 553840
rect 21383 553772 21403 553806
rect 21407 553772 21415 553806
rect 21383 553738 21419 553772
rect 15678 553703 16678 553736
rect 17278 553703 18278 553736
rect 21383 553704 21403 553738
rect 21407 553704 21415 553738
rect 21481 553705 22881 553833
rect 23617 553705 25017 553833
rect 25101 553806 25147 553840
rect 25101 553772 25121 553806
rect 25125 553772 25143 553806
rect 25725 553775 26325 553825
rect 25101 553738 25147 553772
rect 25101 553704 25121 553738
rect 25125 553704 25143 553738
rect 21383 553670 21419 553704
rect 25101 553670 25147 553704
rect 21383 553636 21403 553670
rect 21407 553636 21415 553670
rect 7389 553559 8389 553631
rect 8990 553559 9990 553631
rect 21383 553602 21419 553636
rect 15840 553510 15870 553580
rect 15878 553546 15908 553580
rect 21383 553568 21403 553602
rect 21407 553568 21415 553602
rect 15853 553508 15870 553510
rect 21383 553534 21419 553568
rect 21481 553542 22881 553670
rect 23617 553542 25017 553670
rect 25101 553636 25121 553670
rect 25125 553636 25143 553670
rect 25725 553649 26325 553699
rect 25101 553602 25147 553636
rect 25101 553568 25121 553602
rect 25125 553568 25143 553602
rect 25101 553534 25147 553568
rect 5981 553483 6021 553493
rect 5137 553469 6021 553483
rect 21383 553500 21403 553534
rect 21407 553500 21415 553534
rect 21383 553466 21419 553500
rect 7389 553369 8389 553463
rect 7389 553359 8413 553369
rect 8990 553359 9990 553463
rect 21383 553432 21403 553466
rect 21407 553432 21415 553466
rect 21383 553398 21419 553432
rect 21383 553364 21403 553398
rect 21407 553364 21415 553398
rect 21481 553379 22881 553507
rect 23617 553379 25017 553507
rect 25101 553500 25121 553534
rect 25125 553500 25143 553534
rect 25101 553466 25147 553500
rect 25725 553499 26325 553549
rect 25101 553432 25121 553466
rect 25125 553432 25143 553466
rect 25101 553398 25147 553432
rect 25101 553364 25121 553398
rect 25125 553364 25143 553398
rect 25725 553377 26325 553427
rect 21383 553330 21419 553364
rect 25101 553330 25147 553364
rect 21383 553296 21403 553330
rect 21407 553296 21415 553330
rect 25101 553296 25121 553330
rect 25125 553296 25143 553330
rect 21383 553262 21419 553296
rect 21383 553228 21403 553262
rect 21407 553228 21415 553262
rect 21481 553229 22881 553272
rect 23617 553229 25017 553272
rect 25101 553262 25147 553296
rect 25101 553228 25121 553262
rect 25125 553228 25143 553262
rect 21383 553194 21419 553228
rect 25101 553194 25147 553228
rect 25725 553227 26325 553277
rect 21383 553160 21403 553194
rect 21407 553160 21415 553194
rect 25101 553160 25121 553194
rect 25125 553160 25143 553194
rect 27162 553170 27212 554170
rect 27312 553170 27440 554060
rect 27468 553170 27596 554060
rect 27624 553170 27752 554060
rect 27780 553170 27908 554060
rect 27936 553170 28064 554060
rect 28092 553170 28220 554060
rect 28248 553170 28376 554060
rect 28404 553170 28532 554060
rect 28560 553170 28688 554060
rect 28716 553170 28844 554060
rect 28872 553170 29000 554060
rect 29028 553170 29156 554060
rect 29184 553170 29312 554060
rect 29340 553170 29390 554170
rect 30245 554029 30445 554209
rect 30245 554018 30260 554029
rect 30245 554014 30257 554018
rect 30430 554014 30445 554029
rect 30543 554029 30580 554209
rect 678680 554151 678704 554185
rect 680215 554178 680815 554228
rect 681745 554209 682345 554259
rect 678680 554083 678704 554117
rect 30543 554014 30558 554029
rect 678680 554015 678704 554049
rect 680215 554002 680815 554058
rect 681745 554053 682345 554181
rect 682509 554030 683109 554080
rect 30245 553984 30257 553988
rect 30245 553973 30260 553984
rect 30430 553973 30445 553988
rect 30245 553793 30445 553973
rect 678680 553947 678704 553981
rect 678680 553879 678704 553913
rect 681745 553897 682345 553953
rect 31453 553818 32053 553868
rect 678680 553811 678704 553845
rect 680215 553826 680815 553882
rect 30245 553782 30260 553793
rect 30245 553778 30257 553782
rect 30430 553778 30445 553793
rect 678680 553743 678704 553777
rect 681745 553741 682345 553869
rect 682509 553854 683109 553910
rect 31453 553648 32053 553698
rect 678680 553675 678704 553709
rect 680215 553656 680815 553706
rect 682509 553684 683109 553734
rect 683248 553680 683298 554268
rect 683398 553680 683448 554268
rect 684519 554158 685119 554286
rect 685551 554282 686551 554410
rect 686865 554300 687465 554428
rect 684519 554002 685119 554130
rect 685551 554126 686551 554254
rect 686865 554124 687465 554252
rect 685551 553970 686551 554098
rect 686865 553954 687465 554004
rect 684519 553852 685119 553902
rect 685551 553814 686551 553870
rect 686865 553838 687465 553888
rect 683248 553668 683448 553680
rect 685551 553658 686551 553786
rect 686865 553662 687465 553790
rect 678680 553607 678704 553641
rect 681745 553591 682345 553641
rect 683571 553605 683581 553646
rect 678680 553539 678704 553573
rect 680215 553524 680815 553574
rect 682509 553555 683509 553605
rect 30245 553472 30845 553522
rect 678680 553471 678704 553505
rect 685551 553502 686551 553630
rect 686865 553486 687465 553542
rect 678680 553403 678704 553437
rect 30245 553296 30845 553352
rect 678680 553335 678704 553369
rect 680215 553348 680815 553404
rect 681745 553389 682345 553439
rect 682509 553385 683509 553435
rect 683278 553382 683398 553385
rect 683571 553382 683581 553385
rect 685551 553346 686551 553474
rect 678680 553267 678704 553301
rect 678680 553199 678704 553233
rect 21383 553126 21419 553160
rect 25101 553126 25147 553160
rect 21383 553102 21403 553126
rect 21385 553048 21403 553102
rect 21407 553082 21415 553126
rect 25101 553102 25121 553126
rect 25113 553082 25121 553102
rect 25125 553048 25143 553126
rect 30245 553120 30845 553176
rect 680215 553172 680815 553228
rect 681745 553213 682345 553341
rect 682509 553247 683109 553297
rect 678680 553131 678704 553165
rect 678680 553063 678704 553097
rect 678654 553013 678680 553039
rect 680215 553002 680815 553052
rect 681745 553037 682345 553093
rect 682509 553071 683109 553127
rect 30245 552950 30845 553000
rect 678680 552929 678704 552963
rect 21000 552800 21003 552920
rect 21352 552885 21376 552909
rect 25122 552885 25146 552909
rect 21385 552861 21400 552885
rect 25098 552861 25113 552885
rect 678680 552861 678704 552895
rect 21274 552783 21294 552851
rect 21410 552817 21430 552851
rect 25068 552817 25088 552851
rect 25204 552817 25224 552851
rect 21385 552807 21430 552817
rect 25102 552807 25137 552817
rect 21361 552783 21430 552807
rect 25089 552783 25137 552807
rect 25238 552783 25258 552817
rect 678680 552793 678704 552827
rect 679007 552826 679607 552876
rect 681745 552867 682345 552917
rect 682509 552901 683109 552951
rect 678680 552725 678704 552759
rect 680615 552731 680630 552746
rect 680803 552742 680815 552746
rect 680800 552731 680815 552742
rect 678680 552657 678704 552691
rect 679007 552656 679607 552706
rect 678680 552589 678704 552623
rect 678680 552521 678704 552555
rect 680615 552551 680815 552731
rect 681345 552651 682345 552701
rect 682508 552631 683108 552681
rect 680615 552536 680630 552551
rect 680800 552540 680815 552551
rect 680803 552536 680815 552540
rect 680502 552495 680517 552510
rect 678680 552453 678704 552487
rect 678680 552385 678704 552419
rect 678680 552317 678704 552351
rect 680480 552315 680517 552495
rect 680502 552300 680517 552315
rect 680615 552495 680630 552510
rect 680803 552506 680815 552510
rect 680800 552495 680815 552506
rect 680615 552315 680815 552495
rect 681345 552475 682345 552531
rect 682508 552455 683108 552511
rect 680615 552300 680630 552315
rect 680800 552304 680815 552315
rect 680803 552300 680815 552304
rect 681345 552299 682345 552427
rect 682508 552285 683108 552335
rect 683228 552322 683278 553322
rect 683398 552322 683448 553322
rect 685551 553190 686551 553318
rect 686865 553310 687465 553438
rect 685551 553034 686551 553162
rect 686865 553140 687465 553190
rect 686865 553024 687465 553074
rect 685551 552884 686551 552934
rect 686865 552848 687465 552976
rect 685551 552768 686551 552818
rect 686865 552672 687465 552800
rect 684404 552609 685004 552659
rect 685551 552612 686551 552668
rect 685551 552456 686551 552512
rect 686865 552496 687465 552624
rect 685551 552300 686551 552356
rect 686865 552320 687465 552376
rect 678680 552249 678704 552283
rect 679002 552230 679602 552280
rect 678680 552181 678704 552215
rect 678680 552113 678704 552147
rect 681345 552129 682345 552179
rect 684404 552175 685004 552225
rect 685551 552150 686551 552200
rect 686865 552150 687465 552200
rect 678680 552045 678704 552079
rect 679002 552054 679602 552110
rect 681390 552070 681424 552080
rect 681458 552070 681492 552080
rect 681526 552070 681560 552080
rect 681594 552070 681628 552080
rect 681662 552070 681696 552080
rect 681730 552070 681764 552080
rect 681798 552070 681832 552080
rect 681866 552070 681900 552080
rect 681934 552070 681968 552080
rect 682002 552070 682036 552080
rect 682077 552070 682111 552080
rect 682145 552070 682179 552080
rect 682213 552070 682247 552080
rect 682281 552070 682315 552080
rect 681345 552034 682345 552046
rect 678680 551977 678704 552011
rect 678680 551909 678704 551943
rect 679002 551884 679602 551934
rect 681345 551927 682345 551977
rect 684004 551973 685004 552023
rect 685551 552014 686551 552064
rect 686865 552034 687465 552084
rect 679061 551881 679355 551884
rect 679380 551881 679602 551884
rect 678680 551841 678704 551875
rect 678680 551773 678704 551807
rect 681345 551751 682345 551879
rect 684004 551817 685004 551873
rect 685551 551858 686551 551914
rect 686865 551858 687465 551914
rect 686686 551812 686714 551840
rect 678680 551705 678704 551739
rect 678680 551637 678704 551671
rect 678680 551569 678704 551603
rect 681345 551575 682345 551703
rect 684004 551661 685004 551789
rect 685551 551708 686551 551758
rect 686865 551688 687465 551738
rect 678680 551501 678704 551535
rect 684004 551505 685004 551633
rect 687573 551554 687585 557277
rect 689154 557107 689204 557355
rect 689151 557023 689204 557107
rect 689154 556897 689204 557023
rect 689304 556897 689360 557897
rect 689460 556897 689516 557897
rect 689616 556897 689672 557897
rect 689772 556897 689828 557897
rect 689928 556897 689978 557897
rect 692485 557872 692521 557906
rect 692485 557838 692505 557872
rect 692509 557838 692517 557872
rect 690952 557509 691122 557815
rect 692485 557804 692521 557838
rect 692485 557770 692505 557804
rect 692509 557770 692517 557804
rect 692583 557775 693983 557903
rect 694719 557775 696119 557903
rect 696203 557872 696249 557906
rect 696203 557838 696223 557872
rect 696227 557838 696245 557872
rect 699322 557860 700322 557916
rect 700922 557860 701922 557916
rect 707610 557905 708610 557961
rect 709211 557905 710211 557961
rect 696203 557804 696249 557838
rect 696203 557770 696223 557804
rect 696227 557770 696245 557804
rect 699322 557788 700322 557844
rect 700922 557788 701922 557844
rect 707610 557833 708610 557889
rect 709211 557833 710211 557889
rect 692485 557736 692521 557770
rect 692485 557702 692505 557736
rect 692509 557702 692517 557736
rect 692485 557668 692521 557702
rect 692485 557634 692505 557668
rect 692509 557634 692517 557668
rect 692485 557600 692521 557634
rect 692583 557612 693983 557740
rect 694719 557612 696119 557740
rect 696203 557736 696249 557770
rect 696203 557702 696223 557736
rect 696227 557702 696245 557736
rect 696203 557668 696249 557702
rect 696203 557634 696223 557668
rect 696227 557634 696245 557668
rect 696203 557600 696249 557634
rect 692485 557566 692505 557600
rect 692509 557566 692517 557600
rect 692485 557532 692521 557566
rect 692485 557498 692505 557532
rect 692509 557498 692517 557532
rect 692485 557464 692521 557498
rect 692485 557430 692505 557464
rect 692509 557430 692517 557464
rect 692583 557449 693983 557577
rect 694719 557449 696119 557577
rect 696203 557566 696223 557600
rect 696227 557566 696245 557600
rect 696203 557532 696249 557566
rect 696203 557498 696223 557532
rect 696227 557498 696245 557532
rect 696203 557464 696249 557498
rect 699322 557486 700322 557558
rect 700922 557486 701922 557558
rect 707610 557531 708610 557603
rect 709211 557531 710211 557603
rect 711579 557553 711605 559307
rect 715956 558297 716006 559297
rect 716106 558297 716234 559297
rect 716262 558297 716312 559297
rect 699392 557475 699426 557486
rect 699460 557475 699494 557486
rect 699528 557475 699562 557486
rect 699596 557475 699630 557486
rect 699664 557475 699698 557486
rect 699732 557475 699766 557486
rect 699800 557475 699834 557486
rect 699868 557475 699902 557486
rect 699936 557475 699970 557486
rect 700004 557475 700038 557486
rect 700072 557475 700106 557486
rect 700140 557475 700174 557486
rect 700208 557475 700242 557486
rect 700276 557475 700310 557486
rect 700934 557475 700968 557486
rect 701002 557475 701036 557486
rect 701070 557475 701104 557486
rect 701138 557475 701172 557486
rect 701206 557475 701240 557486
rect 701274 557475 701308 557486
rect 701342 557475 701376 557486
rect 701410 557475 701444 557486
rect 701478 557475 701512 557486
rect 701546 557475 701580 557486
rect 701614 557475 701648 557486
rect 701682 557475 701716 557486
rect 701750 557475 701784 557486
rect 701818 557475 701852 557486
rect 711511 557485 711663 557553
rect 712447 557501 712557 557511
rect 711579 557482 711663 557485
rect 699392 557465 699450 557475
rect 699460 557465 699518 557475
rect 699528 557465 699586 557475
rect 699596 557465 699654 557475
rect 699664 557465 699722 557475
rect 699732 557465 699790 557475
rect 699800 557465 699858 557475
rect 699868 557465 699926 557475
rect 699936 557465 699994 557475
rect 700004 557465 700062 557475
rect 700072 557465 700130 557475
rect 700140 557465 700198 557475
rect 700208 557465 700266 557475
rect 700276 557465 700334 557475
rect 700934 557465 700992 557475
rect 701002 557465 701060 557475
rect 701070 557465 701128 557475
rect 701138 557465 701196 557475
rect 701206 557465 701264 557475
rect 701274 557465 701332 557475
rect 701342 557465 701400 557475
rect 701410 557465 701468 557475
rect 701478 557465 701536 557475
rect 701546 557465 701604 557475
rect 701614 557465 701672 557475
rect 701682 557465 701740 557475
rect 701750 557465 701808 557475
rect 701818 557465 701876 557475
rect 696203 557430 696223 557464
rect 696227 557430 696245 557464
rect 699368 557441 700334 557465
rect 700910 557441 701876 557465
rect 711541 557461 711633 557482
rect 692485 557396 692521 557430
rect 692485 557362 692505 557396
rect 692509 557362 692517 557396
rect 692485 557328 692521 557362
rect 692485 557294 692505 557328
rect 692509 557294 692517 557328
rect 692485 557260 692521 557294
rect 692583 557286 693983 557414
rect 694719 557286 696119 557414
rect 696203 557396 696249 557430
rect 699392 557426 699416 557441
rect 699460 557426 699484 557441
rect 699528 557426 699552 557441
rect 699596 557426 699620 557441
rect 699664 557426 699688 557441
rect 699732 557426 699756 557441
rect 699800 557426 699824 557441
rect 699868 557426 699892 557441
rect 699936 557426 699960 557441
rect 700004 557426 700028 557441
rect 700072 557426 700096 557441
rect 700140 557426 700164 557441
rect 700208 557426 700232 557441
rect 700276 557426 700300 557441
rect 700934 557426 700958 557441
rect 701002 557426 701026 557441
rect 701070 557426 701094 557441
rect 701138 557426 701162 557441
rect 701206 557426 701230 557441
rect 701274 557426 701298 557441
rect 701342 557426 701366 557441
rect 701410 557426 701434 557441
rect 701478 557426 701502 557441
rect 701546 557426 701570 557441
rect 701614 557426 701638 557441
rect 701682 557426 701706 557441
rect 701750 557426 701774 557441
rect 701818 557426 701842 557441
rect 696203 557362 696223 557396
rect 696227 557362 696245 557396
rect 696203 557328 696249 557362
rect 696203 557294 696223 557328
rect 696227 557294 696245 557328
rect 696203 557260 696249 557294
rect 699322 557271 700322 557426
rect 692485 557226 692505 557260
rect 692509 557226 692517 557260
rect 692485 557192 692521 557226
rect 692485 557158 692505 557192
rect 692509 557158 692517 557192
rect 692485 557124 692521 557158
rect 692485 557090 692505 557124
rect 692509 557090 692517 557124
rect 692583 557123 693983 557251
rect 694719 557123 696119 557251
rect 696203 557226 696223 557260
rect 696227 557226 696245 557260
rect 699322 557237 700334 557271
rect 700922 557261 701922 557426
rect 707610 557271 708610 557331
rect 709211 557271 710211 557331
rect 700910 557237 701922 557261
rect 699322 557226 700322 557237
rect 700922 557226 701922 557237
rect 696203 557192 696249 557226
rect 699392 557213 699416 557226
rect 699460 557213 699484 557226
rect 699528 557213 699552 557226
rect 699596 557213 699620 557226
rect 699664 557213 699688 557226
rect 699732 557213 699756 557226
rect 699800 557213 699824 557226
rect 699868 557213 699892 557226
rect 699936 557213 699960 557226
rect 700004 557213 700028 557226
rect 700072 557213 700096 557226
rect 700140 557213 700164 557226
rect 700208 557213 700232 557226
rect 700276 557213 700300 557226
rect 700934 557213 700958 557226
rect 701002 557213 701026 557226
rect 701070 557213 701094 557226
rect 701138 557213 701162 557226
rect 701206 557213 701230 557226
rect 701274 557213 701298 557226
rect 701342 557213 701366 557226
rect 701410 557213 701434 557226
rect 701478 557213 701502 557226
rect 701546 557213 701570 557226
rect 701614 557213 701638 557226
rect 701682 557213 701706 557226
rect 701750 557213 701774 557226
rect 701818 557213 701842 557226
rect 696203 557158 696223 557192
rect 696227 557158 696245 557192
rect 696203 557124 696249 557158
rect 696203 557090 696223 557124
rect 696227 557090 696245 557124
rect 692485 557056 692521 557090
rect 696203 557056 696249 557090
rect 692485 557022 692505 557056
rect 692509 557022 692517 557056
rect 696203 557022 696223 557056
rect 696227 557022 696245 557056
rect 692485 556988 692521 557022
rect 692485 556954 692505 556988
rect 692509 556954 692517 556988
rect 692583 556966 693983 557016
rect 694719 556966 696119 557016
rect 696203 556988 696249 557022
rect 696203 556954 696223 556988
rect 696227 556954 696245 556988
rect 692485 556920 692521 556954
rect 696203 556920 696249 556954
rect 692485 556896 692505 556920
rect 692487 556852 692505 556896
rect 692509 556886 692517 556920
rect 696203 556896 696223 556920
rect 696215 556886 696223 556896
rect 696227 556852 696245 556920
rect 697284 556870 697350 556886
rect 699322 556868 700322 556924
rect 700922 556868 701922 556924
rect 707610 556913 708610 556969
rect 709211 556913 710211 556969
rect 692174 556787 692186 556811
rect 692288 556787 692312 556811
rect 696390 556787 696414 556811
rect 696516 556787 696528 556811
rect 699322 556796 700322 556852
rect 700922 556796 701922 556852
rect 707610 556841 708610 556897
rect 709211 556841 710211 556897
rect 692264 556763 692288 556777
rect 696414 556763 696438 556777
rect 692288 556729 692312 556753
rect 696390 556729 696414 556753
rect 688940 556475 688990 556675
rect 689110 556475 689238 556675
rect 689286 556475 689342 556675
rect 689462 556475 689590 556675
rect 689638 556559 689688 556675
rect 692736 556597 695966 556699
rect 689638 556475 689691 556559
rect 699322 556494 700322 556566
rect 700922 556494 701922 556566
rect 707610 556539 708610 556611
rect 709211 556539 710211 556611
rect 699392 556483 699426 556494
rect 699460 556483 699494 556494
rect 699528 556483 699562 556494
rect 699596 556483 699630 556494
rect 699664 556483 699698 556494
rect 699732 556483 699766 556494
rect 699800 556483 699834 556494
rect 699868 556483 699902 556494
rect 699936 556483 699970 556494
rect 700004 556483 700038 556494
rect 700072 556483 700106 556494
rect 700140 556483 700174 556494
rect 700208 556483 700242 556494
rect 700276 556483 700310 556494
rect 700934 556483 700968 556494
rect 701002 556483 701036 556494
rect 701070 556483 701104 556494
rect 701138 556483 701172 556494
rect 701206 556483 701240 556494
rect 701274 556483 701308 556494
rect 701342 556483 701376 556494
rect 701410 556483 701444 556494
rect 701478 556483 701512 556494
rect 701546 556483 701580 556494
rect 701614 556483 701648 556494
rect 701682 556483 701716 556494
rect 701750 556483 701784 556494
rect 701818 556483 701852 556494
rect 689649 556471 689683 556475
rect 699392 556473 699450 556483
rect 699460 556473 699518 556483
rect 699528 556473 699586 556483
rect 699596 556473 699654 556483
rect 699664 556473 699722 556483
rect 699732 556473 699790 556483
rect 699800 556473 699858 556483
rect 699868 556473 699926 556483
rect 699936 556473 699994 556483
rect 700004 556473 700062 556483
rect 700072 556473 700130 556483
rect 700140 556473 700198 556483
rect 700208 556473 700266 556483
rect 700276 556473 700334 556483
rect 700934 556473 700992 556483
rect 701002 556473 701060 556483
rect 701070 556473 701128 556483
rect 701138 556473 701196 556483
rect 701206 556473 701264 556483
rect 701274 556473 701332 556483
rect 701342 556473 701400 556483
rect 701410 556473 701468 556483
rect 701478 556473 701536 556483
rect 701546 556473 701604 556483
rect 701614 556473 701672 556483
rect 701682 556473 701740 556483
rect 701750 556473 701808 556483
rect 701818 556473 701876 556483
rect 692451 556444 692475 556468
rect 692509 556444 692533 556468
rect 696169 556444 696193 556468
rect 696227 556444 696251 556468
rect 699368 556449 700334 556473
rect 700910 556449 701876 556473
rect 692485 556410 692499 556444
rect 696203 556410 696217 556444
rect 699392 556434 699416 556449
rect 699460 556434 699484 556449
rect 699528 556434 699552 556449
rect 699596 556434 699620 556449
rect 699664 556434 699688 556449
rect 699732 556434 699756 556449
rect 699800 556434 699824 556449
rect 699868 556434 699892 556449
rect 699936 556434 699960 556449
rect 700004 556434 700028 556449
rect 700072 556434 700096 556449
rect 700140 556434 700164 556449
rect 700208 556434 700232 556449
rect 700276 556434 700300 556449
rect 700934 556434 700958 556449
rect 701002 556434 701026 556449
rect 701070 556434 701094 556449
rect 701138 556434 701162 556449
rect 701206 556434 701230 556449
rect 701274 556434 701298 556449
rect 701342 556434 701366 556449
rect 701410 556434 701434 556449
rect 701478 556434 701502 556449
rect 701546 556434 701570 556449
rect 701614 556434 701638 556449
rect 701682 556434 701706 556449
rect 701750 556434 701774 556449
rect 701818 556434 701842 556449
rect 692451 556386 692475 556410
rect 692509 556386 692533 556410
rect 696169 556386 696193 556410
rect 696227 556386 696251 556410
rect 690664 556318 691664 556368
rect 692515 556280 693915 556330
rect 694787 556280 696187 556330
rect 699322 556279 700322 556434
rect 699322 556245 700334 556279
rect 700922 556269 701922 556434
rect 703539 556286 703699 556290
rect 707610 556279 708610 556339
rect 709211 556279 710211 556339
rect 700910 556245 701922 556269
rect 690242 556219 690326 556222
rect 690242 556214 690442 556219
rect 690238 556180 690442 556214
rect 690242 556169 690442 556180
rect 690664 556162 691664 556218
rect 687686 556128 687720 556162
rect 687686 556104 687710 556128
rect 689649 556127 689683 556131
rect 688940 555927 688990 556127
rect 689110 555927 689238 556127
rect 689286 555927 689342 556127
rect 689462 555927 689590 556127
rect 689638 556043 689691 556127
rect 689638 555927 689688 556043
rect 690242 555993 690442 556121
rect 692515 556117 693915 556245
rect 694787 556117 696187 556245
rect 699322 556234 700322 556245
rect 700922 556234 701922 556245
rect 699392 556221 699416 556234
rect 699460 556221 699484 556234
rect 699528 556221 699552 556234
rect 699596 556221 699620 556234
rect 699664 556221 699688 556234
rect 699732 556221 699756 556234
rect 699800 556221 699824 556234
rect 699868 556221 699892 556234
rect 699936 556221 699960 556234
rect 700004 556221 700028 556234
rect 700072 556221 700096 556234
rect 700140 556221 700164 556234
rect 700208 556221 700232 556234
rect 700276 556221 700300 556234
rect 700934 556221 700958 556234
rect 701002 556221 701026 556234
rect 701070 556221 701094 556234
rect 701138 556221 701162 556234
rect 701206 556221 701230 556234
rect 701274 556221 701298 556234
rect 701342 556221 701366 556234
rect 701410 556221 701434 556234
rect 701478 556221 701502 556234
rect 701546 556221 701570 556234
rect 701614 556221 701638 556234
rect 701682 556221 701706 556234
rect 701750 556221 701774 556234
rect 701818 556221 701842 556234
rect 703541 556140 703701 556144
rect 690664 556006 691664 556062
rect 692515 555954 693915 556082
rect 694787 555954 696187 556082
rect 690242 555817 690442 555873
rect 690664 555850 691664 555906
rect 692515 555791 693915 555919
rect 694787 555791 696187 555919
rect 699322 555876 700322 555932
rect 700922 555876 701922 555932
rect 707610 555921 708610 555977
rect 709211 555921 710211 555977
rect 699322 555804 700322 555860
rect 700922 555804 701922 555860
rect 707610 555849 708610 555905
rect 709211 555849 710211 555905
rect 689154 555579 689204 555705
rect 687686 555501 687720 555535
rect 687798 555515 687822 555539
rect 687774 555491 687798 555504
rect 689151 555495 689204 555579
rect 687798 555456 687822 555480
rect 689154 555247 689204 555495
rect 689151 555163 689204 555247
rect 689154 554705 689204 555163
rect 689304 554705 689360 555705
rect 689460 554705 689516 555705
rect 689616 554705 689672 555705
rect 689772 554705 689828 555705
rect 689928 554705 689978 555705
rect 690242 555641 690442 555769
rect 690664 555700 691664 555750
rect 690790 555697 690874 555700
rect 691123 555697 691207 555700
rect 692515 555628 693915 555756
rect 694787 555628 696187 555756
rect 704735 555731 705041 555833
rect 704719 555715 705057 555731
rect 690242 555465 690442 555521
rect 692515 555465 693915 555593
rect 694787 555465 696187 555593
rect 699322 555502 700322 555574
rect 700922 555502 701922 555574
rect 707610 555547 708610 555619
rect 709211 555547 710211 555619
rect 699392 555491 699426 555502
rect 699460 555491 699494 555502
rect 699528 555491 699562 555502
rect 699596 555491 699630 555502
rect 699664 555491 699698 555502
rect 699732 555491 699766 555502
rect 699800 555491 699834 555502
rect 699868 555491 699902 555502
rect 699936 555491 699970 555502
rect 700004 555491 700038 555502
rect 700072 555491 700106 555502
rect 700140 555491 700174 555502
rect 700208 555491 700242 555502
rect 700276 555491 700310 555502
rect 700934 555491 700968 555502
rect 701002 555491 701036 555502
rect 701070 555491 701104 555502
rect 701138 555491 701172 555502
rect 701206 555491 701240 555502
rect 701274 555491 701308 555502
rect 701342 555491 701376 555502
rect 701410 555491 701444 555502
rect 701478 555491 701512 555502
rect 701546 555491 701580 555502
rect 701614 555491 701648 555502
rect 701682 555491 701716 555502
rect 701750 555491 701784 555502
rect 701818 555491 701852 555502
rect 699392 555481 699450 555491
rect 699460 555481 699518 555491
rect 699528 555481 699586 555491
rect 699596 555481 699654 555491
rect 699664 555481 699722 555491
rect 699732 555481 699790 555491
rect 699800 555481 699858 555491
rect 699868 555481 699926 555491
rect 699936 555481 699994 555491
rect 700004 555481 700062 555491
rect 700072 555481 700130 555491
rect 700140 555481 700198 555491
rect 700208 555481 700266 555491
rect 700276 555481 700334 555491
rect 700934 555481 700992 555491
rect 701002 555481 701060 555491
rect 701070 555481 701128 555491
rect 701138 555481 701196 555491
rect 701206 555481 701264 555491
rect 701274 555481 701332 555491
rect 701342 555481 701400 555491
rect 701410 555481 701468 555491
rect 701478 555481 701536 555491
rect 701546 555481 701604 555491
rect 701614 555481 701672 555491
rect 701682 555481 701740 555491
rect 701750 555481 701808 555491
rect 701818 555481 701876 555491
rect 699368 555457 700334 555481
rect 700910 555457 701876 555481
rect 699392 555442 699416 555457
rect 699460 555442 699484 555457
rect 699528 555442 699552 555457
rect 699596 555442 699620 555457
rect 699664 555442 699688 555457
rect 699732 555442 699756 555457
rect 699800 555442 699824 555457
rect 699868 555442 699892 555457
rect 699936 555442 699960 555457
rect 700004 555442 700028 555457
rect 700072 555442 700096 555457
rect 700140 555442 700164 555457
rect 700208 555442 700232 555457
rect 700276 555442 700300 555457
rect 700934 555442 700958 555457
rect 701002 555442 701026 555457
rect 701070 555442 701094 555457
rect 701138 555442 701162 555457
rect 701206 555442 701230 555457
rect 701274 555442 701298 555457
rect 701342 555442 701366 555457
rect 701410 555442 701434 555457
rect 701478 555442 701502 555457
rect 701546 555442 701570 555457
rect 701614 555442 701638 555457
rect 701682 555442 701706 555457
rect 701750 555442 701774 555457
rect 701818 555442 701842 555457
rect 690242 555289 690442 555417
rect 692515 555302 693915 555430
rect 694787 555302 696187 555430
rect 690790 555286 690874 555289
rect 691123 555286 691207 555289
rect 699322 555287 700322 555442
rect 690664 555236 691664 555286
rect 699322 555253 700334 555287
rect 700922 555277 701922 555442
rect 707610 555287 708610 555347
rect 709211 555287 710211 555347
rect 700910 555253 701922 555277
rect 699322 555242 700322 555253
rect 700922 555242 701922 555253
rect 699392 555229 699416 555242
rect 699460 555229 699484 555242
rect 699528 555229 699552 555242
rect 699596 555229 699620 555242
rect 699664 555229 699688 555242
rect 699732 555229 699756 555242
rect 699800 555229 699824 555242
rect 699868 555229 699892 555242
rect 699936 555229 699960 555242
rect 700004 555229 700028 555242
rect 700072 555229 700096 555242
rect 700140 555229 700164 555242
rect 700208 555229 700232 555242
rect 700276 555229 700300 555242
rect 700934 555229 700958 555242
rect 701002 555229 701026 555242
rect 701070 555229 701094 555242
rect 701138 555229 701162 555242
rect 701206 555229 701230 555242
rect 701274 555229 701298 555242
rect 701342 555229 701366 555242
rect 701410 555229 701434 555242
rect 701478 555229 701502 555242
rect 701546 555229 701570 555242
rect 701614 555229 701638 555242
rect 701682 555229 701706 555242
rect 701750 555229 701774 555242
rect 701818 555229 701842 555242
rect 690242 555113 690442 555169
rect 692515 555152 693915 555195
rect 694787 555152 696187 555195
rect 690664 555080 691664 555136
rect 690242 554937 690442 555065
rect 692515 555016 693915 555059
rect 694787 555016 696187 555059
rect 690664 554924 691664 554980
rect 692515 554853 693915 554981
rect 694787 554853 696187 554981
rect 703541 554944 703701 554948
rect 699322 554884 700322 554940
rect 700922 554884 701922 554940
rect 707610 554929 708610 554985
rect 709211 554929 710211 554985
rect 690242 554806 690442 554817
rect 690238 554772 690442 554806
rect 690242 554767 690442 554772
rect 690664 554768 691664 554824
rect 690242 554764 690326 554767
rect 692515 554690 693915 554818
rect 694787 554690 696187 554818
rect 699322 554812 700322 554868
rect 700922 554812 701922 554868
rect 707610 554857 708610 554913
rect 709211 554857 710211 554913
rect 703541 554798 703701 554802
rect 690664 554618 691664 554668
rect 692515 554527 693915 554655
rect 694787 554527 696187 554655
rect 699322 554510 700322 554582
rect 700922 554510 701922 554582
rect 707610 554555 708610 554627
rect 709211 554555 710211 554627
rect 699392 554499 699426 554510
rect 699460 554499 699494 554510
rect 699528 554499 699562 554510
rect 699596 554499 699630 554510
rect 699664 554499 699698 554510
rect 699732 554499 699766 554510
rect 699800 554499 699834 554510
rect 699868 554499 699902 554510
rect 699936 554499 699970 554510
rect 700004 554499 700038 554510
rect 700072 554499 700106 554510
rect 700140 554499 700174 554510
rect 700208 554499 700242 554510
rect 700276 554499 700310 554510
rect 700934 554499 700968 554510
rect 701002 554499 701036 554510
rect 701070 554499 701104 554510
rect 701138 554499 701172 554510
rect 701206 554499 701240 554510
rect 701274 554499 701308 554510
rect 701342 554499 701376 554510
rect 701410 554499 701444 554510
rect 701478 554499 701512 554510
rect 701546 554499 701580 554510
rect 701614 554499 701648 554510
rect 701682 554499 701716 554510
rect 701750 554499 701784 554510
rect 701818 554499 701852 554510
rect 692515 554364 693915 554492
rect 694787 554364 696187 554492
rect 699392 554489 699450 554499
rect 699460 554489 699518 554499
rect 699528 554489 699586 554499
rect 699596 554489 699654 554499
rect 699664 554489 699722 554499
rect 699732 554489 699790 554499
rect 699800 554489 699858 554499
rect 699868 554489 699926 554499
rect 699936 554489 699994 554499
rect 700004 554489 700062 554499
rect 700072 554489 700130 554499
rect 700140 554489 700198 554499
rect 700208 554489 700266 554499
rect 700276 554489 700334 554499
rect 700934 554489 700992 554499
rect 701002 554489 701060 554499
rect 701070 554489 701128 554499
rect 701138 554489 701196 554499
rect 701206 554489 701264 554499
rect 701274 554489 701332 554499
rect 701342 554489 701400 554499
rect 701410 554489 701468 554499
rect 701478 554489 701536 554499
rect 701546 554489 701604 554499
rect 701614 554489 701672 554499
rect 701682 554489 701740 554499
rect 701750 554489 701808 554499
rect 701818 554489 701876 554499
rect 699368 554465 700334 554489
rect 700910 554465 701876 554489
rect 699392 554450 699416 554465
rect 699460 554450 699484 554465
rect 699528 554450 699552 554465
rect 699596 554450 699620 554465
rect 699664 554450 699688 554465
rect 699732 554450 699756 554465
rect 699800 554450 699824 554465
rect 699868 554450 699892 554465
rect 699936 554450 699960 554465
rect 700004 554450 700028 554465
rect 700072 554450 700096 554465
rect 700140 554450 700164 554465
rect 700208 554450 700232 554465
rect 700276 554450 700300 554465
rect 700934 554450 700958 554465
rect 701002 554450 701026 554465
rect 701070 554450 701094 554465
rect 701138 554450 701162 554465
rect 701206 554450 701230 554465
rect 701274 554450 701298 554465
rect 701342 554450 701366 554465
rect 701410 554450 701434 554465
rect 701478 554450 701502 554465
rect 701546 554450 701570 554465
rect 701614 554450 701638 554465
rect 701682 554450 701706 554465
rect 701750 554450 701774 554465
rect 701818 554450 701842 554465
rect 692515 554201 693915 554329
rect 694787 554201 696187 554329
rect 699322 554295 700322 554450
rect 699322 554261 700334 554295
rect 700922 554285 701922 554450
rect 707610 554295 708610 554355
rect 709211 554295 710211 554355
rect 700910 554261 701922 554285
rect 699322 554250 700322 554261
rect 700922 554250 701922 554261
rect 699392 554237 699416 554250
rect 699460 554237 699484 554250
rect 699528 554237 699552 554250
rect 699596 554237 699620 554250
rect 699664 554237 699688 554250
rect 699732 554237 699756 554250
rect 699800 554237 699824 554250
rect 699868 554237 699892 554250
rect 699936 554237 699960 554250
rect 700004 554237 700028 554250
rect 700072 554237 700096 554250
rect 700140 554237 700164 554250
rect 700208 554237 700232 554250
rect 700276 554237 700300 554250
rect 700934 554237 700958 554250
rect 701002 554237 701026 554250
rect 701070 554237 701094 554250
rect 701138 554237 701162 554250
rect 701206 554237 701230 554250
rect 701274 554237 701298 554250
rect 701342 554237 701366 554250
rect 701410 554237 701434 554250
rect 701478 554237 701502 554250
rect 701546 554237 701570 554250
rect 701614 554237 701638 554250
rect 701682 554237 701706 554250
rect 701750 554237 701774 554250
rect 701818 554237 701842 554250
rect 692515 554038 693915 554166
rect 694787 554038 696187 554166
rect 692047 553468 696655 554004
rect 699322 553892 700322 553948
rect 700922 553892 701922 553948
rect 707610 553937 708610 553993
rect 709211 553937 710211 553993
rect 699322 553820 700322 553876
rect 700922 553820 701922 553876
rect 707610 553865 708610 553921
rect 709211 553865 710211 553921
rect 697314 553582 697620 553752
rect 699322 553518 700322 553590
rect 700922 553518 701922 553590
rect 707610 553563 708610 553635
rect 709211 553563 710211 553635
rect 704719 553527 705057 553543
rect 699392 553507 699426 553518
rect 699460 553507 699494 553518
rect 699528 553507 699562 553518
rect 699596 553507 699630 553518
rect 699664 553507 699698 553518
rect 699732 553507 699766 553518
rect 699800 553507 699834 553518
rect 699868 553507 699902 553518
rect 699936 553507 699970 553518
rect 700004 553507 700038 553518
rect 700072 553507 700106 553518
rect 700140 553507 700174 553518
rect 700208 553507 700242 553518
rect 700276 553507 700310 553518
rect 700934 553507 700968 553518
rect 701002 553507 701036 553518
rect 701070 553507 701104 553518
rect 701138 553507 701172 553518
rect 701206 553507 701240 553518
rect 701274 553507 701308 553518
rect 701342 553507 701376 553518
rect 701410 553507 701444 553518
rect 701478 553507 701512 553518
rect 701546 553507 701580 553518
rect 701614 553507 701648 553518
rect 701682 553507 701716 553518
rect 701750 553507 701784 553518
rect 701818 553507 701852 553518
rect 699392 553497 699450 553507
rect 699460 553497 699518 553507
rect 699528 553497 699586 553507
rect 699596 553497 699654 553507
rect 699664 553497 699722 553507
rect 699732 553497 699790 553507
rect 699800 553497 699858 553507
rect 699868 553497 699926 553507
rect 699936 553497 699994 553507
rect 700004 553497 700062 553507
rect 700072 553497 700130 553507
rect 700140 553497 700198 553507
rect 700208 553497 700266 553507
rect 700276 553497 700334 553507
rect 700934 553497 700992 553507
rect 701002 553497 701060 553507
rect 701070 553497 701128 553507
rect 701138 553497 701196 553507
rect 701206 553497 701264 553507
rect 701274 553497 701332 553507
rect 701342 553497 701400 553507
rect 701410 553497 701468 553507
rect 701478 553497 701536 553507
rect 701546 553497 701604 553507
rect 701614 553497 701672 553507
rect 701682 553497 701740 553507
rect 701750 553497 701808 553507
rect 701818 553497 701876 553507
rect 699368 553473 700334 553497
rect 700910 553473 701876 553497
rect 699392 553458 699416 553473
rect 699460 553458 699484 553473
rect 699528 553458 699552 553473
rect 699596 553458 699620 553473
rect 699664 553458 699688 553473
rect 699732 553458 699756 553473
rect 699800 553458 699824 553473
rect 699868 553458 699892 553473
rect 699936 553458 699960 553473
rect 700004 553458 700028 553473
rect 700072 553458 700096 553473
rect 700140 553458 700164 553473
rect 700208 553458 700232 553473
rect 700276 553458 700300 553473
rect 700934 553458 700958 553473
rect 701002 553458 701026 553473
rect 701070 553458 701094 553473
rect 701138 553458 701162 553473
rect 701206 553458 701230 553473
rect 701274 553458 701298 553473
rect 701342 553458 701366 553473
rect 701410 553458 701434 553473
rect 701478 553458 701502 553473
rect 701546 553458 701570 553473
rect 701614 553458 701638 553473
rect 701682 553458 701706 553473
rect 701750 553458 701774 553473
rect 701818 553458 701842 553473
rect 699322 553303 700322 553458
rect 692463 553268 692511 553292
rect 696191 553268 696239 553292
rect 692487 553214 692511 553268
rect 696215 553214 696239 553268
rect 699322 553269 700334 553303
rect 700922 553293 701922 553458
rect 704735 553425 705041 553527
rect 707610 553303 708610 553363
rect 709211 553303 710211 553363
rect 700910 553269 701922 553293
rect 699322 553258 700322 553269
rect 700922 553258 701922 553269
rect 699392 553245 699416 553258
rect 699460 553245 699484 553258
rect 699528 553245 699552 553258
rect 699596 553245 699620 553258
rect 699664 553245 699688 553258
rect 699732 553245 699756 553258
rect 699800 553245 699824 553258
rect 699868 553245 699892 553258
rect 699936 553245 699960 553258
rect 700004 553245 700028 553258
rect 700072 553245 700096 553258
rect 700140 553245 700164 553258
rect 700208 553245 700232 553258
rect 700276 553245 700300 553258
rect 700934 553245 700958 553258
rect 701002 553245 701026 553258
rect 701070 553245 701094 553258
rect 701138 553245 701162 553258
rect 701206 553245 701230 553258
rect 701274 553245 701298 553258
rect 701342 553245 701366 553258
rect 701410 553245 701434 553258
rect 701478 553245 701502 553258
rect 701546 553245 701570 553258
rect 701614 553245 701638 553258
rect 701682 553245 701706 553258
rect 701750 553245 701774 553258
rect 701818 553245 701842 553258
rect 692463 553190 692511 553214
rect 696191 553190 696239 553214
rect 687686 553119 687720 553153
rect 687798 553141 687822 553165
rect 687686 553095 687710 553119
rect 687774 553117 687798 553129
rect 687798 553081 687822 553105
rect 692450 553037 692474 553061
rect 692508 553037 692532 553061
rect 696170 553037 696194 553061
rect 696228 553037 696252 553061
rect 692484 553013 692498 553037
rect 696204 553013 696218 553037
rect 692484 552935 692487 552959
rect 696215 552935 696218 552959
rect 692508 552911 692532 552935
rect 696170 552911 696194 552935
rect 699322 552900 700322 552956
rect 700922 552900 701922 552956
rect 707610 552945 708610 553001
rect 709211 552945 710211 553001
rect 692515 552805 693915 552848
rect 694787 552805 696187 552848
rect 699322 552828 700322 552884
rect 700922 552828 701922 552884
rect 707610 552873 708610 552929
rect 709211 552873 710211 552929
rect 692515 552642 693915 552770
rect 694787 552642 696187 552770
rect 688883 552473 688918 552502
rect 692515 552479 693915 552607
rect 694787 552479 696187 552607
rect 699322 552526 700322 552598
rect 700922 552526 701922 552598
rect 707610 552571 708610 552643
rect 709211 552571 710211 552643
rect 699392 552515 699426 552526
rect 699460 552515 699494 552526
rect 699528 552515 699562 552526
rect 699596 552515 699630 552526
rect 699664 552515 699698 552526
rect 699732 552515 699766 552526
rect 699800 552515 699834 552526
rect 699868 552515 699902 552526
rect 699936 552515 699970 552526
rect 700004 552515 700038 552526
rect 700072 552515 700106 552526
rect 700140 552515 700174 552526
rect 700208 552515 700242 552526
rect 700276 552515 700310 552526
rect 700934 552515 700968 552526
rect 701002 552515 701036 552526
rect 701070 552515 701104 552526
rect 701138 552515 701172 552526
rect 701206 552515 701240 552526
rect 701274 552515 701308 552526
rect 701342 552515 701376 552526
rect 701410 552515 701444 552526
rect 701478 552515 701512 552526
rect 701546 552515 701580 552526
rect 701614 552515 701648 552526
rect 701682 552515 701716 552526
rect 701750 552515 701784 552526
rect 701818 552515 701852 552526
rect 699392 552505 699450 552515
rect 699460 552505 699518 552515
rect 699528 552505 699586 552515
rect 699596 552505 699654 552515
rect 699664 552505 699722 552515
rect 699732 552505 699790 552515
rect 699800 552505 699858 552515
rect 699868 552505 699926 552515
rect 699936 552505 699994 552515
rect 700004 552505 700062 552515
rect 700072 552505 700130 552515
rect 700140 552505 700198 552515
rect 700208 552505 700266 552515
rect 700276 552505 700334 552515
rect 700934 552505 700992 552515
rect 701002 552505 701060 552515
rect 701070 552505 701128 552515
rect 701138 552505 701196 552515
rect 701206 552505 701264 552515
rect 701274 552505 701332 552515
rect 701342 552505 701400 552515
rect 701410 552505 701468 552515
rect 701478 552505 701536 552515
rect 701546 552505 701604 552515
rect 701614 552505 701672 552515
rect 701682 552505 701740 552515
rect 701750 552505 701808 552515
rect 701818 552505 701876 552515
rect 699368 552481 700334 552505
rect 700910 552481 701876 552505
rect 688883 552468 688884 552473
rect 688917 552468 688918 552473
rect 688917 552439 688951 552468
rect 699392 552466 699416 552481
rect 699460 552466 699484 552481
rect 699528 552466 699552 552481
rect 699596 552466 699620 552481
rect 699664 552466 699688 552481
rect 699732 552466 699756 552481
rect 699800 552466 699824 552481
rect 699868 552466 699892 552481
rect 699936 552466 699960 552481
rect 700004 552466 700028 552481
rect 700072 552466 700096 552481
rect 700140 552466 700164 552481
rect 700208 552466 700232 552481
rect 700276 552466 700300 552481
rect 700934 552466 700958 552481
rect 701002 552466 701026 552481
rect 701070 552466 701094 552481
rect 701138 552466 701162 552481
rect 701206 552466 701230 552481
rect 701274 552466 701298 552481
rect 701342 552466 701366 552481
rect 701410 552466 701434 552481
rect 701478 552466 701502 552481
rect 701546 552466 701570 552481
rect 701614 552466 701638 552481
rect 701682 552466 701706 552481
rect 701750 552466 701774 552481
rect 701818 552466 701842 552481
rect 688917 552370 688951 552404
rect 688917 552301 688951 552335
rect 692515 552316 693915 552444
rect 694787 552316 696187 552444
rect 699322 552311 700322 552466
rect 688917 552232 688951 552266
rect 688917 552163 688951 552197
rect 692515 552153 693915 552281
rect 694787 552153 696187 552281
rect 699322 552277 700334 552311
rect 700922 552301 701922 552466
rect 707610 552311 708610 552371
rect 709211 552311 710211 552371
rect 700910 552277 701922 552301
rect 699322 552266 700322 552277
rect 700922 552266 701922 552277
rect 699392 552253 699416 552266
rect 699460 552253 699484 552266
rect 699528 552253 699552 552266
rect 699596 552253 699620 552266
rect 699664 552253 699688 552266
rect 699732 552253 699756 552266
rect 699800 552253 699824 552266
rect 699868 552253 699892 552266
rect 699936 552253 699960 552266
rect 700004 552253 700028 552266
rect 700072 552253 700096 552266
rect 700140 552253 700164 552266
rect 700208 552253 700232 552266
rect 700276 552253 700300 552266
rect 700934 552253 700958 552266
rect 701002 552253 701026 552266
rect 701070 552253 701094 552266
rect 701138 552253 701162 552266
rect 701206 552253 701230 552266
rect 701274 552253 701298 552266
rect 701342 552253 701366 552266
rect 701410 552253 701434 552266
rect 701478 552253 701502 552266
rect 701546 552253 701570 552266
rect 701614 552253 701638 552266
rect 701682 552253 701706 552266
rect 701750 552253 701774 552266
rect 701818 552253 701842 552266
rect 688917 552094 688951 552128
rect 688917 552025 688951 552059
rect 692515 551996 693915 552046
rect 694787 551996 696187 552046
rect 688917 551956 688951 551990
rect 698017 551933 698120 551969
rect 688917 551887 688951 551921
rect 692463 551885 692511 551909
rect 696191 551885 696239 551909
rect 688917 551818 688951 551852
rect 692487 551831 692511 551885
rect 696215 551831 696239 551885
rect 698017 551858 698053 551933
rect 692463 551807 692511 551831
rect 696191 551807 696239 551831
rect 698030 551824 698077 551858
rect 698017 551790 698053 551824
rect 688917 551749 688951 551783
rect 698030 551756 698077 551790
rect 698017 551722 698053 551756
rect 688917 551680 688951 551714
rect 698030 551688 698077 551722
rect 698017 551654 698053 551688
rect 688917 551611 688951 551645
rect 692463 551629 692521 551653
rect 696191 551629 696249 551653
rect 692487 551619 692521 551629
rect 696215 551619 696249 551629
rect 698030 551620 698077 551654
rect 698017 551586 698053 551620
rect 686879 551544 687585 551554
rect 686882 551528 687585 551544
rect 688917 551542 688951 551576
rect 692487 551547 692521 551581
rect 696215 551547 696249 551581
rect 678680 551433 678704 551467
rect 681345 551399 682345 551455
rect 678680 551365 678704 551399
rect 684004 551349 685004 551477
rect 688917 551473 688951 551507
rect 692487 551475 692521 551509
rect 696215 551475 696249 551509
rect 688917 551404 688951 551438
rect 692487 551427 692521 551437
rect 696215 551427 696249 551437
rect 692463 551403 692521 551427
rect 696191 551403 696249 551427
rect 688917 551335 688951 551369
rect 678680 551297 678704 551331
rect 678680 551229 678704 551263
rect 679133 551255 679283 551267
rect 679452 551255 679602 551267
rect 681345 551229 682345 551279
rect 678680 551161 678704 551195
rect 684004 551193 685004 551321
rect 688917 551266 688951 551300
rect 679002 551142 679602 551192
rect 678680 551093 678704 551127
rect 681441 551064 681457 551130
rect 682225 551064 682241 551130
rect 678680 551025 678704 551059
rect 684004 551037 685004 551165
rect 685537 551161 686137 551211
rect 688917 551197 688951 551231
rect 692463 551214 692521 551248
rect 696191 551214 696249 551248
rect 688917 551128 688951 551162
rect 678680 550957 678704 550991
rect 679002 550966 679602 551022
rect 678680 550889 678704 550923
rect 681441 550902 681457 550968
rect 683625 550902 683641 550968
rect 684004 550881 685004 551009
rect 685537 551005 686137 551061
rect 688917 551059 688951 551093
rect 692515 551084 693915 551127
rect 694787 551084 696187 551127
rect 688917 550990 688951 551024
rect 688917 550921 688951 550955
rect 692515 550921 693915 551049
rect 694787 550921 696187 551049
rect 685537 550855 686137 550905
rect 678680 550821 678704 550855
rect 679002 550796 679602 550846
rect 678680 550753 678704 550787
rect 680502 550761 680517 550776
rect 678680 550685 678704 550719
rect 678680 550617 678704 550651
rect 678680 550549 678704 550583
rect 680480 550581 680517 550761
rect 680502 550566 680517 550581
rect 680615 550761 680630 550776
rect 680803 550772 680815 550776
rect 680800 550761 680815 550772
rect 680615 550581 680815 550761
rect 681441 550740 681457 550806
rect 683625 550740 683641 550806
rect 684004 550725 685004 550853
rect 688917 550852 688951 550886
rect 688917 550783 688951 550817
rect 692515 550758 693915 550886
rect 694787 550758 696187 550886
rect 688917 550714 688951 550748
rect 686829 550649 687429 550699
rect 688917 550645 688951 550679
rect 680615 550566 680630 550581
rect 680800 550570 680815 550581
rect 681441 550578 681457 550644
rect 682225 550578 682241 550644
rect 684004 550575 685004 550625
rect 688917 550576 688951 550610
rect 692515 550595 693915 550723
rect 694787 550595 696187 550723
rect 680803 550566 680815 550570
rect 680615 550525 680630 550540
rect 680803 550536 680815 550540
rect 680800 550525 680815 550536
rect 678680 550481 678704 550515
rect 678680 550413 678704 550447
rect 678680 550345 678704 550379
rect 679007 550370 679607 550420
rect 680615 550345 680815 550525
rect 681345 550429 682345 550479
rect 686829 550473 687429 550529
rect 688917 550507 688951 550541
rect 688917 550438 688951 550472
rect 692515 550432 693915 550560
rect 694787 550432 696187 550560
rect 684054 550373 685054 550423
rect 688917 550393 688951 550403
rect 688893 550369 688951 550393
rect 680615 550330 680630 550345
rect 680800 550334 680815 550345
rect 680803 550330 680815 550334
rect 678680 550277 678704 550311
rect 681345 550253 682345 550309
rect 678680 550209 678704 550243
rect 679007 550200 679607 550250
rect 684054 550217 685054 550345
rect 686829 550303 687429 550353
rect 692515 550269 693915 550397
rect 694787 550269 696187 550397
rect 678680 550141 678704 550175
rect 678680 550073 678704 550107
rect 681345 550077 682345 550205
rect 678680 550005 678704 550039
rect 680215 550024 680815 550074
rect 684054 550061 685054 550189
rect 685793 550182 685805 550186
rect 685793 550171 685808 550182
rect 685978 550171 685993 550186
rect 678680 549937 678704 549971
rect 678680 549869 678704 549903
rect 680215 549848 680815 549904
rect 681345 549901 682345 550029
rect 684054 549905 685054 550033
rect 685793 549991 685993 550171
rect 685793 549980 685808 549991
rect 685793 549976 685805 549980
rect 685978 549976 685993 549991
rect 686053 550182 686065 550186
rect 686053 550171 686068 550182
rect 686238 550171 686253 550186
rect 686053 549991 686253 550171
rect 686607 550164 687607 550214
rect 697088 550171 697138 551571
rect 697238 550171 697366 551571
rect 697394 550171 697522 551571
rect 697550 550171 697678 551571
rect 697706 550171 697756 551571
rect 698030 551552 698077 551586
rect 698017 551518 698053 551552
rect 698030 551484 698077 551518
rect 698017 551450 698053 551484
rect 698030 551416 698077 551450
rect 698017 551382 698053 551416
rect 698030 551348 698077 551382
rect 698017 551314 698053 551348
rect 698030 551280 698077 551314
rect 698017 551246 698053 551280
rect 698030 551212 698077 551246
rect 698017 551178 698053 551212
rect 698030 551144 698077 551178
rect 698017 551110 698053 551144
rect 698030 551076 698077 551110
rect 698017 551042 698053 551076
rect 698030 551008 698077 551042
rect 698017 550974 698053 551008
rect 698030 550940 698077 550974
rect 698017 550906 698053 550940
rect 698030 550872 698077 550906
rect 698017 550838 698053 550872
rect 698030 550804 698077 550838
rect 698017 550770 698053 550804
rect 698030 550736 698077 550770
rect 698017 550702 698053 550736
rect 698030 550668 698077 550702
rect 698017 550634 698053 550668
rect 698030 550600 698077 550634
rect 698017 550566 698053 550600
rect 698030 550532 698077 550566
rect 698017 550498 698053 550532
rect 698030 550464 698077 550498
rect 698017 550430 698053 550464
rect 698030 550396 698077 550430
rect 698017 550362 698053 550396
rect 698030 550328 698077 550362
rect 698017 550294 698053 550328
rect 698030 550260 698077 550294
rect 698017 550226 698053 550260
rect 698030 550192 698077 550226
rect 692515 550119 693915 550162
rect 694787 550119 696187 550162
rect 698017 550158 698053 550192
rect 698030 550124 698077 550158
rect 698017 550090 698053 550124
rect 686607 550014 687607 550064
rect 698030 550056 698077 550090
rect 686053 549980 686068 549991
rect 686053 549976 686065 549980
rect 686238 549976 686253 549991
rect 685793 549946 685805 549950
rect 685793 549935 685808 549946
rect 685978 549935 685993 549950
rect 678680 549801 678704 549835
rect 678680 549733 678704 549767
rect 681345 549731 682345 549781
rect 684054 549749 685054 549877
rect 685793 549755 685993 549935
rect 685793 549744 685808 549755
rect 685793 549740 685805 549744
rect 685978 549740 685993 549755
rect 686053 549946 686065 549950
rect 686053 549935 686068 549946
rect 686238 549935 686253 549950
rect 686053 549755 686253 549935
rect 686607 549855 687607 549905
rect 692463 549809 692511 549833
rect 696191 549809 696239 549833
rect 686053 549744 686068 549755
rect 686053 549740 686065 549744
rect 686238 549740 686253 549755
rect 678680 549665 678704 549699
rect 680215 549672 680815 549728
rect 681345 549662 682345 549674
rect 678680 549597 678704 549631
rect 684054 549593 685054 549721
rect 686607 549705 687607 549755
rect 692487 549731 692511 549809
rect 696215 549755 696239 549809
rect 696191 549731 696239 549755
rect 696617 549772 696651 549773
rect 696617 549749 696626 549772
rect 696617 549731 696675 549749
rect 696651 549715 696675 549731
rect 696651 549647 696675 549681
rect 685533 549586 685545 549590
rect 685533 549575 685548 549586
rect 685718 549575 685733 549590
rect 678680 549529 678704 549563
rect 680215 549502 680815 549552
rect 678680 549461 678704 549495
rect 678680 549393 678704 549427
rect 680215 549370 680815 549420
rect 681466 549411 682466 549461
rect 684054 549437 685054 549565
rect 678680 549325 678704 549359
rect 678680 549257 678704 549291
rect 681466 549255 682466 549383
rect 682890 549339 683490 549389
rect 678680 549189 678704 549223
rect 680215 549194 680815 549250
rect 682890 549183 683490 549311
rect 684054 549281 685054 549409
rect 685533 549395 685733 549575
rect 685533 549384 685548 549395
rect 685533 549380 685545 549384
rect 685718 549380 685733 549395
rect 685793 549586 685805 549590
rect 685793 549575 685808 549586
rect 685978 549575 685993 549590
rect 685793 549395 685993 549575
rect 685793 549384 685808 549395
rect 685793 549380 685805 549384
rect 685978 549380 685993 549395
rect 686053 549586 686065 549590
rect 686053 549575 686068 549586
rect 686238 549575 686253 549590
rect 686053 549395 686253 549575
rect 686053 549384 686068 549395
rect 686053 549380 686065 549384
rect 686238 549380 686253 549395
rect 686313 549586 686325 549590
rect 686313 549575 686328 549586
rect 686498 549575 686513 549590
rect 686313 549395 686513 549575
rect 686313 549384 686328 549395
rect 686313 549380 686325 549384
rect 686498 549380 686513 549395
rect 686627 549586 686639 549590
rect 686627 549575 686642 549586
rect 686812 549575 686827 549590
rect 686627 549395 686827 549575
rect 686627 549384 686642 549395
rect 686627 549380 686639 549384
rect 686812 549380 686827 549395
rect 686887 549586 686899 549590
rect 686887 549575 686902 549586
rect 687072 549575 687087 549590
rect 686887 549395 687087 549575
rect 686887 549384 686902 549395
rect 686887 549380 686899 549384
rect 687072 549380 687087 549395
rect 687147 549586 687159 549590
rect 687147 549575 687162 549586
rect 687332 549575 687347 549590
rect 696651 549579 696675 549613
rect 687147 549395 687347 549575
rect 696651 549511 696675 549545
rect 696651 549443 696675 549477
rect 687147 549384 687162 549395
rect 687147 549380 687159 549384
rect 687332 549380 687347 549395
rect 696651 549375 696675 549409
rect 696651 549307 696675 549341
rect 685718 549215 685733 549230
rect 685679 549185 685733 549215
rect 678680 549121 678704 549155
rect 681466 549105 682466 549155
rect 684054 549131 685054 549181
rect 685718 549170 685733 549185
rect 685793 549226 685805 549230
rect 685793 549215 685808 549226
rect 685978 549215 685993 549230
rect 685793 549185 685993 549215
rect 685793 549174 685808 549185
rect 685793 549170 685805 549174
rect 685978 549170 685993 549185
rect 686053 549226 686065 549230
rect 686053 549215 686068 549226
rect 686238 549215 686253 549230
rect 686812 549215 686827 549230
rect 686053 549185 686253 549215
rect 686807 549185 686827 549215
rect 686053 549174 686068 549185
rect 686053 549170 686065 549174
rect 686238 549170 686253 549185
rect 686812 549170 686827 549185
rect 686887 549226 686899 549230
rect 686887 549215 686902 549226
rect 687072 549215 687087 549230
rect 686887 549185 687087 549215
rect 686887 549174 686902 549185
rect 686887 549170 686899 549174
rect 687072 549170 687087 549185
rect 687147 549226 687159 549230
rect 687147 549215 687162 549226
rect 687332 549215 687347 549230
rect 687147 549185 687347 549215
rect 687147 549174 687162 549185
rect 687147 549170 687159 549174
rect 687332 549170 687347 549185
rect 685718 549129 685733 549144
rect 681794 549102 682466 549105
rect 685679 549099 685733 549129
rect 678680 549053 678704 549087
rect 685718 549084 685733 549099
rect 685793 549140 685805 549144
rect 685793 549129 685808 549140
rect 685978 549129 685993 549144
rect 685793 549099 685993 549129
rect 685793 549088 685808 549099
rect 685793 549084 685805 549088
rect 685978 549084 685993 549099
rect 686053 549140 686065 549144
rect 686053 549129 686068 549140
rect 686238 549129 686253 549144
rect 686812 549129 686827 549144
rect 686053 549099 686253 549129
rect 686807 549099 686827 549129
rect 686053 549088 686068 549099
rect 686053 549084 686065 549088
rect 686238 549084 686253 549099
rect 686812 549084 686827 549099
rect 686887 549140 686899 549144
rect 686887 549129 686902 549140
rect 687072 549129 687087 549144
rect 686887 549099 687087 549129
rect 686887 549088 686902 549099
rect 686887 549084 686899 549088
rect 687072 549084 687087 549099
rect 687147 549140 687159 549144
rect 687147 549129 687162 549140
rect 687332 549129 687347 549144
rect 687147 549099 687347 549129
rect 687147 549088 687162 549099
rect 687147 549084 687159 549088
rect 687332 549084 687347 549099
rect 678680 548985 678704 549019
rect 680215 549018 680815 549074
rect 682890 549027 683490 549083
rect 678680 548917 678704 548951
rect 678680 548849 678704 548883
rect 680215 548848 680815 548898
rect 678680 548781 678704 548815
rect 678680 548713 678704 548747
rect 678680 548645 678704 548679
rect 679007 548672 679607 548722
rect 678680 548577 678704 548611
rect 680615 548577 680630 548592
rect 680803 548588 680815 548592
rect 680800 548577 680815 548588
rect 678680 548509 678704 548543
rect 679007 548502 679607 548552
rect 678680 548441 678704 548475
rect 678680 548373 678704 548407
rect 680615 548397 680815 548577
rect 681502 548505 681529 548995
rect 681866 548896 682466 549024
rect 682890 548871 683490 548999
rect 684004 548929 685004 548979
rect 685539 548940 685777 548972
rect 685803 548920 686119 548938
rect 681866 548740 682466 548868
rect 684004 548773 685004 548901
rect 682890 548721 683490 548771
rect 681866 548584 682466 548712
rect 682890 548605 683490 548655
rect 684004 548617 685004 548745
rect 681866 548434 682466 548484
rect 682890 548449 683490 548505
rect 684004 548461 685004 548589
rect 692427 548522 693027 548572
rect 680615 548382 680630 548397
rect 680800 548386 680815 548397
rect 680803 548382 680815 548386
rect 680502 548341 680517 548356
rect 678680 548305 678704 548339
rect 678680 548237 678704 548271
rect 678680 548169 678704 548203
rect 680480 548161 680517 548341
rect 680502 548146 680517 548161
rect 680615 548341 680630 548356
rect 680803 548352 680815 548356
rect 680800 548341 680815 548352
rect 680615 548161 680815 548341
rect 681866 548318 682466 548368
rect 682890 548293 683490 548349
rect 684004 548305 685004 548433
rect 692427 548366 693027 548494
rect 693888 548375 694194 548545
rect 694388 548375 694694 548545
rect 689309 548278 689909 548328
rect 681866 548168 682466 548218
rect 682041 548165 682385 548168
rect 680615 548146 680630 548161
rect 680800 548150 680815 548161
rect 680803 548146 680815 548150
rect 682890 548137 683490 548193
rect 684004 548149 685004 548277
rect 678680 548101 678704 548135
rect 679002 548076 679602 548126
rect 689309 548122 689909 548250
rect 692427 548210 693027 548338
rect 678680 548033 678704 548067
rect 678680 547965 678704 547999
rect 682890 547981 683490 548109
rect 684004 547993 685004 548121
rect 689309 547966 689909 548094
rect 692427 548054 693027 548110
rect 678680 547897 678704 547931
rect 679002 547900 679602 547956
rect 678680 547829 678704 547863
rect 682890 547825 683490 547953
rect 684004 547837 685004 547965
rect 692427 547898 693027 548026
rect 689309 547810 689909 547866
rect 678680 547761 678704 547795
rect 679002 547730 679602 547780
rect 679061 547727 679355 547730
rect 679380 547727 679602 547730
rect 678680 547693 678704 547727
rect 682890 547669 683490 547797
rect 684004 547687 685004 547737
rect 685803 547720 686119 547732
rect 685539 547716 686119 547720
rect 685513 547682 685537 547716
rect 685539 547682 685777 547716
rect 678680 547625 678704 547659
rect 689309 547654 689909 547782
rect 690910 547754 691110 547765
rect 692427 547742 693027 547870
rect 690910 547640 691110 547690
rect 678680 547557 678704 547591
rect 678680 547489 678704 547523
rect 682890 547513 683490 547569
rect 685718 547555 685733 547570
rect 684004 547485 685004 547535
rect 685679 547525 685733 547555
rect 685718 547510 685733 547525
rect 685793 547566 685805 547570
rect 685793 547555 685808 547566
rect 685978 547555 685993 547570
rect 685793 547525 685993 547555
rect 685793 547514 685808 547525
rect 685793 547510 685805 547514
rect 685978 547510 685993 547525
rect 686053 547566 686065 547570
rect 686053 547555 686068 547566
rect 686238 547555 686253 547570
rect 686812 547555 686827 547570
rect 686053 547525 686253 547555
rect 686807 547525 686827 547555
rect 686053 547514 686068 547525
rect 686053 547510 686065 547514
rect 686238 547510 686253 547525
rect 686812 547510 686827 547525
rect 686887 547566 686899 547570
rect 686887 547555 686902 547566
rect 687072 547555 687087 547570
rect 686887 547525 687087 547555
rect 686887 547514 686902 547525
rect 686887 547510 686899 547514
rect 687072 547510 687087 547525
rect 687147 547566 687159 547570
rect 687147 547555 687162 547566
rect 687332 547555 687347 547570
rect 687147 547525 687347 547555
rect 687147 547514 687162 547525
rect 687147 547510 687159 547514
rect 687332 547510 687347 547525
rect 689309 547498 689909 547626
rect 692427 547592 693027 547642
rect 693888 547575 694194 547745
rect 694388 547575 694694 547745
rect 678680 547421 678704 547455
rect 678680 547353 678704 547387
rect 682890 547357 683490 547485
rect 690910 547484 691110 547540
rect 685718 547469 685733 547484
rect 684004 547329 685004 547457
rect 685679 547439 685733 547469
rect 685718 547424 685733 547439
rect 685793 547480 685805 547484
rect 685793 547469 685808 547480
rect 685978 547469 685993 547484
rect 685793 547439 685993 547469
rect 685793 547428 685808 547439
rect 685793 547424 685805 547428
rect 685978 547424 685993 547439
rect 686053 547480 686065 547484
rect 686053 547469 686068 547480
rect 686238 547469 686253 547484
rect 686812 547469 686827 547484
rect 686053 547439 686253 547469
rect 686807 547439 686827 547469
rect 686053 547428 686068 547439
rect 686053 547424 686065 547428
rect 686238 547424 686253 547439
rect 686812 547424 686827 547439
rect 686887 547480 686899 547484
rect 686887 547469 686902 547480
rect 687072 547469 687087 547484
rect 686887 547439 687087 547469
rect 686887 547428 686902 547439
rect 686887 547424 686899 547428
rect 687072 547424 687087 547439
rect 687147 547480 687159 547484
rect 687147 547469 687162 547480
rect 687332 547469 687347 547484
rect 687147 547439 687347 547469
rect 692427 547462 693027 547512
rect 687147 547428 687162 547439
rect 687147 547424 687159 547428
rect 687332 547424 687347 547439
rect 689309 547348 689909 547398
rect 690910 547334 691110 547384
rect 678680 547285 678704 547319
rect 678680 547217 678704 547251
rect 682890 547201 683490 547329
rect 692427 547312 693027 547362
rect 678680 547149 678704 547183
rect 684004 547173 685004 547301
rect 685533 547270 685545 547274
rect 685533 547259 685548 547270
rect 685718 547259 685733 547274
rect 678680 547081 678704 547115
rect 679133 547101 679283 547113
rect 679452 547101 679602 547113
rect 678680 547013 678704 547047
rect 682890 547045 683490 547173
rect 679002 546988 679602 547038
rect 684004 547017 685004 547145
rect 685533 547079 685733 547259
rect 685533 547068 685548 547079
rect 685533 547064 685545 547068
rect 685718 547064 685733 547079
rect 685793 547270 685805 547274
rect 685793 547259 685808 547270
rect 685978 547259 685993 547274
rect 685793 547079 685993 547259
rect 685793 547068 685808 547079
rect 685793 547064 685805 547068
rect 685978 547064 685993 547079
rect 686053 547270 686065 547274
rect 686053 547259 686068 547270
rect 686238 547259 686253 547274
rect 686053 547079 686253 547259
rect 686053 547068 686068 547079
rect 686053 547064 686065 547068
rect 686238 547064 686253 547079
rect 686313 547270 686325 547274
rect 686313 547259 686328 547270
rect 686498 547259 686513 547274
rect 686313 547079 686513 547259
rect 686313 547068 686328 547079
rect 686313 547064 686325 547068
rect 686498 547064 686513 547079
rect 686627 547270 686639 547274
rect 686627 547259 686642 547270
rect 686812 547259 686827 547274
rect 686627 547079 686827 547259
rect 686627 547068 686642 547079
rect 686627 547064 686639 547068
rect 686812 547064 686827 547079
rect 686887 547270 686899 547274
rect 686887 547259 686902 547270
rect 687072 547259 687087 547274
rect 686887 547079 687087 547259
rect 686887 547068 686902 547079
rect 686887 547064 686899 547068
rect 687072 547064 687087 547079
rect 687147 547270 687159 547274
rect 687147 547259 687162 547270
rect 687332 547259 687347 547274
rect 687147 547079 687347 547259
rect 689309 547218 689909 547268
rect 692427 547140 693027 547190
rect 687147 547068 687162 547079
rect 687147 547064 687159 547068
rect 687332 547064 687347 547079
rect 689309 547068 689909 547118
rect 692427 546990 693027 547040
rect 678680 546945 678704 546979
rect 678680 546877 678704 546911
rect 682890 546895 683490 546945
rect 678680 546809 678704 546843
rect 679002 546812 679602 546868
rect 684004 546861 685004 546917
rect 685793 546910 685805 546914
rect 685793 546899 685808 546910
rect 685978 546899 685993 546914
rect 682890 546779 683490 546829
rect 678680 546741 678704 546775
rect 678680 546673 678704 546707
rect 679002 546642 679602 546692
rect 678680 546605 678704 546639
rect 682890 546623 683490 546751
rect 684004 546705 685004 546833
rect 685793 546719 685993 546899
rect 685793 546708 685808 546719
rect 685793 546704 685805 546708
rect 685978 546704 685993 546719
rect 686053 546910 686065 546914
rect 686053 546899 686068 546910
rect 686238 546899 686253 546914
rect 686607 546899 687607 546949
rect 690910 546934 691110 546984
rect 686053 546719 686253 546899
rect 692427 546860 693027 546910
rect 686607 546749 687607 546799
rect 690910 546778 691110 546834
rect 686053 546708 686068 546719
rect 686053 546704 686065 546708
rect 686238 546704 686253 546719
rect 692427 546704 693027 546832
rect 693888 546775 694194 546945
rect 694388 546775 694694 546945
rect 680502 546607 680517 546622
rect 678680 546537 678704 546571
rect 678680 546469 678704 546503
rect 678680 546401 678704 546435
rect 680480 546427 680517 546607
rect 680502 546412 680517 546427
rect 680615 546607 680630 546622
rect 680803 546618 680815 546622
rect 680800 546607 680815 546618
rect 680615 546427 680815 546607
rect 682890 546467 683490 546595
rect 684004 546549 685004 546677
rect 685793 546674 685805 546678
rect 685793 546663 685808 546674
rect 685978 546663 685993 546678
rect 680615 546412 680630 546427
rect 680800 546416 680815 546427
rect 680803 546412 680815 546416
rect 680615 546371 680630 546386
rect 680803 546382 680815 546386
rect 680800 546371 680815 546382
rect 678680 546333 678704 546367
rect 678680 546265 678704 546299
rect 678680 546197 678704 546231
rect 679007 546216 679607 546266
rect 680615 546191 680815 546371
rect 682890 546311 683490 546439
rect 684004 546393 685004 546521
rect 685793 546483 685993 546663
rect 685793 546472 685808 546483
rect 685793 546468 685805 546472
rect 685978 546468 685993 546483
rect 686053 546674 686065 546678
rect 686053 546663 686068 546674
rect 686238 546663 686253 546678
rect 686053 546483 686253 546663
rect 686607 546590 687607 546640
rect 690910 546628 691110 546678
rect 692427 546548 693027 546676
rect 686053 546472 686068 546483
rect 686053 546468 686065 546472
rect 686238 546468 686253 546483
rect 686607 546440 687607 546490
rect 692427 546392 693027 546448
rect 686829 546301 687429 546351
rect 684004 546243 685004 546293
rect 692427 546236 693027 546364
rect 695201 546282 695251 549282
rect 695351 546282 695479 549282
rect 695507 546282 695635 549282
rect 695663 546282 695791 549282
rect 695819 546282 695947 549282
rect 695975 546282 696103 549282
rect 696131 546282 696259 549282
rect 696287 546282 696337 549282
rect 696651 549239 696675 549273
rect 696651 549171 696675 549205
rect 696651 549103 696675 549137
rect 696651 549035 696675 549069
rect 696651 548967 696675 549001
rect 696651 548899 696675 548933
rect 696651 548831 696675 548865
rect 696651 548763 696675 548797
rect 696651 548695 696675 548729
rect 696651 548627 696675 548661
rect 697088 548641 697138 550041
rect 697238 548641 697366 550041
rect 697394 548641 697522 550041
rect 697550 548641 697678 550041
rect 697706 548641 697756 550041
rect 698017 550022 698053 550056
rect 698030 549988 698077 550022
rect 698017 549954 698053 549988
rect 698030 549920 698077 549954
rect 698017 549886 698053 549920
rect 698030 549852 698077 549886
rect 698017 549818 698053 549852
rect 698030 549784 698077 549818
rect 698017 549750 698053 549784
rect 698030 549716 698077 549750
rect 698017 549682 698053 549716
rect 698030 549648 698077 549682
rect 698017 549614 698053 549648
rect 698030 549580 698077 549614
rect 698017 549546 698053 549580
rect 698030 549512 698077 549546
rect 698017 549478 698053 549512
rect 698030 549444 698077 549478
rect 698017 549410 698053 549444
rect 698030 549376 698077 549410
rect 698017 549342 698053 549376
rect 698030 549308 698077 549342
rect 698017 549274 698053 549308
rect 698030 549240 698077 549274
rect 698017 549206 698053 549240
rect 698030 549172 698077 549206
rect 698017 549138 698053 549172
rect 698030 549104 698077 549138
rect 698017 549070 698053 549104
rect 698030 549036 698077 549070
rect 698017 549002 698053 549036
rect 698030 548968 698077 549002
rect 698017 548934 698053 548968
rect 698030 548900 698077 548934
rect 698017 548866 698053 548900
rect 698030 548832 698077 548866
rect 698017 548798 698053 548832
rect 698030 548764 698077 548798
rect 698017 548730 698053 548764
rect 698030 548696 698077 548730
rect 698017 548662 698053 548696
rect 698030 548628 698077 548662
rect 698017 548594 698053 548628
rect 696651 548559 696675 548593
rect 698030 548560 698077 548594
rect 698017 548526 698053 548560
rect 696651 548491 696675 548525
rect 698030 548492 698077 548526
rect 696651 548423 696675 548457
rect 698017 548428 698053 548492
rect 698030 548394 698077 548428
rect 696651 548355 696675 548389
rect 698017 548360 698053 548394
rect 698030 548326 698077 548360
rect 696651 548287 696675 548321
rect 698017 548292 698053 548326
rect 696651 548219 696675 548253
rect 696651 548151 696675 548185
rect 696651 548083 696675 548117
rect 696651 548015 696675 548049
rect 696651 547947 696675 547981
rect 696651 547879 696675 547913
rect 696651 547811 696675 547845
rect 696651 547743 696675 547777
rect 696651 547675 696675 547709
rect 696651 547607 696675 547641
rect 696651 547539 696675 547573
rect 696651 547471 696675 547505
rect 696651 547403 696675 547437
rect 696651 547335 696675 547369
rect 696651 547267 696675 547301
rect 696651 547199 696675 547233
rect 696651 547131 696675 547165
rect 696651 547063 696675 547097
rect 696651 546995 696675 547029
rect 696651 546927 696675 546961
rect 696651 546859 696675 546893
rect 697088 546879 697138 548279
rect 697238 546879 697366 548279
rect 697394 546879 697522 548279
rect 697550 546879 697678 548279
rect 697706 546879 697756 548279
rect 698030 548258 698077 548292
rect 698017 548224 698053 548258
rect 698030 548190 698077 548224
rect 698017 548156 698053 548190
rect 698030 548122 698077 548156
rect 698017 548088 698053 548122
rect 698030 548054 698077 548088
rect 698017 548020 698053 548054
rect 698030 547986 698077 548020
rect 698017 547952 698053 547986
rect 698030 547918 698077 547952
rect 698017 547884 698053 547918
rect 698030 547850 698077 547884
rect 698017 547816 698053 547850
rect 698030 547782 698077 547816
rect 698017 547748 698053 547782
rect 698030 547714 698077 547748
rect 698017 547680 698053 547714
rect 698030 547646 698077 547680
rect 698017 547612 698053 547646
rect 698030 547578 698077 547612
rect 698017 547544 698053 547578
rect 698030 547510 698077 547544
rect 698017 547476 698053 547510
rect 698030 547442 698077 547476
rect 698017 547408 698053 547442
rect 698030 547374 698077 547408
rect 698017 547340 698053 547374
rect 698030 547306 698077 547340
rect 698017 547272 698053 547306
rect 698030 547238 698077 547272
rect 698017 547204 698053 547238
rect 698030 547170 698077 547204
rect 698017 547136 698053 547170
rect 698030 547102 698077 547136
rect 698017 547068 698053 547102
rect 698030 547034 698077 547068
rect 698017 547000 698053 547034
rect 698030 546966 698077 547000
rect 698017 546932 698053 546966
rect 698030 546898 698077 546932
rect 698017 546864 698053 546898
rect 698030 546830 698077 546864
rect 696651 546791 696675 546825
rect 698017 546796 698053 546830
rect 698030 546762 698077 546796
rect 696651 546723 696675 546757
rect 696651 546655 696675 546689
rect 696651 546587 696675 546621
rect 696651 546519 696675 546553
rect 696651 546451 696675 546485
rect 696651 546383 696675 546417
rect 696651 546315 696675 546349
rect 696651 546247 696675 546281
rect 680615 546176 680630 546191
rect 680800 546180 680815 546191
rect 680803 546176 680815 546180
rect 678680 546129 678704 546163
rect 682890 546161 683490 546211
rect 684004 546127 685004 546177
rect 686829 546125 687429 546181
rect 678680 546061 678704 546095
rect 679007 546046 679607 546096
rect 692427 546080 693027 546208
rect 696651 546179 696675 546213
rect 696651 546111 696675 546145
rect 696651 546043 696675 546077
rect 678680 545993 678704 546027
rect 681664 546002 681812 546006
rect 681641 545994 681812 546002
rect 682113 545994 682313 546006
rect 684004 545971 685004 546027
rect 678680 545925 678704 545959
rect 686829 545955 687429 546005
rect 678680 545857 678704 545891
rect 680215 545870 680815 545920
rect 681713 545881 682313 545931
rect 682921 545899 683521 545949
rect 692427 545930 693027 545980
rect 696651 545975 696675 546009
rect 696651 545907 696675 545941
rect 678680 545789 678704 545823
rect 684004 545821 685004 545871
rect 678680 545721 678704 545755
rect 680215 545694 680815 545750
rect 681713 545705 682313 545761
rect 682921 545743 683521 545799
rect 685537 545749 686137 545799
rect 697088 545749 697138 546749
rect 697238 545749 697366 546749
rect 697394 545749 697522 546749
rect 697550 545749 697678 546749
rect 697706 545749 697756 546749
rect 698017 546728 698053 546762
rect 698030 546694 698077 546728
rect 698017 546660 698053 546694
rect 698030 546626 698077 546660
rect 698017 546592 698053 546626
rect 698030 546558 698077 546592
rect 698017 546524 698053 546558
rect 698030 546490 698077 546524
rect 698017 546456 698053 546490
rect 698030 546422 698077 546456
rect 698017 546388 698053 546422
rect 698030 546354 698077 546388
rect 698017 546320 698053 546354
rect 698030 546286 698077 546320
rect 698017 546252 698053 546286
rect 698030 546218 698077 546252
rect 698017 546184 698053 546218
rect 698030 546150 698077 546184
rect 698017 546116 698053 546150
rect 698030 546082 698077 546116
rect 698017 546048 698053 546082
rect 698030 546014 698077 546048
rect 698017 545980 698053 546014
rect 698030 545946 698077 545980
rect 698017 545912 698053 545946
rect 698030 545878 698077 545912
rect 698017 545844 698053 545878
rect 698030 545810 698077 545844
rect 698017 545776 698053 545810
rect 698030 545742 698077 545776
rect 698017 545708 698053 545742
rect 678680 545653 678704 545687
rect 698030 545674 698077 545708
rect 678680 545585 678704 545619
rect 680215 545518 680815 545574
rect 681713 545529 682313 545657
rect 682921 545593 683521 545643
rect 684070 545599 684670 545649
rect 685537 545593 686137 545649
rect 698017 545640 698053 545674
rect 698030 545606 698077 545640
rect 698017 545572 698053 545606
rect 698030 545538 698077 545572
rect 698017 545504 698053 545538
rect 684070 545443 684670 545499
rect 685537 545443 686137 545493
rect 692428 545442 693028 545492
rect 698030 545470 698077 545504
rect 698017 545436 698053 545470
rect 680215 545348 680815 545398
rect 681713 545359 682313 545409
rect 698030 545402 698077 545436
rect 698017 545368 698053 545402
rect 684070 545293 684670 545343
rect 692428 545292 693028 545342
rect 698030 545334 698077 545368
rect 698017 545300 698053 545334
rect 680215 545232 680815 545282
rect 698030 545266 698077 545300
rect 698017 545232 698053 545266
rect 692428 545162 693028 545212
rect 698030 545198 698077 545232
rect 698017 545164 698053 545198
rect 680215 545056 680815 545112
rect 692428 545006 693028 545134
rect 698030 545130 698077 545164
rect 698017 545096 698053 545130
rect 698030 545062 698077 545096
rect 698017 544983 698053 545062
rect 698084 544983 698120 551933
rect 699322 551908 700322 551964
rect 700922 551908 701922 551964
rect 707610 551953 708610 552009
rect 709211 551953 710211 552009
rect 699322 551836 700322 551892
rect 700922 551836 701922 551892
rect 707610 551881 708610 551937
rect 709211 551881 710211 551937
rect 699322 551534 700322 551606
rect 700922 551534 701922 551606
rect 707610 551579 708610 551651
rect 709211 551579 710211 551651
rect 699392 551523 699426 551534
rect 699460 551523 699494 551534
rect 699528 551523 699562 551534
rect 699596 551523 699630 551534
rect 699664 551523 699698 551534
rect 699732 551523 699766 551534
rect 699800 551523 699834 551534
rect 699868 551523 699902 551534
rect 699936 551523 699970 551534
rect 700004 551523 700038 551534
rect 700072 551523 700106 551534
rect 700140 551523 700174 551534
rect 700208 551523 700242 551534
rect 700276 551523 700310 551534
rect 700934 551523 700968 551534
rect 701002 551523 701036 551534
rect 701070 551523 701104 551534
rect 701138 551523 701172 551534
rect 701206 551523 701240 551534
rect 701274 551523 701308 551534
rect 701342 551523 701376 551534
rect 701410 551523 701444 551534
rect 701478 551523 701512 551534
rect 701546 551523 701580 551534
rect 701614 551523 701648 551534
rect 701682 551523 701716 551534
rect 701750 551523 701784 551534
rect 701818 551523 701852 551534
rect 699392 551513 699450 551523
rect 699460 551513 699518 551523
rect 699528 551513 699586 551523
rect 699596 551513 699654 551523
rect 699664 551513 699722 551523
rect 699732 551513 699790 551523
rect 699800 551513 699858 551523
rect 699868 551513 699926 551523
rect 699936 551513 699994 551523
rect 700004 551513 700062 551523
rect 700072 551513 700130 551523
rect 700140 551513 700198 551523
rect 700208 551513 700266 551523
rect 700276 551513 700334 551523
rect 700934 551513 700992 551523
rect 701002 551513 701060 551523
rect 701070 551513 701128 551523
rect 701138 551513 701196 551523
rect 701206 551513 701264 551523
rect 701274 551513 701332 551523
rect 701342 551513 701400 551523
rect 701410 551513 701468 551523
rect 701478 551513 701536 551523
rect 701546 551513 701604 551523
rect 701614 551513 701672 551523
rect 701682 551513 701740 551523
rect 701750 551513 701808 551523
rect 701818 551513 701876 551523
rect 699368 551489 700334 551513
rect 700910 551489 701876 551513
rect 699392 551474 699416 551489
rect 699460 551474 699484 551489
rect 699528 551474 699552 551489
rect 699596 551474 699620 551489
rect 699664 551474 699688 551489
rect 699732 551474 699756 551489
rect 699800 551474 699824 551489
rect 699868 551474 699892 551489
rect 699936 551474 699960 551489
rect 700004 551474 700028 551489
rect 700072 551474 700096 551489
rect 700140 551474 700164 551489
rect 700208 551474 700232 551489
rect 700276 551474 700300 551489
rect 700934 551474 700958 551489
rect 701002 551474 701026 551489
rect 701070 551474 701094 551489
rect 701138 551474 701162 551489
rect 701206 551474 701230 551489
rect 701274 551474 701298 551489
rect 701342 551474 701366 551489
rect 701410 551474 701434 551489
rect 701478 551474 701502 551489
rect 701546 551474 701570 551489
rect 701614 551474 701638 551489
rect 701682 551474 701706 551489
rect 701750 551474 701774 551489
rect 701818 551474 701842 551489
rect 699322 551319 700322 551474
rect 699322 551285 700334 551319
rect 700922 551309 701922 551474
rect 707610 551319 708610 551379
rect 709211 551319 710211 551379
rect 700910 551285 701922 551309
rect 699322 551274 700322 551285
rect 700922 551274 701922 551285
rect 699392 551261 699416 551274
rect 699460 551261 699484 551274
rect 699528 551261 699552 551274
rect 699596 551261 699620 551274
rect 699664 551261 699688 551274
rect 699732 551261 699756 551274
rect 699800 551261 699824 551274
rect 699868 551261 699892 551274
rect 699936 551261 699960 551274
rect 700004 551261 700028 551274
rect 700072 551261 700096 551274
rect 700140 551261 700164 551274
rect 700208 551261 700232 551274
rect 700276 551261 700300 551274
rect 700934 551261 700958 551274
rect 701002 551261 701026 551274
rect 701070 551261 701094 551274
rect 701138 551261 701162 551274
rect 701206 551261 701230 551274
rect 701274 551261 701298 551274
rect 701342 551261 701366 551274
rect 701410 551261 701434 551274
rect 701478 551261 701502 551274
rect 701546 551261 701570 551274
rect 701614 551261 701638 551274
rect 701682 551261 701706 551274
rect 701750 551261 701774 551274
rect 701818 551261 701842 551274
rect 699322 550916 700322 550972
rect 700922 550916 701922 550972
rect 707610 550961 708610 551017
rect 709211 550961 710211 551017
rect 699322 550844 700322 550900
rect 700922 550844 701922 550900
rect 707610 550889 708610 550945
rect 709211 550889 710211 550945
rect 699322 550542 700322 550614
rect 700922 550542 701922 550614
rect 707610 550587 708610 550659
rect 709211 550587 710211 550659
rect 699392 550531 699426 550542
rect 699460 550531 699494 550542
rect 699528 550531 699562 550542
rect 699596 550531 699630 550542
rect 699664 550531 699698 550542
rect 699732 550531 699766 550542
rect 699800 550531 699834 550542
rect 699868 550531 699902 550542
rect 699936 550531 699970 550542
rect 700004 550531 700038 550542
rect 700072 550531 700106 550542
rect 700140 550531 700174 550542
rect 700208 550531 700242 550542
rect 700276 550531 700310 550542
rect 700934 550531 700968 550542
rect 701002 550531 701036 550542
rect 701070 550531 701104 550542
rect 701138 550531 701172 550542
rect 701206 550531 701240 550542
rect 701274 550531 701308 550542
rect 701342 550531 701376 550542
rect 701410 550531 701444 550542
rect 701478 550531 701512 550542
rect 701546 550531 701580 550542
rect 701614 550531 701648 550542
rect 701682 550531 701716 550542
rect 701750 550531 701784 550542
rect 701818 550531 701852 550542
rect 699392 550521 699450 550531
rect 699460 550521 699518 550531
rect 699528 550521 699586 550531
rect 699596 550521 699654 550531
rect 699664 550521 699722 550531
rect 699732 550521 699790 550531
rect 699800 550521 699858 550531
rect 699868 550521 699926 550531
rect 699936 550521 699994 550531
rect 700004 550521 700062 550531
rect 700072 550521 700130 550531
rect 700140 550521 700198 550531
rect 700208 550521 700266 550531
rect 700276 550521 700334 550531
rect 700934 550521 700992 550531
rect 701002 550521 701060 550531
rect 701070 550521 701128 550531
rect 701138 550521 701196 550531
rect 701206 550521 701264 550531
rect 701274 550521 701332 550531
rect 701342 550521 701400 550531
rect 701410 550521 701468 550531
rect 701478 550521 701536 550531
rect 701546 550521 701604 550531
rect 701614 550521 701672 550531
rect 701682 550521 701740 550531
rect 701750 550521 701808 550531
rect 701818 550521 701876 550531
rect 699368 550497 700334 550521
rect 700910 550497 701876 550521
rect 699392 550482 699416 550497
rect 699460 550482 699484 550497
rect 699528 550482 699552 550497
rect 699596 550482 699620 550497
rect 699664 550482 699688 550497
rect 699732 550482 699756 550497
rect 699800 550482 699824 550497
rect 699868 550482 699892 550497
rect 699936 550482 699960 550497
rect 700004 550482 700028 550497
rect 700072 550482 700096 550497
rect 700140 550482 700164 550497
rect 700208 550482 700232 550497
rect 700276 550482 700300 550497
rect 700934 550482 700958 550497
rect 701002 550482 701026 550497
rect 701070 550482 701094 550497
rect 701138 550482 701162 550497
rect 701206 550482 701230 550497
rect 701274 550482 701298 550497
rect 701342 550482 701366 550497
rect 701410 550482 701434 550497
rect 701478 550482 701502 550497
rect 701546 550482 701570 550497
rect 701614 550482 701638 550497
rect 701682 550482 701706 550497
rect 701750 550482 701774 550497
rect 701818 550482 701842 550497
rect 699322 550327 700322 550482
rect 699322 550293 700334 550327
rect 700922 550317 701922 550482
rect 707610 550327 708610 550387
rect 709211 550327 710211 550387
rect 711541 550345 711629 557461
rect 711892 556200 711942 557200
rect 712062 556200 712112 557200
rect 711892 555079 711942 556079
rect 712062 555079 712112 556079
rect 711892 553958 711942 554958
rect 712062 553958 712112 554958
rect 711892 552848 711942 553848
rect 712062 552848 712112 553848
rect 711892 551727 711942 552727
rect 712062 551727 712112 552727
rect 711892 550606 711942 551606
rect 712062 550606 712112 551606
rect 712409 550371 712431 557485
rect 712469 557459 712487 557501
rect 712499 557459 712505 557467
rect 712499 557455 712511 557459
rect 712539 557455 712557 557501
rect 713640 555461 713674 557785
rect 713750 557772 714750 557822
rect 717367 557820 717413 557853
rect 717367 557819 717379 557820
rect 717401 557819 717413 557820
rect 717401 557809 717600 557819
rect 717401 557786 717413 557809
rect 713750 557562 714750 557612
rect 713750 557446 714750 557496
rect 713750 557230 714750 557358
rect 713750 557014 714750 557070
rect 713750 556798 714750 556926
rect 713750 556588 714750 556638
rect 714478 556585 714750 556588
rect 715486 555931 715536 556931
rect 715696 555931 715824 556931
rect 715912 555931 715962 556931
rect 713641 555345 713663 555461
rect 713640 555309 713674 555345
rect 713750 555314 714750 555364
rect 713750 555158 714750 555214
rect 713750 555002 714750 555130
rect 713750 554846 714750 554974
rect 713750 554690 714750 554746
rect 716425 554709 716725 554721
rect 713750 554534 714750 554662
rect 716425 554596 717425 554646
rect 713750 554378 714750 554506
rect 716425 554440 717425 554568
rect 713750 554222 714750 554350
rect 716425 554284 717425 554340
rect 713750 554072 714750 554122
rect 713750 553956 714750 554006
rect 713750 553800 714750 553928
rect 713750 553644 714750 553772
rect 713750 553488 714750 553616
rect 715354 553587 715404 554187
rect 715504 553587 715560 554187
rect 715660 553587 715716 554187
rect 715816 553587 715872 554187
rect 715972 553587 716022 554187
rect 716425 554128 717425 554256
rect 716425 553978 717425 554028
rect 716425 553862 717425 553912
rect 716425 553706 717425 553834
rect 716425 553550 717425 553606
rect 716425 553394 717425 553522
rect 713750 553332 714750 553388
rect 713750 553176 714750 553304
rect 716425 553244 717425 553294
rect 713750 553020 714750 553148
rect 713750 552870 714750 552920
rect 713750 552742 714750 552792
rect 713750 552586 714750 552642
rect 713750 552436 714750 552486
rect 713750 552320 714350 552370
rect 713750 552164 714350 552292
rect 715510 552191 715560 553191
rect 715660 552191 715788 553191
rect 715816 552191 715944 553191
rect 715972 552191 716022 553191
rect 716425 553128 717425 553178
rect 716425 552972 717425 553028
rect 716425 552822 717425 552872
rect 716425 552706 717425 552756
rect 716425 552550 717425 552678
rect 716425 552394 717425 552522
rect 716425 552238 717425 552366
rect 716425 552082 717425 552210
rect 713750 552008 714350 552064
rect 713750 551852 714350 551980
rect 716425 551932 717425 551982
rect 713750 551696 714350 551752
rect 713750 551446 714350 551496
rect 714565 551443 714765 551455
rect 713750 551330 714750 551380
rect 713750 551120 714750 551170
rect 716413 551092 716447 551150
rect 713750 551004 714750 551054
rect 713750 550794 714750 550844
rect 713750 550678 714750 550728
rect 713750 550468 714750 550518
rect 713750 550352 714750 550402
rect 700910 550293 701922 550317
rect 699322 550282 700322 550293
rect 700922 550282 701922 550293
rect 711541 550311 711633 550345
rect 699392 550269 699416 550282
rect 699460 550269 699484 550282
rect 699528 550269 699552 550282
rect 699596 550269 699620 550282
rect 699664 550269 699688 550282
rect 699732 550269 699756 550282
rect 699800 550269 699824 550282
rect 699868 550269 699892 550282
rect 699936 550269 699960 550282
rect 700004 550269 700028 550282
rect 700072 550269 700096 550282
rect 700140 550269 700164 550282
rect 700208 550269 700232 550282
rect 700276 550269 700300 550282
rect 700934 550269 700958 550282
rect 701002 550269 701026 550282
rect 701070 550269 701094 550282
rect 701138 550269 701162 550282
rect 701206 550269 701230 550282
rect 701274 550269 701298 550282
rect 701342 550269 701366 550282
rect 701410 550269 701434 550282
rect 701478 550269 701502 550282
rect 701546 550269 701570 550282
rect 701614 550269 701638 550282
rect 701682 550269 701706 550282
rect 701750 550269 701774 550282
rect 701818 550269 701842 550282
rect 699322 549924 700322 549980
rect 700922 549924 701922 549980
rect 707610 549969 708610 550025
rect 709211 549969 710211 550025
rect 699322 549852 700322 549908
rect 700922 549852 701922 549908
rect 707610 549897 708610 549953
rect 709211 549897 710211 549953
rect 699322 549550 700322 549622
rect 700922 549550 701922 549622
rect 707610 549595 708610 549667
rect 709211 549595 710211 549667
rect 699392 549539 699426 549550
rect 699460 549539 699494 549550
rect 699528 549539 699562 549550
rect 699596 549539 699630 549550
rect 699664 549539 699698 549550
rect 699732 549539 699766 549550
rect 699800 549539 699834 549550
rect 699868 549539 699902 549550
rect 699936 549539 699970 549550
rect 700004 549539 700038 549550
rect 700072 549539 700106 549550
rect 700140 549539 700174 549550
rect 700208 549539 700242 549550
rect 700276 549539 700310 549550
rect 700934 549539 700968 549550
rect 701002 549539 701036 549550
rect 701070 549539 701104 549550
rect 701138 549539 701172 549550
rect 701206 549539 701240 549550
rect 701274 549539 701308 549550
rect 701342 549539 701376 549550
rect 701410 549539 701444 549550
rect 701478 549539 701512 549550
rect 701546 549539 701580 549550
rect 701614 549539 701648 549550
rect 701682 549539 701716 549550
rect 701750 549539 701784 549550
rect 701818 549539 701852 549550
rect 699392 549529 699450 549539
rect 699460 549529 699518 549539
rect 699528 549529 699586 549539
rect 699596 549529 699654 549539
rect 699664 549529 699722 549539
rect 699732 549529 699790 549539
rect 699800 549529 699858 549539
rect 699868 549529 699926 549539
rect 699936 549529 699994 549539
rect 700004 549529 700062 549539
rect 700072 549529 700130 549539
rect 700140 549529 700198 549539
rect 700208 549529 700266 549539
rect 700276 549529 700334 549539
rect 700934 549529 700992 549539
rect 701002 549529 701060 549539
rect 701070 549529 701128 549539
rect 701138 549529 701196 549539
rect 701206 549529 701264 549539
rect 701274 549529 701332 549539
rect 701342 549529 701400 549539
rect 701410 549529 701468 549539
rect 701478 549529 701536 549539
rect 701546 549529 701604 549539
rect 701614 549529 701672 549539
rect 701682 549529 701740 549539
rect 701750 549529 701808 549539
rect 701818 549529 701876 549539
rect 699368 549505 700334 549529
rect 700910 549505 701876 549529
rect 699392 549490 699416 549505
rect 699460 549490 699484 549505
rect 699528 549490 699552 549505
rect 699596 549490 699620 549505
rect 699664 549490 699688 549505
rect 699732 549490 699756 549505
rect 699800 549490 699824 549505
rect 699868 549490 699892 549505
rect 699936 549490 699960 549505
rect 700004 549490 700028 549505
rect 700072 549490 700096 549505
rect 700140 549490 700164 549505
rect 700208 549490 700232 549505
rect 700276 549490 700300 549505
rect 700934 549490 700958 549505
rect 701002 549490 701026 549505
rect 701070 549490 701094 549505
rect 701138 549490 701162 549505
rect 701206 549490 701230 549505
rect 701274 549490 701298 549505
rect 701342 549490 701366 549505
rect 701410 549490 701434 549505
rect 701478 549490 701502 549505
rect 701546 549490 701570 549505
rect 701614 549490 701638 549505
rect 701682 549490 701706 549505
rect 701750 549490 701774 549505
rect 701818 549490 701842 549505
rect 699322 549335 700322 549490
rect 699322 549301 700334 549335
rect 700922 549325 701922 549490
rect 707610 549335 708610 549395
rect 709211 549335 710211 549395
rect 700910 549301 701922 549325
rect 699322 549290 700322 549301
rect 700922 549290 701922 549301
rect 699392 549277 699416 549290
rect 699460 549277 699484 549290
rect 699528 549277 699552 549290
rect 699596 549277 699620 549290
rect 699664 549277 699688 549290
rect 699732 549277 699756 549290
rect 699800 549277 699824 549290
rect 699868 549277 699892 549290
rect 699936 549277 699960 549290
rect 700004 549277 700028 549290
rect 700072 549277 700096 549290
rect 700140 549277 700164 549290
rect 700208 549277 700232 549290
rect 700276 549277 700300 549290
rect 700934 549277 700958 549290
rect 701002 549277 701026 549290
rect 701070 549277 701094 549290
rect 701138 549277 701162 549290
rect 701206 549277 701230 549290
rect 701274 549277 701298 549290
rect 701342 549277 701366 549290
rect 701410 549277 701434 549290
rect 701478 549277 701502 549290
rect 701546 549277 701570 549290
rect 701614 549277 701638 549290
rect 701682 549277 701706 549290
rect 701750 549277 701774 549290
rect 701818 549277 701842 549290
rect 699322 548932 700322 548988
rect 700922 548932 701922 548988
rect 707610 548977 708610 549033
rect 709211 548977 710211 549033
rect 699322 548860 700322 548916
rect 700922 548860 701922 548916
rect 707610 548905 708610 548961
rect 709211 548905 710211 548961
rect 699322 548558 700322 548630
rect 700922 548558 701922 548630
rect 707610 548603 708610 548675
rect 709211 548603 710211 548675
rect 699392 548547 699426 548558
rect 699460 548547 699494 548558
rect 699528 548547 699562 548558
rect 699596 548547 699630 548558
rect 699664 548547 699698 548558
rect 699732 548547 699766 548558
rect 699800 548547 699834 548558
rect 699868 548547 699902 548558
rect 699936 548547 699970 548558
rect 700004 548547 700038 548558
rect 700072 548547 700106 548558
rect 700140 548547 700174 548558
rect 700208 548547 700242 548558
rect 700276 548547 700310 548558
rect 700934 548547 700968 548558
rect 701002 548547 701036 548558
rect 701070 548547 701104 548558
rect 701138 548547 701172 548558
rect 701206 548547 701240 548558
rect 701274 548547 701308 548558
rect 701342 548547 701376 548558
rect 701410 548547 701444 548558
rect 701478 548547 701512 548558
rect 701546 548547 701580 548558
rect 701614 548547 701648 548558
rect 701682 548547 701716 548558
rect 701750 548547 701784 548558
rect 701818 548547 701852 548558
rect 699392 548537 699450 548547
rect 699460 548537 699518 548547
rect 699528 548537 699586 548547
rect 699596 548537 699654 548547
rect 699664 548537 699722 548547
rect 699732 548537 699790 548547
rect 699800 548537 699858 548547
rect 699868 548537 699926 548547
rect 699936 548537 699994 548547
rect 700004 548537 700062 548547
rect 700072 548537 700130 548547
rect 700140 548537 700198 548547
rect 700208 548537 700266 548547
rect 700276 548537 700334 548547
rect 700934 548537 700992 548547
rect 701002 548537 701060 548547
rect 701070 548537 701128 548547
rect 701138 548537 701196 548547
rect 701206 548537 701264 548547
rect 701274 548537 701332 548547
rect 701342 548537 701400 548547
rect 701410 548537 701468 548547
rect 701478 548537 701536 548547
rect 701546 548537 701604 548547
rect 701614 548537 701672 548547
rect 701682 548537 701740 548547
rect 701750 548537 701808 548547
rect 701818 548537 701876 548547
rect 699368 548513 700334 548537
rect 700910 548513 701876 548537
rect 699392 548498 699416 548513
rect 699460 548498 699484 548513
rect 699528 548498 699552 548513
rect 699596 548498 699620 548513
rect 699664 548498 699688 548513
rect 699732 548498 699756 548513
rect 699800 548498 699824 548513
rect 699868 548498 699892 548513
rect 699936 548498 699960 548513
rect 700004 548498 700028 548513
rect 700072 548498 700096 548513
rect 700140 548498 700164 548513
rect 700208 548498 700232 548513
rect 700276 548498 700300 548513
rect 700934 548498 700958 548513
rect 701002 548498 701026 548513
rect 701070 548498 701094 548513
rect 701138 548498 701162 548513
rect 701206 548498 701230 548513
rect 701274 548498 701298 548513
rect 701342 548498 701366 548513
rect 701410 548498 701434 548513
rect 701478 548498 701502 548513
rect 701546 548498 701570 548513
rect 701614 548498 701638 548513
rect 701682 548498 701706 548513
rect 701750 548498 701774 548513
rect 701818 548498 701842 548513
rect 699322 548343 700322 548498
rect 699322 548309 700334 548343
rect 700922 548333 701922 548498
rect 707610 548343 708610 548403
rect 709211 548343 710211 548403
rect 700910 548309 701922 548333
rect 699322 548298 700322 548309
rect 700922 548298 701922 548309
rect 699392 548285 699416 548298
rect 699460 548285 699484 548298
rect 699528 548285 699552 548298
rect 699596 548285 699620 548298
rect 699664 548285 699688 548298
rect 699732 548285 699756 548298
rect 699800 548285 699824 548298
rect 699868 548285 699892 548298
rect 699936 548285 699960 548298
rect 700004 548285 700028 548298
rect 700072 548285 700096 548298
rect 700140 548285 700164 548298
rect 700208 548285 700232 548298
rect 700276 548285 700300 548298
rect 700934 548285 700958 548298
rect 701002 548285 701026 548298
rect 701070 548285 701094 548298
rect 701138 548285 701162 548298
rect 701206 548285 701230 548298
rect 701274 548285 701298 548298
rect 701342 548285 701366 548298
rect 701410 548285 701434 548298
rect 701478 548285 701502 548298
rect 701546 548285 701570 548298
rect 701614 548285 701638 548298
rect 701682 548285 701706 548298
rect 701750 548285 701774 548298
rect 701818 548285 701842 548298
rect 699322 547940 700322 547996
rect 700922 547940 701922 547996
rect 707610 547985 708610 548041
rect 709211 547985 710211 548041
rect 699322 547868 700322 547924
rect 700922 547868 701922 547924
rect 707610 547913 708610 547969
rect 709211 547913 710211 547969
rect 699322 547566 700322 547638
rect 700922 547566 701922 547638
rect 707610 547611 708610 547683
rect 709211 547611 710211 547683
rect 699392 547555 699426 547566
rect 699460 547555 699494 547566
rect 699528 547555 699562 547566
rect 699596 547555 699630 547566
rect 699664 547555 699698 547566
rect 699732 547555 699766 547566
rect 699800 547555 699834 547566
rect 699868 547555 699902 547566
rect 699936 547555 699970 547566
rect 700004 547555 700038 547566
rect 700072 547555 700106 547566
rect 700140 547555 700174 547566
rect 700208 547555 700242 547566
rect 700276 547555 700310 547566
rect 700934 547555 700968 547566
rect 701002 547555 701036 547566
rect 701070 547555 701104 547566
rect 701138 547555 701172 547566
rect 701206 547555 701240 547566
rect 701274 547555 701308 547566
rect 701342 547555 701376 547566
rect 701410 547555 701444 547566
rect 701478 547555 701512 547566
rect 701546 547555 701580 547566
rect 701614 547555 701648 547566
rect 701682 547555 701716 547566
rect 701750 547555 701784 547566
rect 701818 547555 701852 547566
rect 699392 547545 699450 547555
rect 699460 547545 699518 547555
rect 699528 547545 699586 547555
rect 699596 547545 699654 547555
rect 699664 547545 699722 547555
rect 699732 547545 699790 547555
rect 699800 547545 699858 547555
rect 699868 547545 699926 547555
rect 699936 547545 699994 547555
rect 700004 547545 700062 547555
rect 700072 547545 700130 547555
rect 700140 547545 700198 547555
rect 700208 547545 700266 547555
rect 700276 547545 700334 547555
rect 700934 547545 700992 547555
rect 701002 547545 701060 547555
rect 701070 547545 701128 547555
rect 701138 547545 701196 547555
rect 701206 547545 701264 547555
rect 701274 547545 701332 547555
rect 701342 547545 701400 547555
rect 701410 547545 701468 547555
rect 701478 547545 701536 547555
rect 701546 547545 701604 547555
rect 701614 547545 701672 547555
rect 701682 547545 701740 547555
rect 701750 547545 701808 547555
rect 701818 547545 701876 547555
rect 699368 547521 700334 547545
rect 700910 547521 701876 547545
rect 699392 547506 699416 547521
rect 699460 547506 699484 547521
rect 699528 547506 699552 547521
rect 699596 547506 699620 547521
rect 699664 547506 699688 547521
rect 699732 547506 699756 547521
rect 699800 547506 699824 547521
rect 699868 547506 699892 547521
rect 699936 547506 699960 547521
rect 700004 547506 700028 547521
rect 700072 547506 700096 547521
rect 700140 547506 700164 547521
rect 700208 547506 700232 547521
rect 700276 547506 700300 547521
rect 700934 547506 700958 547521
rect 701002 547506 701026 547521
rect 701070 547506 701094 547521
rect 701138 547506 701162 547521
rect 701206 547506 701230 547521
rect 701274 547506 701298 547521
rect 701342 547506 701366 547521
rect 701410 547506 701434 547521
rect 701478 547506 701502 547521
rect 701546 547506 701570 547521
rect 701614 547506 701638 547521
rect 701682 547506 701706 547521
rect 701750 547506 701774 547521
rect 701818 547506 701842 547521
rect 699322 547351 700322 547506
rect 699322 547317 700334 547351
rect 700922 547341 701922 547506
rect 705107 547360 705173 547376
rect 707610 547351 708610 547411
rect 709211 547351 710211 547411
rect 700910 547317 701922 547341
rect 699322 547306 700322 547317
rect 700922 547306 701922 547317
rect 699392 547293 699416 547306
rect 699460 547293 699484 547306
rect 699528 547293 699552 547306
rect 699596 547293 699620 547306
rect 699664 547293 699688 547306
rect 699732 547293 699756 547306
rect 699800 547293 699824 547306
rect 699868 547293 699892 547306
rect 699936 547293 699960 547306
rect 700004 547293 700028 547306
rect 700072 547293 700096 547306
rect 700140 547293 700164 547306
rect 700208 547293 700232 547306
rect 700276 547293 700300 547306
rect 700934 547293 700958 547306
rect 701002 547293 701026 547306
rect 701070 547293 701094 547306
rect 701138 547293 701162 547306
rect 701206 547293 701230 547306
rect 701274 547293 701298 547306
rect 701342 547293 701366 547306
rect 701410 547293 701434 547306
rect 701478 547293 701502 547306
rect 701546 547293 701570 547306
rect 701614 547293 701638 547306
rect 701682 547293 701706 547306
rect 701750 547293 701774 547306
rect 701818 547293 701842 547306
rect 699322 546948 700322 547004
rect 700922 546948 701922 547004
rect 707610 546993 708610 547049
rect 709211 546993 710211 547049
rect 699322 546876 700322 546932
rect 700922 546876 701922 546932
rect 707610 546921 708610 546977
rect 709211 546921 710211 546977
rect 699322 546574 700322 546646
rect 700922 546574 701922 546646
rect 707610 546619 708610 546691
rect 709211 546619 710211 546691
rect 699392 546563 699426 546574
rect 699460 546563 699494 546574
rect 699528 546563 699562 546574
rect 699596 546563 699630 546574
rect 699664 546563 699698 546574
rect 699732 546563 699766 546574
rect 699800 546563 699834 546574
rect 699868 546563 699902 546574
rect 699936 546563 699970 546574
rect 700004 546563 700038 546574
rect 700072 546563 700106 546574
rect 700140 546563 700174 546574
rect 700208 546563 700242 546574
rect 700276 546563 700310 546574
rect 700934 546563 700968 546574
rect 701002 546563 701036 546574
rect 701070 546563 701104 546574
rect 701138 546563 701172 546574
rect 701206 546563 701240 546574
rect 701274 546563 701308 546574
rect 701342 546563 701376 546574
rect 701410 546563 701444 546574
rect 701478 546563 701512 546574
rect 701546 546563 701580 546574
rect 701614 546563 701648 546574
rect 701682 546563 701716 546574
rect 701750 546563 701784 546574
rect 701818 546563 701852 546574
rect 699392 546553 699450 546563
rect 699460 546553 699518 546563
rect 699528 546553 699586 546563
rect 699596 546553 699654 546563
rect 699664 546553 699722 546563
rect 699732 546553 699790 546563
rect 699800 546553 699858 546563
rect 699868 546553 699926 546563
rect 699936 546553 699994 546563
rect 700004 546553 700062 546563
rect 700072 546553 700130 546563
rect 700140 546553 700198 546563
rect 700208 546553 700266 546563
rect 700276 546553 700334 546563
rect 700934 546553 700992 546563
rect 701002 546553 701060 546563
rect 701070 546553 701128 546563
rect 701138 546553 701196 546563
rect 701206 546553 701264 546563
rect 701274 546553 701332 546563
rect 701342 546553 701400 546563
rect 701410 546553 701468 546563
rect 701478 546553 701536 546563
rect 701546 546553 701604 546563
rect 701614 546553 701672 546563
rect 701682 546553 701740 546563
rect 701750 546553 701808 546563
rect 701818 546553 701876 546563
rect 699368 546529 700334 546553
rect 700910 546529 701876 546553
rect 699392 546514 699416 546529
rect 699460 546514 699484 546529
rect 699528 546514 699552 546529
rect 699596 546514 699620 546529
rect 699664 546514 699688 546529
rect 699732 546514 699756 546529
rect 699800 546514 699824 546529
rect 699868 546514 699892 546529
rect 699936 546514 699960 546529
rect 700004 546514 700028 546529
rect 700072 546514 700096 546529
rect 700140 546514 700164 546529
rect 700208 546514 700232 546529
rect 700276 546514 700300 546529
rect 700934 546514 700958 546529
rect 701002 546514 701026 546529
rect 701070 546514 701094 546529
rect 701138 546514 701162 546529
rect 701206 546514 701230 546529
rect 701274 546514 701298 546529
rect 701342 546514 701366 546529
rect 701410 546514 701434 546529
rect 701478 546514 701502 546529
rect 701546 546514 701570 546529
rect 701614 546514 701638 546529
rect 701682 546514 701706 546529
rect 701750 546514 701774 546529
rect 701818 546514 701842 546529
rect 699322 546359 700322 546514
rect 699322 546325 700334 546359
rect 700922 546349 701922 546514
rect 707610 546359 708610 546419
rect 709211 546359 710211 546419
rect 700910 546325 701922 546349
rect 699322 546314 700322 546325
rect 700922 546314 701922 546325
rect 699392 546301 699416 546314
rect 699460 546301 699484 546314
rect 699528 546301 699552 546314
rect 699596 546301 699620 546314
rect 699664 546301 699688 546314
rect 699732 546301 699756 546314
rect 699800 546301 699824 546314
rect 699868 546301 699892 546314
rect 699936 546301 699960 546314
rect 700004 546301 700028 546314
rect 700072 546301 700096 546314
rect 700140 546301 700164 546314
rect 700208 546301 700232 546314
rect 700276 546301 700300 546314
rect 700934 546301 700958 546314
rect 701002 546301 701026 546314
rect 701070 546301 701094 546314
rect 701138 546301 701162 546314
rect 701206 546301 701230 546314
rect 701274 546301 701298 546314
rect 701342 546301 701366 546314
rect 701410 546301 701434 546314
rect 701478 546301 701502 546314
rect 701546 546301 701570 546314
rect 701614 546301 701638 546314
rect 701682 546301 701706 546314
rect 701750 546301 701774 546314
rect 701818 546301 701842 546314
rect 709211 546148 710211 546152
rect 707574 546099 707610 546134
rect 708610 546099 708646 546134
rect 707574 546098 708646 546099
rect 707574 546057 707610 546098
rect 708610 546057 708646 546098
rect 699322 545956 700322 546012
rect 700922 545956 701922 546012
rect 707574 546001 708646 546057
rect 707574 545964 707610 546001
rect 708610 545964 708646 546001
rect 707574 545959 708646 545964
rect 699322 545884 700322 545940
rect 700922 545884 701922 545940
rect 707574 545924 707610 545959
rect 708610 545924 708646 545959
rect 709175 546098 710247 546134
rect 709175 546057 709211 546098
rect 710211 546057 710247 546098
rect 709175 546001 710247 546057
rect 709175 545964 709211 546001
rect 710211 545964 710247 546001
rect 709175 545936 710247 545964
rect 709175 545924 709211 545936
rect 710211 545924 710247 545936
rect 707610 545713 708610 545785
rect 709211 545713 710211 545785
rect 699322 545623 700322 545673
rect 700922 545623 701922 545673
rect 707610 545523 708610 545617
rect 707610 545513 708644 545523
rect 709211 545513 710211 545591
rect 711541 545437 711629 550311
rect 713750 550136 714750 550264
rect 716417 550152 717417 550202
rect 711892 549049 711942 550049
rect 712062 549049 712112 550049
rect 713750 549920 714750 550048
rect 716417 549996 717417 550052
rect 716417 549846 717417 549896
rect 713750 549704 714750 549832
rect 716417 549730 717017 549780
rect 716417 549580 717017 549630
rect 713750 549488 714750 549544
rect 716417 549464 717417 549514
rect 713750 549272 714750 549400
rect 716417 549308 717417 549364
rect 713750 549056 714750 549184
rect 716417 549152 717417 549280
rect 716417 548996 717417 549052
rect 711892 547928 711942 548928
rect 712062 547928 712112 548928
rect 713750 548840 714750 548968
rect 716417 548840 717417 548968
rect 713750 548624 714750 548752
rect 716417 548684 717417 548740
rect 716417 548474 717417 548524
rect 713750 548408 714750 548464
rect 716417 548308 717417 548358
rect 713750 548192 714750 548248
rect 716417 548152 717417 548280
rect 713750 547976 714750 548104
rect 716417 547996 717417 548052
rect 711892 546807 711942 547807
rect 712062 546807 712112 547807
rect 713750 547760 714750 547888
rect 716417 547780 717417 547836
rect 713750 547544 714750 547672
rect 716417 547570 717417 547620
rect 713750 547328 714750 547456
rect 716417 547454 717417 547504
rect 716417 547298 717417 547426
rect 713750 547118 714750 547168
rect 716417 547148 717417 547198
rect 711892 545697 711942 546697
rect 712062 545697 712112 546697
rect 714686 546357 714794 546424
rect 714645 546323 714794 546357
rect 716071 546357 716074 546358
rect 716071 546356 716072 546357
rect 716073 546356 716074 546357
rect 716071 546355 716074 546356
rect 716208 546357 716211 546358
rect 716208 546356 716209 546357
rect 716210 546356 716211 546357
rect 716208 546355 716211 546356
rect 714964 546247 715998 546329
rect 716284 546247 717318 546329
rect 705107 545336 705173 545352
rect 711541 545302 711633 545437
rect 714175 545398 714225 545998
rect 714425 545398 714475 545998
rect 711579 545301 711595 545302
rect 714781 545191 714863 546226
rect 715134 545955 715828 546037
rect 714686 545123 714863 545191
rect 714645 545089 714863 545123
rect 680215 544880 680815 544936
rect 686719 544893 686739 544917
rect 686743 544893 686753 544917
rect 686719 544859 686757 544893
rect 686719 544822 686739 544859
rect 686743 544822 686753 544859
rect 692428 544850 693028 544978
rect 698017 544947 698210 544983
rect 698084 544935 698210 544947
rect 702756 544959 703645 544983
rect 702756 544935 702853 544959
rect 698084 544828 702853 544935
rect 686719 544788 686757 544822
rect 680215 544704 680815 544760
rect 686719 544751 686739 544788
rect 686743 544751 686753 544788
rect 686719 544741 686757 544751
rect 686699 544717 686767 544741
rect 686719 544704 686739 544717
rect 686743 544704 686753 544717
rect 686719 544695 686753 544704
rect 686719 544693 686743 544695
rect 692428 544694 693028 544750
rect 686685 544656 686709 544680
rect 686743 544656 686767 544680
rect 678799 544503 679399 544553
rect 680215 544534 680815 544584
rect 692428 544538 693028 544666
rect 680593 544531 680815 544534
rect 682009 544501 682069 544516
rect 682024 544465 682054 544501
rect 683708 544387 684308 544437
rect 678799 544327 679399 544383
rect 692428 544382 693028 544510
rect 683708 544237 684308 544287
rect 678799 544157 679399 544207
rect 685242 544187 686142 544320
rect 714781 544308 714863 545089
rect 715063 544609 715145 545915
rect 715342 545752 715382 545792
rect 715582 545752 715622 545792
rect 715289 544777 715339 545719
rect 715382 545668 715422 545752
rect 715542 545668 715582 545752
rect 715633 544777 715683 545719
rect 715382 544672 715422 544756
rect 715542 544672 715582 544756
rect 715342 544632 715382 544672
rect 715582 544632 715622 544672
rect 715815 544609 715897 545915
rect 715134 544387 715828 544469
rect 716100 544308 716182 546226
rect 716454 545955 717148 546037
rect 716385 544609 716467 545915
rect 716660 545752 716700 545792
rect 716900 545752 716940 545792
rect 716599 544777 716649 545719
rect 716700 545668 716740 545752
rect 716860 545668 716900 545752
rect 716943 544777 716993 545719
rect 716700 544672 716740 544756
rect 716860 544672 716900 544756
rect 716660 544632 716700 544672
rect 716900 544632 716940 544672
rect 717137 544609 717219 545915
rect 716454 544387 717148 544469
rect 717419 544308 717501 546226
rect 692428 544232 693028 544282
rect 684565 544160 684790 544168
rect 685242 544144 685808 544187
rect 696597 544000 696600 544120
rect 714964 544095 715998 544177
rect 716284 544095 717318 544177
rect 21000 517000 21003 517120
rect 282 516623 1316 516705
rect 1602 516623 2636 516705
rect 32810 516662 33035 516670
rect 38201 516593 38801 516643
rect 24572 516518 25172 516568
rect 33292 516513 33892 516563
rect 99 514574 181 516492
rect 452 516331 1146 516413
rect 381 514885 463 516191
rect 660 516128 700 516168
rect 900 516128 940 516168
rect 700 516044 740 516128
rect 860 516044 900 516128
rect 607 515081 657 516023
rect 951 515081 1001 516023
rect 1133 514885 1215 516191
rect 452 514763 1146 514845
rect 1418 514574 1500 516492
rect 1772 516331 2466 516413
rect 1703 514885 1785 516191
rect 1978 516128 2018 516168
rect 2218 516128 2258 516168
rect 2018 516044 2058 516128
rect 2178 516044 2218 516128
rect 1917 515081 1967 516023
rect 2261 515081 2311 516023
rect 2455 514885 2537 516191
rect 2737 515779 2819 516492
rect 24572 516362 25172 516490
rect 38201 516417 38801 516473
rect 33292 516363 33892 516413
rect 24572 516206 25172 516334
rect 35546 516299 35576 516335
rect 36785 516329 36935 516341
rect 35531 516284 35591 516299
rect 36785 516216 37385 516266
rect 38201 516247 38801 516297
rect 30833 516120 30857 516144
rect 30891 516120 30915 516144
rect 24572 516050 25172 516106
rect 30857 516105 30881 516107
rect 30857 516096 30887 516105
rect 30867 516083 30887 516096
rect 30891 516083 30907 516120
rect 30833 516059 30857 516083
rect 30867 516049 30911 516083
rect 14747 515865 19516 515972
rect 24572 515894 25172 516022
rect 30867 516012 30887 516049
rect 30891 516012 30907 516049
rect 36785 516040 37385 516096
rect 30867 515978 30911 516012
rect 30867 515941 30887 515978
rect 30891 515941 30907 515978
rect 30867 515907 30911 515941
rect 30867 515883 30887 515907
rect 30891 515883 30907 515907
rect 14747 515841 14844 515865
rect 13955 515817 14844 515841
rect 19390 515853 19516 515865
rect 19390 515841 19583 515853
rect 19390 515817 19605 515841
rect 19639 515817 19673 515841
rect 19707 515817 19741 515841
rect 19775 515817 19809 515841
rect 19843 515817 19877 515841
rect 19911 515817 19945 515841
rect 19979 515817 20013 515841
rect 20047 515817 20081 515841
rect 20115 515817 20149 515841
rect 20183 515817 20217 515841
rect 20251 515817 20285 515841
rect 20319 515817 20353 515841
rect 20387 515817 20421 515841
rect 20455 515817 20489 515841
rect 20523 515817 20557 515841
rect 20591 515817 20625 515841
rect 20659 515817 20693 515841
rect 2737 515711 2914 515779
rect 1772 514763 2466 514845
rect 2737 514574 2819 515711
rect 2848 515677 2955 515711
rect 19480 515540 19516 515817
rect 19547 515540 19583 515817
rect 24572 515738 25172 515866
rect 36785 515864 37385 515920
rect 36785 515688 37385 515744
rect 20809 515650 20833 515684
rect 20809 515582 20833 515616
rect 24572 515588 25172 515638
rect 20809 515540 20833 515548
rect 36785 515518 37385 515568
rect 3125 514802 3175 515402
rect 3375 514802 3425 515402
rect 282 514471 1316 514553
rect 1602 514471 2636 514553
rect 1389 514444 1392 514445
rect 1389 514443 1390 514444
rect 1391 514443 1392 514444
rect 1389 514442 1392 514443
rect 1526 514444 1529 514445
rect 1526 514443 1527 514444
rect 1528 514443 1529 514444
rect 2848 514443 2955 514477
rect 1526 514442 1529 514443
rect 5488 514280 5538 515103
rect 5658 514280 5708 515103
rect 6005 514280 6021 515499
rect 12427 515448 12493 515464
rect 24572 515458 25172 515508
rect 32930 515457 33530 515507
rect 35287 515391 35887 515441
rect 36785 515402 37385 515452
rect 24572 515308 25172 515358
rect 31463 515307 32063 515357
rect 32930 515301 33530 515357
rect 7389 515277 7406 515287
rect 7440 515277 7477 515287
rect 7511 515277 7551 515287
rect 7585 515277 7622 515287
rect 7656 515277 7696 515287
rect 7730 515277 7767 515287
rect 7801 515277 7841 515287
rect 7875 515277 7912 515287
rect 7946 515277 7986 515287
rect 8020 515277 8057 515287
rect 8091 515277 8131 515287
rect 8165 515277 8202 515287
rect 8236 515277 8296 515287
rect 8330 515277 8381 515287
rect 8996 515277 9044 515287
rect 9078 515277 9120 515287
rect 9154 515277 9197 515287
rect 9231 515277 9291 515287
rect 9325 515277 9362 515287
rect 9396 515277 9436 515287
rect 9470 515277 9507 515287
rect 9541 515277 9581 515287
rect 9615 515277 9652 515287
rect 9686 515277 9726 515287
rect 9760 515277 9797 515287
rect 9831 515277 9871 515287
rect 9905 515277 9942 515287
rect 9976 515277 9990 515287
rect 7389 515209 8389 515277
rect 8990 515183 9990 515277
rect 36785 515226 37385 515282
rect 15678 515127 16678 515177
rect 17278 515127 18278 515177
rect 31463 515151 32063 515207
rect 32930 515151 33530 515201
rect 34079 515157 34679 515207
rect 7389 514840 8389 514864
rect 15678 514860 16678 514916
rect 17278 514860 18278 514916
rect 8990 514840 9990 514841
rect 7389 514743 8389 514799
rect 8990 514743 9990 514799
rect 15678 514788 16678 514844
rect 17278 514788 18278 514844
rect 8990 514701 9990 514702
rect 15678 514286 16678 514426
rect 17278 514286 18278 514426
rect 19844 514280 19894 515051
rect 20462 514280 20512 515051
rect 31463 515001 32063 515051
rect 34079 515001 34679 515057
rect 35287 515039 35887 515095
rect 36785 515050 37385 515106
rect 32596 514929 33596 514979
rect 24573 514820 25173 514870
rect 34079 514851 34679 514901
rect 35287 514869 35887 514919
rect 36785 514880 37385 514930
rect 30171 514795 30771 514845
rect 32596 514773 33596 514829
rect 37993 514704 38593 514754
rect 30171 514619 30771 514675
rect 32596 514623 33596 514673
rect 34110 514589 34710 514639
rect 21263 514280 21313 514518
rect 22349 514280 22399 514518
rect 32596 514507 33596 514557
rect 30171 514449 30771 514499
rect 36785 514429 36985 514609
rect 37993 514534 38593 514584
rect 24573 514352 25173 514408
rect 29993 514310 30993 514360
rect 31347 514280 31547 514317
rect 31607 514280 31807 514317
rect 36785 514280 36985 514373
rect 37083 514280 37120 514373
rect 696597 508200 696600 508320
rect 692376 507983 692396 508017
rect 692463 507993 692532 508017
rect 696191 507993 696239 508017
rect 692487 507983 692532 507993
rect 696204 507983 696239 507993
rect 696340 507983 696360 508017
rect 692487 507915 692502 507939
rect 696200 507915 696215 507939
rect 692454 507891 692478 507915
rect 696224 507891 696248 507915
rect 686755 507800 687355 507850
rect 692487 507748 692505 507752
rect 692479 507718 692505 507748
rect 692487 507698 692505 507718
rect 686755 507624 687355 507680
rect 692485 507674 692505 507698
rect 692509 507674 692517 507718
rect 696215 507698 696223 507748
rect 696203 507674 696223 507698
rect 696227 507674 696245 507752
rect 692485 507640 692521 507674
rect 696203 507640 696249 507674
rect 686755 507448 687355 507504
rect 686755 507278 687355 507328
rect 685547 507102 686147 507152
rect 687155 507007 687170 507022
rect 687343 507018 687355 507022
rect 687340 507007 687355 507018
rect 685547 506932 686147 506982
rect 687155 506827 687355 507007
rect 687155 506812 687170 506827
rect 687340 506816 687355 506827
rect 687343 506812 687355 506816
rect 687042 506771 687057 506786
rect 687020 506591 687057 506771
rect 687155 506771 687170 506786
rect 687343 506782 687355 506786
rect 687340 506771 687355 506782
rect 687155 506591 687355 506771
rect 688210 506630 688260 507630
rect 688360 506740 688488 507630
rect 688516 506740 688644 507630
rect 688672 506740 688800 507630
rect 688828 506740 688956 507630
rect 688984 506740 689112 507630
rect 689140 506740 689268 507630
rect 689296 506740 689424 507630
rect 689452 506740 689580 507630
rect 689608 506740 689736 507630
rect 689764 506740 689892 507630
rect 689920 506740 690048 507630
rect 690076 506740 690204 507630
rect 690232 506740 690360 507630
rect 690388 506630 690438 507630
rect 692485 507606 692505 507640
rect 692509 507606 692517 507640
rect 696203 507606 696223 507640
rect 696227 507606 696245 507640
rect 691275 507523 691875 507573
rect 692485 507572 692521 507606
rect 696203 507572 696249 507606
rect 692485 507538 692505 507572
rect 692509 507538 692517 507572
rect 692485 507504 692521 507538
rect 692583 507528 693983 507571
rect 694719 507528 696119 507571
rect 696203 507538 696223 507572
rect 696227 507538 696245 507572
rect 696203 507504 696249 507538
rect 692485 507470 692505 507504
rect 692509 507470 692517 507504
rect 692485 507436 692521 507470
rect 691275 507373 691875 507423
rect 692485 507402 692505 507436
rect 692509 507402 692517 507436
rect 692485 507368 692521 507402
rect 692485 507334 692505 507368
rect 692509 507334 692517 507368
rect 692583 507365 693983 507493
rect 694719 507365 696119 507493
rect 696203 507470 696223 507504
rect 696227 507470 696245 507504
rect 696203 507436 696249 507470
rect 707624 507441 707658 507475
rect 707695 507441 707729 507475
rect 707769 507441 707803 507475
rect 707840 507441 707874 507475
rect 707914 507441 707948 507475
rect 707985 507441 708019 507475
rect 708059 507441 708093 507475
rect 708130 507441 708164 507475
rect 708204 507441 708238 507475
rect 708275 507441 708309 507475
rect 708369 507441 708403 507475
rect 708446 507441 708480 507475
rect 708520 507441 708554 507465
rect 708588 507441 708610 507465
rect 709211 507441 709234 507465
rect 709270 507441 709304 507475
rect 709364 507441 709398 507475
rect 709435 507441 709469 507475
rect 709509 507441 709543 507475
rect 709580 507441 709614 507475
rect 709654 507441 709688 507475
rect 709725 507441 709759 507475
rect 709799 507441 709833 507475
rect 709870 507441 709904 507475
rect 709944 507441 709978 507475
rect 710015 507441 710049 507475
rect 710089 507441 710123 507475
rect 710160 507441 710194 507475
rect 696203 507402 696223 507436
rect 696227 507402 696245 507436
rect 707610 507431 707624 507441
rect 707658 507431 707695 507441
rect 707729 507431 707769 507441
rect 707803 507431 707840 507441
rect 707874 507431 707914 507441
rect 707948 507431 707985 507441
rect 708019 507431 708059 507441
rect 708093 507431 708130 507441
rect 708164 507431 708204 507441
rect 708238 507431 708275 507441
rect 708309 507431 708369 507441
rect 708403 507431 708446 507441
rect 708480 507431 708520 507441
rect 708554 507431 708588 507441
rect 708610 507431 708634 507441
rect 709211 507431 709270 507441
rect 709304 507431 709364 507441
rect 709398 507431 709435 507441
rect 709469 507431 709509 507441
rect 709543 507431 709580 507441
rect 709614 507431 709654 507441
rect 709688 507431 709725 507441
rect 709759 507431 709799 507441
rect 709833 507431 709870 507441
rect 709904 507431 709944 507441
rect 709978 507431 710015 507441
rect 710049 507431 710089 507441
rect 710123 507431 710160 507441
rect 710194 507431 710211 507441
rect 696203 507368 696249 507402
rect 696203 507334 696223 507368
rect 696227 507334 696245 507368
rect 707610 507337 708610 507431
rect 709211 507337 710211 507431
rect 691275 507251 691875 507301
rect 692485 507300 692521 507334
rect 692485 507266 692505 507300
rect 692509 507266 692517 507300
rect 692485 507232 692521 507266
rect 692485 507198 692505 507232
rect 692509 507198 692517 507232
rect 692583 507202 693983 507330
rect 694719 507202 696119 507330
rect 696203 507300 696249 507334
rect 711579 507317 712463 507331
rect 711579 507307 711619 507317
rect 696203 507266 696223 507300
rect 696227 507266 696245 507300
rect 701730 507290 701747 507292
rect 696203 507232 696249 507266
rect 696203 507198 696223 507232
rect 696227 507198 696245 507232
rect 701692 507220 701722 507254
rect 701730 507220 701760 507290
rect 707610 507241 708610 507301
rect 709211 507241 710211 507301
rect 692485 507164 692521 507198
rect 691275 507101 691875 507151
rect 692485 507130 692505 507164
rect 692509 507130 692517 507164
rect 692485 507096 692521 507130
rect 692485 507062 692505 507096
rect 692509 507062 692517 507096
rect 692485 507028 692521 507062
rect 692583 507039 693983 507167
rect 694719 507039 696119 507167
rect 696203 507164 696249 507198
rect 696203 507130 696223 507164
rect 696227 507130 696245 507164
rect 696203 507096 696249 507130
rect 696203 507062 696223 507096
rect 696227 507062 696245 507096
rect 699322 507064 700322 507097
rect 700922 507064 701922 507097
rect 696203 507028 696249 507062
rect 707610 507044 708610 507048
rect 709211 507044 710211 507048
rect 691275 506975 691875 507025
rect 692485 506994 692505 507028
rect 692509 506994 692517 507028
rect 692485 506960 692521 506994
rect 692485 506926 692505 506960
rect 692509 506926 692517 506960
rect 692485 506892 692521 506926
rect 691275 506825 691875 506875
rect 692485 506858 692505 506892
rect 692509 506858 692517 506892
rect 692583 506876 693983 507004
rect 694719 506876 696119 507004
rect 696203 506994 696223 507028
rect 696227 506994 696245 507028
rect 707574 506994 708646 507030
rect 696203 506960 696249 506994
rect 696203 506926 696223 506960
rect 696227 506926 696245 506960
rect 707574 506953 707610 506994
rect 708610 506953 708646 506994
rect 696203 506892 696249 506926
rect 697284 506894 697350 506910
rect 707574 506897 708646 506953
rect 696203 506858 696223 506892
rect 696227 506858 696245 506892
rect 699322 506877 700322 506894
rect 700922 506877 701922 506894
rect 707574 506881 707610 506897
rect 708610 506881 708646 506897
rect 692485 506824 692521 506858
rect 692485 506790 692505 506824
rect 692509 506790 692517 506824
rect 692485 506756 692521 506790
rect 691275 506703 691875 506753
rect 692485 506740 692505 506756
rect 692509 506740 692517 506756
rect 692583 506740 693983 506841
rect 694719 506740 696119 506841
rect 696203 506824 696249 506858
rect 707574 506825 708646 506881
rect 696203 506790 696223 506824
rect 696227 506790 696245 506824
rect 696203 506756 696249 506790
rect 696203 506740 696223 506756
rect 696227 506740 696245 506756
rect 699322 506740 700322 506811
rect 700922 506740 701922 506811
rect 707574 506788 707610 506825
rect 708610 506788 708646 506825
rect 707574 506748 708646 506788
rect 709175 506994 710247 507030
rect 709175 506953 709211 506994
rect 710211 506953 710247 506994
rect 709175 506897 710247 506953
rect 709175 506881 709211 506897
rect 710211 506881 710247 506897
rect 709175 506825 710247 506881
rect 709175 506788 709211 506825
rect 710211 506788 710247 506825
rect 709175 506748 710247 506788
rect 685542 506506 686142 506556
rect 691275 506553 691875 506603
rect 685542 506330 686142 506386
rect 692583 506237 693983 506280
rect 694719 506237 696119 506280
rect 699322 506278 700322 506418
rect 700922 506278 701922 506418
rect 685542 506160 686142 506210
rect 692583 506101 693983 506144
rect 694719 506101 696119 506144
rect 680215 505678 680815 505728
rect 680215 505502 680815 505558
rect 685551 505516 686551 505566
rect 689154 505480 689204 505897
rect 689304 505480 689360 505897
rect 689460 505480 689516 505897
rect 689616 505480 689672 505897
rect 689772 505480 689828 505897
rect 689928 505480 689978 505897
rect 699322 505860 700322 505916
rect 700922 505860 701922 505916
rect 707610 505905 708610 505961
rect 709211 505905 710211 505961
rect 699322 505788 700322 505844
rect 700922 505788 701922 505844
rect 707610 505833 708610 505889
rect 709211 505833 710211 505889
rect 711579 505525 711605 507307
rect 715956 506297 716006 507297
rect 716106 506740 716234 507297
rect 716262 506297 716312 507297
rect 711579 505480 711595 505495
rect 712409 505480 712431 505485
rect 713640 505480 713641 505785
rect 713750 505772 714750 505822
rect 713750 505562 714750 505612
rect 713750 505480 714750 505496
rect 2850 503304 3850 503320
rect 2850 503188 3850 503238
rect 2850 502978 3850 503028
rect 3959 503015 3960 503320
rect 5169 503315 5191 503320
rect 6005 503305 6021 503320
rect 1288 501503 1338 502503
rect 1438 501503 1566 502060
rect 1594 501503 1644 502503
rect 5995 501493 6021 503275
rect 7389 502911 8389 502967
rect 8990 502911 9990 502967
rect 15678 502956 16678 503012
rect 17278 502956 18278 503012
rect 7389 502839 8389 502895
rect 8990 502839 9990 502895
rect 15678 502884 16678 502940
rect 17278 502884 18278 502940
rect 27622 502903 27672 503320
rect 27772 502903 27828 503320
rect 27928 502903 27984 503320
rect 28084 502903 28140 503320
rect 28240 502903 28296 503320
rect 28396 502903 28446 503320
rect 31049 503234 32049 503284
rect 36785 503242 37385 503298
rect 36785 503072 37385 503122
rect 21481 502656 22881 502699
rect 23617 502656 25017 502699
rect 31458 502590 32058 502640
rect 15678 502382 16678 502522
rect 17278 502382 18278 502522
rect 21481 502520 22881 502563
rect 23617 502520 25017 502563
rect 31458 502414 32058 502470
rect 25725 502197 26325 502247
rect 31458 502244 32058 502294
rect 7353 502016 8425 502052
rect 7353 501975 7389 502016
rect 8389 501975 8425 502016
rect 7353 501919 8425 501975
rect 7353 501903 7389 501919
rect 8389 501903 8425 501919
rect 7353 501847 8425 501903
rect 7353 501810 7389 501847
rect 8389 501810 8425 501847
rect 7353 501770 8425 501810
rect 8954 502016 10026 502052
rect 8954 501975 8990 502016
rect 9990 501975 10026 502016
rect 8954 501919 10026 501975
rect 21383 502044 21403 502060
rect 21407 502044 21415 502060
rect 21383 502010 21419 502044
rect 21481 502031 22881 502060
rect 23617 502031 25017 502060
rect 25101 502044 25121 502060
rect 25125 502044 25143 502060
rect 25725 502047 26325 502097
rect 25101 502010 25147 502044
rect 21383 501976 21403 502010
rect 21407 501976 21415 502010
rect 21383 501942 21419 501976
rect 8954 501903 8990 501919
rect 9990 501903 10026 501919
rect 15678 501906 16678 501923
rect 17278 501906 18278 501923
rect 21383 501908 21403 501942
rect 21407 501908 21415 501942
rect 8954 501847 10026 501903
rect 20250 501890 20316 501906
rect 8954 501810 8990 501847
rect 9990 501810 10026 501847
rect 8954 501770 10026 501810
rect 21383 501874 21419 501908
rect 21383 501840 21403 501874
rect 21407 501840 21415 501874
rect 21481 501868 22881 501996
rect 23617 501868 25017 501996
rect 25101 501976 25121 502010
rect 25125 501976 25143 502010
rect 25101 501942 25147 501976
rect 25101 501908 25121 501942
rect 25125 501908 25143 501942
rect 25725 501925 26325 501975
rect 25101 501874 25147 501908
rect 25101 501840 25121 501874
rect 25125 501840 25143 501874
rect 21383 501806 21419 501840
rect 21383 501772 21403 501806
rect 21407 501772 21415 501806
rect 21383 501738 21419 501772
rect 15678 501703 16678 501736
rect 17278 501703 18278 501736
rect 21383 501704 21403 501738
rect 21407 501704 21415 501738
rect 21481 501705 22881 501833
rect 23617 501705 25017 501833
rect 25101 501806 25147 501840
rect 25101 501772 25121 501806
rect 25125 501772 25143 501806
rect 25725 501775 26325 501825
rect 25101 501738 25147 501772
rect 25101 501704 25121 501738
rect 25125 501704 25143 501738
rect 21383 501670 21419 501704
rect 25101 501670 25147 501704
rect 21383 501636 21403 501670
rect 21407 501636 21415 501670
rect 7389 501559 8389 501631
rect 8990 501559 9990 501631
rect 21383 501602 21419 501636
rect 15840 501510 15870 501580
rect 15878 501546 15908 501580
rect 21383 501568 21403 501602
rect 21407 501568 21415 501602
rect 15853 501508 15870 501510
rect 21383 501534 21419 501568
rect 21481 501542 22881 501670
rect 23617 501542 25017 501670
rect 25101 501636 25121 501670
rect 25125 501636 25143 501670
rect 25725 501649 26325 501699
rect 25101 501602 25147 501636
rect 25101 501568 25121 501602
rect 25125 501568 25143 501602
rect 25101 501534 25147 501568
rect 5981 501483 6021 501493
rect 5137 501469 6021 501483
rect 21383 501500 21403 501534
rect 21407 501500 21415 501534
rect 21383 501466 21419 501500
rect 7389 501369 8389 501463
rect 7389 501359 8413 501369
rect 8990 501359 9990 501463
rect 21383 501432 21403 501466
rect 21407 501432 21415 501466
rect 21383 501398 21419 501432
rect 21383 501364 21403 501398
rect 21407 501364 21415 501398
rect 21481 501379 22881 501507
rect 23617 501379 25017 501507
rect 25101 501500 25121 501534
rect 25125 501500 25143 501534
rect 25101 501466 25147 501500
rect 25725 501499 26325 501549
rect 25101 501432 25121 501466
rect 25125 501432 25143 501466
rect 25101 501398 25147 501432
rect 25101 501364 25121 501398
rect 25125 501364 25143 501398
rect 25725 501377 26325 501427
rect 21383 501330 21419 501364
rect 25101 501330 25147 501364
rect 21383 501296 21403 501330
rect 21407 501296 21415 501330
rect 25101 501296 25121 501330
rect 25125 501296 25143 501330
rect 21383 501262 21419 501296
rect 21383 501228 21403 501262
rect 21407 501228 21415 501262
rect 21481 501229 22881 501272
rect 23617 501229 25017 501272
rect 25101 501262 25147 501296
rect 25101 501228 25121 501262
rect 25125 501228 25143 501262
rect 21383 501194 21419 501228
rect 25101 501194 25147 501228
rect 25725 501227 26325 501277
rect 21383 501160 21403 501194
rect 21407 501160 21415 501194
rect 25101 501160 25121 501194
rect 25125 501160 25143 501194
rect 27162 501170 27212 502170
rect 27312 501170 27440 502060
rect 27468 501170 27596 502060
rect 27624 501170 27752 502060
rect 27780 501170 27908 502060
rect 27936 501170 28064 502060
rect 28092 501170 28220 502060
rect 28248 501170 28376 502060
rect 28404 501170 28532 502060
rect 28560 501170 28688 502060
rect 28716 501170 28844 502060
rect 28872 501170 29000 502060
rect 29028 501170 29156 502060
rect 29184 501170 29312 502060
rect 29340 501170 29390 502170
rect 30245 502029 30445 502209
rect 30245 502018 30260 502029
rect 30245 502014 30257 502018
rect 30430 502014 30445 502029
rect 30543 502029 30580 502209
rect 30543 502014 30558 502029
rect 30245 501984 30257 501988
rect 30245 501973 30260 501984
rect 30430 501973 30445 501988
rect 30245 501793 30445 501973
rect 31453 501818 32053 501868
rect 30245 501782 30260 501793
rect 30245 501778 30257 501782
rect 30430 501778 30445 501793
rect 31453 501648 32053 501698
rect 30245 501472 30845 501522
rect 30245 501296 30845 501352
rect 21383 501126 21419 501160
rect 25101 501126 25147 501160
rect 21383 501102 21403 501126
rect 21385 501048 21403 501102
rect 21407 501082 21415 501126
rect 25101 501102 25121 501126
rect 25113 501082 25121 501102
rect 25125 501048 25143 501126
rect 30245 501120 30845 501176
rect 30245 500950 30845 501000
rect 21000 500800 21003 500920
rect 21352 500885 21376 500909
rect 25122 500885 25146 500909
rect 21385 500861 21400 500885
rect 25098 500861 25113 500885
rect 21274 500783 21294 500851
rect 21410 500817 21430 500851
rect 25068 500817 25088 500851
rect 25204 500817 25224 500851
rect 21385 500807 21430 500817
rect 25102 500807 25137 500817
rect 21361 500783 21430 500807
rect 25089 500783 25137 500807
rect 25238 500783 25258 500817
rect 680480 494427 680517 494520
rect 680615 494427 680815 494520
rect 685793 494483 685993 494520
rect 686053 494483 686253 494520
rect 686607 494440 687607 494490
rect 692427 494392 693027 494448
rect 679007 494216 679607 494266
rect 680615 494191 680815 494371
rect 686829 494301 687429 494351
rect 684004 494243 685004 494293
rect 695201 494282 695251 494520
rect 696287 494282 696337 494520
rect 682890 494161 683490 494211
rect 684004 494127 685004 494177
rect 686829 494125 687429 494181
rect 679007 494046 679607 494096
rect 684004 493971 685004 494027
rect 686829 493955 687429 494005
rect 680215 493870 680815 493920
rect 681713 493881 682313 493931
rect 682921 493899 683521 493949
rect 692427 493930 693027 493980
rect 684004 493821 685004 493871
rect 680215 493694 680815 493750
rect 681713 493705 682313 493761
rect 682921 493743 683521 493799
rect 685537 493749 686137 493799
rect 697088 493749 697138 494520
rect 697706 493749 697756 494520
rect 699322 494374 700322 494514
rect 700922 494374 701922 494514
rect 707610 494098 708610 494099
rect 699322 493956 700322 494012
rect 700922 493956 701922 494012
rect 707610 494001 708610 494057
rect 709211 494001 710211 494057
rect 707610 493959 708610 493960
rect 699322 493884 700322 493940
rect 700922 493884 701922 493940
rect 709211 493936 710211 493960
rect 682921 493593 683521 493643
rect 684070 493599 684670 493649
rect 685537 493593 686137 493649
rect 699322 493623 700322 493673
rect 700922 493623 701922 493673
rect 680215 493518 680815 493574
rect 707610 493523 708610 493617
rect 709211 493523 710211 493591
rect 707610 493513 707624 493523
rect 707658 493513 707695 493523
rect 707729 493513 707769 493523
rect 707803 493513 707840 493523
rect 707874 493513 707914 493523
rect 707948 493513 707985 493523
rect 708019 493513 708059 493523
rect 708093 493513 708130 493523
rect 708164 493513 708204 493523
rect 708238 493513 708275 493523
rect 708309 493513 708369 493523
rect 708403 493513 708446 493523
rect 708480 493513 708522 493523
rect 708556 493513 708604 493523
rect 709219 493513 709270 493523
rect 709304 493513 709364 493523
rect 709398 493513 709435 493523
rect 709469 493513 709509 493523
rect 709543 493513 709580 493523
rect 709614 493513 709654 493523
rect 709688 493513 709725 493523
rect 709759 493513 709799 493523
rect 709833 493513 709870 493523
rect 709904 493513 709944 493523
rect 709978 493513 710015 493523
rect 710049 493513 710089 493523
rect 710123 493513 710160 493523
rect 710194 493513 710211 493523
rect 684070 493443 684670 493499
rect 685537 493443 686137 493493
rect 692428 493442 693028 493492
rect 680215 493348 680815 493398
rect 681713 493359 682313 493409
rect 684070 493293 684670 493343
rect 692428 493292 693028 493342
rect 705107 493336 705173 493352
rect 711579 493301 711595 494520
rect 711892 493697 711942 494520
rect 712062 493697 712112 494520
rect 716071 494357 716074 494358
rect 714645 494323 714752 494357
rect 716071 494356 716072 494357
rect 716073 494356 716074 494357
rect 716071 494355 716074 494356
rect 716208 494357 716211 494358
rect 716208 494356 716209 494357
rect 716210 494356 716211 494357
rect 716208 494355 716211 494356
rect 714964 494247 715998 494329
rect 716284 494247 717318 494329
rect 714175 493398 714225 493998
rect 714425 493398 714475 493998
rect 680215 493232 680815 493282
rect 698017 493232 698053 493260
rect 692428 493162 693028 493212
rect 698030 493198 698077 493232
rect 698017 493164 698053 493198
rect 680215 493056 680815 493112
rect 692428 493006 693028 493134
rect 698030 493130 698077 493164
rect 698017 493096 698053 493130
rect 698030 493062 698077 493096
rect 698017 492983 698053 493062
rect 698084 492983 698120 493260
rect 714781 493191 714863 494226
rect 715134 493955 715828 494037
rect 714686 493123 714863 493191
rect 714645 493089 714863 493123
rect 680215 492880 680815 492936
rect 686719 492893 686739 492917
rect 686743 492893 686753 492917
rect 686719 492859 686757 492893
rect 686719 492822 686739 492859
rect 686743 492822 686753 492859
rect 692428 492850 693028 492978
rect 698017 492947 698210 492983
rect 698084 492935 698210 492947
rect 702756 492959 703645 492983
rect 702756 492935 702853 492959
rect 698084 492828 702853 492935
rect 686719 492788 686757 492822
rect 680215 492704 680815 492760
rect 686719 492751 686739 492788
rect 686743 492751 686753 492788
rect 686719 492741 686757 492751
rect 686699 492717 686767 492741
rect 686719 492704 686739 492717
rect 686743 492704 686753 492717
rect 686719 492695 686753 492704
rect 686719 492693 686743 492695
rect 692428 492694 693028 492750
rect 686685 492656 686709 492680
rect 686743 492656 686767 492680
rect 678799 492503 679399 492553
rect 680215 492534 680815 492584
rect 692428 492538 693028 492666
rect 680593 492531 680815 492534
rect 682009 492501 682069 492516
rect 682024 492465 682054 492501
rect 683708 492387 684308 492437
rect 678799 492327 679399 492383
rect 692428 492382 693028 492510
rect 714781 492308 714863 493089
rect 715063 492609 715145 493915
rect 715289 492777 715339 493719
rect 715633 492777 715683 493719
rect 715382 492672 715422 492756
rect 715542 492672 715582 492756
rect 715342 492632 715382 492672
rect 715582 492632 715622 492672
rect 715815 492609 715897 493915
rect 715134 492387 715828 492469
rect 716100 492308 716182 494226
rect 716454 493955 717148 494037
rect 716385 492609 716467 493915
rect 716599 492777 716649 493719
rect 716943 492777 716993 493719
rect 716700 492672 716740 492756
rect 716860 492672 716900 492756
rect 716660 492632 716700 492672
rect 716900 492632 716940 492672
rect 717137 492609 717219 493915
rect 716454 492387 717148 492469
rect 717419 492308 717501 494226
rect 683708 492237 684308 492287
rect 692428 492232 693028 492282
rect 678799 492157 679399 492207
rect 684565 492160 684790 492168
rect 696597 492000 696600 492120
rect 714964 492095 715998 492177
rect 716284 492095 717318 492177
rect 21000 465000 21003 465120
rect 282 464623 1316 464705
rect 1602 464623 2636 464705
rect 32810 464662 33035 464670
rect 38201 464593 38801 464643
rect 24572 464518 25172 464568
rect 33292 464513 33892 464563
rect 99 462574 181 464492
rect 452 464331 1146 464413
rect 381 462885 463 464191
rect 660 464128 700 464168
rect 900 464128 940 464168
rect 700 464044 740 464128
rect 860 464044 900 464128
rect 607 463081 657 464023
rect 700 463048 740 463132
rect 860 463048 900 463132
rect 951 463081 1001 464023
rect 660 463008 700 463048
rect 900 463008 940 463048
rect 1133 462885 1215 464191
rect 452 462763 1146 462845
rect 1418 462574 1500 464492
rect 1772 464331 2466 464413
rect 1703 462885 1785 464191
rect 1978 464128 2018 464168
rect 2218 464128 2258 464168
rect 2018 464044 2058 464128
rect 2178 464044 2218 464128
rect 1917 463081 1967 464023
rect 2018 463048 2058 463132
rect 2178 463048 2218 463132
rect 2261 463081 2311 464023
rect 1978 463008 2018 463048
rect 2218 463008 2258 463048
rect 2455 462885 2537 464191
rect 2737 463779 2819 464492
rect 24572 464362 25172 464490
rect 38201 464417 38801 464473
rect 33292 464363 33892 464413
rect 24572 464206 25172 464334
rect 35546 464299 35576 464335
rect 36785 464329 36935 464341
rect 35531 464284 35591 464299
rect 36785 464216 37385 464266
rect 38201 464247 38801 464297
rect 30833 464120 30857 464144
rect 30891 464120 30915 464144
rect 24572 464050 25172 464106
rect 30857 464105 30881 464107
rect 30857 464096 30887 464105
rect 30867 464083 30887 464096
rect 30891 464083 30907 464120
rect 30833 464059 30857 464083
rect 30867 464049 30911 464083
rect 14747 463865 19516 463972
rect 24572 463894 25172 464022
rect 30867 464012 30887 464049
rect 30891 464012 30907 464049
rect 36785 464040 37385 464096
rect 30867 463978 30911 464012
rect 30867 463941 30887 463978
rect 30891 463941 30907 463978
rect 30867 463907 30911 463941
rect 30867 463883 30887 463907
rect 30891 463883 30907 463907
rect 14747 463841 14844 463865
rect 13955 463817 14844 463841
rect 19390 463853 19516 463865
rect 19390 463841 19583 463853
rect 19390 463817 19605 463841
rect 19639 463817 19673 463841
rect 19707 463817 19741 463841
rect 19775 463817 19809 463841
rect 19843 463817 19877 463841
rect 19911 463817 19945 463841
rect 19979 463817 20013 463841
rect 20047 463817 20081 463841
rect 20115 463817 20149 463841
rect 20183 463817 20217 463841
rect 20251 463817 20285 463841
rect 20319 463817 20353 463841
rect 20387 463817 20421 463841
rect 20455 463817 20489 463841
rect 20523 463817 20557 463841
rect 20591 463817 20625 463841
rect 20659 463817 20693 463841
rect 2737 463711 2914 463779
rect 1772 462763 2466 462845
rect 2737 462574 2819 463711
rect 2848 463677 2955 463711
rect 6005 463498 6021 463499
rect 3125 462802 3175 463402
rect 3375 462802 3425 463402
rect 5967 463363 6059 463498
rect 12427 463448 12493 463464
rect 282 462471 1316 462553
rect 1602 462471 2636 462553
rect 2806 462477 2914 462545
rect 1389 462444 1392 462445
rect 1389 462443 1390 462444
rect 1391 462443 1392 462444
rect 1389 462442 1392 462443
rect 1526 462444 1529 462445
rect 1526 462443 1527 462444
rect 1528 462443 1529 462444
rect 2848 462443 2955 462477
rect 1526 462442 1529 462443
rect 5488 462103 5538 463103
rect 5658 462103 5708 463103
rect 183 461602 1183 461652
rect 2850 461632 3850 461682
rect 183 461446 1183 461574
rect 2850 461416 3850 461544
rect 183 461296 1183 461346
rect 183 461180 1183 461230
rect 2850 461200 3850 461328
rect 183 460964 1183 461020
rect 2850 460984 3850 461112
rect 5488 460993 5538 461993
rect 5658 460993 5708 461993
rect 183 460748 1183 460804
rect 2850 460768 3850 460896
rect 183 460592 1183 460720
rect 2850 460552 3850 460608
rect 183 460442 1183 460492
rect 2850 460336 3850 460392
rect 183 460276 1183 460326
rect 2850 460120 3850 460248
rect 183 460060 1183 460116
rect 183 459904 1183 460032
rect 2850 459904 3850 460032
rect 5488 459872 5538 460872
rect 5658 459872 5708 460872
rect 183 459748 1183 459804
rect 183 459592 1183 459720
rect 2850 459688 3850 459816
rect 183 459436 1183 459492
rect 2850 459472 3850 459600
rect 183 459286 1183 459336
rect 2850 459256 3850 459312
rect 583 459170 1183 459220
rect 583 459020 1183 459070
rect 2850 459040 3850 459168
rect 183 458904 1183 458954
rect 2850 458824 3850 458952
rect 183 458748 1183 458804
rect 5488 458751 5538 459751
rect 5658 458751 5708 459751
rect 183 458598 1183 458648
rect 2850 458608 3850 458736
rect 5971 458489 6059 463363
rect 7406 463287 7440 463321
rect 7477 463287 7511 463321
rect 7551 463287 7585 463321
rect 7622 463287 7656 463321
rect 7696 463287 7730 463321
rect 7767 463287 7801 463321
rect 7841 463287 7875 463321
rect 7912 463287 7946 463321
rect 7986 463287 8020 463321
rect 8057 463287 8091 463321
rect 8131 463287 8165 463321
rect 8202 463287 8236 463321
rect 8296 463287 8330 463321
rect 8381 463311 8423 463321
rect 8381 463287 8389 463311
rect 8415 463287 8423 463311
rect 8956 463311 8996 463321
rect 8956 463287 8962 463311
rect 8990 463287 8996 463311
rect 9044 463287 9078 463321
rect 9120 463287 9154 463321
rect 9197 463287 9231 463321
rect 9291 463287 9325 463321
rect 9362 463287 9396 463321
rect 9436 463287 9470 463321
rect 9507 463287 9541 463321
rect 9581 463287 9615 463321
rect 9652 463287 9686 463321
rect 9726 463287 9760 463321
rect 9797 463287 9831 463321
rect 9871 463287 9905 463321
rect 9942 463287 9976 463321
rect 7389 463277 7406 463287
rect 7440 463277 7477 463287
rect 7511 463277 7551 463287
rect 7585 463277 7622 463287
rect 7656 463277 7696 463287
rect 7730 463277 7767 463287
rect 7801 463277 7841 463287
rect 7875 463277 7912 463287
rect 7946 463277 7986 463287
rect 8020 463277 8057 463287
rect 8091 463277 8131 463287
rect 8165 463277 8202 463287
rect 8236 463277 8296 463287
rect 8330 463277 8381 463287
rect 8389 463277 8423 463287
rect 8990 463277 9044 463287
rect 9078 463277 9120 463287
rect 9154 463277 9197 463287
rect 9231 463277 9291 463287
rect 9325 463277 9362 463287
rect 9396 463277 9436 463287
rect 9470 463277 9507 463287
rect 9541 463277 9581 463287
rect 9615 463277 9652 463287
rect 9686 463277 9726 463287
rect 9760 463277 9797 463287
rect 9831 463277 9871 463287
rect 9905 463277 9942 463287
rect 9976 463277 9990 463287
rect 7389 463209 8389 463277
rect 8990 463183 9990 463277
rect 7389 463087 8389 463147
rect 8990 463087 9990 463147
rect 15678 463127 16678 463177
rect 17278 463127 18278 463177
rect 7353 462864 7389 462876
rect 8389 462864 8425 462876
rect 7353 462840 8425 462864
rect 7353 462799 7389 462840
rect 8389 462799 8425 462840
rect 7353 462743 8425 462799
rect 7353 462706 7389 462743
rect 8389 462706 8425 462743
rect 7353 462666 8425 462706
rect 8954 462841 8990 462876
rect 9990 462841 10026 462876
rect 15678 462860 16678 462916
rect 17278 462860 18278 462916
rect 8954 462840 10026 462841
rect 8954 462799 8990 462840
rect 9990 462799 10026 462840
rect 8954 462743 10026 462799
rect 15678 462788 16678 462844
rect 17278 462788 18278 462844
rect 8954 462706 8990 462743
rect 9990 462706 10026 462743
rect 8954 462701 10026 462706
rect 8954 462666 8990 462701
rect 9990 462666 10026 462701
rect 7389 462441 8389 462513
rect 8990 462441 9990 462513
rect 15678 462486 16678 462558
rect 17278 462486 18278 462558
rect 15748 462475 15782 462486
rect 15816 462475 15850 462486
rect 15884 462475 15918 462486
rect 15952 462475 15986 462486
rect 16020 462475 16054 462486
rect 16088 462475 16122 462486
rect 16156 462475 16190 462486
rect 16224 462475 16258 462486
rect 16292 462475 16326 462486
rect 16360 462475 16394 462486
rect 16428 462475 16462 462486
rect 16496 462475 16530 462486
rect 16564 462475 16598 462486
rect 16632 462475 16666 462486
rect 17290 462475 17324 462486
rect 17358 462475 17392 462486
rect 17426 462475 17460 462486
rect 17494 462475 17528 462486
rect 17562 462475 17596 462486
rect 17630 462475 17664 462486
rect 17698 462475 17732 462486
rect 17766 462475 17800 462486
rect 17834 462475 17868 462486
rect 17902 462475 17936 462486
rect 17970 462475 18004 462486
rect 18038 462475 18072 462486
rect 18106 462475 18140 462486
rect 18174 462475 18208 462486
rect 15748 462465 15806 462475
rect 15816 462465 15874 462475
rect 15884 462465 15942 462475
rect 15952 462465 16010 462475
rect 16020 462465 16078 462475
rect 16088 462465 16146 462475
rect 16156 462465 16214 462475
rect 16224 462465 16282 462475
rect 16292 462465 16350 462475
rect 16360 462465 16418 462475
rect 16428 462465 16486 462475
rect 16496 462465 16554 462475
rect 16564 462465 16622 462475
rect 16632 462465 16690 462475
rect 17290 462465 17348 462475
rect 17358 462465 17416 462475
rect 17426 462465 17484 462475
rect 17494 462465 17552 462475
rect 17562 462465 17620 462475
rect 17630 462465 17688 462475
rect 17698 462465 17756 462475
rect 17766 462465 17824 462475
rect 17834 462465 17892 462475
rect 17902 462465 17960 462475
rect 17970 462465 18028 462475
rect 18038 462465 18096 462475
rect 18106 462465 18164 462475
rect 18174 462465 18232 462475
rect 15724 462441 16690 462465
rect 17266 462441 18232 462465
rect 15748 462426 15772 462441
rect 15816 462426 15840 462441
rect 15884 462426 15908 462441
rect 15952 462426 15976 462441
rect 16020 462426 16044 462441
rect 16088 462426 16112 462441
rect 16156 462426 16180 462441
rect 16224 462426 16248 462441
rect 16292 462426 16316 462441
rect 16360 462426 16384 462441
rect 16428 462426 16452 462441
rect 16496 462426 16520 462441
rect 16564 462426 16588 462441
rect 16632 462426 16656 462441
rect 17290 462426 17314 462441
rect 17358 462426 17382 462441
rect 17426 462426 17450 462441
rect 17494 462426 17518 462441
rect 17562 462426 17586 462441
rect 17630 462426 17654 462441
rect 17698 462426 17722 462441
rect 17766 462426 17790 462441
rect 17834 462426 17858 462441
rect 17902 462426 17926 462441
rect 17970 462426 17994 462441
rect 18038 462426 18062 462441
rect 18106 462426 18130 462441
rect 18174 462426 18198 462441
rect 15678 462271 16678 462426
rect 7389 462181 8389 462241
rect 8990 462181 9990 462241
rect 15678 462237 16690 462271
rect 17278 462261 18278 462426
rect 17266 462237 18278 462261
rect 15678 462226 16678 462237
rect 17278 462226 18278 462237
rect 15748 462213 15772 462226
rect 15816 462213 15840 462226
rect 15884 462213 15908 462226
rect 15952 462213 15976 462226
rect 16020 462213 16044 462226
rect 16088 462213 16112 462226
rect 16156 462213 16180 462226
rect 16224 462213 16248 462226
rect 16292 462213 16316 462226
rect 16360 462213 16384 462226
rect 16428 462213 16452 462226
rect 16496 462213 16520 462226
rect 16564 462213 16588 462226
rect 16632 462213 16656 462226
rect 17290 462213 17314 462226
rect 17358 462213 17382 462226
rect 17426 462213 17450 462226
rect 17494 462213 17518 462226
rect 17562 462213 17586 462226
rect 17630 462213 17654 462226
rect 17698 462213 17722 462226
rect 17766 462213 17790 462226
rect 17834 462213 17858 462226
rect 17902 462213 17926 462226
rect 17970 462213 17994 462226
rect 18038 462213 18062 462226
rect 18106 462213 18130 462226
rect 18174 462213 18198 462226
rect 7389 461823 8389 461879
rect 8990 461823 9990 461879
rect 15678 461868 16678 461924
rect 17278 461868 18278 461924
rect 7389 461751 8389 461807
rect 8990 461751 9990 461807
rect 15678 461796 16678 461852
rect 17278 461796 18278 461852
rect 7389 461449 8389 461521
rect 8990 461449 9990 461521
rect 15678 461494 16678 461566
rect 17278 461494 18278 461566
rect 15748 461483 15782 461494
rect 15816 461483 15850 461494
rect 15884 461483 15918 461494
rect 15952 461483 15986 461494
rect 16020 461483 16054 461494
rect 16088 461483 16122 461494
rect 16156 461483 16190 461494
rect 16224 461483 16258 461494
rect 16292 461483 16326 461494
rect 16360 461483 16394 461494
rect 16428 461483 16462 461494
rect 16496 461483 16530 461494
rect 16564 461483 16598 461494
rect 16632 461483 16666 461494
rect 17290 461483 17324 461494
rect 17358 461483 17392 461494
rect 17426 461483 17460 461494
rect 17494 461483 17528 461494
rect 17562 461483 17596 461494
rect 17630 461483 17664 461494
rect 17698 461483 17732 461494
rect 17766 461483 17800 461494
rect 17834 461483 17868 461494
rect 17902 461483 17936 461494
rect 17970 461483 18004 461494
rect 18038 461483 18072 461494
rect 18106 461483 18140 461494
rect 18174 461483 18208 461494
rect 15748 461473 15806 461483
rect 15816 461473 15874 461483
rect 15884 461473 15942 461483
rect 15952 461473 16010 461483
rect 16020 461473 16078 461483
rect 16088 461473 16146 461483
rect 16156 461473 16214 461483
rect 16224 461473 16282 461483
rect 16292 461473 16350 461483
rect 16360 461473 16418 461483
rect 16428 461473 16486 461483
rect 16496 461473 16554 461483
rect 16564 461473 16622 461483
rect 16632 461473 16690 461483
rect 17290 461473 17348 461483
rect 17358 461473 17416 461483
rect 17426 461473 17484 461483
rect 17494 461473 17552 461483
rect 17562 461473 17620 461483
rect 17630 461473 17688 461483
rect 17698 461473 17756 461483
rect 17766 461473 17824 461483
rect 17834 461473 17892 461483
rect 17902 461473 17960 461483
rect 17970 461473 18028 461483
rect 18038 461473 18096 461483
rect 18106 461473 18164 461483
rect 18174 461473 18232 461483
rect 15724 461449 16690 461473
rect 17266 461449 18232 461473
rect 12427 461424 12493 461440
rect 15748 461434 15772 461449
rect 15816 461434 15840 461449
rect 15884 461434 15908 461449
rect 15952 461434 15976 461449
rect 16020 461434 16044 461449
rect 16088 461434 16112 461449
rect 16156 461434 16180 461449
rect 16224 461434 16248 461449
rect 16292 461434 16316 461449
rect 16360 461434 16384 461449
rect 16428 461434 16452 461449
rect 16496 461434 16520 461449
rect 16564 461434 16588 461449
rect 16632 461434 16656 461449
rect 17290 461434 17314 461449
rect 17358 461434 17382 461449
rect 17426 461434 17450 461449
rect 17494 461434 17518 461449
rect 17562 461434 17586 461449
rect 17630 461434 17654 461449
rect 17698 461434 17722 461449
rect 17766 461434 17790 461449
rect 17834 461434 17858 461449
rect 17902 461434 17926 461449
rect 17970 461434 17994 461449
rect 18038 461434 18062 461449
rect 18106 461434 18130 461449
rect 18174 461434 18198 461449
rect 15678 461279 16678 461434
rect 7389 461189 8389 461249
rect 8990 461189 9990 461249
rect 15678 461245 16690 461279
rect 17278 461269 18278 461434
rect 17266 461245 18278 461269
rect 15678 461234 16678 461245
rect 17278 461234 18278 461245
rect 15748 461221 15772 461234
rect 15816 461221 15840 461234
rect 15884 461221 15908 461234
rect 15952 461221 15976 461234
rect 16020 461221 16044 461234
rect 16088 461221 16112 461234
rect 16156 461221 16180 461234
rect 16224 461221 16248 461234
rect 16292 461221 16316 461234
rect 16360 461221 16384 461234
rect 16428 461221 16452 461234
rect 16496 461221 16520 461234
rect 16564 461221 16588 461234
rect 16632 461221 16656 461234
rect 17290 461221 17314 461234
rect 17358 461221 17382 461234
rect 17426 461221 17450 461234
rect 17494 461221 17518 461234
rect 17562 461221 17586 461234
rect 17630 461221 17654 461234
rect 17698 461221 17722 461234
rect 17766 461221 17790 461234
rect 17834 461221 17858 461234
rect 17902 461221 17926 461234
rect 17970 461221 17994 461234
rect 18038 461221 18062 461234
rect 18106 461221 18130 461234
rect 18174 461221 18198 461234
rect 7389 460831 8389 460887
rect 8990 460831 9990 460887
rect 15678 460876 16678 460932
rect 17278 460876 18278 460932
rect 7389 460759 8389 460815
rect 8990 460759 9990 460815
rect 15678 460804 16678 460860
rect 17278 460804 18278 460860
rect 7389 460457 8389 460529
rect 8990 460457 9990 460529
rect 15678 460502 16678 460574
rect 17278 460502 18278 460574
rect 15748 460491 15782 460502
rect 15816 460491 15850 460502
rect 15884 460491 15918 460502
rect 15952 460491 15986 460502
rect 16020 460491 16054 460502
rect 16088 460491 16122 460502
rect 16156 460491 16190 460502
rect 16224 460491 16258 460502
rect 16292 460491 16326 460502
rect 16360 460491 16394 460502
rect 16428 460491 16462 460502
rect 16496 460491 16530 460502
rect 16564 460491 16598 460502
rect 16632 460491 16666 460502
rect 17290 460491 17324 460502
rect 17358 460491 17392 460502
rect 17426 460491 17460 460502
rect 17494 460491 17528 460502
rect 17562 460491 17596 460502
rect 17630 460491 17664 460502
rect 17698 460491 17732 460502
rect 17766 460491 17800 460502
rect 17834 460491 17868 460502
rect 17902 460491 17936 460502
rect 17970 460491 18004 460502
rect 18038 460491 18072 460502
rect 18106 460491 18140 460502
rect 18174 460491 18208 460502
rect 15748 460481 15806 460491
rect 15816 460481 15874 460491
rect 15884 460481 15942 460491
rect 15952 460481 16010 460491
rect 16020 460481 16078 460491
rect 16088 460481 16146 460491
rect 16156 460481 16214 460491
rect 16224 460481 16282 460491
rect 16292 460481 16350 460491
rect 16360 460481 16418 460491
rect 16428 460481 16486 460491
rect 16496 460481 16554 460491
rect 16564 460481 16622 460491
rect 16632 460481 16690 460491
rect 17290 460481 17348 460491
rect 17358 460481 17416 460491
rect 17426 460481 17484 460491
rect 17494 460481 17552 460491
rect 17562 460481 17620 460491
rect 17630 460481 17688 460491
rect 17698 460481 17756 460491
rect 17766 460481 17824 460491
rect 17834 460481 17892 460491
rect 17902 460481 17960 460491
rect 17970 460481 18028 460491
rect 18038 460481 18096 460491
rect 18106 460481 18164 460491
rect 18174 460481 18232 460491
rect 15724 460457 16690 460481
rect 17266 460457 18232 460481
rect 15748 460442 15772 460457
rect 15816 460442 15840 460457
rect 15884 460442 15908 460457
rect 15952 460442 15976 460457
rect 16020 460442 16044 460457
rect 16088 460442 16112 460457
rect 16156 460442 16180 460457
rect 16224 460442 16248 460457
rect 16292 460442 16316 460457
rect 16360 460442 16384 460457
rect 16428 460442 16452 460457
rect 16496 460442 16520 460457
rect 16564 460442 16588 460457
rect 16632 460442 16656 460457
rect 17290 460442 17314 460457
rect 17358 460442 17382 460457
rect 17426 460442 17450 460457
rect 17494 460442 17518 460457
rect 17562 460442 17586 460457
rect 17630 460442 17654 460457
rect 17698 460442 17722 460457
rect 17766 460442 17790 460457
rect 17834 460442 17858 460457
rect 17902 460442 17926 460457
rect 17970 460442 17994 460457
rect 18038 460442 18062 460457
rect 18106 460442 18130 460457
rect 18174 460442 18198 460457
rect 15678 460287 16678 460442
rect 7389 460197 8389 460257
rect 8990 460197 9990 460257
rect 15678 460253 16690 460287
rect 17278 460277 18278 460442
rect 17266 460253 18278 460277
rect 15678 460242 16678 460253
rect 17278 460242 18278 460253
rect 15748 460229 15772 460242
rect 15816 460229 15840 460242
rect 15884 460229 15908 460242
rect 15952 460229 15976 460242
rect 16020 460229 16044 460242
rect 16088 460229 16112 460242
rect 16156 460229 16180 460242
rect 16224 460229 16248 460242
rect 16292 460229 16316 460242
rect 16360 460229 16384 460242
rect 16428 460229 16452 460242
rect 16496 460229 16520 460242
rect 16564 460229 16588 460242
rect 16632 460229 16656 460242
rect 17290 460229 17314 460242
rect 17358 460229 17382 460242
rect 17426 460229 17450 460242
rect 17494 460229 17518 460242
rect 17562 460229 17586 460242
rect 17630 460229 17654 460242
rect 17698 460229 17722 460242
rect 17766 460229 17790 460242
rect 17834 460229 17858 460242
rect 17902 460229 17926 460242
rect 17970 460229 17994 460242
rect 18038 460229 18062 460242
rect 18106 460229 18130 460242
rect 18174 460229 18198 460242
rect 7389 459839 8389 459895
rect 8990 459839 9990 459895
rect 15678 459884 16678 459940
rect 17278 459884 18278 459940
rect 7389 459767 8389 459823
rect 8990 459767 9990 459823
rect 15678 459812 16678 459868
rect 17278 459812 18278 459868
rect 7389 459465 8389 459537
rect 8990 459465 9990 459537
rect 15678 459510 16678 459582
rect 17278 459510 18278 459582
rect 15748 459499 15782 459510
rect 15816 459499 15850 459510
rect 15884 459499 15918 459510
rect 15952 459499 15986 459510
rect 16020 459499 16054 459510
rect 16088 459499 16122 459510
rect 16156 459499 16190 459510
rect 16224 459499 16258 459510
rect 16292 459499 16326 459510
rect 16360 459499 16394 459510
rect 16428 459499 16462 459510
rect 16496 459499 16530 459510
rect 16564 459499 16598 459510
rect 16632 459499 16666 459510
rect 17290 459499 17324 459510
rect 17358 459499 17392 459510
rect 17426 459499 17460 459510
rect 17494 459499 17528 459510
rect 17562 459499 17596 459510
rect 17630 459499 17664 459510
rect 17698 459499 17732 459510
rect 17766 459499 17800 459510
rect 17834 459499 17868 459510
rect 17902 459499 17936 459510
rect 17970 459499 18004 459510
rect 18038 459499 18072 459510
rect 18106 459499 18140 459510
rect 18174 459499 18208 459510
rect 15748 459489 15806 459499
rect 15816 459489 15874 459499
rect 15884 459489 15942 459499
rect 15952 459489 16010 459499
rect 16020 459489 16078 459499
rect 16088 459489 16146 459499
rect 16156 459489 16214 459499
rect 16224 459489 16282 459499
rect 16292 459489 16350 459499
rect 16360 459489 16418 459499
rect 16428 459489 16486 459499
rect 16496 459489 16554 459499
rect 16564 459489 16622 459499
rect 16632 459489 16690 459499
rect 17290 459489 17348 459499
rect 17358 459489 17416 459499
rect 17426 459489 17484 459499
rect 17494 459489 17552 459499
rect 17562 459489 17620 459499
rect 17630 459489 17688 459499
rect 17698 459489 17756 459499
rect 17766 459489 17824 459499
rect 17834 459489 17892 459499
rect 17902 459489 17960 459499
rect 17970 459489 18028 459499
rect 18038 459489 18096 459499
rect 18106 459489 18164 459499
rect 18174 459489 18232 459499
rect 15724 459465 16690 459489
rect 17266 459465 18232 459489
rect 15748 459450 15772 459465
rect 15816 459450 15840 459465
rect 15884 459450 15908 459465
rect 15952 459450 15976 459465
rect 16020 459450 16044 459465
rect 16088 459450 16112 459465
rect 16156 459450 16180 459465
rect 16224 459450 16248 459465
rect 16292 459450 16316 459465
rect 16360 459450 16384 459465
rect 16428 459450 16452 459465
rect 16496 459450 16520 459465
rect 16564 459450 16588 459465
rect 16632 459450 16656 459465
rect 17290 459450 17314 459465
rect 17358 459450 17382 459465
rect 17426 459450 17450 459465
rect 17494 459450 17518 459465
rect 17562 459450 17586 459465
rect 17630 459450 17654 459465
rect 17698 459450 17722 459465
rect 17766 459450 17790 459465
rect 17834 459450 17858 459465
rect 17902 459450 17926 459465
rect 17970 459450 17994 459465
rect 18038 459450 18062 459465
rect 18106 459450 18130 459465
rect 18174 459450 18198 459465
rect 15678 459295 16678 459450
rect 7389 459205 8389 459265
rect 8990 459205 9990 459265
rect 15678 459261 16690 459295
rect 17278 459285 18278 459450
rect 17266 459261 18278 459285
rect 15678 459250 16678 459261
rect 17278 459250 18278 459261
rect 15748 459237 15772 459250
rect 15816 459237 15840 459250
rect 15884 459237 15908 459250
rect 15952 459237 15976 459250
rect 16020 459237 16044 459250
rect 16088 459237 16112 459250
rect 16156 459237 16180 459250
rect 16224 459237 16248 459250
rect 16292 459237 16316 459250
rect 16360 459237 16384 459250
rect 16428 459237 16452 459250
rect 16496 459237 16520 459250
rect 16564 459237 16588 459250
rect 16632 459237 16656 459250
rect 17290 459237 17314 459250
rect 17358 459237 17382 459250
rect 17426 459237 17450 459250
rect 17494 459237 17518 459250
rect 17562 459237 17586 459250
rect 17630 459237 17654 459250
rect 17698 459237 17722 459250
rect 17766 459237 17790 459250
rect 17834 459237 17858 459250
rect 17902 459237 17926 459250
rect 17970 459237 17994 459250
rect 18038 459237 18062 459250
rect 18106 459237 18130 459250
rect 18174 459237 18198 459250
rect 7389 458847 8389 458903
rect 8990 458847 9990 458903
rect 15678 458892 16678 458948
rect 17278 458892 18278 458948
rect 7389 458775 8389 458831
rect 8990 458775 9990 458831
rect 15678 458820 16678 458876
rect 17278 458820 18278 458876
rect 5967 458455 6059 458489
rect 7389 458473 8389 458545
rect 8990 458473 9990 458545
rect 15678 458518 16678 458590
rect 17278 458518 18278 458590
rect 15748 458507 15782 458518
rect 15816 458507 15850 458518
rect 15884 458507 15918 458518
rect 15952 458507 15986 458518
rect 16020 458507 16054 458518
rect 16088 458507 16122 458518
rect 16156 458507 16190 458518
rect 16224 458507 16258 458518
rect 16292 458507 16326 458518
rect 16360 458507 16394 458518
rect 16428 458507 16462 458518
rect 16496 458507 16530 458518
rect 16564 458507 16598 458518
rect 16632 458507 16666 458518
rect 17290 458507 17324 458518
rect 17358 458507 17392 458518
rect 17426 458507 17460 458518
rect 17494 458507 17528 458518
rect 17562 458507 17596 458518
rect 17630 458507 17664 458518
rect 17698 458507 17732 458518
rect 17766 458507 17800 458518
rect 17834 458507 17868 458518
rect 17902 458507 17936 458518
rect 17970 458507 18004 458518
rect 18038 458507 18072 458518
rect 18106 458507 18140 458518
rect 18174 458507 18208 458518
rect 15748 458497 15806 458507
rect 15816 458497 15874 458507
rect 15884 458497 15942 458507
rect 15952 458497 16010 458507
rect 16020 458497 16078 458507
rect 16088 458497 16146 458507
rect 16156 458497 16214 458507
rect 16224 458497 16282 458507
rect 16292 458497 16350 458507
rect 16360 458497 16418 458507
rect 16428 458497 16486 458507
rect 16496 458497 16554 458507
rect 16564 458497 16622 458507
rect 16632 458497 16690 458507
rect 17290 458497 17348 458507
rect 17358 458497 17416 458507
rect 17426 458497 17484 458507
rect 17494 458497 17552 458507
rect 17562 458497 17620 458507
rect 17630 458497 17688 458507
rect 17698 458497 17756 458507
rect 17766 458497 17824 458507
rect 17834 458497 17892 458507
rect 17902 458497 17960 458507
rect 17970 458497 18028 458507
rect 18038 458497 18096 458507
rect 18106 458497 18164 458507
rect 18174 458497 18232 458507
rect 15724 458473 16690 458497
rect 17266 458473 18232 458497
rect 15748 458458 15772 458473
rect 15816 458458 15840 458473
rect 15884 458458 15908 458473
rect 15952 458458 15976 458473
rect 16020 458458 16044 458473
rect 16088 458458 16112 458473
rect 16156 458458 16180 458473
rect 16224 458458 16248 458473
rect 16292 458458 16316 458473
rect 16360 458458 16384 458473
rect 16428 458458 16452 458473
rect 16496 458458 16520 458473
rect 16564 458458 16588 458473
rect 16632 458458 16656 458473
rect 17290 458458 17314 458473
rect 17358 458458 17382 458473
rect 17426 458458 17450 458473
rect 17494 458458 17518 458473
rect 17562 458458 17586 458473
rect 17630 458458 17654 458473
rect 17698 458458 17722 458473
rect 17766 458458 17790 458473
rect 17834 458458 17858 458473
rect 17902 458458 17926 458473
rect 17970 458458 17994 458473
rect 18038 458458 18062 458473
rect 18106 458458 18130 458473
rect 18174 458458 18198 458473
rect 2850 458398 3850 458448
rect 2850 458282 3850 458332
rect 2850 458072 3850 458122
rect 2850 457956 3850 458006
rect 2850 457746 3850 457796
rect 1153 457660 1187 457718
rect 2850 457630 3850 457680
rect 2850 457420 3850 457470
rect 2850 457417 3107 457420
rect 3250 457304 3850 457354
rect 3250 457048 3850 457104
rect 3250 456892 3850 457020
rect 175 456818 1175 456868
rect 175 456662 1175 456790
rect 3250 456736 3850 456792
rect 175 456506 1175 456634
rect 175 456350 1175 456478
rect 175 456194 1175 456322
rect 175 456044 1175 456094
rect 175 455928 1175 455978
rect 175 455772 1175 455828
rect 175 455622 1175 455672
rect 1578 455609 1628 456609
rect 1728 455609 1856 456609
rect 1884 455609 2012 456609
rect 2040 455609 2090 456609
rect 3250 456580 3850 456708
rect 3250 456430 3850 456480
rect 2850 456314 3850 456364
rect 2850 456158 3850 456214
rect 2850 456008 3850 456058
rect 2850 455880 3850 455930
rect 2850 455724 3850 455852
rect 2850 455568 3850 455696
rect 175 455506 1175 455556
rect 175 455350 1175 455478
rect 2850 455412 3850 455468
rect 2850 455256 3850 455384
rect 175 455194 1175 455250
rect 175 455038 1175 455166
rect 175 454888 1175 454938
rect 175 454772 1175 454822
rect 175 454616 1175 454744
rect 1578 454613 1628 455213
rect 1728 454613 1784 455213
rect 1884 454613 1940 455213
rect 2040 454613 2096 455213
rect 2196 454613 2246 455213
rect 2850 455100 3850 455228
rect 2850 454944 3850 455072
rect 2850 454794 3850 454844
rect 2850 454678 3850 454728
rect 2850 454522 3850 454650
rect 175 454460 1175 454516
rect 175 454304 1175 454432
rect 2850 454366 3850 454494
rect 2850 454210 3850 454338
rect 175 454154 1175 454204
rect 803 454151 1175 454154
rect 2850 454054 3850 454110
rect 2850 453898 3850 454026
rect 2850 453742 3850 453870
rect 2850 453586 3850 453642
rect 2850 453436 3850 453486
rect 3926 453455 3960 453491
rect 3967 453339 3989 453455
rect 1638 451869 1688 452869
rect 1848 451869 1976 452869
rect 2064 451869 2114 452869
rect 2850 452275 3050 452287
rect 2850 452162 3850 452212
rect 2850 451946 3850 452074
rect 2850 451730 3850 451786
rect 2850 451514 3850 451642
rect 2850 451304 3850 451354
rect 2850 451188 3850 451238
rect 2850 450978 3850 451028
rect 3926 451015 3960 453339
rect 5169 451315 5191 458429
rect 5488 457194 5538 458194
rect 5658 457194 5708 458194
rect 5488 456073 5538 457073
rect 5658 456073 5708 457073
rect 5488 454952 5538 455952
rect 5658 454952 5708 455952
rect 5488 453842 5538 454842
rect 5658 453842 5708 454842
rect 5488 452721 5538 453721
rect 5658 452721 5708 453721
rect 5488 451600 5538 452600
rect 5658 451600 5708 452600
rect 5971 451386 6059 458455
rect 15678 458303 16678 458458
rect 7389 458213 8389 458273
rect 8990 458213 9990 458273
rect 15678 458269 16690 458303
rect 17278 458293 18278 458458
rect 17266 458269 18278 458293
rect 15678 458258 16678 458269
rect 17278 458258 18278 458269
rect 15748 458245 15772 458258
rect 15816 458245 15840 458258
rect 15884 458245 15908 458258
rect 15952 458245 15976 458258
rect 16020 458245 16044 458258
rect 16088 458245 16112 458258
rect 16156 458245 16180 458258
rect 16224 458245 16248 458258
rect 16292 458245 16316 458258
rect 16360 458245 16384 458258
rect 16428 458245 16452 458258
rect 16496 458245 16520 458258
rect 16564 458245 16588 458258
rect 16632 458245 16656 458258
rect 17290 458245 17314 458258
rect 17358 458245 17382 458258
rect 17426 458245 17450 458258
rect 17494 458245 17518 458258
rect 17562 458245 17586 458258
rect 17630 458245 17654 458258
rect 17698 458245 17722 458258
rect 17766 458245 17790 458258
rect 17834 458245 17858 458258
rect 17902 458245 17926 458258
rect 17970 458245 17994 458258
rect 18038 458245 18062 458258
rect 18106 458245 18130 458258
rect 18174 458245 18198 458258
rect 7389 457855 8389 457911
rect 8990 457855 9990 457911
rect 15678 457900 16678 457956
rect 17278 457900 18278 457956
rect 7389 457783 8389 457839
rect 8990 457783 9990 457839
rect 15678 457828 16678 457884
rect 17278 457828 18278 457884
rect 7389 457481 8389 457553
rect 8990 457481 9990 457553
rect 15678 457526 16678 457598
rect 17278 457526 18278 457598
rect 15748 457515 15782 457526
rect 15816 457515 15850 457526
rect 15884 457515 15918 457526
rect 15952 457515 15986 457526
rect 16020 457515 16054 457526
rect 16088 457515 16122 457526
rect 16156 457515 16190 457526
rect 16224 457515 16258 457526
rect 16292 457515 16326 457526
rect 16360 457515 16394 457526
rect 16428 457515 16462 457526
rect 16496 457515 16530 457526
rect 16564 457515 16598 457526
rect 16632 457515 16666 457526
rect 17290 457515 17324 457526
rect 17358 457515 17392 457526
rect 17426 457515 17460 457526
rect 17494 457515 17528 457526
rect 17562 457515 17596 457526
rect 17630 457515 17664 457526
rect 17698 457515 17732 457526
rect 17766 457515 17800 457526
rect 17834 457515 17868 457526
rect 17902 457515 17936 457526
rect 17970 457515 18004 457526
rect 18038 457515 18072 457526
rect 18106 457515 18140 457526
rect 18174 457515 18208 457526
rect 15748 457505 15806 457515
rect 15816 457505 15874 457515
rect 15884 457505 15942 457515
rect 15952 457505 16010 457515
rect 16020 457505 16078 457515
rect 16088 457505 16146 457515
rect 16156 457505 16214 457515
rect 16224 457505 16282 457515
rect 16292 457505 16350 457515
rect 16360 457505 16418 457515
rect 16428 457505 16486 457515
rect 16496 457505 16554 457515
rect 16564 457505 16622 457515
rect 16632 457505 16690 457515
rect 17290 457505 17348 457515
rect 17358 457505 17416 457515
rect 17426 457505 17484 457515
rect 17494 457505 17552 457515
rect 17562 457505 17620 457515
rect 17630 457505 17688 457515
rect 17698 457505 17756 457515
rect 17766 457505 17824 457515
rect 17834 457505 17892 457515
rect 17902 457505 17960 457515
rect 17970 457505 18028 457515
rect 18038 457505 18096 457515
rect 18106 457505 18164 457515
rect 18174 457505 18232 457515
rect 15724 457481 16690 457505
rect 17266 457481 18232 457505
rect 15748 457466 15772 457481
rect 15816 457466 15840 457481
rect 15884 457466 15908 457481
rect 15952 457466 15976 457481
rect 16020 457466 16044 457481
rect 16088 457466 16112 457481
rect 16156 457466 16180 457481
rect 16224 457466 16248 457481
rect 16292 457466 16316 457481
rect 16360 457466 16384 457481
rect 16428 457466 16452 457481
rect 16496 457466 16520 457481
rect 16564 457466 16588 457481
rect 16632 457466 16656 457481
rect 17290 457466 17314 457481
rect 17358 457466 17382 457481
rect 17426 457466 17450 457481
rect 17494 457466 17518 457481
rect 17562 457466 17586 457481
rect 17630 457466 17654 457481
rect 17698 457466 17722 457481
rect 17766 457466 17790 457481
rect 17834 457466 17858 457481
rect 17902 457466 17926 457481
rect 17970 457466 17994 457481
rect 18038 457466 18062 457481
rect 18106 457466 18130 457481
rect 18174 457466 18198 457481
rect 15678 457311 16678 457466
rect 7389 457221 8389 457281
rect 8990 457221 9990 457281
rect 15678 457277 16690 457311
rect 17278 457301 18278 457466
rect 17266 457277 18278 457301
rect 15678 457266 16678 457277
rect 17278 457266 18278 457277
rect 15748 457253 15772 457266
rect 15816 457253 15840 457266
rect 15884 457253 15908 457266
rect 15952 457253 15976 457266
rect 16020 457253 16044 457266
rect 16088 457253 16112 457266
rect 16156 457253 16180 457266
rect 16224 457253 16248 457266
rect 16292 457253 16316 457266
rect 16360 457253 16384 457266
rect 16428 457253 16452 457266
rect 16496 457253 16520 457266
rect 16564 457253 16588 457266
rect 16632 457253 16656 457266
rect 17290 457253 17314 457266
rect 17358 457253 17382 457266
rect 17426 457253 17450 457266
rect 17494 457253 17518 457266
rect 17562 457253 17586 457266
rect 17630 457253 17654 457266
rect 17698 457253 17722 457266
rect 17766 457253 17790 457266
rect 17834 457253 17858 457266
rect 17902 457253 17926 457266
rect 17970 457253 17994 457266
rect 18038 457253 18062 457266
rect 18106 457253 18130 457266
rect 18174 457253 18198 457266
rect 7389 456863 8389 456919
rect 8990 456863 9990 456919
rect 15678 456908 16678 456964
rect 17278 456908 18278 456964
rect 7389 456791 8389 456847
rect 8990 456791 9990 456847
rect 15678 456836 16678 456892
rect 17278 456836 18278 456892
rect 19480 456867 19516 463817
rect 19547 456867 19583 463817
rect 24572 463738 25172 463866
rect 36785 463864 37385 463920
rect 36785 463688 37385 463744
rect 20809 463650 20833 463684
rect 20809 463582 20833 463616
rect 24572 463588 25172 463638
rect 20809 463514 20833 463548
rect 36785 463518 37385 463568
rect 20809 463446 20833 463480
rect 24572 463458 25172 463508
rect 32930 463457 33530 463507
rect 20809 463378 20833 463412
rect 35287 463391 35887 463441
rect 36785 463402 37385 463452
rect 20809 463310 20833 463344
rect 24572 463308 25172 463358
rect 31463 463307 32063 463357
rect 32930 463301 33530 463357
rect 20809 463242 20833 463276
rect 35287 463215 35887 463343
rect 36785 463226 37385 463282
rect 20809 463174 20833 463208
rect 31463 463151 32063 463207
rect 32930 463151 33530 463201
rect 34079 463157 34679 463207
rect 20809 463106 20833 463140
rect 19844 462051 19894 463051
rect 19994 462051 20122 463051
rect 20150 462051 20278 463051
rect 20306 462051 20434 463051
rect 20462 462051 20512 463051
rect 20809 463038 20833 463072
rect 20809 462970 20833 463004
rect 20973 463000 21007 463024
rect 21041 463000 21075 463024
rect 21109 463000 21143 463024
rect 21177 463000 21211 463024
rect 21245 463000 21279 463024
rect 21313 463000 21347 463024
rect 21381 463000 21415 463024
rect 21449 463000 21483 463024
rect 21517 463000 21551 463024
rect 21585 463000 21619 463024
rect 21653 463000 21687 463024
rect 21721 463000 21755 463024
rect 21789 463000 21823 463024
rect 21857 463000 21891 463024
rect 21925 463000 21959 463024
rect 21993 463000 22027 463024
rect 22061 463000 22095 463024
rect 22129 463000 22163 463024
rect 22197 463000 22210 463024
rect 31463 463001 32063 463051
rect 34079 463001 34679 463057
rect 35287 463039 35887 463095
rect 36785 463050 37385 463106
rect 20809 462902 20833 462936
rect 32596 462929 33596 462979
rect 20809 462834 20833 462868
rect 24573 462820 25173 462870
rect 34079 462851 34679 462901
rect 35287 462869 35887 462919
rect 36785 462880 37385 462930
rect 35287 462866 35559 462869
rect 35716 462866 35887 462869
rect 20809 462766 20833 462800
rect 30171 462795 30771 462845
rect 20809 462698 20833 462732
rect 24573 462664 25173 462792
rect 32596 462773 33596 462829
rect 37993 462704 38593 462754
rect 19844 460521 19894 461921
rect 19994 460521 20122 461921
rect 20150 460521 20278 461921
rect 20306 460521 20434 461921
rect 20462 460521 20512 461921
rect 20809 460219 20833 460253
rect 19844 458759 19894 460159
rect 19994 458759 20122 460159
rect 20150 458759 20278 460159
rect 20306 458759 20434 460159
rect 20462 458759 20512 460159
rect 20809 460151 20833 460185
rect 20809 460083 20833 460117
rect 20809 460015 20833 460049
rect 20809 459947 20833 459981
rect 20809 459879 20833 459913
rect 20809 459811 20833 459845
rect 20809 459743 20833 459777
rect 20809 459675 20833 459709
rect 20809 459607 20833 459641
rect 20809 459539 20833 459573
rect 21263 459518 21313 462518
rect 21413 459518 21541 462518
rect 21569 459518 21697 462518
rect 21725 459518 21853 462518
rect 21881 459518 22009 462518
rect 22037 459518 22165 462518
rect 22193 459518 22321 462518
rect 22349 459518 22399 462518
rect 24573 462508 25173 462636
rect 30171 462619 30771 462675
rect 32596 462623 33596 462673
rect 34110 462589 34710 462639
rect 36785 462620 36797 462624
rect 36785 462609 36800 462620
rect 36970 462609 36985 462624
rect 26348 462530 26372 462564
rect 32596 462507 33596 462557
rect 26348 462461 26372 462495
rect 30171 462449 30771 462499
rect 24573 462352 25173 462408
rect 24573 462196 25173 462324
rect 29993 462310 30993 462360
rect 32596 462351 33596 462479
rect 34110 462433 34710 462561
rect 36785 462429 36985 462609
rect 37993 462534 38593 462584
rect 36785 462418 36800 462429
rect 36785 462414 36797 462418
rect 36970 462414 36985 462429
rect 31347 462317 31362 462332
rect 31535 462328 31547 462332
rect 31532 462317 31547 462328
rect 24573 462040 25173 462168
rect 26490 462122 26690 462172
rect 29993 462160 30993 462210
rect 31347 462137 31547 462317
rect 31347 462122 31362 462137
rect 31532 462126 31547 462137
rect 31535 462122 31547 462126
rect 31607 462317 31622 462332
rect 31795 462328 31807 462332
rect 31792 462317 31807 462328
rect 31607 462137 31807 462317
rect 32596 462195 33596 462323
rect 34110 462277 34710 462405
rect 36785 462384 36797 462388
rect 36785 462373 36800 462384
rect 36970 462373 36985 462388
rect 31607 462122 31622 462137
rect 31792 462126 31807 462137
rect 31795 462122 31807 462126
rect 31347 462081 31362 462096
rect 31535 462092 31547 462096
rect 31532 462081 31547 462092
rect 22906 461855 23212 462025
rect 23406 461855 23712 462025
rect 26490 461966 26690 462022
rect 29993 462001 30993 462051
rect 24573 461890 25173 461940
rect 31347 461901 31547 462081
rect 26490 461816 26690 461866
rect 29993 461851 30993 461901
rect 31347 461886 31362 461901
rect 31532 461890 31547 461901
rect 31535 461886 31547 461890
rect 31607 462081 31622 462096
rect 31795 462092 31807 462096
rect 31792 462081 31807 462092
rect 31607 461901 31807 462081
rect 32596 462039 33596 462167
rect 34110 462121 34710 462249
rect 36785 462193 36985 462373
rect 36785 462182 36800 462193
rect 36785 462178 36797 462182
rect 36970 462178 36985 462193
rect 37083 462373 37098 462388
rect 37083 462193 37120 462373
rect 37083 462178 37098 462193
rect 37998 462108 38598 462158
rect 34110 461971 34710 462021
rect 31607 461886 31622 461901
rect 31792 461890 31807 461901
rect 31795 461886 31807 461890
rect 32596 461883 33596 461939
rect 37998 461932 38598 461988
rect 34110 461855 34710 461905
rect 24573 461760 25173 461810
rect 27691 461682 28291 461732
rect 30253 461721 30268 461736
rect 30441 461732 30453 461736
rect 30438 461721 30453 461732
rect 24573 461610 25173 461660
rect 27691 461532 28291 461582
rect 30253 461541 30453 461721
rect 30253 461526 30268 461541
rect 30438 461530 30453 461541
rect 30441 461526 30453 461530
rect 30513 461721 30528 461736
rect 30701 461732 30713 461736
rect 30698 461721 30713 461732
rect 30513 461541 30713 461721
rect 30513 461526 30528 461541
rect 30698 461530 30713 461541
rect 30701 461526 30713 461530
rect 30773 461721 30788 461736
rect 30961 461732 30973 461736
rect 30958 461721 30973 461732
rect 30773 461541 30973 461721
rect 30773 461526 30788 461541
rect 30958 461530 30973 461541
rect 30961 461526 30973 461530
rect 31087 461721 31102 461736
rect 31275 461732 31287 461736
rect 31272 461721 31287 461732
rect 31087 461541 31287 461721
rect 31087 461526 31102 461541
rect 31272 461530 31287 461541
rect 31275 461526 31287 461530
rect 31347 461721 31362 461736
rect 31535 461732 31547 461736
rect 31532 461721 31547 461732
rect 31347 461541 31547 461721
rect 31347 461526 31362 461541
rect 31532 461530 31547 461541
rect 31535 461526 31547 461530
rect 31607 461721 31622 461736
rect 31795 461732 31807 461736
rect 31792 461721 31807 461732
rect 31607 461541 31807 461721
rect 31607 461526 31622 461541
rect 31792 461530 31807 461541
rect 31795 461526 31807 461530
rect 31867 461721 31882 461736
rect 32055 461732 32067 461736
rect 32052 461721 32067 461732
rect 32596 461727 33596 461855
rect 31867 461541 32067 461721
rect 34110 461699 34710 461827
rect 37998 461762 38598 461812
rect 37998 461759 38220 461762
rect 38245 461759 38539 461762
rect 32596 461571 33596 461699
rect 34110 461543 34710 461671
rect 31867 461526 31882 461541
rect 32052 461530 32067 461541
rect 32055 461526 32067 461530
rect 22619 461446 22647 461474
rect 24573 461438 25173 461488
rect 26490 461416 26690 461466
rect 27691 461402 28291 461452
rect 32596 461415 33596 461543
rect 34110 461387 34710 461515
rect 24573 461288 25173 461338
rect 26490 461260 26690 461316
rect 27691 461246 28291 461374
rect 30253 461361 30268 461376
rect 30441 461372 30453 461376
rect 30438 461361 30453 461372
rect 30253 461331 30453 461361
rect 30253 461316 30268 461331
rect 30438 461320 30453 461331
rect 30441 461316 30453 461320
rect 30513 461361 30528 461376
rect 30701 461372 30713 461376
rect 30698 461361 30713 461372
rect 30513 461331 30713 461361
rect 30513 461316 30528 461331
rect 30698 461320 30713 461331
rect 30701 461316 30713 461320
rect 30773 461361 30788 461376
rect 31347 461361 31362 461376
rect 31535 461372 31547 461376
rect 31532 461361 31547 461372
rect 30773 461331 30793 461361
rect 31347 461331 31547 461361
rect 30773 461316 30788 461331
rect 31347 461316 31362 461331
rect 31532 461320 31547 461331
rect 31535 461316 31547 461320
rect 31607 461361 31622 461376
rect 31795 461372 31807 461376
rect 31792 461361 31807 461372
rect 31607 461331 31807 461361
rect 31607 461316 31622 461331
rect 31792 461320 31807 461331
rect 31795 461316 31807 461320
rect 31867 461361 31882 461376
rect 31867 461331 31921 461361
rect 31867 461316 31882 461331
rect 30253 461275 30268 461290
rect 30441 461286 30453 461290
rect 30438 461275 30453 461286
rect 30253 461245 30453 461275
rect 30253 461230 30268 461245
rect 30438 461234 30453 461245
rect 30441 461230 30453 461234
rect 30513 461275 30528 461290
rect 30701 461286 30713 461290
rect 30698 461275 30713 461286
rect 30513 461245 30713 461275
rect 30513 461230 30528 461245
rect 30698 461234 30713 461245
rect 30701 461230 30713 461234
rect 30773 461275 30788 461290
rect 31347 461275 31362 461290
rect 31535 461286 31547 461290
rect 31532 461275 31547 461286
rect 30773 461245 30793 461275
rect 31347 461245 31547 461275
rect 30773 461230 30788 461245
rect 31347 461230 31362 461245
rect 31532 461234 31547 461245
rect 31535 461230 31547 461234
rect 31607 461275 31622 461290
rect 31795 461286 31807 461290
rect 31792 461275 31807 461286
rect 31607 461245 31807 461275
rect 31607 461230 31622 461245
rect 31792 461234 31807 461245
rect 31795 461230 31807 461234
rect 31867 461275 31882 461290
rect 31867 461245 31921 461275
rect 32596 461265 33596 461315
rect 31867 461230 31882 461245
rect 34110 461231 34710 461287
rect 22906 461055 23212 461225
rect 23406 461055 23712 461225
rect 24573 461158 25173 461208
rect 24573 461002 25173 461130
rect 26490 461107 26690 461160
rect 27691 461090 28291 461218
rect 31823 461084 32061 461118
rect 31481 461080 32061 461084
rect 31481 461068 31797 461080
rect 32596 461063 33596 461113
rect 34110 461075 34710 461203
rect 37998 461133 38148 461145
rect 38317 461133 38467 461145
rect 24573 460846 25173 460974
rect 27691 460934 28291 460990
rect 32596 460907 33596 461035
rect 34110 460919 34710 461047
rect 37998 461020 38598 461070
rect 27691 460778 28291 460906
rect 25286 460758 25310 460762
rect 32596 460751 33596 460879
rect 34110 460763 34710 460891
rect 37998 460844 38598 460900
rect 24573 460690 25173 460746
rect 25286 460687 25310 460721
rect 24573 460534 25173 460662
rect 25286 460615 25310 460649
rect 27691 460622 28291 460750
rect 32596 460595 33596 460723
rect 35287 460695 35487 460707
rect 37998 460674 38598 460724
rect 34110 460607 34710 460663
rect 36785 460650 36797 460654
rect 36785 460639 36800 460650
rect 36970 460639 36985 460654
rect 35134 460582 35734 460632
rect 25286 460543 25310 460577
rect 22906 460255 23212 460425
rect 23406 460255 23712 460425
rect 24573 460378 25173 460506
rect 25286 460471 25310 460505
rect 27691 460472 28291 460522
rect 32596 460439 33596 460567
rect 34110 460451 34710 460507
rect 35134 460432 35734 460482
rect 36785 460459 36985 460639
rect 36785 460448 36800 460459
rect 36785 460444 36797 460448
rect 36970 460444 36985 460459
rect 37083 460639 37098 460654
rect 37083 460459 37120 460639
rect 37083 460444 37098 460459
rect 36785 460414 36797 460418
rect 32596 460283 33596 460411
rect 36785 460403 36800 460414
rect 36970 460403 36985 460418
rect 34110 460295 34710 460351
rect 35134 460316 35734 460366
rect 24573 460228 25173 460278
rect 32596 460127 33596 460255
rect 34110 460145 34710 460195
rect 35134 460160 35734 460288
rect 32596 459971 33596 460099
rect 34110 460029 34710 460079
rect 35134 460004 35734 460132
rect 31481 459862 31797 459880
rect 34110 459873 34710 460001
rect 31823 459828 32061 459860
rect 32596 459821 33596 459871
rect 35134 459848 35734 459976
rect 36071 459805 36098 460295
rect 36785 460223 36985 460403
rect 37993 460248 38593 460298
rect 36785 460212 36800 460223
rect 36785 460208 36797 460212
rect 36970 460208 36985 460223
rect 696597 460200 696600 460320
rect 37993 460078 38593 460128
rect 692376 459983 692396 460017
rect 692463 459993 692532 460017
rect 696191 459993 696239 460017
rect 692487 459983 692532 459993
rect 696204 459983 696239 459993
rect 696340 459983 696360 460017
rect 36785 459902 37385 459952
rect 692487 459915 692502 459939
rect 696200 459915 696215 459939
rect 692454 459891 692478 459915
rect 696224 459891 696248 459915
rect 686755 459800 687355 459850
rect 34110 459717 34710 459773
rect 30253 459701 30268 459716
rect 30441 459712 30453 459716
rect 30438 459701 30453 459712
rect 30253 459671 30453 459701
rect 30253 459656 30268 459671
rect 30438 459660 30453 459671
rect 30441 459656 30453 459660
rect 30513 459701 30528 459716
rect 30701 459712 30713 459716
rect 30698 459701 30713 459712
rect 30513 459671 30713 459701
rect 30513 459656 30528 459671
rect 30698 459660 30713 459671
rect 30701 459656 30713 459660
rect 30773 459701 30788 459716
rect 31347 459701 31362 459716
rect 31535 459712 31547 459716
rect 31532 459701 31547 459712
rect 30773 459671 30793 459701
rect 31347 459671 31547 459701
rect 30773 459656 30788 459671
rect 31347 459656 31362 459671
rect 31532 459660 31547 459671
rect 31535 459656 31547 459660
rect 31607 459701 31622 459716
rect 31795 459712 31807 459716
rect 31792 459701 31807 459712
rect 31607 459671 31807 459701
rect 31607 459656 31622 459671
rect 31792 459660 31807 459671
rect 31795 459656 31807 459660
rect 31867 459701 31882 459716
rect 31867 459671 31921 459701
rect 35134 459698 35734 459770
rect 36785 459726 37385 459782
rect 692487 459748 692505 459752
rect 692479 459718 692505 459748
rect 692487 459698 692505 459718
rect 31867 459656 31882 459671
rect 30253 459615 30268 459630
rect 30441 459626 30453 459630
rect 30438 459615 30453 459626
rect 30253 459585 30453 459615
rect 30253 459570 30268 459585
rect 30438 459574 30453 459585
rect 30441 459570 30453 459574
rect 30513 459615 30528 459630
rect 30701 459626 30713 459630
rect 30698 459615 30713 459626
rect 30513 459585 30713 459615
rect 30513 459570 30528 459585
rect 30698 459574 30713 459585
rect 30701 459570 30713 459574
rect 30773 459615 30788 459630
rect 31347 459615 31362 459630
rect 31535 459626 31547 459630
rect 31532 459615 31547 459626
rect 30773 459585 30793 459615
rect 31347 459585 31547 459615
rect 30773 459570 30788 459585
rect 31347 459570 31362 459585
rect 31532 459574 31547 459585
rect 31535 459570 31547 459574
rect 31607 459615 31622 459630
rect 31795 459626 31807 459630
rect 31792 459615 31807 459626
rect 31607 459585 31807 459615
rect 31607 459570 31622 459585
rect 31792 459574 31807 459585
rect 31795 459570 31807 459574
rect 31867 459615 31882 459630
rect 32546 459619 33546 459669
rect 31867 459585 31921 459615
rect 31867 459570 31882 459585
rect 20809 459471 20833 459505
rect 32546 459463 33546 459591
rect 34110 459561 34710 459689
rect 35134 459645 36134 459695
rect 686755 459624 687355 459680
rect 692485 459674 692505 459698
rect 692509 459674 692517 459718
rect 696215 459698 696223 459748
rect 696203 459674 696223 459698
rect 696227 459674 696245 459752
rect 692485 459640 692521 459674
rect 696203 459640 696249 459674
rect 35134 459489 36134 459617
rect 36785 459550 37385 459606
rect 20809 459403 20833 459437
rect 30253 459405 30268 459420
rect 30441 459416 30453 459420
rect 30438 459405 30453 459416
rect 20809 459335 20833 459369
rect 20809 459267 20833 459301
rect 20809 459199 20833 459233
rect 30253 459225 30453 459405
rect 30253 459210 30268 459225
rect 30438 459214 30453 459225
rect 30441 459210 30453 459214
rect 30513 459405 30528 459420
rect 30701 459416 30713 459420
rect 30698 459405 30713 459416
rect 30513 459225 30713 459405
rect 30513 459210 30528 459225
rect 30698 459214 30713 459225
rect 30701 459210 30713 459214
rect 30773 459405 30788 459420
rect 30961 459416 30973 459420
rect 30958 459405 30973 459416
rect 30773 459225 30973 459405
rect 30773 459210 30788 459225
rect 30958 459214 30973 459225
rect 30961 459210 30973 459214
rect 31087 459405 31102 459420
rect 31275 459416 31287 459420
rect 31272 459405 31287 459416
rect 31087 459225 31287 459405
rect 31087 459210 31102 459225
rect 31272 459214 31287 459225
rect 31275 459210 31287 459214
rect 31347 459405 31362 459420
rect 31535 459416 31547 459420
rect 31532 459405 31547 459416
rect 31347 459225 31547 459405
rect 31347 459210 31362 459225
rect 31532 459214 31547 459225
rect 31535 459210 31547 459214
rect 31607 459405 31622 459420
rect 31795 459416 31807 459420
rect 31792 459405 31807 459416
rect 31607 459225 31807 459405
rect 31607 459210 31622 459225
rect 31792 459214 31807 459225
rect 31795 459210 31807 459214
rect 31867 459405 31882 459420
rect 32055 459416 32067 459420
rect 32052 459405 32067 459416
rect 31867 459225 32067 459405
rect 32546 459307 33546 459435
rect 34110 459411 34710 459461
rect 686755 459448 687355 459504
rect 35134 459339 36134 459389
rect 36785 459380 37385 459430
rect 31867 459210 31882 459225
rect 32052 459214 32067 459225
rect 32055 459210 32067 459214
rect 20809 459131 20833 459165
rect 32546 459151 33546 459279
rect 36785 459248 37385 459298
rect 686755 459278 687355 459328
rect 35285 459162 35319 459172
rect 35353 459162 35387 459172
rect 35421 459162 35455 459172
rect 35489 459162 35523 459172
rect 35564 459162 35598 459172
rect 35632 459162 35666 459172
rect 35700 459162 35734 459172
rect 35768 459162 35802 459172
rect 35836 459162 35870 459172
rect 35904 459162 35938 459172
rect 35972 459162 36006 459172
rect 36040 459162 36074 459172
rect 36108 459162 36142 459172
rect 36176 459162 36210 459172
rect 35255 459126 36255 459138
rect 20809 459063 20833 459097
rect 20940 459085 20983 459103
rect 20940 459069 20949 459085
rect 20974 459069 20983 459085
rect 25113 459069 25349 459093
rect 25383 459069 25417 459093
rect 20974 459051 21008 459069
rect 20809 458995 20833 459029
rect 20974 459028 21003 459051
rect 21361 459045 21409 459069
rect 20949 459027 20983 459028
rect 21385 458991 21409 459045
rect 25113 458991 25137 459069
rect 29993 459045 30993 459095
rect 31347 459045 31362 459060
rect 31535 459056 31547 459060
rect 31532 459045 31547 459056
rect 21361 458967 21409 458991
rect 25089 458967 25137 458991
rect 20809 458927 20833 458961
rect 20809 458859 20833 458893
rect 20809 458791 20833 458825
rect 20809 458723 20833 458757
rect 20809 458655 20833 458689
rect 21413 458638 22813 458681
rect 23685 458638 25085 458681
rect 19844 457229 19894 458629
rect 19994 457229 20122 458629
rect 20150 457229 20278 458629
rect 20306 457229 20434 458629
rect 20462 457229 20512 458629
rect 20809 458587 20833 458621
rect 20809 458519 20833 458553
rect 20809 458451 20833 458485
rect 21413 458475 22813 458603
rect 23685 458475 25085 458603
rect 20809 458383 20833 458417
rect 20809 458315 20833 458349
rect 21413 458312 22813 458440
rect 23685 458312 25085 458440
rect 20809 458247 20833 458281
rect 20809 458179 20833 458213
rect 21413 458149 22813 458277
rect 23685 458149 25085 458277
rect 20809 458111 20833 458145
rect 20809 458043 20833 458077
rect 20809 457975 20833 458009
rect 21413 457986 22813 458114
rect 23685 457986 25085 458114
rect 20809 457907 20833 457941
rect 20809 457839 20833 457873
rect 21413 457823 22813 457951
rect 23685 457823 25085 457951
rect 20809 457771 20833 457805
rect 20809 457703 20833 457737
rect 21413 457673 22813 457716
rect 23685 457673 25085 457716
rect 20809 457635 20833 457669
rect 20809 457567 20833 457601
rect 21361 457552 21419 457586
rect 25089 457552 25147 457586
rect 20809 457499 20833 457533
rect 20809 457431 20833 457465
rect 20809 457363 20833 457397
rect 21361 457373 21419 457397
rect 25089 457373 25147 457397
rect 21385 457363 21419 457373
rect 25113 457363 25147 457373
rect 20809 457295 20833 457329
rect 21385 457291 21419 457325
rect 25113 457291 25147 457325
rect 20809 457227 20833 457261
rect 21385 457219 21419 457253
rect 25113 457219 25147 457253
rect 20809 457159 20833 457193
rect 21385 457171 21419 457181
rect 25113 457171 25147 457181
rect 21361 457147 21419 457171
rect 25089 457147 25147 457171
rect 20809 457091 20833 457125
rect 20809 457023 20833 457057
rect 20809 456955 20833 456989
rect 21361 456969 21409 456993
rect 25089 456969 25137 456993
rect 20809 456887 20833 456921
rect 21385 456915 21409 456969
rect 25113 456915 25137 456969
rect 21361 456891 21409 456915
rect 25089 456891 25137 456915
rect 19480 456831 19583 456867
rect 21413 456754 22813 456804
rect 23685 456754 25085 456804
rect 7389 456489 8389 456561
rect 8990 456489 9990 456561
rect 15678 456534 16678 456606
rect 17278 456534 18278 456606
rect 21413 456591 22813 456719
rect 23685 456591 25085 456719
rect 15748 456523 15782 456534
rect 15816 456523 15850 456534
rect 15884 456523 15918 456534
rect 15952 456523 15986 456534
rect 16020 456523 16054 456534
rect 16088 456523 16122 456534
rect 16156 456523 16190 456534
rect 16224 456523 16258 456534
rect 16292 456523 16326 456534
rect 16360 456523 16394 456534
rect 16428 456523 16462 456534
rect 16496 456523 16530 456534
rect 16564 456523 16598 456534
rect 16632 456523 16666 456534
rect 17290 456523 17324 456534
rect 17358 456523 17392 456534
rect 17426 456523 17460 456534
rect 17494 456523 17528 456534
rect 17562 456523 17596 456534
rect 17630 456523 17664 456534
rect 17698 456523 17732 456534
rect 17766 456523 17800 456534
rect 17834 456523 17868 456534
rect 17902 456523 17936 456534
rect 17970 456523 18004 456534
rect 18038 456523 18072 456534
rect 18106 456523 18140 456534
rect 18174 456523 18208 456534
rect 15748 456513 15806 456523
rect 15816 456513 15874 456523
rect 15884 456513 15942 456523
rect 15952 456513 16010 456523
rect 16020 456513 16078 456523
rect 16088 456513 16146 456523
rect 16156 456513 16214 456523
rect 16224 456513 16282 456523
rect 16292 456513 16350 456523
rect 16360 456513 16418 456523
rect 16428 456513 16486 456523
rect 16496 456513 16554 456523
rect 16564 456513 16622 456523
rect 16632 456513 16690 456523
rect 17290 456513 17348 456523
rect 17358 456513 17416 456523
rect 17426 456513 17484 456523
rect 17494 456513 17552 456523
rect 17562 456513 17620 456523
rect 17630 456513 17688 456523
rect 17698 456513 17756 456523
rect 17766 456513 17824 456523
rect 17834 456513 17892 456523
rect 17902 456513 17960 456523
rect 17970 456513 18028 456523
rect 18038 456513 18096 456523
rect 18106 456513 18164 456523
rect 18174 456513 18232 456523
rect 15724 456489 16690 456513
rect 17266 456489 18232 456513
rect 15748 456474 15772 456489
rect 15816 456474 15840 456489
rect 15884 456474 15908 456489
rect 15952 456474 15976 456489
rect 16020 456474 16044 456489
rect 16088 456474 16112 456489
rect 16156 456474 16180 456489
rect 16224 456474 16248 456489
rect 16292 456474 16316 456489
rect 16360 456474 16384 456489
rect 16428 456474 16452 456489
rect 16496 456474 16520 456489
rect 16564 456474 16588 456489
rect 16632 456474 16656 456489
rect 17290 456474 17314 456489
rect 17358 456474 17382 456489
rect 17426 456474 17450 456489
rect 17494 456474 17518 456489
rect 17562 456474 17586 456489
rect 17630 456474 17654 456489
rect 17698 456474 17722 456489
rect 17766 456474 17790 456489
rect 17834 456474 17858 456489
rect 17902 456474 17926 456489
rect 17970 456474 17994 456489
rect 18038 456474 18062 456489
rect 18106 456474 18130 456489
rect 18174 456474 18198 456489
rect 15678 456319 16678 456474
rect 7389 456229 8389 456289
rect 8990 456229 9990 456289
rect 15678 456285 16690 456319
rect 17278 456309 18278 456474
rect 21413 456428 22813 456556
rect 23685 456428 25085 456556
rect 17266 456285 18278 456309
rect 15678 456274 16678 456285
rect 17278 456274 18278 456285
rect 15748 456261 15772 456274
rect 15816 456261 15840 456274
rect 15884 456261 15908 456274
rect 15952 456261 15976 456274
rect 16020 456261 16044 456274
rect 16088 456261 16112 456274
rect 16156 456261 16180 456274
rect 16224 456261 16248 456274
rect 16292 456261 16316 456274
rect 16360 456261 16384 456274
rect 16428 456261 16452 456274
rect 16496 456261 16520 456274
rect 16564 456261 16588 456274
rect 16632 456261 16656 456274
rect 17290 456261 17314 456274
rect 17358 456261 17382 456274
rect 17426 456261 17450 456274
rect 17494 456261 17518 456274
rect 17562 456261 17586 456274
rect 17630 456261 17654 456274
rect 17698 456261 17722 456274
rect 17766 456261 17790 456274
rect 17834 456261 17858 456274
rect 17902 456261 17926 456274
rect 17970 456261 17994 456274
rect 18038 456261 18062 456274
rect 18106 456261 18130 456274
rect 18174 456261 18198 456274
rect 21413 456265 22813 456393
rect 23685 456265 25085 456393
rect 21413 456102 22813 456230
rect 23685 456102 25085 456230
rect 7389 455871 8389 455927
rect 8990 455871 9990 455927
rect 15678 455916 16678 455972
rect 17278 455916 18278 455972
rect 21413 455952 22813 455995
rect 23685 455952 25085 455995
rect 7389 455799 8389 455855
rect 8990 455799 9990 455855
rect 15678 455844 16678 455900
rect 17278 455844 18278 455900
rect 21406 455865 21430 455889
rect 25068 455865 25092 455889
rect 21382 455841 21385 455865
rect 25113 455841 25116 455865
rect 21382 455763 21396 455787
rect 25102 455763 25116 455787
rect 21348 455739 21372 455763
rect 21406 455739 21430 455763
rect 25068 455739 25092 455763
rect 25126 455739 25150 455763
rect 25524 455703 25548 459001
rect 29993 458895 30993 458945
rect 31347 458865 31547 459045
rect 31347 458850 31362 458865
rect 31532 458854 31547 458865
rect 31535 458850 31547 458854
rect 31607 459045 31622 459060
rect 31795 459056 31807 459060
rect 31792 459045 31807 459056
rect 31607 458865 31807 459045
rect 32546 458995 33546 459123
rect 36785 459072 37385 459128
rect 685547 459102 686147 459152
rect 35255 459019 36255 459069
rect 687155 459007 687170 459022
rect 687343 459018 687355 459022
rect 687340 459007 687355 459018
rect 31607 458850 31622 458865
rect 31792 458854 31807 458865
rect 31795 458850 31807 458854
rect 32546 458839 33546 458967
rect 35255 458843 36255 458971
rect 36785 458896 37385 458952
rect 685547 458932 686147 458982
rect 687155 458827 687355 459007
rect 31347 458809 31362 458824
rect 31535 458820 31547 458824
rect 31532 458809 31547 458820
rect 29993 458736 30993 458786
rect 29993 458586 30993 458636
rect 31347 458629 31547 458809
rect 31347 458614 31362 458629
rect 31532 458618 31547 458629
rect 31535 458614 31547 458618
rect 31607 458809 31622 458824
rect 31795 458820 31807 458824
rect 31792 458809 31807 458820
rect 687155 458812 687170 458827
rect 687340 458816 687355 458827
rect 687343 458812 687355 458816
rect 31607 458629 31807 458809
rect 32546 458683 33546 458811
rect 35255 458667 36255 458795
rect 36785 458726 37385 458776
rect 687042 458771 687057 458786
rect 31607 458614 31622 458629
rect 31792 458618 31807 458629
rect 31795 458614 31807 458618
rect 32546 458527 33546 458655
rect 37993 458550 38593 458600
rect 687020 458591 687057 458771
rect 687042 458576 687057 458591
rect 687155 458771 687170 458786
rect 687343 458782 687355 458786
rect 687340 458771 687355 458782
rect 687155 458591 687355 458771
rect 688210 458630 688260 459630
rect 688360 458630 688488 459630
rect 688516 458630 688644 459630
rect 688672 458630 688800 459630
rect 688828 458630 688956 459630
rect 688984 458630 689112 459630
rect 689140 458630 689268 459630
rect 689296 458630 689424 459630
rect 689452 458630 689580 459630
rect 689608 458630 689736 459630
rect 689764 458630 689892 459630
rect 689920 458630 690048 459630
rect 690076 458630 690204 459630
rect 690232 458630 690360 459630
rect 690388 458630 690438 459630
rect 692485 459606 692505 459640
rect 692509 459606 692517 459640
rect 696203 459606 696223 459640
rect 696227 459606 696245 459640
rect 691275 459523 691875 459573
rect 692485 459572 692521 459606
rect 696203 459572 696249 459606
rect 692485 459538 692505 459572
rect 692509 459538 692517 459572
rect 692485 459504 692521 459538
rect 692583 459528 693983 459571
rect 694719 459528 696119 459571
rect 696203 459538 696223 459572
rect 696227 459538 696245 459572
rect 696203 459504 696249 459538
rect 692485 459470 692505 459504
rect 692509 459470 692517 459504
rect 692485 459436 692521 459470
rect 691275 459373 691875 459423
rect 692485 459402 692505 459436
rect 692509 459402 692517 459436
rect 692485 459368 692521 459402
rect 692485 459334 692505 459368
rect 692509 459334 692517 459368
rect 692583 459365 693983 459493
rect 694719 459365 696119 459493
rect 696203 459470 696223 459504
rect 696227 459470 696245 459504
rect 696203 459436 696249 459470
rect 707624 459441 707658 459475
rect 707695 459441 707729 459475
rect 707769 459441 707803 459475
rect 707840 459441 707874 459475
rect 707914 459441 707948 459475
rect 707985 459441 708019 459475
rect 708059 459441 708093 459475
rect 708130 459441 708164 459475
rect 708204 459441 708238 459475
rect 708275 459441 708309 459475
rect 708369 459441 708403 459475
rect 708446 459441 708480 459475
rect 708520 459441 708554 459465
rect 708588 459441 708610 459465
rect 709211 459441 709234 459465
rect 709270 459441 709304 459475
rect 709364 459441 709398 459475
rect 709435 459441 709469 459475
rect 709509 459441 709543 459475
rect 709580 459441 709614 459475
rect 709654 459441 709688 459475
rect 709725 459441 709759 459475
rect 709799 459441 709833 459475
rect 709870 459441 709904 459475
rect 709944 459441 709978 459475
rect 710015 459441 710049 459475
rect 710089 459441 710123 459475
rect 710160 459441 710194 459475
rect 696203 459402 696223 459436
rect 696227 459402 696245 459436
rect 707610 459431 707624 459441
rect 707658 459431 707695 459441
rect 707729 459431 707769 459441
rect 707803 459431 707840 459441
rect 707874 459431 707914 459441
rect 707948 459431 707985 459441
rect 708019 459431 708059 459441
rect 708093 459431 708130 459441
rect 708164 459431 708204 459441
rect 708238 459431 708275 459441
rect 708309 459431 708369 459441
rect 708403 459431 708446 459441
rect 708480 459431 708520 459441
rect 708554 459431 708588 459441
rect 708610 459431 708634 459441
rect 709211 459431 709270 459441
rect 709304 459431 709364 459441
rect 709398 459431 709435 459441
rect 709469 459431 709509 459441
rect 709543 459431 709580 459441
rect 709614 459431 709654 459441
rect 709688 459431 709725 459441
rect 709759 459431 709799 459441
rect 709833 459431 709870 459441
rect 709904 459431 709944 459441
rect 709978 459431 710015 459441
rect 710049 459431 710089 459441
rect 710123 459431 710160 459441
rect 710194 459431 710211 459441
rect 696203 459368 696249 459402
rect 696203 459334 696223 459368
rect 696227 459334 696245 459368
rect 707610 459337 708610 459431
rect 709211 459337 710211 459431
rect 691275 459251 691875 459301
rect 692485 459300 692521 459334
rect 692485 459266 692505 459300
rect 692509 459266 692517 459300
rect 692485 459232 692521 459266
rect 692485 459198 692505 459232
rect 692509 459198 692517 459232
rect 692583 459202 693983 459330
rect 694719 459202 696119 459330
rect 696203 459300 696249 459334
rect 711579 459317 712463 459331
rect 711579 459307 711619 459317
rect 696203 459266 696223 459300
rect 696227 459266 696245 459300
rect 701730 459290 701747 459292
rect 696203 459232 696249 459266
rect 696203 459198 696223 459232
rect 696227 459198 696245 459232
rect 701692 459220 701722 459254
rect 701730 459220 701760 459290
rect 707610 459241 708610 459301
rect 709211 459241 710211 459301
rect 692485 459164 692521 459198
rect 691275 459101 691875 459151
rect 692485 459130 692505 459164
rect 692509 459130 692517 459164
rect 692485 459096 692521 459130
rect 692485 459062 692505 459096
rect 692509 459062 692517 459096
rect 692485 459028 692521 459062
rect 692583 459039 693983 459167
rect 694719 459039 696119 459167
rect 696203 459164 696249 459198
rect 696203 459130 696223 459164
rect 696227 459130 696245 459164
rect 696203 459096 696249 459130
rect 696203 459062 696223 459096
rect 696227 459062 696245 459096
rect 699322 459064 700322 459097
rect 700922 459064 701922 459097
rect 696203 459028 696249 459062
rect 707610 459044 708610 459048
rect 709211 459044 710211 459048
rect 691275 458975 691875 459025
rect 692485 458994 692505 459028
rect 692509 458994 692517 459028
rect 692485 458960 692521 458994
rect 692485 458926 692505 458960
rect 692509 458926 692517 458960
rect 692485 458892 692521 458926
rect 691275 458825 691875 458875
rect 692485 458858 692505 458892
rect 692509 458858 692517 458892
rect 692583 458876 693983 459004
rect 694719 458876 696119 459004
rect 696203 458994 696223 459028
rect 696227 458994 696245 459028
rect 707574 458994 708646 459030
rect 696203 458960 696249 458994
rect 696203 458926 696223 458960
rect 696227 458926 696245 458960
rect 707574 458953 707610 458994
rect 708610 458953 708646 458994
rect 696203 458892 696249 458926
rect 697284 458894 697350 458910
rect 707574 458897 708646 458953
rect 696203 458858 696223 458892
rect 696227 458858 696245 458892
rect 699322 458877 700322 458894
rect 700922 458877 701922 458894
rect 707574 458881 707610 458897
rect 708610 458881 708646 458897
rect 692485 458824 692521 458858
rect 692485 458790 692505 458824
rect 692509 458790 692517 458824
rect 692485 458756 692521 458790
rect 691275 458703 691875 458753
rect 692485 458722 692505 458756
rect 692509 458722 692517 458756
rect 692485 458688 692521 458722
rect 692583 458713 693983 458841
rect 694719 458713 696119 458841
rect 696203 458824 696249 458858
rect 707574 458825 708646 458881
rect 696203 458790 696223 458824
rect 696227 458790 696245 458824
rect 696203 458756 696249 458790
rect 696203 458722 696223 458756
rect 696227 458722 696245 458756
rect 699322 458739 700322 458811
rect 700922 458739 701922 458811
rect 707574 458788 707610 458825
rect 708610 458788 708646 458825
rect 707574 458748 708646 458788
rect 709175 458994 710247 459030
rect 709175 458953 709211 458994
rect 710211 458953 710247 458994
rect 709175 458897 710247 458953
rect 709175 458881 709211 458897
rect 710211 458881 710247 458897
rect 709175 458825 710247 458881
rect 709175 458788 709211 458825
rect 710211 458788 710247 458825
rect 709175 458748 710247 458788
rect 696203 458688 696249 458722
rect 692485 458654 692505 458688
rect 692509 458654 692517 458688
rect 692485 458620 692521 458654
rect 687155 458576 687170 458591
rect 687340 458580 687355 458591
rect 687343 458576 687355 458580
rect 28647 458450 28671 458477
rect 30171 458447 30771 458497
rect 35255 458491 36255 458547
rect 685542 458506 686142 458556
rect 691275 458553 691875 458603
rect 692485 458586 692505 458620
rect 692509 458586 692517 458620
rect 692485 458552 692521 458586
rect 692485 458518 692505 458552
rect 692509 458518 692517 458552
rect 692583 458550 693983 458678
rect 694719 458550 696119 458678
rect 696203 458654 696223 458688
rect 696227 458654 696245 458688
rect 696203 458620 696249 458654
rect 696203 458586 696223 458620
rect 696227 458586 696245 458620
rect 696203 458552 696249 458586
rect 696203 458518 696223 458552
rect 696227 458518 696245 458552
rect 692485 458484 692521 458518
rect 36785 458466 36797 458470
rect 36785 458455 36800 458466
rect 36970 458455 36985 458470
rect 28683 458397 28717 458431
rect 32546 458377 33546 458427
rect 28683 458328 28717 458362
rect 28683 458259 28717 458293
rect 30171 458271 30771 458327
rect 35255 458321 36255 458371
rect 36785 458275 36985 458455
rect 692485 458450 692505 458484
rect 692509 458450 692517 458484
rect 37993 458380 38593 458430
rect 692485 458416 692521 458450
rect 679817 458330 679841 458354
rect 685542 458330 686142 458386
rect 692485 458382 692505 458416
rect 692509 458382 692517 458416
rect 692583 458387 693983 458515
rect 694719 458387 696119 458515
rect 696203 458484 696249 458518
rect 696203 458450 696223 458484
rect 696227 458450 696245 458484
rect 699322 458478 700322 458550
rect 700922 458478 701922 458550
rect 707610 458523 708610 458595
rect 709211 458523 710211 458595
rect 699392 458467 699426 458478
rect 699460 458467 699494 458478
rect 699528 458467 699562 458478
rect 699596 458467 699630 458478
rect 699664 458467 699698 458478
rect 699732 458467 699766 458478
rect 699800 458467 699834 458478
rect 699868 458467 699902 458478
rect 699936 458467 699970 458478
rect 700004 458467 700038 458478
rect 700072 458467 700106 458478
rect 700140 458467 700174 458478
rect 700208 458467 700242 458478
rect 700276 458467 700310 458478
rect 700934 458467 700968 458478
rect 701002 458467 701036 458478
rect 701070 458467 701104 458478
rect 701138 458467 701172 458478
rect 701206 458467 701240 458478
rect 701274 458467 701308 458478
rect 701342 458467 701376 458478
rect 701410 458467 701444 458478
rect 701478 458467 701512 458478
rect 701546 458467 701580 458478
rect 701614 458467 701648 458478
rect 701682 458467 701716 458478
rect 701750 458467 701784 458478
rect 701818 458467 701852 458478
rect 699392 458457 699450 458467
rect 699460 458457 699518 458467
rect 699528 458457 699586 458467
rect 699596 458457 699654 458467
rect 699664 458457 699722 458467
rect 699732 458457 699790 458467
rect 699800 458457 699858 458467
rect 699868 458457 699926 458467
rect 699936 458457 699994 458467
rect 700004 458457 700062 458467
rect 700072 458457 700130 458467
rect 700140 458457 700198 458467
rect 700208 458457 700266 458467
rect 700276 458457 700334 458467
rect 700934 458457 700992 458467
rect 701002 458457 701060 458467
rect 701070 458457 701128 458467
rect 701138 458457 701196 458467
rect 701206 458457 701264 458467
rect 701274 458457 701332 458467
rect 701342 458457 701400 458467
rect 701410 458457 701468 458467
rect 701478 458457 701536 458467
rect 701546 458457 701604 458467
rect 701614 458457 701672 458467
rect 701682 458457 701740 458467
rect 701750 458457 701808 458467
rect 701818 458457 701876 458467
rect 696203 458416 696249 458450
rect 699368 458433 700334 458457
rect 700910 458433 701876 458457
rect 699392 458418 699416 458433
rect 699460 458418 699484 458433
rect 699528 458418 699552 458433
rect 699596 458418 699620 458433
rect 699664 458418 699688 458433
rect 699732 458418 699756 458433
rect 699800 458418 699824 458433
rect 699868 458418 699892 458433
rect 699936 458418 699960 458433
rect 700004 458418 700028 458433
rect 700072 458418 700096 458433
rect 700140 458418 700164 458433
rect 700208 458418 700232 458433
rect 700276 458418 700300 458433
rect 700934 458418 700958 458433
rect 701002 458418 701026 458433
rect 701070 458418 701094 458433
rect 701138 458418 701162 458433
rect 701206 458418 701230 458433
rect 701274 458418 701298 458433
rect 701342 458418 701366 458433
rect 701410 458418 701434 458433
rect 701478 458418 701502 458433
rect 701546 458418 701570 458433
rect 701614 458418 701638 458433
rect 701682 458418 701706 458433
rect 701750 458418 701774 458433
rect 701818 458418 701842 458433
rect 696203 458382 696223 458416
rect 696227 458382 696245 458416
rect 692485 458348 692521 458382
rect 696203 458348 696249 458382
rect 679549 458307 679573 458330
rect 679793 458306 679808 458330
rect 692485 458314 692505 458348
rect 692509 458314 692517 458348
rect 696203 458314 696223 458348
rect 696227 458314 696245 458348
rect 36785 458264 36800 458275
rect 36785 458260 36797 458264
rect 36970 458260 36985 458275
rect 692485 458280 692521 458314
rect 696203 458280 696249 458314
rect 679549 458237 679573 458271
rect 692485 458246 692505 458280
rect 692509 458246 692517 458280
rect 36785 458230 36797 458234
rect 28683 458190 28717 458224
rect 32596 458175 33596 458225
rect 35359 458156 35375 458222
rect 36143 458156 36159 458222
rect 36785 458219 36800 458230
rect 36970 458219 36985 458234
rect 28683 458121 28717 458155
rect 30171 458101 30771 458151
rect 28683 458052 28717 458086
rect 32596 458019 33596 458147
rect 28683 457983 28717 458017
rect 33959 457994 33975 458060
rect 36143 457994 36159 458060
rect 36785 458039 36985 458219
rect 36785 458028 36800 458039
rect 36785 458024 36797 458028
rect 36970 458024 36985 458039
rect 37083 458219 37098 458234
rect 37083 458039 37120 458219
rect 692485 458212 692521 458246
rect 692583 458237 693983 458280
rect 694719 458237 696119 458280
rect 696203 458246 696223 458280
rect 696227 458246 696245 458280
rect 699322 458263 700322 458418
rect 696203 458212 696249 458246
rect 699322 458229 700334 458263
rect 700922 458253 701922 458418
rect 700910 458229 701922 458253
rect 699322 458218 700322 458229
rect 700922 458218 701922 458229
rect 707574 458263 708646 458299
rect 707574 458226 707610 458263
rect 708610 458226 708646 458263
rect 679549 458167 679573 458201
rect 685542 458160 686142 458210
rect 685601 458157 685895 458160
rect 685920 458157 686142 458160
rect 692485 458178 692505 458212
rect 692509 458178 692517 458212
rect 696203 458178 696223 458212
rect 696227 458178 696245 458212
rect 699392 458205 699416 458218
rect 699460 458205 699484 458218
rect 699528 458205 699552 458218
rect 699596 458205 699620 458218
rect 699664 458205 699688 458218
rect 699732 458205 699756 458218
rect 699800 458205 699824 458218
rect 699868 458205 699892 458218
rect 699936 458205 699960 458218
rect 700004 458205 700028 458218
rect 700072 458205 700096 458218
rect 700140 458205 700164 458218
rect 700208 458205 700232 458218
rect 700276 458205 700300 458218
rect 700934 458205 700958 458218
rect 701002 458205 701026 458218
rect 701070 458205 701094 458218
rect 701138 458205 701162 458218
rect 701206 458205 701230 458218
rect 701274 458205 701298 458218
rect 701342 458205 701366 458218
rect 701410 458205 701434 458218
rect 701478 458205 701502 458218
rect 701546 458205 701570 458218
rect 701614 458205 701638 458218
rect 701682 458205 701706 458218
rect 701750 458205 701774 458218
rect 701818 458205 701842 458218
rect 707574 458186 708646 458226
rect 709175 458263 710247 458299
rect 709175 458226 709211 458263
rect 710211 458226 710247 458263
rect 709175 458186 710247 458226
rect 692485 458144 692521 458178
rect 696203 458144 696249 458178
rect 679549 458097 679573 458131
rect 692485 458110 692505 458144
rect 692509 458110 692517 458144
rect 692485 458076 692521 458110
rect 692583 458101 693983 458144
rect 694719 458101 696119 458144
rect 696203 458110 696223 458144
rect 696227 458110 696245 458144
rect 696203 458076 696249 458110
rect 37083 458024 37098 458039
rect 679549 458027 679573 458061
rect 692485 458042 692505 458076
rect 692509 458042 692517 458076
rect 692485 458008 692521 458042
rect 28683 457914 28717 457948
rect 31463 457895 32063 457945
rect 28683 457845 28717 457879
rect 32596 457863 33596 457991
rect 37998 457954 38598 458004
rect 679549 457957 679573 457991
rect 692485 457974 692505 458008
rect 692509 457974 692517 458008
rect 679793 457933 679808 457957
rect 692485 457940 692521 457974
rect 679817 457909 679841 457933
rect 692485 457906 692505 457940
rect 692509 457906 692517 457940
rect 692583 457938 693983 458066
rect 694719 457938 696119 458066
rect 696203 458042 696223 458076
rect 696227 458042 696245 458076
rect 696203 458008 696249 458042
rect 696203 457974 696223 458008
rect 696227 457974 696245 458008
rect 696203 457940 696249 457974
rect 696203 457906 696223 457940
rect 696227 457906 696245 457940
rect 28683 457776 28717 457810
rect 28683 457707 28717 457741
rect 31463 457739 32063 457795
rect 32596 457707 33596 457835
rect 33959 457832 33975 457898
rect 36143 457832 36159 457898
rect 687685 457838 687709 457862
rect 37998 457778 38598 457834
rect 687661 457814 687675 457838
rect 687669 457797 687675 457814
rect 679515 457762 679539 457785
rect 679613 457762 679637 457785
rect 679491 457737 679515 457761
rect 679637 457737 679661 457761
rect 28683 457638 28717 457672
rect 28683 457569 28717 457603
rect 31463 457589 32063 457639
rect 32596 457551 33596 457679
rect 35359 457670 35375 457736
rect 36143 457670 36159 457736
rect 680215 457678 680815 457728
rect 37998 457608 38598 457658
rect 37998 457605 38220 457608
rect 38245 457605 38539 457608
rect 28683 457500 28717 457534
rect 28683 457431 28717 457465
rect 28683 457362 28717 457396
rect 32596 457395 33596 457523
rect 35255 457521 36255 457571
rect 680215 457502 680815 457558
rect 685551 457516 686551 457566
rect 28683 457293 28717 457327
rect 28683 457224 28717 457258
rect 30015 457256 30718 457272
rect 30015 457246 30721 457256
rect 28683 457155 28717 457189
rect 28683 457086 28717 457120
rect 28683 457017 28717 457051
rect 28683 456948 28717 456982
rect 28683 456879 28717 456913
rect 28683 456810 28717 456844
rect 28683 456741 28717 456775
rect 28683 456672 28717 456706
rect 28683 456603 28717 456637
rect 28683 456534 28717 456568
rect 28683 456465 28717 456499
rect 28683 456396 28717 456430
rect 28682 456361 28683 456366
rect 28682 456332 28717 456361
rect 28647 456303 28671 456332
rect 28647 456234 28671 456268
rect 28647 456165 28671 456199
rect 28647 456096 28671 456130
rect 28647 456027 28671 456061
rect 28647 455958 28671 455992
rect 28647 455889 28671 455923
rect 28647 455820 28671 455854
rect 28647 455751 28671 455785
rect 28647 455682 28671 455716
rect 29778 455695 29802 455719
rect 29802 455671 29826 455683
rect 29880 455681 29914 455715
rect 25524 455635 25548 455669
rect 7389 455497 8389 455569
rect 8990 455497 9990 455569
rect 15678 455542 16678 455614
rect 17278 455542 18278 455614
rect 28647 455613 28671 455647
rect 29778 455635 29802 455659
rect 21361 455586 21409 455610
rect 25089 455586 25137 455610
rect 15748 455531 15782 455542
rect 15816 455531 15850 455542
rect 15884 455531 15918 455542
rect 15952 455531 15986 455542
rect 16020 455531 16054 455542
rect 16088 455531 16122 455542
rect 16156 455531 16190 455542
rect 16224 455531 16258 455542
rect 16292 455531 16326 455542
rect 16360 455531 16394 455542
rect 16428 455531 16462 455542
rect 16496 455531 16530 455542
rect 16564 455531 16598 455542
rect 16632 455531 16666 455542
rect 17290 455531 17324 455542
rect 17358 455531 17392 455542
rect 17426 455531 17460 455542
rect 17494 455531 17528 455542
rect 17562 455531 17596 455542
rect 17630 455531 17664 455542
rect 17698 455531 17732 455542
rect 17766 455531 17800 455542
rect 17834 455531 17868 455542
rect 17902 455531 17936 455542
rect 17970 455531 18004 455542
rect 18038 455531 18072 455542
rect 18106 455531 18140 455542
rect 18174 455531 18208 455542
rect 21385 455532 21409 455586
rect 25113 455532 25137 455586
rect 28647 455544 28671 455578
rect 15748 455521 15806 455531
rect 15816 455521 15874 455531
rect 15884 455521 15942 455531
rect 15952 455521 16010 455531
rect 16020 455521 16078 455531
rect 16088 455521 16146 455531
rect 16156 455521 16214 455531
rect 16224 455521 16282 455531
rect 16292 455521 16350 455531
rect 16360 455521 16418 455531
rect 16428 455521 16486 455531
rect 16496 455521 16554 455531
rect 16564 455521 16622 455531
rect 16632 455521 16690 455531
rect 17290 455521 17348 455531
rect 17358 455521 17416 455531
rect 17426 455521 17484 455531
rect 17494 455521 17552 455531
rect 17562 455521 17620 455531
rect 17630 455521 17688 455531
rect 17698 455521 17756 455531
rect 17766 455521 17824 455531
rect 17834 455521 17892 455531
rect 17902 455521 17960 455531
rect 17970 455521 18028 455531
rect 18038 455521 18096 455531
rect 18106 455521 18164 455531
rect 18174 455521 18232 455531
rect 15724 455497 16690 455521
rect 17266 455497 18232 455521
rect 21361 455508 21409 455532
rect 25089 455508 25137 455532
rect 15748 455482 15772 455497
rect 15816 455482 15840 455497
rect 15884 455482 15908 455497
rect 15952 455482 15976 455497
rect 16020 455482 16044 455497
rect 16088 455482 16112 455497
rect 16156 455482 16180 455497
rect 16224 455482 16248 455497
rect 16292 455482 16316 455497
rect 16360 455482 16384 455497
rect 16428 455482 16452 455497
rect 16496 455482 16520 455497
rect 16564 455482 16588 455497
rect 16632 455482 16656 455497
rect 17290 455482 17314 455497
rect 17358 455482 17382 455497
rect 17426 455482 17450 455497
rect 17494 455482 17518 455497
rect 17562 455482 17586 455497
rect 17630 455482 17654 455497
rect 17698 455482 17722 455497
rect 17766 455482 17790 455497
rect 17834 455482 17858 455497
rect 17902 455482 17926 455497
rect 17970 455482 17994 455497
rect 18038 455482 18062 455497
rect 18106 455482 18130 455497
rect 18174 455482 18198 455497
rect 7389 455237 8389 455297
rect 8990 455237 9990 455297
rect 12559 455273 12865 455375
rect 15678 455327 16678 455482
rect 15678 455293 16690 455327
rect 17278 455317 18278 455482
rect 28647 455475 28671 455509
rect 28647 455406 28671 455440
rect 28647 455337 28671 455371
rect 17266 455293 18278 455317
rect 15678 455282 16678 455293
rect 17278 455282 18278 455293
rect 12543 455257 12881 455273
rect 15748 455269 15772 455282
rect 15816 455269 15840 455282
rect 15884 455269 15908 455282
rect 15952 455269 15976 455282
rect 16020 455269 16044 455282
rect 16088 455269 16112 455282
rect 16156 455269 16180 455282
rect 16224 455269 16248 455282
rect 16292 455269 16316 455282
rect 16360 455269 16384 455282
rect 16428 455269 16452 455282
rect 16496 455269 16520 455282
rect 16564 455269 16588 455282
rect 16632 455269 16656 455282
rect 17290 455269 17314 455282
rect 17358 455269 17382 455282
rect 17426 455269 17450 455282
rect 17494 455269 17518 455282
rect 17562 455269 17586 455282
rect 17630 455269 17654 455282
rect 17698 455269 17722 455282
rect 17766 455269 17790 455282
rect 17834 455269 17858 455282
rect 17902 455269 17926 455282
rect 17970 455269 17994 455282
rect 18038 455269 18062 455282
rect 18106 455269 18130 455282
rect 18174 455269 18198 455282
rect 19980 455048 20286 455218
rect 7389 454879 8389 454935
rect 8990 454879 9990 454935
rect 15678 454924 16678 454980
rect 17278 454924 18278 454980
rect 7389 454807 8389 454863
rect 8990 454807 9990 454863
rect 15678 454852 16678 454908
rect 17278 454852 18278 454908
rect 20945 454796 25553 455332
rect 28647 455268 28671 455302
rect 28647 455199 28671 455233
rect 28647 455154 28671 455164
rect 21413 454706 22813 454796
rect 23685 454706 25085 454796
rect 7389 454505 8389 454577
rect 8990 454505 9990 454577
rect 15678 454550 16678 454622
rect 17278 454550 18278 454622
rect 15748 454539 15782 454550
rect 15816 454539 15850 454550
rect 15884 454539 15918 454550
rect 15952 454539 15986 454550
rect 16020 454539 16054 454550
rect 16088 454539 16122 454550
rect 16156 454539 16190 454550
rect 16224 454539 16258 454550
rect 16292 454539 16326 454550
rect 16360 454539 16394 454550
rect 16428 454539 16462 454550
rect 16496 454539 16530 454550
rect 16564 454539 16598 454550
rect 16632 454539 16666 454550
rect 17290 454539 17324 454550
rect 17358 454539 17392 454550
rect 17426 454539 17460 454550
rect 17494 454539 17528 454550
rect 17562 454539 17596 454550
rect 17630 454539 17664 454550
rect 17698 454539 17732 454550
rect 17766 454539 17800 454550
rect 17834 454539 17868 454550
rect 17902 454539 17936 454550
rect 17970 454539 18004 454550
rect 18038 454539 18072 454550
rect 18106 454539 18140 454550
rect 18174 454539 18208 454550
rect 21413 454543 22813 454671
rect 23685 454543 25085 454671
rect 15748 454529 15806 454539
rect 15816 454529 15874 454539
rect 15884 454529 15942 454539
rect 15952 454529 16010 454539
rect 16020 454529 16078 454539
rect 16088 454529 16146 454539
rect 16156 454529 16214 454539
rect 16224 454529 16282 454539
rect 16292 454529 16350 454539
rect 16360 454529 16418 454539
rect 16428 454529 16486 454539
rect 16496 454529 16554 454539
rect 16564 454529 16622 454539
rect 16632 454529 16690 454539
rect 17290 454529 17348 454539
rect 17358 454529 17416 454539
rect 17426 454529 17484 454539
rect 17494 454529 17552 454539
rect 17562 454529 17620 454539
rect 17630 454529 17688 454539
rect 17698 454529 17756 454539
rect 17766 454529 17824 454539
rect 17834 454529 17892 454539
rect 17902 454529 17960 454539
rect 17970 454529 18028 454539
rect 18038 454529 18096 454539
rect 18106 454529 18164 454539
rect 18174 454529 18232 454539
rect 15724 454505 16690 454529
rect 17266 454505 18232 454529
rect 15748 454490 15772 454505
rect 15816 454490 15840 454505
rect 15884 454490 15908 454505
rect 15952 454490 15976 454505
rect 16020 454490 16044 454505
rect 16088 454490 16112 454505
rect 16156 454490 16180 454505
rect 16224 454490 16248 454505
rect 16292 454490 16316 454505
rect 16360 454490 16384 454505
rect 16428 454490 16452 454505
rect 16496 454490 16520 454505
rect 16564 454490 16588 454505
rect 16632 454490 16656 454505
rect 17290 454490 17314 454505
rect 17358 454490 17382 454505
rect 17426 454490 17450 454505
rect 17494 454490 17518 454505
rect 17562 454490 17586 454505
rect 17630 454490 17654 454505
rect 17698 454490 17722 454505
rect 17766 454490 17790 454505
rect 17834 454490 17858 454505
rect 17902 454490 17926 454505
rect 17970 454490 17994 454505
rect 18038 454490 18062 454505
rect 18106 454490 18130 454505
rect 18174 454490 18198 454505
rect 15678 454335 16678 454490
rect 7389 454245 8389 454305
rect 8990 454245 9990 454305
rect 15678 454301 16690 454335
rect 17278 454325 18278 454490
rect 21413 454380 22813 454508
rect 23685 454380 25085 454508
rect 17266 454301 18278 454325
rect 15678 454290 16678 454301
rect 17278 454290 18278 454301
rect 15748 454277 15772 454290
rect 15816 454277 15840 454290
rect 15884 454277 15908 454290
rect 15952 454277 15976 454290
rect 16020 454277 16044 454290
rect 16088 454277 16112 454290
rect 16156 454277 16180 454290
rect 16224 454277 16248 454290
rect 16292 454277 16316 454290
rect 16360 454277 16384 454290
rect 16428 454277 16452 454290
rect 16496 454277 16520 454290
rect 16564 454277 16588 454290
rect 16632 454277 16656 454290
rect 17290 454277 17314 454290
rect 17358 454277 17382 454290
rect 17426 454277 17450 454290
rect 17494 454277 17518 454290
rect 17562 454277 17586 454290
rect 17630 454277 17654 454290
rect 17698 454277 17722 454290
rect 17766 454277 17790 454290
rect 17834 454277 17858 454290
rect 17902 454277 17926 454290
rect 17970 454277 17994 454290
rect 18038 454277 18062 454290
rect 18106 454277 18130 454290
rect 18174 454277 18198 454290
rect 21413 454217 22813 454345
rect 23685 454217 25085 454345
rect 21413 454054 22813 454182
rect 23685 454054 25085 454182
rect 25936 454132 26936 454182
rect 27274 454033 27358 454036
rect 13899 453998 14059 454002
rect 7389 453887 8389 453943
rect 8990 453887 9990 453943
rect 15678 453932 16678 453988
rect 17278 453932 18278 453988
rect 7389 453815 8389 453871
rect 8990 453815 9990 453871
rect 15678 453860 16678 453916
rect 17278 453860 18278 453916
rect 21413 453891 22813 454019
rect 23685 453891 25085 454019
rect 25936 453976 26936 454032
rect 27158 453983 27358 454033
rect 13899 453852 14059 453856
rect 25936 453820 26936 453876
rect 27158 453807 27358 453935
rect 21413 453741 22813 453784
rect 23685 453741 25085 453784
rect 25936 453664 26936 453720
rect 7389 453513 8389 453585
rect 8990 453513 9990 453585
rect 15678 453558 16678 453630
rect 17278 453558 18278 453630
rect 21413 453605 22813 453648
rect 23685 453605 25085 453648
rect 27158 453631 27358 453687
rect 15748 453547 15782 453558
rect 15816 453547 15850 453558
rect 15884 453547 15918 453558
rect 15952 453547 15986 453558
rect 16020 453547 16054 453558
rect 16088 453547 16122 453558
rect 16156 453547 16190 453558
rect 16224 453547 16258 453558
rect 16292 453547 16326 453558
rect 16360 453547 16394 453558
rect 16428 453547 16462 453558
rect 16496 453547 16530 453558
rect 16564 453547 16598 453558
rect 16632 453547 16666 453558
rect 17290 453547 17324 453558
rect 17358 453547 17392 453558
rect 17426 453547 17460 453558
rect 17494 453547 17528 453558
rect 17562 453547 17596 453558
rect 17630 453547 17664 453558
rect 17698 453547 17732 453558
rect 17766 453547 17800 453558
rect 17834 453547 17868 453558
rect 17902 453547 17936 453558
rect 17970 453547 18004 453558
rect 18038 453547 18072 453558
rect 18106 453547 18140 453558
rect 18174 453547 18208 453558
rect 15748 453537 15806 453547
rect 15816 453537 15874 453547
rect 15884 453537 15942 453547
rect 15952 453537 16010 453547
rect 16020 453537 16078 453547
rect 16088 453537 16146 453547
rect 16156 453537 16214 453547
rect 16224 453537 16282 453547
rect 16292 453537 16350 453547
rect 16360 453537 16418 453547
rect 16428 453537 16486 453547
rect 16496 453537 16554 453547
rect 16564 453537 16622 453547
rect 16632 453537 16690 453547
rect 17290 453537 17348 453547
rect 17358 453537 17416 453547
rect 17426 453537 17484 453547
rect 17494 453537 17552 453547
rect 17562 453537 17620 453547
rect 17630 453537 17688 453547
rect 17698 453537 17756 453547
rect 17766 453537 17824 453547
rect 17834 453537 17892 453547
rect 17902 453537 17960 453547
rect 17970 453537 18028 453547
rect 18038 453537 18096 453547
rect 18106 453537 18164 453547
rect 18174 453537 18232 453547
rect 15724 453513 16690 453537
rect 17266 453513 18232 453537
rect 15748 453498 15772 453513
rect 15816 453498 15840 453513
rect 15884 453498 15908 453513
rect 15952 453498 15976 453513
rect 16020 453498 16044 453513
rect 16088 453498 16112 453513
rect 16156 453498 16180 453513
rect 16224 453498 16248 453513
rect 16292 453498 16316 453513
rect 16360 453498 16384 453513
rect 16428 453498 16452 453513
rect 16496 453498 16520 453513
rect 16564 453498 16588 453513
rect 16632 453498 16656 453513
rect 17290 453498 17314 453513
rect 17358 453498 17382 453513
rect 17426 453498 17450 453513
rect 17494 453498 17518 453513
rect 17562 453498 17586 453513
rect 17630 453498 17654 453513
rect 17698 453498 17722 453513
rect 17766 453498 17790 453513
rect 17834 453498 17858 453513
rect 17902 453498 17926 453513
rect 17970 453498 17994 453513
rect 18038 453498 18062 453513
rect 18106 453498 18130 453513
rect 18174 453498 18198 453513
rect 15678 453343 16678 453498
rect 7389 453253 8389 453313
rect 8990 453253 9990 453313
rect 15678 453309 16690 453343
rect 17278 453333 18278 453498
rect 21413 453442 22813 453570
rect 23685 453442 25085 453570
rect 25936 453514 26936 453564
rect 26393 453511 26477 453514
rect 26726 453511 26810 453514
rect 27158 453455 27358 453583
rect 17266 453309 18278 453333
rect 15678 453298 16678 453309
rect 17278 453298 18278 453309
rect 15748 453285 15772 453298
rect 15816 453285 15840 453298
rect 15884 453285 15908 453298
rect 15952 453285 15976 453298
rect 16020 453285 16044 453298
rect 16088 453285 16112 453298
rect 16156 453285 16180 453298
rect 16224 453285 16248 453298
rect 16292 453285 16316 453298
rect 16360 453285 16384 453298
rect 16428 453285 16452 453298
rect 16496 453285 16520 453298
rect 16564 453285 16588 453298
rect 16632 453285 16656 453298
rect 17290 453285 17314 453298
rect 17358 453285 17382 453298
rect 17426 453285 17450 453298
rect 17494 453285 17518 453298
rect 17562 453285 17586 453298
rect 17630 453285 17654 453298
rect 17698 453285 17722 453298
rect 17766 453285 17790 453298
rect 17834 453285 17858 453298
rect 17902 453285 17926 453298
rect 17970 453285 17994 453298
rect 18038 453285 18062 453298
rect 18106 453285 18130 453298
rect 18174 453285 18198 453298
rect 21413 453279 22813 453407
rect 23685 453279 25085 453407
rect 27158 453279 27358 453335
rect 21413 453116 22813 453244
rect 23685 453116 25085 453244
rect 27158 453103 27358 453231
rect 26393 453100 26477 453103
rect 26726 453100 26810 453103
rect 12543 453069 12881 453085
rect 12559 452967 12865 453069
rect 7389 452895 8389 452951
rect 8990 452895 9990 452951
rect 15678 452940 16678 452996
rect 17278 452940 18278 452996
rect 21413 452953 22813 453081
rect 23685 452953 25085 453081
rect 25936 453050 26936 453100
rect 27622 453095 27672 454095
rect 27772 453095 27828 454095
rect 27928 453095 27984 454095
rect 28084 453095 28140 454095
rect 28240 453095 28296 454095
rect 28396 453637 28446 454095
rect 28396 453553 28449 453637
rect 28396 453305 28446 453553
rect 29778 453320 29802 453344
rect 28396 453221 28449 453305
rect 29802 453296 29826 453309
rect 29880 453299 29914 453333
rect 29778 453261 29802 453285
rect 29890 453275 29914 453299
rect 28396 453095 28446 453221
rect 7389 452823 8389 452879
rect 8990 452823 9990 452879
rect 15678 452868 16678 452924
rect 17278 452868 18278 452924
rect 21413 452790 22813 452918
rect 23685 452790 25085 452918
rect 25936 452894 26936 452950
rect 27158 452927 27358 452983
rect 13899 452656 14059 452660
rect 7389 452521 8389 452593
rect 8990 452521 9990 452593
rect 15678 452566 16678 452638
rect 17278 452566 18278 452638
rect 21413 452627 22813 452755
rect 23685 452627 25085 452755
rect 25936 452738 26936 452794
rect 27158 452751 27358 452879
rect 27912 452757 27962 452873
rect 27909 452673 27962 452757
rect 28082 452673 28210 452873
rect 28258 452673 28314 452873
rect 28434 452673 28562 452873
rect 28610 452673 28660 452873
rect 27917 452669 27951 452673
rect 29880 452672 29914 452706
rect 25936 452582 26936 452638
rect 27158 452581 27358 452631
rect 27274 452578 27358 452581
rect 15748 452555 15782 452566
rect 15816 452555 15850 452566
rect 15884 452555 15918 452566
rect 15952 452555 15986 452566
rect 16020 452555 16054 452566
rect 16088 452555 16122 452566
rect 16156 452555 16190 452566
rect 16224 452555 16258 452566
rect 16292 452555 16326 452566
rect 16360 452555 16394 452566
rect 16428 452555 16462 452566
rect 16496 452555 16530 452566
rect 16564 452555 16598 452566
rect 16632 452555 16666 452566
rect 17290 452555 17324 452566
rect 17358 452555 17392 452566
rect 17426 452555 17460 452566
rect 17494 452555 17528 452566
rect 17562 452555 17596 452566
rect 17630 452555 17664 452566
rect 17698 452555 17732 452566
rect 17766 452555 17800 452566
rect 17834 452555 17868 452566
rect 17902 452555 17936 452566
rect 17970 452555 18004 452566
rect 18038 452555 18072 452566
rect 18106 452555 18140 452566
rect 18174 452555 18208 452566
rect 15748 452545 15806 452555
rect 15816 452545 15874 452555
rect 15884 452545 15942 452555
rect 15952 452545 16010 452555
rect 16020 452545 16078 452555
rect 16088 452545 16146 452555
rect 16156 452545 16214 452555
rect 16224 452545 16282 452555
rect 16292 452545 16350 452555
rect 16360 452545 16418 452555
rect 16428 452545 16486 452555
rect 16496 452545 16554 452555
rect 16564 452545 16622 452555
rect 16632 452545 16690 452555
rect 17290 452545 17348 452555
rect 17358 452545 17416 452555
rect 17426 452545 17484 452555
rect 17494 452545 17552 452555
rect 17562 452545 17620 452555
rect 17630 452545 17688 452555
rect 17698 452545 17756 452555
rect 17766 452545 17824 452555
rect 17834 452545 17892 452555
rect 17902 452545 17960 452555
rect 17970 452545 18028 452555
rect 18038 452545 18096 452555
rect 18106 452545 18164 452555
rect 18174 452545 18232 452555
rect 15724 452521 16690 452545
rect 17266 452521 18232 452545
rect 13901 452510 14061 452514
rect 15748 452506 15772 452521
rect 15816 452506 15840 452521
rect 15884 452506 15908 452521
rect 15952 452506 15976 452521
rect 16020 452506 16044 452521
rect 16088 452506 16112 452521
rect 16156 452506 16180 452521
rect 16224 452506 16248 452521
rect 16292 452506 16316 452521
rect 16360 452506 16384 452521
rect 16428 452506 16452 452521
rect 16496 452506 16520 452521
rect 16564 452506 16588 452521
rect 16632 452506 16656 452521
rect 17290 452506 17314 452521
rect 17358 452506 17382 452521
rect 17426 452506 17450 452521
rect 17494 452506 17518 452521
rect 17562 452506 17586 452521
rect 17630 452506 17654 452521
rect 17698 452506 17722 452521
rect 17766 452506 17790 452521
rect 17834 452506 17858 452521
rect 17902 452506 17926 452521
rect 17970 452506 17994 452521
rect 18038 452506 18062 452521
rect 18106 452506 18130 452521
rect 18174 452506 18198 452521
rect 15678 452351 16678 452506
rect 7389 452261 8389 452321
rect 8990 452261 9990 452321
rect 15678 452317 16690 452351
rect 17278 452341 18278 452506
rect 21413 452470 22813 452520
rect 23685 452470 25085 452520
rect 25936 452432 26936 452482
rect 21349 452390 21373 452414
rect 21407 452390 21431 452414
rect 25067 452390 25091 452414
rect 25125 452390 25149 452414
rect 21383 452356 21397 452390
rect 25101 452356 25115 452390
rect 17266 452317 18278 452341
rect 21349 452332 21373 452356
rect 21407 452332 21431 452356
rect 25067 452332 25091 452356
rect 25125 452332 25149 452356
rect 27917 452325 27951 452329
rect 15678 452306 16678 452317
rect 17278 452306 18278 452317
rect 15748 452293 15772 452306
rect 15816 452293 15840 452306
rect 15884 452293 15908 452306
rect 15952 452293 15976 452306
rect 16020 452293 16044 452306
rect 16088 452293 16112 452306
rect 16156 452293 16180 452306
rect 16224 452293 16248 452306
rect 16292 452293 16316 452306
rect 16360 452293 16384 452306
rect 16428 452293 16452 452306
rect 16496 452293 16520 452306
rect 16564 452293 16588 452306
rect 16632 452293 16656 452306
rect 17290 452293 17314 452306
rect 17358 452293 17382 452306
rect 17426 452293 17450 452306
rect 17494 452293 17518 452306
rect 17562 452293 17586 452306
rect 17630 452293 17654 452306
rect 17698 452293 17722 452306
rect 17766 452293 17790 452306
rect 17834 452293 17858 452306
rect 17902 452293 17926 452306
rect 17970 452293 17994 452306
rect 18038 452293 18062 452306
rect 18106 452293 18130 452306
rect 18174 452293 18198 452306
rect 27909 452241 27962 452325
rect 21634 452101 24864 452203
rect 27912 452125 27962 452241
rect 28082 452125 28210 452325
rect 28258 452125 28314 452325
rect 28434 452125 28562 452325
rect 28610 452125 28660 452325
rect 21186 452047 21210 452071
rect 25288 452047 25312 452071
rect 21162 452023 21186 452037
rect 25312 452023 25336 452037
rect 7389 451903 8389 451959
rect 8990 451903 9990 451959
rect 15678 451948 16678 452004
rect 17278 451948 18278 452004
rect 21072 451989 21084 452013
rect 21186 451989 21210 452013
rect 25288 451989 25312 452013
rect 25414 451989 25426 452013
rect 21385 451944 21403 451948
rect 7389 451831 8389 451887
rect 8990 451831 9990 451887
rect 15678 451876 16678 451932
rect 17278 451876 18278 451932
rect 20250 451914 20316 451930
rect 21377 451914 21403 451944
rect 21385 451904 21403 451914
rect 21383 451880 21403 451904
rect 21407 451880 21415 451914
rect 25113 451904 25121 451944
rect 25101 451880 25121 451904
rect 25125 451880 25143 451948
rect 21383 451846 21419 451880
rect 25101 451846 25147 451880
rect 21383 451812 21403 451846
rect 21407 451812 21415 451846
rect 21383 451778 21419 451812
rect 21481 451784 22881 451834
rect 23617 451784 25017 451834
rect 25101 451812 25121 451846
rect 25125 451812 25143 451846
rect 25101 451778 25147 451812
rect 21383 451744 21403 451778
rect 21407 451744 21415 451778
rect 21383 451710 21419 451744
rect 21383 451676 21403 451710
rect 21407 451676 21415 451710
rect 7389 451529 8389 451601
rect 8990 451529 9990 451601
rect 15678 451574 16678 451646
rect 17278 451574 18278 451646
rect 21383 451642 21419 451676
rect 21383 451608 21403 451642
rect 21407 451608 21415 451642
rect 21481 451621 22881 451749
rect 23617 451621 25017 451749
rect 25101 451744 25121 451778
rect 25125 451744 25143 451778
rect 25101 451710 25147 451744
rect 25101 451676 25121 451710
rect 25125 451676 25143 451710
rect 25101 451642 25147 451676
rect 25101 451608 25121 451642
rect 25125 451608 25143 451642
rect 21383 451574 21419 451608
rect 15748 451563 15782 451574
rect 15816 451563 15850 451574
rect 15884 451563 15918 451574
rect 15952 451563 15986 451574
rect 16020 451563 16054 451574
rect 16088 451563 16122 451574
rect 16156 451563 16190 451574
rect 16224 451563 16258 451574
rect 16292 451563 16326 451574
rect 16360 451563 16394 451574
rect 16428 451563 16462 451574
rect 16496 451563 16530 451574
rect 16564 451563 16598 451574
rect 16632 451563 16666 451574
rect 17290 451563 17324 451574
rect 17358 451563 17392 451574
rect 17426 451563 17460 451574
rect 17494 451563 17528 451574
rect 17562 451563 17596 451574
rect 17630 451563 17664 451574
rect 17698 451563 17732 451574
rect 17766 451563 17800 451574
rect 17834 451563 17868 451574
rect 17902 451563 17936 451574
rect 17970 451563 18004 451574
rect 18038 451563 18072 451574
rect 18106 451563 18140 451574
rect 18174 451563 18208 451574
rect 15748 451553 15806 451563
rect 15816 451553 15874 451563
rect 15884 451553 15942 451563
rect 15952 451553 16010 451563
rect 16020 451553 16078 451563
rect 16088 451553 16146 451563
rect 16156 451553 16214 451563
rect 16224 451553 16282 451563
rect 16292 451553 16350 451563
rect 16360 451553 16418 451563
rect 16428 451553 16486 451563
rect 16496 451553 16554 451563
rect 16564 451553 16622 451563
rect 16632 451553 16690 451563
rect 17290 451553 17348 451563
rect 17358 451553 17416 451563
rect 17426 451553 17484 451563
rect 17494 451553 17552 451563
rect 17562 451553 17620 451563
rect 17630 451553 17688 451563
rect 17698 451553 17756 451563
rect 17766 451553 17824 451563
rect 17834 451553 17892 451563
rect 17902 451553 17960 451563
rect 17970 451553 18028 451563
rect 18038 451553 18096 451563
rect 18106 451553 18164 451563
rect 18174 451553 18232 451563
rect 15724 451529 16690 451553
rect 17266 451529 18232 451553
rect 21383 451540 21403 451574
rect 21407 451540 21415 451574
rect 15748 451514 15772 451529
rect 15816 451514 15840 451529
rect 15884 451514 15908 451529
rect 15952 451514 15976 451529
rect 16020 451514 16044 451529
rect 16088 451514 16112 451529
rect 16156 451514 16180 451529
rect 16224 451514 16248 451529
rect 16292 451514 16316 451529
rect 16360 451514 16384 451529
rect 16428 451514 16452 451529
rect 16496 451514 16520 451529
rect 16564 451514 16588 451529
rect 16632 451514 16656 451529
rect 17290 451514 17314 451529
rect 17358 451514 17382 451529
rect 17426 451514 17450 451529
rect 17494 451514 17518 451529
rect 17562 451514 17586 451529
rect 17630 451514 17654 451529
rect 17698 451514 17722 451529
rect 17766 451514 17790 451529
rect 17834 451514 17858 451529
rect 17902 451514 17926 451529
rect 17970 451514 17994 451529
rect 18038 451514 18062 451529
rect 18106 451514 18130 451529
rect 18174 451514 18198 451529
rect 5937 451318 6089 451386
rect 15678 451359 16678 451514
rect 6005 451315 6089 451318
rect 5967 451305 6059 451315
rect 6005 451275 6021 451305
rect 1288 449503 1338 450503
rect 1438 449503 1566 450503
rect 1594 449503 1644 450503
rect 5995 449493 6021 451275
rect 7389 451269 8389 451329
rect 8990 451269 9990 451329
rect 15678 451325 16690 451359
rect 17278 451349 18278 451514
rect 17266 451325 18278 451349
rect 15678 451314 16678 451325
rect 17278 451314 18278 451325
rect 21383 451506 21419 451540
rect 21383 451472 21403 451506
rect 21407 451472 21415 451506
rect 21383 451438 21419 451472
rect 21481 451458 22881 451586
rect 23617 451458 25017 451586
rect 25101 451574 25147 451608
rect 25101 451540 25121 451574
rect 25125 451540 25143 451574
rect 25101 451506 25147 451540
rect 25101 451472 25121 451506
rect 25125 451472 25143 451506
rect 25101 451438 25147 451472
rect 21383 451404 21403 451438
rect 21407 451404 21415 451438
rect 21383 451370 21419 451404
rect 21383 451336 21403 451370
rect 21407 451336 21415 451370
rect 15748 451301 15772 451314
rect 15816 451301 15840 451314
rect 15884 451301 15908 451314
rect 15952 451301 15976 451314
rect 16020 451301 16044 451314
rect 16088 451301 16112 451314
rect 16156 451301 16180 451314
rect 16224 451301 16248 451314
rect 16292 451301 16316 451314
rect 16360 451301 16384 451314
rect 16428 451301 16452 451314
rect 16496 451301 16520 451314
rect 16564 451301 16588 451314
rect 16632 451301 16656 451314
rect 17290 451301 17314 451314
rect 17358 451301 17382 451314
rect 17426 451301 17450 451314
rect 17494 451301 17518 451314
rect 17562 451301 17586 451314
rect 17630 451301 17654 451314
rect 17698 451301 17722 451314
rect 17766 451301 17790 451314
rect 17834 451301 17858 451314
rect 17902 451301 17926 451314
rect 17970 451301 17994 451314
rect 18038 451301 18062 451314
rect 18106 451301 18130 451314
rect 18174 451301 18198 451314
rect 21383 451302 21419 451336
rect 21383 451268 21403 451302
rect 21407 451268 21415 451302
rect 21481 451295 22881 451423
rect 23617 451295 25017 451423
rect 25101 451404 25121 451438
rect 25125 451404 25143 451438
rect 25101 451370 25147 451404
rect 25101 451336 25121 451370
rect 25125 451336 25143 451370
rect 25101 451302 25147 451336
rect 25101 451268 25121 451302
rect 25125 451268 25143 451302
rect 21383 451234 21419 451268
rect 21383 451200 21403 451234
rect 21407 451200 21415 451234
rect 21383 451166 21419 451200
rect 21383 451132 21403 451166
rect 21407 451132 21415 451166
rect 21481 451132 22881 451260
rect 23617 451132 25017 451260
rect 25101 451234 25147 451268
rect 25101 451200 25121 451234
rect 25125 451200 25143 451234
rect 25101 451166 25147 451200
rect 25101 451132 25121 451166
rect 25125 451132 25143 451166
rect 21383 451098 21419 451132
rect 25101 451098 25147 451132
rect 21383 451064 21403 451098
rect 21407 451064 21415 451098
rect 21383 451030 21419 451064
rect 7389 450911 8389 450967
rect 8990 450911 9990 450967
rect 15678 450956 16678 451012
rect 17278 450956 18278 451012
rect 21383 450996 21403 451030
rect 21407 450996 21415 451030
rect 21383 450962 21419 450996
rect 21481 450969 22881 451097
rect 23617 450969 25017 451097
rect 25101 451064 25121 451098
rect 25125 451064 25143 451098
rect 25101 451030 25147 451064
rect 25101 450996 25121 451030
rect 25125 450996 25143 451030
rect 25101 450962 25147 450996
rect 26478 450985 26648 451291
rect 7389 450839 8389 450895
rect 8990 450839 9990 450895
rect 15678 450884 16678 450940
rect 17278 450884 18278 450940
rect 21383 450928 21403 450962
rect 21407 450928 21415 450962
rect 21383 450894 21419 450928
rect 21383 450860 21403 450894
rect 21407 450860 21415 450894
rect 21383 450826 21419 450860
rect 21383 450792 21403 450826
rect 21407 450792 21415 450826
rect 21481 450806 22881 450934
rect 23617 450806 25017 450934
rect 25101 450928 25121 450962
rect 25125 450928 25143 450962
rect 25101 450894 25147 450928
rect 27622 450903 27672 451903
rect 27772 450903 27828 451903
rect 27928 450903 27984 451903
rect 28084 450903 28140 451903
rect 28240 450903 28296 451903
rect 28396 451777 28446 451903
rect 28396 451693 28449 451777
rect 28396 451445 28446 451693
rect 30015 451523 30027 457246
rect 32596 457239 33596 457367
rect 35255 457345 36255 457401
rect 680215 457326 680815 457382
rect 685551 457360 686551 457488
rect 689154 457439 689204 457897
rect 689151 457355 689204 457439
rect 30135 457062 30735 457112
rect 31049 457042 32049 457092
rect 32596 457083 33596 457211
rect 35255 457169 36255 457297
rect 680215 457156 680815 457206
rect 685551 457204 686551 457332
rect 35255 456993 36255 457121
rect 685551 457048 686551 457176
rect 686865 457116 687465 457166
rect 30135 456886 30735 456942
rect 31049 456886 32049 456942
rect 32596 456927 33596 456983
rect 37998 456979 38148 456991
rect 38317 456979 38467 456991
rect 679007 456980 679607 457030
rect 30135 456716 30735 456766
rect 31049 456736 32049 456786
rect 32596 456777 33596 456827
rect 35255 456823 36255 456873
rect 37998 456866 38598 456916
rect 680615 456885 680630 456900
rect 680803 456896 680815 456900
rect 680800 456885 680815 456896
rect 685551 456892 686551 456948
rect 686865 456940 687465 457068
rect 679007 456810 679607 456860
rect 35255 456754 36255 456766
rect 37998 456690 38598 456746
rect 680615 456705 680815 456885
rect 683328 456793 683928 456843
rect 682573 456717 683173 456767
rect 680615 456690 680630 456705
rect 680800 456694 680815 456705
rect 680803 456690 680815 456694
rect 30135 456600 30735 456650
rect 31049 456600 32049 456650
rect 32596 456575 33196 456625
rect 35255 456621 36255 456671
rect 680502 456649 680517 456664
rect 30135 456424 30735 456480
rect 31049 456444 32049 456500
rect 30135 456248 30735 456376
rect 31049 456288 32049 456344
rect 30135 456072 30735 456200
rect 31049 456132 32049 456188
rect 32596 456141 33196 456191
rect 30135 455896 30735 456024
rect 31049 455982 32049 456032
rect 31049 455866 32049 455916
rect 30135 455726 30735 455776
rect 31049 455710 32049 455838
rect 30135 455610 30735 455660
rect 30135 455434 30735 455562
rect 31049 455554 32049 455682
rect 31049 455398 32049 455526
rect 34152 455490 34202 456478
rect 34322 455490 34372 456478
rect 34492 456465 35092 456515
rect 35255 456445 36255 456573
rect 37998 456520 38598 456570
rect 36785 456496 36797 456500
rect 36785 456485 36800 456496
rect 36970 456485 36985 456500
rect 34492 456289 35092 456345
rect 35255 456269 36255 456325
rect 36785 456305 36985 456485
rect 36785 456294 36800 456305
rect 36785 456290 36797 456294
rect 36970 456290 36985 456305
rect 37083 456485 37098 456500
rect 37083 456305 37120 456485
rect 680480 456469 680517 456649
rect 680502 456454 680517 456469
rect 680615 456649 680630 456664
rect 680803 456660 680815 456664
rect 680800 456649 680815 456660
rect 680615 456469 680815 456649
rect 682573 456541 683173 456669
rect 683328 456617 683928 456745
rect 685551 456736 686551 456864
rect 686865 456764 687465 456820
rect 685551 456580 686551 456708
rect 686865 456588 687465 456716
rect 680615 456454 680630 456469
rect 680800 456458 680815 456469
rect 680803 456454 680815 456458
rect 683328 456441 683928 456497
rect 679002 456384 679602 456434
rect 685551 456424 686551 456552
rect 682573 456365 683173 456421
rect 686865 456412 687465 456468
rect 37083 456290 37098 456305
rect 36785 456260 36797 456264
rect 36785 456249 36800 456260
rect 36970 456249 36985 456264
rect 34492 456119 35092 456169
rect 35255 456099 36255 456149
rect 36785 456069 36985 456249
rect 679002 456208 679602 456264
rect 682573 456189 683173 456317
rect 683328 456265 683928 456321
rect 685551 456274 686551 456324
rect 686865 456236 687465 456364
rect 685551 456158 686551 456208
rect 37993 456094 38593 456144
rect 678680 456123 678704 456157
rect 36785 456058 36800 456069
rect 36785 456054 36797 456058
rect 36970 456054 36985 456069
rect 678680 456055 678704 456089
rect 679002 456038 679602 456088
rect 679061 456035 679355 456038
rect 679380 456035 679602 456038
rect 678680 455987 678704 456021
rect 682573 456013 683173 456141
rect 683328 456089 683928 456145
rect 34491 455849 35091 455899
rect 35255 455883 35855 455933
rect 37993 455924 38593 455974
rect 678680 455919 678704 455953
rect 678680 455851 678704 455885
rect 682573 455837 683173 455965
rect 683328 455913 683928 456041
rect 685551 455982 686551 456110
rect 686865 456060 687465 456116
rect 34491 455673 35091 455729
rect 35255 455707 35855 455763
rect 36785 455748 37385 455798
rect 38920 455761 38946 455787
rect 678680 455783 678704 455817
rect 685551 455806 686551 455934
rect 686865 455884 687465 456012
rect 678680 455715 678704 455749
rect 34491 455503 35091 455553
rect 35255 455531 35855 455659
rect 678680 455647 678704 455681
rect 682573 455661 683173 455789
rect 683328 455737 683928 455793
rect 685551 455630 686551 455758
rect 686865 455708 687465 455836
rect 36785 455572 37385 455628
rect 678680 455579 678704 455613
rect 683328 455567 683928 455617
rect 678680 455511 678704 455545
rect 682573 455491 683173 455541
rect 684519 455498 685119 455548
rect 34019 455418 34029 455490
rect 34152 455478 34372 455490
rect 34091 455415 34101 455418
rect 30135 455258 30735 455314
rect 31049 455242 32049 455370
rect 34091 455365 35091 455415
rect 35255 455361 35855 455411
rect 36785 455396 37385 455452
rect 678680 455443 678704 455477
rect 685551 455454 686551 455582
rect 686865 455532 687465 455660
rect 679133 455409 679283 455421
rect 679452 455409 679602 455421
rect 678680 455375 678704 455409
rect 678680 455307 678704 455341
rect 679002 455296 679602 455346
rect 684519 455342 685119 455398
rect 685551 455278 686551 455406
rect 686865 455356 687465 455484
rect 30135 455082 30735 455210
rect 31049 455086 32049 455214
rect 34091 455195 35091 455245
rect 36785 455226 37385 455276
rect 678680 455239 678704 455273
rect 34091 455192 34101 455195
rect 34202 455192 34302 455195
rect 35255 455159 35855 455209
rect 678680 455171 678704 455205
rect 684519 455192 685119 455242
rect 30135 454912 30735 454962
rect 31049 454930 32049 454986
rect 30135 454796 30735 454846
rect 31049 454774 32049 454902
rect 32481 454898 33081 454948
rect 30135 454620 30735 454748
rect 31049 454618 32049 454746
rect 32481 454742 33081 454870
rect 30135 454444 30735 454572
rect 31049 454462 32049 454590
rect 32481 454586 33081 454714
rect 34152 454532 34202 455132
rect 34302 454532 34352 455132
rect 34491 455066 35091 455116
rect 35255 455003 35855 455131
rect 36785 455094 37385 455144
rect 678680 455103 678704 455137
rect 679002 455120 679602 455176
rect 681745 455081 682345 455131
rect 682509 455069 683109 455119
rect 678680 455035 678704 455069
rect 683739 455027 684339 455077
rect 684519 455062 685119 455112
rect 685551 455102 686551 455230
rect 686865 455180 687465 455308
rect 34491 454890 35091 454946
rect 36785 454918 37385 454974
rect 678680 454967 678704 455001
rect 679002 454950 679602 455000
rect 35255 454847 35855 454903
rect 678680 454899 678704 454933
rect 680502 454915 680517 454930
rect 678680 454831 678704 454865
rect 34491 454720 35091 454770
rect 35255 454691 35855 454819
rect 36785 454742 37385 454798
rect 678680 454763 678704 454797
rect 680480 454735 680517 454915
rect 678680 454695 678704 454729
rect 680502 454720 680517 454735
rect 680615 454915 680630 454930
rect 680803 454926 680815 454930
rect 680800 454915 680815 454926
rect 681745 454925 682345 454981
rect 680615 454735 680815 454915
rect 681745 454769 682345 454897
rect 682509 454893 683109 455021
rect 684519 454906 685119 455034
rect 685551 454926 686551 455054
rect 686865 455004 687465 455060
rect 683739 454837 684339 454893
rect 686865 454828 687465 454956
rect 680615 454720 680630 454735
rect 680800 454724 680815 454735
rect 680803 454720 680815 454724
rect 680615 454679 680630 454694
rect 680803 454690 680815 454694
rect 680800 454679 680815 454690
rect 678680 454627 678704 454661
rect 35255 454541 35855 454591
rect 36785 454572 37385 454622
rect 678680 454559 678704 454593
rect 678680 454491 678704 454525
rect 679007 454524 679607 454574
rect 680615 454499 680815 454679
rect 681745 454613 682345 454741
rect 682509 454717 683109 454773
rect 684519 454750 685119 454806
rect 685551 454750 686551 454806
rect 682509 454541 683109 454669
rect 684519 454594 685119 454722
rect 685551 454594 686551 454722
rect 686865 454652 687465 454780
rect 32481 454436 33081 454486
rect 680615 454484 680630 454499
rect 680800 454488 680815 454499
rect 680803 454484 680815 454488
rect 681745 454463 682345 454513
rect 683739 454477 684339 454513
rect 30135 454268 30735 454396
rect 31049 454306 32049 454434
rect 34491 454379 35091 454429
rect 37993 454396 38593 454446
rect 678680 454423 678704 454457
rect 684519 454444 685119 454494
rect 685551 454438 686551 454566
rect 686865 454476 687465 454604
rect 32481 454306 33081 454356
rect 678680 454355 678704 454389
rect 679007 454354 679607 454404
rect 682509 454371 683109 454421
rect 33261 454287 33861 454323
rect 30135 454092 30735 454220
rect 31049 454150 32049 454278
rect 32481 454150 33081 454278
rect 34491 454203 35091 454331
rect 35255 454287 35855 454337
rect 36785 454312 36797 454316
rect 36785 454301 36800 454312
rect 36970 454301 36985 454316
rect 35255 454131 35855 454259
rect 36785 454121 36985 454301
rect 678680 454287 678704 454321
rect 684519 454314 685119 454364
rect 37993 454226 38593 454276
rect 678680 454219 678704 454253
rect 678680 454151 678704 454185
rect 680215 454178 680815 454228
rect 681745 454209 682345 454259
rect 36785 454110 36800 454121
rect 36785 454106 36797 454110
rect 36970 454106 36985 454121
rect 30135 453916 30735 454044
rect 31049 453994 32049 454050
rect 32481 453994 33081 454050
rect 34491 454027 35091 454083
rect 31049 453818 32049 453946
rect 32481 453838 33081 453966
rect 33261 453907 33861 453963
rect 34491 453851 35091 453979
rect 35255 453975 35855 454103
rect 678680 454083 678704 454117
rect 36785 454076 36797 454080
rect 36785 454065 36800 454076
rect 36970 454065 36985 454080
rect 36785 453885 36985 454065
rect 35255 453819 35855 453875
rect 36785 453874 36800 453885
rect 36785 453870 36797 453874
rect 36970 453870 36985 453885
rect 37083 454065 37098 454080
rect 37083 453885 37120 454065
rect 678680 454015 678704 454049
rect 680215 454002 680815 454058
rect 681745 454053 682345 454181
rect 682509 454030 683109 454080
rect 678680 453947 678704 453981
rect 37083 453870 37098 453885
rect 678680 453879 678704 453913
rect 681745 453897 682345 453953
rect 37998 453800 38598 453850
rect 678680 453811 678704 453845
rect 680215 453826 680815 453882
rect 30135 453740 30735 453796
rect 30135 453564 30735 453692
rect 31049 453642 32049 453770
rect 32481 453688 33081 453738
rect 33261 453723 33861 453773
rect 678680 453743 678704 453777
rect 681745 453741 682345 453869
rect 682509 453854 683109 453910
rect 34491 453681 35091 453731
rect 35255 453669 35855 453719
rect 37998 453624 38598 453680
rect 678680 453675 678704 453709
rect 680215 453656 680815 453706
rect 682509 453684 683109 453734
rect 683248 453680 683298 454268
rect 683398 453680 683448 454268
rect 684519 454158 685119 454286
rect 685551 454282 686551 454410
rect 686865 454300 687465 454428
rect 684519 454002 685119 454130
rect 685551 454126 686551 454254
rect 686865 454124 687465 454252
rect 685551 453970 686551 454098
rect 686865 453954 687465 454004
rect 684519 453852 685119 453902
rect 685551 453814 686551 453870
rect 686865 453838 687465 453888
rect 683248 453668 683448 453680
rect 685551 453658 686551 453786
rect 686865 453662 687465 453790
rect 30135 453388 30735 453516
rect 31049 453466 32049 453594
rect 32481 453558 33081 453608
rect 678680 453607 678704 453641
rect 681745 453591 682345 453641
rect 683571 453605 683581 453646
rect 678680 453539 678704 453573
rect 680215 453524 680815 453574
rect 682509 453555 683509 453605
rect 30135 453212 30735 453340
rect 31049 453290 32049 453418
rect 32481 453402 33081 453458
rect 37998 453454 38598 453504
rect 678680 453471 678704 453505
rect 685551 453502 686551 453630
rect 686865 453486 687465 453542
rect 37998 453451 38220 453454
rect 38245 453451 38539 453454
rect 678680 453403 678704 453437
rect 678680 453335 678704 453369
rect 680215 453348 680815 453404
rect 681745 453389 682345 453439
rect 682509 453385 683509 453435
rect 683278 453382 683398 453385
rect 683571 453382 683581 453385
rect 685551 453346 686551 453474
rect 32481 453252 33081 453302
rect 34427 453259 35027 453309
rect 678680 453267 678704 453301
rect 30135 453036 30735 453164
rect 31049 453114 32049 453242
rect 33672 453183 34272 453233
rect 34427 453083 35027 453211
rect 678680 453199 678704 453233
rect 680215 453172 680815 453228
rect 681745 453213 682345 453341
rect 682509 453247 683109 453297
rect 678680 453131 678704 453165
rect 30135 452860 30735 452988
rect 31049 452938 32049 453066
rect 678680 453063 678704 453097
rect 33672 453007 34272 453063
rect 31049 452762 32049 452890
rect 33672 452831 34272 452959
rect 34427 452907 35027 453035
rect 678654 453013 678680 453039
rect 680215 453002 680815 453052
rect 681745 453037 682345 453093
rect 682509 453071 683109 453127
rect 678680 452929 678704 452963
rect 678680 452861 678704 452895
rect 30135 452684 30735 452740
rect 34427 452731 35027 452859
rect 37998 452825 38148 452837
rect 38317 452825 38467 452837
rect 678680 452793 678704 452827
rect 679007 452826 679607 452876
rect 681745 452867 682345 452917
rect 682509 452901 683109 452951
rect 37998 452712 38598 452762
rect 678680 452725 678704 452759
rect 680615 452731 680630 452746
rect 680803 452742 680815 452746
rect 680800 452731 680815 452742
rect 33672 452655 34272 452711
rect 30135 452508 30735 452636
rect 31049 452592 32049 452642
rect 34427 452555 35027 452683
rect 678680 452657 678704 452691
rect 679007 452656 679607 452706
rect 37998 452536 38598 452592
rect 678680 452589 678704 452623
rect 31049 452476 32049 452526
rect 33672 452479 34272 452535
rect 678680 452521 678704 452555
rect 680615 452551 680815 452731
rect 681345 452651 682345 452701
rect 682508 452631 683108 452681
rect 680615 452536 680630 452551
rect 680800 452540 680815 452551
rect 680803 452536 680815 452540
rect 680502 452495 680517 452510
rect 678680 452453 678704 452487
rect 30135 452332 30735 452388
rect 31049 452320 32049 452448
rect 34427 452379 35027 452435
rect 37998 452366 38598 452416
rect 678680 452385 678704 452419
rect 33672 452303 34272 452359
rect 36785 452342 36797 452346
rect 36785 452331 36800 452342
rect 36970 452331 36985 452346
rect 30135 452156 30735 452284
rect 31049 452164 32049 452292
rect 30135 451980 30735 452036
rect 31049 452008 32049 452136
rect 33672 452127 34272 452255
rect 34427 452203 35027 452331
rect 36785 452151 36985 452331
rect 36785 452140 36800 452151
rect 36785 452136 36797 452140
rect 36970 452136 36985 452151
rect 37083 452331 37098 452346
rect 37083 452151 37120 452331
rect 678680 452317 678704 452351
rect 680480 452315 680517 452495
rect 680502 452300 680517 452315
rect 680615 452495 680630 452510
rect 680803 452506 680815 452510
rect 680800 452495 680815 452506
rect 680615 452315 680815 452495
rect 681345 452475 682345 452531
rect 682508 452455 683108 452511
rect 680615 452300 680630 452315
rect 680800 452304 680815 452315
rect 680803 452300 680815 452304
rect 681345 452299 682345 452427
rect 682508 452285 683108 452335
rect 683228 452322 683278 453322
rect 683398 452322 683448 453322
rect 685551 453190 686551 453318
rect 686865 453310 687465 453438
rect 685551 453034 686551 453162
rect 686865 453140 687465 453190
rect 686865 453024 687465 453074
rect 685551 452884 686551 452934
rect 686865 452848 687465 452976
rect 685551 452768 686551 452818
rect 686865 452672 687465 452800
rect 684404 452609 685004 452659
rect 685551 452612 686551 452668
rect 685551 452456 686551 452512
rect 686865 452496 687465 452624
rect 685551 452300 686551 452356
rect 686865 452320 687465 452376
rect 678680 452249 678704 452283
rect 679002 452230 679602 452280
rect 678680 452181 678704 452215
rect 37083 452136 37098 452151
rect 678680 452113 678704 452147
rect 681345 452129 682345 452179
rect 684404 452175 685004 452225
rect 685551 452150 686551 452200
rect 686865 452150 687465 452200
rect 36785 452106 36797 452110
rect 36785 452095 36800 452106
rect 36970 452095 36985 452110
rect 34427 452033 35027 452083
rect 33672 451957 34272 452007
rect 30135 451804 30735 451932
rect 36785 451915 36985 452095
rect 678680 452045 678704 452079
rect 679002 452054 679602 452110
rect 681390 452070 681424 452080
rect 681458 452070 681492 452080
rect 681526 452070 681560 452080
rect 681594 452070 681628 452080
rect 681662 452070 681696 452080
rect 681730 452070 681764 452080
rect 681798 452070 681832 452080
rect 681866 452070 681900 452080
rect 681934 452070 681968 452080
rect 682002 452070 682036 452080
rect 682077 452070 682111 452080
rect 682145 452070 682179 452080
rect 682213 452070 682247 452080
rect 682281 452070 682315 452080
rect 681345 452034 682345 452046
rect 37993 451940 38593 451990
rect 678680 451977 678704 452011
rect 31049 451852 32049 451908
rect 36785 451904 36800 451915
rect 36785 451900 36797 451904
rect 36970 451900 36985 451915
rect 678680 451909 678704 451943
rect 679002 451884 679602 451934
rect 681345 451927 682345 451977
rect 684004 451973 685004 452023
rect 685551 452014 686551 452064
rect 686865 452034 687465 452084
rect 679061 451881 679355 451884
rect 679380 451881 679602 451884
rect 678680 451841 678704 451875
rect 31049 451696 32049 451824
rect 37993 451770 38593 451820
rect 678680 451773 678704 451807
rect 681345 451751 682345 451879
rect 684004 451817 685004 451873
rect 685551 451858 686551 451914
rect 686865 451858 687465 451914
rect 686686 451812 686714 451840
rect 678680 451705 678704 451739
rect 30135 451634 30735 451684
rect 31049 451540 32049 451668
rect 36785 451594 37385 451644
rect 678680 451637 678704 451671
rect 678680 451569 678704 451603
rect 681345 451575 682345 451703
rect 684004 451661 685004 451789
rect 685551 451708 686551 451758
rect 686865 451688 687465 451738
rect 28396 451361 28449 451445
rect 31049 451384 32049 451512
rect 678680 451501 678704 451535
rect 684004 451505 685004 451633
rect 687573 451554 687585 457277
rect 689154 457107 689204 457355
rect 689151 457023 689204 457107
rect 689154 456897 689204 457023
rect 689304 456897 689360 457897
rect 689460 456897 689516 457897
rect 689616 456897 689672 457897
rect 689772 456897 689828 457897
rect 689928 456897 689978 457897
rect 692485 457872 692521 457906
rect 692485 457838 692505 457872
rect 692509 457838 692517 457872
rect 690952 457509 691122 457815
rect 692485 457804 692521 457838
rect 692485 457770 692505 457804
rect 692509 457770 692517 457804
rect 692583 457775 693983 457903
rect 694719 457775 696119 457903
rect 696203 457872 696249 457906
rect 696203 457838 696223 457872
rect 696227 457838 696245 457872
rect 699322 457860 700322 457916
rect 700922 457860 701922 457916
rect 707610 457905 708610 457961
rect 709211 457905 710211 457961
rect 696203 457804 696249 457838
rect 696203 457770 696223 457804
rect 696227 457770 696245 457804
rect 699322 457788 700322 457844
rect 700922 457788 701922 457844
rect 707610 457833 708610 457889
rect 709211 457833 710211 457889
rect 692485 457736 692521 457770
rect 692485 457702 692505 457736
rect 692509 457702 692517 457736
rect 692485 457668 692521 457702
rect 692485 457634 692505 457668
rect 692509 457634 692517 457668
rect 692485 457600 692521 457634
rect 692583 457612 693983 457740
rect 694719 457612 696119 457740
rect 696203 457736 696249 457770
rect 696203 457702 696223 457736
rect 696227 457702 696245 457736
rect 696203 457668 696249 457702
rect 696203 457634 696223 457668
rect 696227 457634 696245 457668
rect 696203 457600 696249 457634
rect 692485 457566 692505 457600
rect 692509 457566 692517 457600
rect 692485 457532 692521 457566
rect 692485 457498 692505 457532
rect 692509 457498 692517 457532
rect 692485 457464 692521 457498
rect 692485 457430 692505 457464
rect 692509 457430 692517 457464
rect 692583 457449 693983 457577
rect 694719 457449 696119 457577
rect 696203 457566 696223 457600
rect 696227 457566 696245 457600
rect 696203 457532 696249 457566
rect 696203 457498 696223 457532
rect 696227 457498 696245 457532
rect 696203 457464 696249 457498
rect 699322 457486 700322 457558
rect 700922 457486 701922 457558
rect 707610 457531 708610 457603
rect 709211 457531 710211 457603
rect 711579 457553 711605 459307
rect 715956 458297 716006 459297
rect 716106 458297 716234 459297
rect 716262 458297 716312 459297
rect 699392 457475 699426 457486
rect 699460 457475 699494 457486
rect 699528 457475 699562 457486
rect 699596 457475 699630 457486
rect 699664 457475 699698 457486
rect 699732 457475 699766 457486
rect 699800 457475 699834 457486
rect 699868 457475 699902 457486
rect 699936 457475 699970 457486
rect 700004 457475 700038 457486
rect 700072 457475 700106 457486
rect 700140 457475 700174 457486
rect 700208 457475 700242 457486
rect 700276 457475 700310 457486
rect 700934 457475 700968 457486
rect 701002 457475 701036 457486
rect 701070 457475 701104 457486
rect 701138 457475 701172 457486
rect 701206 457475 701240 457486
rect 701274 457475 701308 457486
rect 701342 457475 701376 457486
rect 701410 457475 701444 457486
rect 701478 457475 701512 457486
rect 701546 457475 701580 457486
rect 701614 457475 701648 457486
rect 701682 457475 701716 457486
rect 701750 457475 701784 457486
rect 701818 457475 701852 457486
rect 711511 457485 711663 457553
rect 712447 457501 712557 457511
rect 711579 457482 711663 457485
rect 699392 457465 699450 457475
rect 699460 457465 699518 457475
rect 699528 457465 699586 457475
rect 699596 457465 699654 457475
rect 699664 457465 699722 457475
rect 699732 457465 699790 457475
rect 699800 457465 699858 457475
rect 699868 457465 699926 457475
rect 699936 457465 699994 457475
rect 700004 457465 700062 457475
rect 700072 457465 700130 457475
rect 700140 457465 700198 457475
rect 700208 457465 700266 457475
rect 700276 457465 700334 457475
rect 700934 457465 700992 457475
rect 701002 457465 701060 457475
rect 701070 457465 701128 457475
rect 701138 457465 701196 457475
rect 701206 457465 701264 457475
rect 701274 457465 701332 457475
rect 701342 457465 701400 457475
rect 701410 457465 701468 457475
rect 701478 457465 701536 457475
rect 701546 457465 701604 457475
rect 701614 457465 701672 457475
rect 701682 457465 701740 457475
rect 701750 457465 701808 457475
rect 701818 457465 701876 457475
rect 696203 457430 696223 457464
rect 696227 457430 696245 457464
rect 699368 457441 700334 457465
rect 700910 457441 701876 457465
rect 711541 457461 711633 457482
rect 692485 457396 692521 457430
rect 692485 457362 692505 457396
rect 692509 457362 692517 457396
rect 692485 457328 692521 457362
rect 692485 457294 692505 457328
rect 692509 457294 692517 457328
rect 692485 457260 692521 457294
rect 692583 457286 693983 457414
rect 694719 457286 696119 457414
rect 696203 457396 696249 457430
rect 699392 457426 699416 457441
rect 699460 457426 699484 457441
rect 699528 457426 699552 457441
rect 699596 457426 699620 457441
rect 699664 457426 699688 457441
rect 699732 457426 699756 457441
rect 699800 457426 699824 457441
rect 699868 457426 699892 457441
rect 699936 457426 699960 457441
rect 700004 457426 700028 457441
rect 700072 457426 700096 457441
rect 700140 457426 700164 457441
rect 700208 457426 700232 457441
rect 700276 457426 700300 457441
rect 700934 457426 700958 457441
rect 701002 457426 701026 457441
rect 701070 457426 701094 457441
rect 701138 457426 701162 457441
rect 701206 457426 701230 457441
rect 701274 457426 701298 457441
rect 701342 457426 701366 457441
rect 701410 457426 701434 457441
rect 701478 457426 701502 457441
rect 701546 457426 701570 457441
rect 701614 457426 701638 457441
rect 701682 457426 701706 457441
rect 701750 457426 701774 457441
rect 701818 457426 701842 457441
rect 696203 457362 696223 457396
rect 696227 457362 696245 457396
rect 696203 457328 696249 457362
rect 696203 457294 696223 457328
rect 696227 457294 696245 457328
rect 696203 457260 696249 457294
rect 699322 457271 700322 457426
rect 692485 457226 692505 457260
rect 692509 457226 692517 457260
rect 692485 457192 692521 457226
rect 692485 457158 692505 457192
rect 692509 457158 692517 457192
rect 692485 457124 692521 457158
rect 692485 457090 692505 457124
rect 692509 457090 692517 457124
rect 692583 457123 693983 457251
rect 694719 457123 696119 457251
rect 696203 457226 696223 457260
rect 696227 457226 696245 457260
rect 699322 457237 700334 457271
rect 700922 457261 701922 457426
rect 707610 457271 708610 457331
rect 709211 457271 710211 457331
rect 700910 457237 701922 457261
rect 699322 457226 700322 457237
rect 700922 457226 701922 457237
rect 696203 457192 696249 457226
rect 699392 457213 699416 457226
rect 699460 457213 699484 457226
rect 699528 457213 699552 457226
rect 699596 457213 699620 457226
rect 699664 457213 699688 457226
rect 699732 457213 699756 457226
rect 699800 457213 699824 457226
rect 699868 457213 699892 457226
rect 699936 457213 699960 457226
rect 700004 457213 700028 457226
rect 700072 457213 700096 457226
rect 700140 457213 700164 457226
rect 700208 457213 700232 457226
rect 700276 457213 700300 457226
rect 700934 457213 700958 457226
rect 701002 457213 701026 457226
rect 701070 457213 701094 457226
rect 701138 457213 701162 457226
rect 701206 457213 701230 457226
rect 701274 457213 701298 457226
rect 701342 457213 701366 457226
rect 701410 457213 701434 457226
rect 701478 457213 701502 457226
rect 701546 457213 701570 457226
rect 701614 457213 701638 457226
rect 701682 457213 701706 457226
rect 701750 457213 701774 457226
rect 701818 457213 701842 457226
rect 696203 457158 696223 457192
rect 696227 457158 696245 457192
rect 696203 457124 696249 457158
rect 696203 457090 696223 457124
rect 696227 457090 696245 457124
rect 692485 457056 692521 457090
rect 696203 457056 696249 457090
rect 692485 457022 692505 457056
rect 692509 457022 692517 457056
rect 696203 457022 696223 457056
rect 696227 457022 696245 457056
rect 692485 456988 692521 457022
rect 692485 456954 692505 456988
rect 692509 456954 692517 456988
rect 692583 456966 693983 457016
rect 694719 456966 696119 457016
rect 696203 456988 696249 457022
rect 696203 456954 696223 456988
rect 696227 456954 696245 456988
rect 692485 456920 692521 456954
rect 696203 456920 696249 456954
rect 692485 456896 692505 456920
rect 692487 456852 692505 456896
rect 692509 456886 692517 456920
rect 696203 456896 696223 456920
rect 696215 456886 696223 456896
rect 696227 456852 696245 456920
rect 697284 456870 697350 456886
rect 699322 456868 700322 456924
rect 700922 456868 701922 456924
rect 707610 456913 708610 456969
rect 709211 456913 710211 456969
rect 692174 456787 692186 456811
rect 692288 456787 692312 456811
rect 696390 456787 696414 456811
rect 696516 456787 696528 456811
rect 699322 456796 700322 456852
rect 700922 456796 701922 456852
rect 707610 456841 708610 456897
rect 709211 456841 710211 456897
rect 692264 456763 692288 456777
rect 696414 456763 696438 456777
rect 692288 456729 692312 456753
rect 696390 456729 696414 456753
rect 688940 456475 688990 456675
rect 689110 456475 689238 456675
rect 689286 456475 689342 456675
rect 689462 456475 689590 456675
rect 689638 456559 689688 456675
rect 692736 456597 695966 456699
rect 689638 456475 689691 456559
rect 699322 456494 700322 456566
rect 700922 456494 701922 456566
rect 707610 456539 708610 456611
rect 709211 456539 710211 456611
rect 699392 456483 699426 456494
rect 699460 456483 699494 456494
rect 699528 456483 699562 456494
rect 699596 456483 699630 456494
rect 699664 456483 699698 456494
rect 699732 456483 699766 456494
rect 699800 456483 699834 456494
rect 699868 456483 699902 456494
rect 699936 456483 699970 456494
rect 700004 456483 700038 456494
rect 700072 456483 700106 456494
rect 700140 456483 700174 456494
rect 700208 456483 700242 456494
rect 700276 456483 700310 456494
rect 700934 456483 700968 456494
rect 701002 456483 701036 456494
rect 701070 456483 701104 456494
rect 701138 456483 701172 456494
rect 701206 456483 701240 456494
rect 701274 456483 701308 456494
rect 701342 456483 701376 456494
rect 701410 456483 701444 456494
rect 701478 456483 701512 456494
rect 701546 456483 701580 456494
rect 701614 456483 701648 456494
rect 701682 456483 701716 456494
rect 701750 456483 701784 456494
rect 701818 456483 701852 456494
rect 689649 456471 689683 456475
rect 699392 456473 699450 456483
rect 699460 456473 699518 456483
rect 699528 456473 699586 456483
rect 699596 456473 699654 456483
rect 699664 456473 699722 456483
rect 699732 456473 699790 456483
rect 699800 456473 699858 456483
rect 699868 456473 699926 456483
rect 699936 456473 699994 456483
rect 700004 456473 700062 456483
rect 700072 456473 700130 456483
rect 700140 456473 700198 456483
rect 700208 456473 700266 456483
rect 700276 456473 700334 456483
rect 700934 456473 700992 456483
rect 701002 456473 701060 456483
rect 701070 456473 701128 456483
rect 701138 456473 701196 456483
rect 701206 456473 701264 456483
rect 701274 456473 701332 456483
rect 701342 456473 701400 456483
rect 701410 456473 701468 456483
rect 701478 456473 701536 456483
rect 701546 456473 701604 456483
rect 701614 456473 701672 456483
rect 701682 456473 701740 456483
rect 701750 456473 701808 456483
rect 701818 456473 701876 456483
rect 692451 456444 692475 456468
rect 692509 456444 692533 456468
rect 696169 456444 696193 456468
rect 696227 456444 696251 456468
rect 699368 456449 700334 456473
rect 700910 456449 701876 456473
rect 692485 456410 692499 456444
rect 696203 456410 696217 456444
rect 699392 456434 699416 456449
rect 699460 456434 699484 456449
rect 699528 456434 699552 456449
rect 699596 456434 699620 456449
rect 699664 456434 699688 456449
rect 699732 456434 699756 456449
rect 699800 456434 699824 456449
rect 699868 456434 699892 456449
rect 699936 456434 699960 456449
rect 700004 456434 700028 456449
rect 700072 456434 700096 456449
rect 700140 456434 700164 456449
rect 700208 456434 700232 456449
rect 700276 456434 700300 456449
rect 700934 456434 700958 456449
rect 701002 456434 701026 456449
rect 701070 456434 701094 456449
rect 701138 456434 701162 456449
rect 701206 456434 701230 456449
rect 701274 456434 701298 456449
rect 701342 456434 701366 456449
rect 701410 456434 701434 456449
rect 701478 456434 701502 456449
rect 701546 456434 701570 456449
rect 701614 456434 701638 456449
rect 701682 456434 701706 456449
rect 701750 456434 701774 456449
rect 701818 456434 701842 456449
rect 692451 456386 692475 456410
rect 692509 456386 692533 456410
rect 696169 456386 696193 456410
rect 696227 456386 696251 456410
rect 690664 456318 691664 456368
rect 692515 456280 693915 456330
rect 694787 456280 696187 456330
rect 699322 456279 700322 456434
rect 699322 456245 700334 456279
rect 700922 456269 701922 456434
rect 703539 456286 703699 456290
rect 707610 456279 708610 456339
rect 709211 456279 710211 456339
rect 700910 456245 701922 456269
rect 690242 456219 690326 456222
rect 690242 456214 690442 456219
rect 690238 456180 690442 456214
rect 690242 456169 690442 456180
rect 690664 456162 691664 456218
rect 687686 456128 687720 456162
rect 687686 456104 687710 456128
rect 689649 456127 689683 456131
rect 688940 455927 688990 456127
rect 689110 455927 689238 456127
rect 689286 455927 689342 456127
rect 689462 455927 689590 456127
rect 689638 456043 689691 456127
rect 689638 455927 689688 456043
rect 690242 455993 690442 456121
rect 692515 456117 693915 456245
rect 694787 456117 696187 456245
rect 699322 456234 700322 456245
rect 700922 456234 701922 456245
rect 699392 456221 699416 456234
rect 699460 456221 699484 456234
rect 699528 456221 699552 456234
rect 699596 456221 699620 456234
rect 699664 456221 699688 456234
rect 699732 456221 699756 456234
rect 699800 456221 699824 456234
rect 699868 456221 699892 456234
rect 699936 456221 699960 456234
rect 700004 456221 700028 456234
rect 700072 456221 700096 456234
rect 700140 456221 700164 456234
rect 700208 456221 700232 456234
rect 700276 456221 700300 456234
rect 700934 456221 700958 456234
rect 701002 456221 701026 456234
rect 701070 456221 701094 456234
rect 701138 456221 701162 456234
rect 701206 456221 701230 456234
rect 701274 456221 701298 456234
rect 701342 456221 701366 456234
rect 701410 456221 701434 456234
rect 701478 456221 701502 456234
rect 701546 456221 701570 456234
rect 701614 456221 701638 456234
rect 701682 456221 701706 456234
rect 701750 456221 701774 456234
rect 701818 456221 701842 456234
rect 703541 456140 703701 456144
rect 690664 456006 691664 456062
rect 692515 455954 693915 456082
rect 694787 455954 696187 456082
rect 690242 455817 690442 455873
rect 690664 455850 691664 455906
rect 692515 455791 693915 455919
rect 694787 455791 696187 455919
rect 699322 455876 700322 455932
rect 700922 455876 701922 455932
rect 707610 455921 708610 455977
rect 709211 455921 710211 455977
rect 699322 455804 700322 455860
rect 700922 455804 701922 455860
rect 707610 455849 708610 455905
rect 709211 455849 710211 455905
rect 689154 455579 689204 455705
rect 687686 455501 687720 455535
rect 687798 455515 687822 455539
rect 687774 455491 687798 455504
rect 689151 455495 689204 455579
rect 687798 455456 687822 455480
rect 689154 455247 689204 455495
rect 689151 455163 689204 455247
rect 689154 454705 689204 455163
rect 689304 454705 689360 455705
rect 689460 454705 689516 455705
rect 689616 454705 689672 455705
rect 689772 454705 689828 455705
rect 689928 454705 689978 455705
rect 690242 455641 690442 455769
rect 690664 455700 691664 455750
rect 690790 455697 690874 455700
rect 691123 455697 691207 455700
rect 692515 455628 693915 455756
rect 694787 455628 696187 455756
rect 704735 455731 705041 455833
rect 704719 455715 705057 455731
rect 690242 455465 690442 455521
rect 692515 455465 693915 455593
rect 694787 455465 696187 455593
rect 699322 455502 700322 455574
rect 700922 455502 701922 455574
rect 707610 455547 708610 455619
rect 709211 455547 710211 455619
rect 699392 455491 699426 455502
rect 699460 455491 699494 455502
rect 699528 455491 699562 455502
rect 699596 455491 699630 455502
rect 699664 455491 699698 455502
rect 699732 455491 699766 455502
rect 699800 455491 699834 455502
rect 699868 455491 699902 455502
rect 699936 455491 699970 455502
rect 700004 455491 700038 455502
rect 700072 455491 700106 455502
rect 700140 455491 700174 455502
rect 700208 455491 700242 455502
rect 700276 455491 700310 455502
rect 700934 455491 700968 455502
rect 701002 455491 701036 455502
rect 701070 455491 701104 455502
rect 701138 455491 701172 455502
rect 701206 455491 701240 455502
rect 701274 455491 701308 455502
rect 701342 455491 701376 455502
rect 701410 455491 701444 455502
rect 701478 455491 701512 455502
rect 701546 455491 701580 455502
rect 701614 455491 701648 455502
rect 701682 455491 701716 455502
rect 701750 455491 701784 455502
rect 701818 455491 701852 455502
rect 699392 455481 699450 455491
rect 699460 455481 699518 455491
rect 699528 455481 699586 455491
rect 699596 455481 699654 455491
rect 699664 455481 699722 455491
rect 699732 455481 699790 455491
rect 699800 455481 699858 455491
rect 699868 455481 699926 455491
rect 699936 455481 699994 455491
rect 700004 455481 700062 455491
rect 700072 455481 700130 455491
rect 700140 455481 700198 455491
rect 700208 455481 700266 455491
rect 700276 455481 700334 455491
rect 700934 455481 700992 455491
rect 701002 455481 701060 455491
rect 701070 455481 701128 455491
rect 701138 455481 701196 455491
rect 701206 455481 701264 455491
rect 701274 455481 701332 455491
rect 701342 455481 701400 455491
rect 701410 455481 701468 455491
rect 701478 455481 701536 455491
rect 701546 455481 701604 455491
rect 701614 455481 701672 455491
rect 701682 455481 701740 455491
rect 701750 455481 701808 455491
rect 701818 455481 701876 455491
rect 699368 455457 700334 455481
rect 700910 455457 701876 455481
rect 699392 455442 699416 455457
rect 699460 455442 699484 455457
rect 699528 455442 699552 455457
rect 699596 455442 699620 455457
rect 699664 455442 699688 455457
rect 699732 455442 699756 455457
rect 699800 455442 699824 455457
rect 699868 455442 699892 455457
rect 699936 455442 699960 455457
rect 700004 455442 700028 455457
rect 700072 455442 700096 455457
rect 700140 455442 700164 455457
rect 700208 455442 700232 455457
rect 700276 455442 700300 455457
rect 700934 455442 700958 455457
rect 701002 455442 701026 455457
rect 701070 455442 701094 455457
rect 701138 455442 701162 455457
rect 701206 455442 701230 455457
rect 701274 455442 701298 455457
rect 701342 455442 701366 455457
rect 701410 455442 701434 455457
rect 701478 455442 701502 455457
rect 701546 455442 701570 455457
rect 701614 455442 701638 455457
rect 701682 455442 701706 455457
rect 701750 455442 701774 455457
rect 701818 455442 701842 455457
rect 690242 455289 690442 455417
rect 692515 455302 693915 455430
rect 694787 455302 696187 455430
rect 690790 455286 690874 455289
rect 691123 455286 691207 455289
rect 699322 455287 700322 455442
rect 690664 455236 691664 455286
rect 699322 455253 700334 455287
rect 700922 455277 701922 455442
rect 707610 455287 708610 455347
rect 709211 455287 710211 455347
rect 700910 455253 701922 455277
rect 699322 455242 700322 455253
rect 700922 455242 701922 455253
rect 699392 455229 699416 455242
rect 699460 455229 699484 455242
rect 699528 455229 699552 455242
rect 699596 455229 699620 455242
rect 699664 455229 699688 455242
rect 699732 455229 699756 455242
rect 699800 455229 699824 455242
rect 699868 455229 699892 455242
rect 699936 455229 699960 455242
rect 700004 455229 700028 455242
rect 700072 455229 700096 455242
rect 700140 455229 700164 455242
rect 700208 455229 700232 455242
rect 700276 455229 700300 455242
rect 700934 455229 700958 455242
rect 701002 455229 701026 455242
rect 701070 455229 701094 455242
rect 701138 455229 701162 455242
rect 701206 455229 701230 455242
rect 701274 455229 701298 455242
rect 701342 455229 701366 455242
rect 701410 455229 701434 455242
rect 701478 455229 701502 455242
rect 701546 455229 701570 455242
rect 701614 455229 701638 455242
rect 701682 455229 701706 455242
rect 701750 455229 701774 455242
rect 701818 455229 701842 455242
rect 690242 455113 690442 455169
rect 692515 455152 693915 455195
rect 694787 455152 696187 455195
rect 690664 455080 691664 455136
rect 690242 454937 690442 455065
rect 692515 455016 693915 455059
rect 694787 455016 696187 455059
rect 690664 454924 691664 454980
rect 692515 454853 693915 454981
rect 694787 454853 696187 454981
rect 703541 454944 703701 454948
rect 699322 454884 700322 454940
rect 700922 454884 701922 454940
rect 707610 454929 708610 454985
rect 709211 454929 710211 454985
rect 690242 454806 690442 454817
rect 690238 454772 690442 454806
rect 690242 454767 690442 454772
rect 690664 454768 691664 454824
rect 690242 454764 690326 454767
rect 692515 454690 693915 454818
rect 694787 454690 696187 454818
rect 699322 454812 700322 454868
rect 700922 454812 701922 454868
rect 707610 454857 708610 454913
rect 709211 454857 710211 454913
rect 703541 454798 703701 454802
rect 690664 454618 691664 454668
rect 692515 454527 693915 454655
rect 694787 454527 696187 454655
rect 699322 454510 700322 454582
rect 700922 454510 701922 454582
rect 707610 454555 708610 454627
rect 709211 454555 710211 454627
rect 699392 454499 699426 454510
rect 699460 454499 699494 454510
rect 699528 454499 699562 454510
rect 699596 454499 699630 454510
rect 699664 454499 699698 454510
rect 699732 454499 699766 454510
rect 699800 454499 699834 454510
rect 699868 454499 699902 454510
rect 699936 454499 699970 454510
rect 700004 454499 700038 454510
rect 700072 454499 700106 454510
rect 700140 454499 700174 454510
rect 700208 454499 700242 454510
rect 700276 454499 700310 454510
rect 700934 454499 700968 454510
rect 701002 454499 701036 454510
rect 701070 454499 701104 454510
rect 701138 454499 701172 454510
rect 701206 454499 701240 454510
rect 701274 454499 701308 454510
rect 701342 454499 701376 454510
rect 701410 454499 701444 454510
rect 701478 454499 701512 454510
rect 701546 454499 701580 454510
rect 701614 454499 701648 454510
rect 701682 454499 701716 454510
rect 701750 454499 701784 454510
rect 701818 454499 701852 454510
rect 692515 454364 693915 454492
rect 694787 454364 696187 454492
rect 699392 454489 699450 454499
rect 699460 454489 699518 454499
rect 699528 454489 699586 454499
rect 699596 454489 699654 454499
rect 699664 454489 699722 454499
rect 699732 454489 699790 454499
rect 699800 454489 699858 454499
rect 699868 454489 699926 454499
rect 699936 454489 699994 454499
rect 700004 454489 700062 454499
rect 700072 454489 700130 454499
rect 700140 454489 700198 454499
rect 700208 454489 700266 454499
rect 700276 454489 700334 454499
rect 700934 454489 700992 454499
rect 701002 454489 701060 454499
rect 701070 454489 701128 454499
rect 701138 454489 701196 454499
rect 701206 454489 701264 454499
rect 701274 454489 701332 454499
rect 701342 454489 701400 454499
rect 701410 454489 701468 454499
rect 701478 454489 701536 454499
rect 701546 454489 701604 454499
rect 701614 454489 701672 454499
rect 701682 454489 701740 454499
rect 701750 454489 701808 454499
rect 701818 454489 701876 454499
rect 699368 454465 700334 454489
rect 700910 454465 701876 454489
rect 699392 454450 699416 454465
rect 699460 454450 699484 454465
rect 699528 454450 699552 454465
rect 699596 454450 699620 454465
rect 699664 454450 699688 454465
rect 699732 454450 699756 454465
rect 699800 454450 699824 454465
rect 699868 454450 699892 454465
rect 699936 454450 699960 454465
rect 700004 454450 700028 454465
rect 700072 454450 700096 454465
rect 700140 454450 700164 454465
rect 700208 454450 700232 454465
rect 700276 454450 700300 454465
rect 700934 454450 700958 454465
rect 701002 454450 701026 454465
rect 701070 454450 701094 454465
rect 701138 454450 701162 454465
rect 701206 454450 701230 454465
rect 701274 454450 701298 454465
rect 701342 454450 701366 454465
rect 701410 454450 701434 454465
rect 701478 454450 701502 454465
rect 701546 454450 701570 454465
rect 701614 454450 701638 454465
rect 701682 454450 701706 454465
rect 701750 454450 701774 454465
rect 701818 454450 701842 454465
rect 692515 454201 693915 454329
rect 694787 454201 696187 454329
rect 699322 454295 700322 454450
rect 699322 454261 700334 454295
rect 700922 454285 701922 454450
rect 707610 454295 708610 454355
rect 709211 454295 710211 454355
rect 700910 454261 701922 454285
rect 699322 454250 700322 454261
rect 700922 454250 701922 454261
rect 699392 454237 699416 454250
rect 699460 454237 699484 454250
rect 699528 454237 699552 454250
rect 699596 454237 699620 454250
rect 699664 454237 699688 454250
rect 699732 454237 699756 454250
rect 699800 454237 699824 454250
rect 699868 454237 699892 454250
rect 699936 454237 699960 454250
rect 700004 454237 700028 454250
rect 700072 454237 700096 454250
rect 700140 454237 700164 454250
rect 700208 454237 700232 454250
rect 700276 454237 700300 454250
rect 700934 454237 700958 454250
rect 701002 454237 701026 454250
rect 701070 454237 701094 454250
rect 701138 454237 701162 454250
rect 701206 454237 701230 454250
rect 701274 454237 701298 454250
rect 701342 454237 701366 454250
rect 701410 454237 701434 454250
rect 701478 454237 701502 454250
rect 701546 454237 701570 454250
rect 701614 454237 701638 454250
rect 701682 454237 701706 454250
rect 701750 454237 701774 454250
rect 701818 454237 701842 454250
rect 692515 454038 693915 454166
rect 694787 454038 696187 454166
rect 692047 453468 696655 454004
rect 699322 453892 700322 453948
rect 700922 453892 701922 453948
rect 707610 453937 708610 453993
rect 709211 453937 710211 453993
rect 699322 453820 700322 453876
rect 700922 453820 701922 453876
rect 707610 453865 708610 453921
rect 709211 453865 710211 453921
rect 697314 453582 697620 453752
rect 699322 453518 700322 453590
rect 700922 453518 701922 453590
rect 707610 453563 708610 453635
rect 709211 453563 710211 453635
rect 704719 453527 705057 453543
rect 699392 453507 699426 453518
rect 699460 453507 699494 453518
rect 699528 453507 699562 453518
rect 699596 453507 699630 453518
rect 699664 453507 699698 453518
rect 699732 453507 699766 453518
rect 699800 453507 699834 453518
rect 699868 453507 699902 453518
rect 699936 453507 699970 453518
rect 700004 453507 700038 453518
rect 700072 453507 700106 453518
rect 700140 453507 700174 453518
rect 700208 453507 700242 453518
rect 700276 453507 700310 453518
rect 700934 453507 700968 453518
rect 701002 453507 701036 453518
rect 701070 453507 701104 453518
rect 701138 453507 701172 453518
rect 701206 453507 701240 453518
rect 701274 453507 701308 453518
rect 701342 453507 701376 453518
rect 701410 453507 701444 453518
rect 701478 453507 701512 453518
rect 701546 453507 701580 453518
rect 701614 453507 701648 453518
rect 701682 453507 701716 453518
rect 701750 453507 701784 453518
rect 701818 453507 701852 453518
rect 699392 453497 699450 453507
rect 699460 453497 699518 453507
rect 699528 453497 699586 453507
rect 699596 453497 699654 453507
rect 699664 453497 699722 453507
rect 699732 453497 699790 453507
rect 699800 453497 699858 453507
rect 699868 453497 699926 453507
rect 699936 453497 699994 453507
rect 700004 453497 700062 453507
rect 700072 453497 700130 453507
rect 700140 453497 700198 453507
rect 700208 453497 700266 453507
rect 700276 453497 700334 453507
rect 700934 453497 700992 453507
rect 701002 453497 701060 453507
rect 701070 453497 701128 453507
rect 701138 453497 701196 453507
rect 701206 453497 701264 453507
rect 701274 453497 701332 453507
rect 701342 453497 701400 453507
rect 701410 453497 701468 453507
rect 701478 453497 701536 453507
rect 701546 453497 701604 453507
rect 701614 453497 701672 453507
rect 701682 453497 701740 453507
rect 701750 453497 701808 453507
rect 701818 453497 701876 453507
rect 699368 453473 700334 453497
rect 700910 453473 701876 453497
rect 699392 453458 699416 453473
rect 699460 453458 699484 453473
rect 699528 453458 699552 453473
rect 699596 453458 699620 453473
rect 699664 453458 699688 453473
rect 699732 453458 699756 453473
rect 699800 453458 699824 453473
rect 699868 453458 699892 453473
rect 699936 453458 699960 453473
rect 700004 453458 700028 453473
rect 700072 453458 700096 453473
rect 700140 453458 700164 453473
rect 700208 453458 700232 453473
rect 700276 453458 700300 453473
rect 700934 453458 700958 453473
rect 701002 453458 701026 453473
rect 701070 453458 701094 453473
rect 701138 453458 701162 453473
rect 701206 453458 701230 453473
rect 701274 453458 701298 453473
rect 701342 453458 701366 453473
rect 701410 453458 701434 453473
rect 701478 453458 701502 453473
rect 701546 453458 701570 453473
rect 701614 453458 701638 453473
rect 701682 453458 701706 453473
rect 701750 453458 701774 453473
rect 701818 453458 701842 453473
rect 699322 453303 700322 453458
rect 692463 453268 692511 453292
rect 696191 453268 696239 453292
rect 692487 453214 692511 453268
rect 696215 453214 696239 453268
rect 699322 453269 700334 453303
rect 700922 453293 701922 453458
rect 704735 453425 705041 453527
rect 707610 453303 708610 453363
rect 709211 453303 710211 453363
rect 700910 453269 701922 453293
rect 699322 453258 700322 453269
rect 700922 453258 701922 453269
rect 699392 453245 699416 453258
rect 699460 453245 699484 453258
rect 699528 453245 699552 453258
rect 699596 453245 699620 453258
rect 699664 453245 699688 453258
rect 699732 453245 699756 453258
rect 699800 453245 699824 453258
rect 699868 453245 699892 453258
rect 699936 453245 699960 453258
rect 700004 453245 700028 453258
rect 700072 453245 700096 453258
rect 700140 453245 700164 453258
rect 700208 453245 700232 453258
rect 700276 453245 700300 453258
rect 700934 453245 700958 453258
rect 701002 453245 701026 453258
rect 701070 453245 701094 453258
rect 701138 453245 701162 453258
rect 701206 453245 701230 453258
rect 701274 453245 701298 453258
rect 701342 453245 701366 453258
rect 701410 453245 701434 453258
rect 701478 453245 701502 453258
rect 701546 453245 701570 453258
rect 701614 453245 701638 453258
rect 701682 453245 701706 453258
rect 701750 453245 701774 453258
rect 701818 453245 701842 453258
rect 692463 453190 692511 453214
rect 696191 453190 696239 453214
rect 687686 453119 687720 453153
rect 687798 453141 687822 453165
rect 687686 453095 687710 453119
rect 687774 453117 687798 453129
rect 687798 453081 687822 453105
rect 692450 453037 692474 453061
rect 692508 453037 692532 453061
rect 696170 453037 696194 453061
rect 696228 453037 696252 453061
rect 692484 453013 692498 453037
rect 696204 453013 696218 453037
rect 692484 452935 692487 452959
rect 696215 452935 696218 452959
rect 692508 452911 692532 452935
rect 696170 452911 696194 452935
rect 699322 452900 700322 452956
rect 700922 452900 701922 452956
rect 707610 452945 708610 453001
rect 709211 452945 710211 453001
rect 692515 452805 693915 452848
rect 694787 452805 696187 452848
rect 699322 452828 700322 452884
rect 700922 452828 701922 452884
rect 707610 452873 708610 452929
rect 709211 452873 710211 452929
rect 692515 452642 693915 452770
rect 694787 452642 696187 452770
rect 688883 452473 688918 452502
rect 692515 452479 693915 452607
rect 694787 452479 696187 452607
rect 699322 452526 700322 452598
rect 700922 452526 701922 452598
rect 707610 452571 708610 452643
rect 709211 452571 710211 452643
rect 699392 452515 699426 452526
rect 699460 452515 699494 452526
rect 699528 452515 699562 452526
rect 699596 452515 699630 452526
rect 699664 452515 699698 452526
rect 699732 452515 699766 452526
rect 699800 452515 699834 452526
rect 699868 452515 699902 452526
rect 699936 452515 699970 452526
rect 700004 452515 700038 452526
rect 700072 452515 700106 452526
rect 700140 452515 700174 452526
rect 700208 452515 700242 452526
rect 700276 452515 700310 452526
rect 700934 452515 700968 452526
rect 701002 452515 701036 452526
rect 701070 452515 701104 452526
rect 701138 452515 701172 452526
rect 701206 452515 701240 452526
rect 701274 452515 701308 452526
rect 701342 452515 701376 452526
rect 701410 452515 701444 452526
rect 701478 452515 701512 452526
rect 701546 452515 701580 452526
rect 701614 452515 701648 452526
rect 701682 452515 701716 452526
rect 701750 452515 701784 452526
rect 701818 452515 701852 452526
rect 699392 452505 699450 452515
rect 699460 452505 699518 452515
rect 699528 452505 699586 452515
rect 699596 452505 699654 452515
rect 699664 452505 699722 452515
rect 699732 452505 699790 452515
rect 699800 452505 699858 452515
rect 699868 452505 699926 452515
rect 699936 452505 699994 452515
rect 700004 452505 700062 452515
rect 700072 452505 700130 452515
rect 700140 452505 700198 452515
rect 700208 452505 700266 452515
rect 700276 452505 700334 452515
rect 700934 452505 700992 452515
rect 701002 452505 701060 452515
rect 701070 452505 701128 452515
rect 701138 452505 701196 452515
rect 701206 452505 701264 452515
rect 701274 452505 701332 452515
rect 701342 452505 701400 452515
rect 701410 452505 701468 452515
rect 701478 452505 701536 452515
rect 701546 452505 701604 452515
rect 701614 452505 701672 452515
rect 701682 452505 701740 452515
rect 701750 452505 701808 452515
rect 701818 452505 701876 452515
rect 699368 452481 700334 452505
rect 700910 452481 701876 452505
rect 688883 452468 688884 452473
rect 688917 452468 688918 452473
rect 688917 452439 688951 452468
rect 699392 452466 699416 452481
rect 699460 452466 699484 452481
rect 699528 452466 699552 452481
rect 699596 452466 699620 452481
rect 699664 452466 699688 452481
rect 699732 452466 699756 452481
rect 699800 452466 699824 452481
rect 699868 452466 699892 452481
rect 699936 452466 699960 452481
rect 700004 452466 700028 452481
rect 700072 452466 700096 452481
rect 700140 452466 700164 452481
rect 700208 452466 700232 452481
rect 700276 452466 700300 452481
rect 700934 452466 700958 452481
rect 701002 452466 701026 452481
rect 701070 452466 701094 452481
rect 701138 452466 701162 452481
rect 701206 452466 701230 452481
rect 701274 452466 701298 452481
rect 701342 452466 701366 452481
rect 701410 452466 701434 452481
rect 701478 452466 701502 452481
rect 701546 452466 701570 452481
rect 701614 452466 701638 452481
rect 701682 452466 701706 452481
rect 701750 452466 701774 452481
rect 701818 452466 701842 452481
rect 688917 452370 688951 452404
rect 688917 452301 688951 452335
rect 692515 452316 693915 452444
rect 694787 452316 696187 452444
rect 699322 452311 700322 452466
rect 688917 452232 688951 452266
rect 688917 452163 688951 452197
rect 692515 452153 693915 452281
rect 694787 452153 696187 452281
rect 699322 452277 700334 452311
rect 700922 452301 701922 452466
rect 707610 452311 708610 452371
rect 709211 452311 710211 452371
rect 700910 452277 701922 452301
rect 699322 452266 700322 452277
rect 700922 452266 701922 452277
rect 699392 452253 699416 452266
rect 699460 452253 699484 452266
rect 699528 452253 699552 452266
rect 699596 452253 699620 452266
rect 699664 452253 699688 452266
rect 699732 452253 699756 452266
rect 699800 452253 699824 452266
rect 699868 452253 699892 452266
rect 699936 452253 699960 452266
rect 700004 452253 700028 452266
rect 700072 452253 700096 452266
rect 700140 452253 700164 452266
rect 700208 452253 700232 452266
rect 700276 452253 700300 452266
rect 700934 452253 700958 452266
rect 701002 452253 701026 452266
rect 701070 452253 701094 452266
rect 701138 452253 701162 452266
rect 701206 452253 701230 452266
rect 701274 452253 701298 452266
rect 701342 452253 701366 452266
rect 701410 452253 701434 452266
rect 701478 452253 701502 452266
rect 701546 452253 701570 452266
rect 701614 452253 701638 452266
rect 701682 452253 701706 452266
rect 701750 452253 701774 452266
rect 701818 452253 701842 452266
rect 688917 452094 688951 452128
rect 688917 452025 688951 452059
rect 692515 451996 693915 452046
rect 694787 451996 696187 452046
rect 688917 451956 688951 451990
rect 698017 451933 698120 451969
rect 688917 451887 688951 451921
rect 692463 451885 692511 451909
rect 696191 451885 696239 451909
rect 688917 451818 688951 451852
rect 692487 451831 692511 451885
rect 696215 451831 696239 451885
rect 698017 451858 698053 451933
rect 692463 451807 692511 451831
rect 696191 451807 696239 451831
rect 698030 451824 698077 451858
rect 698017 451790 698053 451824
rect 688917 451749 688951 451783
rect 698030 451756 698077 451790
rect 698017 451722 698053 451756
rect 688917 451680 688951 451714
rect 698030 451688 698077 451722
rect 698017 451654 698053 451688
rect 688917 451611 688951 451645
rect 692463 451629 692521 451653
rect 696191 451629 696249 451653
rect 692487 451619 692521 451629
rect 696215 451619 696249 451629
rect 698030 451620 698077 451654
rect 698017 451586 698053 451620
rect 686879 451544 687585 451554
rect 686882 451528 687585 451544
rect 688917 451542 688951 451576
rect 692487 451547 692521 451581
rect 696215 451547 696249 451581
rect 36785 451418 37385 451474
rect 678680 451433 678704 451467
rect 681345 451399 682345 451455
rect 678680 451365 678704 451399
rect 28396 450903 28446 451361
rect 684004 451349 685004 451477
rect 688917 451473 688951 451507
rect 692487 451475 692521 451509
rect 696215 451475 696249 451509
rect 688917 451404 688951 451438
rect 692487 451427 692521 451437
rect 696215 451427 696249 451437
rect 692463 451403 692521 451427
rect 696191 451403 696249 451427
rect 688917 451335 688951 451369
rect 31049 451234 32049 451284
rect 36785 451242 37385 451298
rect 678680 451297 678704 451331
rect 678680 451229 678704 451263
rect 679133 451255 679283 451267
rect 679452 451255 679602 451267
rect 681345 451229 682345 451279
rect 678680 451161 678704 451195
rect 684004 451193 685004 451321
rect 688917 451266 688951 451300
rect 679002 451142 679602 451192
rect 36785 451072 37385 451122
rect 678680 451093 678704 451127
rect 681441 451064 681457 451130
rect 682225 451064 682241 451130
rect 37939 451039 37963 451063
rect 38085 451039 38109 451063
rect 29925 451003 29931 451032
rect 30271 451003 30305 451027
rect 30342 451003 30376 451027
rect 30413 451003 30447 451027
rect 30484 451003 30518 451027
rect 30555 451003 30589 451027
rect 30626 451003 30660 451027
rect 30697 451003 30731 451027
rect 37963 451015 37987 451038
rect 38061 451015 38085 451038
rect 678680 451025 678704 451059
rect 684004 451037 685004 451165
rect 685537 451161 686137 451211
rect 688917 451197 688951 451231
rect 692463 451214 692521 451248
rect 696191 451214 696249 451248
rect 688917 451128 688951 451162
rect 29931 450962 29939 450986
rect 29955 450962 29961 451003
rect 29891 450938 29915 450962
rect 678680 450957 678704 450991
rect 679002 450966 679602 451022
rect 25101 450860 25121 450894
rect 25125 450860 25143 450894
rect 37759 450867 37783 450891
rect 678680 450889 678704 450923
rect 681441 450902 681457 450968
rect 683625 450902 683641 450968
rect 684004 450881 685004 451009
rect 685537 451005 686137 451061
rect 688917 451059 688951 451093
rect 692515 451084 693915 451127
rect 694787 451084 696187 451127
rect 688917 450990 688951 451024
rect 688917 450921 688951 450955
rect 692515 450921 693915 451049
rect 694787 450921 696187 451049
rect 25101 450826 25147 450860
rect 37792 450843 37807 450867
rect 685537 450855 686137 450905
rect 25101 450792 25121 450826
rect 25125 450792 25143 450826
rect 678680 450821 678704 450855
rect 679002 450796 679602 450846
rect 21383 450758 21419 450792
rect 25101 450758 25147 450792
rect 21383 450724 21403 450758
rect 21407 450724 21415 450758
rect 25101 450724 25121 450758
rect 25125 450724 25143 450758
rect 678680 450753 678704 450787
rect 680502 450761 680517 450776
rect 21383 450690 21419 450724
rect 21383 450656 21403 450690
rect 21407 450656 21415 450690
rect 21481 450656 22881 450699
rect 22892 450675 22920 450703
rect 23617 450656 25017 450699
rect 25101 450690 25147 450724
rect 31458 450703 31608 450715
rect 31777 450703 31927 450715
rect 25101 450656 25121 450690
rect 25125 450656 25143 450690
rect 678680 450685 678704 450719
rect 7389 450628 8389 450632
rect 8990 450628 9990 450632
rect 7353 450578 8425 450614
rect 7353 450537 7389 450578
rect 8389 450537 8425 450578
rect 7353 450501 8425 450537
rect 8954 450578 10026 450614
rect 15678 450582 16678 450654
rect 17278 450582 18278 450654
rect 21383 450622 21419 450656
rect 25101 450622 25147 450656
rect 21383 450588 21403 450622
rect 21407 450588 21415 450622
rect 25101 450588 25121 450622
rect 25125 450588 25143 450622
rect 8954 450537 8990 450578
rect 9990 450537 10026 450578
rect 15748 450571 15782 450582
rect 15816 450571 15850 450582
rect 15884 450571 15918 450582
rect 15952 450571 15986 450582
rect 16020 450571 16054 450582
rect 16088 450571 16122 450582
rect 16156 450571 16190 450582
rect 16224 450571 16258 450582
rect 16292 450571 16326 450582
rect 16360 450571 16394 450582
rect 16428 450571 16462 450582
rect 16496 450571 16530 450582
rect 16564 450571 16598 450582
rect 16632 450571 16666 450582
rect 17290 450571 17324 450582
rect 17358 450571 17392 450582
rect 17426 450571 17460 450582
rect 17494 450571 17528 450582
rect 17562 450571 17596 450582
rect 17630 450571 17664 450582
rect 17698 450571 17732 450582
rect 17766 450571 17800 450582
rect 17834 450571 17868 450582
rect 17902 450571 17936 450582
rect 17970 450571 18004 450582
rect 18038 450571 18072 450582
rect 18106 450571 18140 450582
rect 18174 450571 18208 450582
rect 15748 450561 15806 450571
rect 15816 450561 15874 450571
rect 15884 450561 15942 450571
rect 15952 450561 16010 450571
rect 16020 450561 16078 450571
rect 16088 450561 16146 450571
rect 16156 450561 16214 450571
rect 16224 450561 16282 450571
rect 16292 450561 16350 450571
rect 16360 450561 16418 450571
rect 16428 450561 16486 450571
rect 16496 450561 16554 450571
rect 16564 450561 16622 450571
rect 16632 450561 16690 450571
rect 17290 450561 17348 450571
rect 17358 450561 17416 450571
rect 17426 450561 17484 450571
rect 17494 450561 17552 450571
rect 17562 450561 17620 450571
rect 17630 450561 17688 450571
rect 17698 450561 17756 450571
rect 17766 450561 17824 450571
rect 17834 450561 17892 450571
rect 17902 450561 17960 450571
rect 17970 450561 18028 450571
rect 18038 450561 18096 450571
rect 18106 450561 18164 450571
rect 18174 450561 18232 450571
rect 15724 450537 16690 450561
rect 17266 450537 18232 450561
rect 21383 450554 21419 450588
rect 8954 450501 10026 450537
rect 15748 450522 15772 450537
rect 15816 450522 15840 450537
rect 15884 450522 15908 450537
rect 15952 450522 15976 450537
rect 16020 450522 16044 450537
rect 16088 450522 16112 450537
rect 16156 450522 16180 450537
rect 16224 450522 16248 450537
rect 16292 450522 16316 450537
rect 16360 450522 16384 450537
rect 16428 450522 16452 450537
rect 16496 450522 16520 450537
rect 16564 450522 16588 450537
rect 16632 450522 16656 450537
rect 17290 450522 17314 450537
rect 17358 450522 17382 450537
rect 17426 450522 17450 450537
rect 17494 450522 17518 450537
rect 17562 450522 17586 450537
rect 17630 450522 17654 450537
rect 17698 450522 17722 450537
rect 17766 450522 17790 450537
rect 17834 450522 17858 450537
rect 17902 450522 17926 450537
rect 17970 450522 17994 450537
rect 18038 450522 18062 450537
rect 18106 450522 18130 450537
rect 18174 450522 18198 450537
rect 15678 450367 16678 450522
rect 7389 450277 8389 450337
rect 8990 450277 9990 450337
rect 15678 450333 16690 450367
rect 17278 450357 18278 450522
rect 17266 450333 18278 450357
rect 15678 450322 16678 450333
rect 17278 450322 18278 450333
rect 21383 450520 21403 450554
rect 21407 450520 21415 450554
rect 21481 450520 22881 450563
rect 23617 450520 25017 450563
rect 25101 450554 25147 450588
rect 25414 450573 25438 450607
rect 31458 450590 32058 450640
rect 678680 450617 678704 450651
rect 25101 450520 25121 450554
rect 25125 450520 25143 450554
rect 678680 450549 678704 450583
rect 680480 450581 680517 450761
rect 680502 450566 680517 450581
rect 680615 450761 680630 450776
rect 680803 450772 680815 450776
rect 680800 450761 680815 450772
rect 680615 450581 680815 450761
rect 681441 450740 681457 450806
rect 683625 450740 683641 450806
rect 684004 450725 685004 450853
rect 688917 450852 688951 450886
rect 688917 450783 688951 450817
rect 692515 450758 693915 450886
rect 694787 450758 696187 450886
rect 688917 450714 688951 450748
rect 686829 450649 687429 450699
rect 688917 450645 688951 450679
rect 680615 450566 680630 450581
rect 680800 450570 680815 450581
rect 681441 450578 681457 450644
rect 682225 450578 682241 450644
rect 684004 450575 685004 450625
rect 688917 450576 688951 450610
rect 692515 450595 693915 450723
rect 694787 450595 696187 450723
rect 680803 450566 680815 450570
rect 680615 450525 680630 450540
rect 680803 450536 680815 450540
rect 680800 450525 680815 450536
rect 21383 450486 21419 450520
rect 25101 450486 25147 450520
rect 21383 450452 21403 450486
rect 21407 450452 21415 450486
rect 21383 450418 21419 450452
rect 21383 450384 21403 450418
rect 21407 450384 21415 450418
rect 21383 450350 21419 450384
rect 21481 450357 22881 450485
rect 23617 450357 25017 450485
rect 25101 450452 25121 450486
rect 25125 450452 25143 450486
rect 37792 450470 37807 450494
rect 678680 450481 678704 450515
rect 25101 450418 25147 450452
rect 25101 450384 25121 450418
rect 25125 450384 25143 450418
rect 31458 450414 32058 450470
rect 37759 450446 37783 450470
rect 678680 450413 678704 450447
rect 25101 450350 25147 450384
rect 15748 450309 15772 450322
rect 15816 450309 15840 450322
rect 15884 450309 15908 450322
rect 15952 450309 15976 450322
rect 16020 450309 16044 450322
rect 16088 450309 16112 450322
rect 16156 450309 16180 450322
rect 16224 450309 16248 450322
rect 16292 450309 16316 450322
rect 16360 450309 16384 450322
rect 16428 450309 16452 450322
rect 16496 450309 16520 450322
rect 16564 450309 16588 450322
rect 16632 450309 16656 450322
rect 17290 450309 17314 450322
rect 17358 450309 17382 450322
rect 17426 450309 17450 450322
rect 17494 450309 17518 450322
rect 17562 450309 17586 450322
rect 17630 450309 17654 450322
rect 17698 450309 17722 450322
rect 17766 450309 17790 450322
rect 17834 450309 17858 450322
rect 17902 450309 17926 450322
rect 17970 450309 17994 450322
rect 18038 450309 18062 450322
rect 18106 450309 18130 450322
rect 18174 450309 18198 450322
rect 21383 450316 21403 450350
rect 21407 450316 21415 450350
rect 21383 450282 21419 450316
rect 21383 450248 21403 450282
rect 21407 450248 21415 450282
rect 21383 450214 21419 450248
rect 21383 450180 21403 450214
rect 21407 450180 21415 450214
rect 21481 450194 22881 450322
rect 23617 450194 25017 450322
rect 25101 450316 25121 450350
rect 25125 450316 25143 450350
rect 678680 450345 678704 450379
rect 679007 450370 679607 450420
rect 680615 450345 680815 450525
rect 681345 450429 682345 450479
rect 686829 450473 687429 450529
rect 688917 450507 688951 450541
rect 688917 450438 688951 450472
rect 692515 450432 693915 450560
rect 694787 450432 696187 450560
rect 684054 450373 685054 450423
rect 688917 450393 688951 450403
rect 688893 450369 688951 450393
rect 680615 450330 680630 450345
rect 680800 450334 680815 450345
rect 680803 450330 680815 450334
rect 25101 450282 25147 450316
rect 25101 450248 25121 450282
rect 25125 450248 25143 450282
rect 25101 450214 25147 450248
rect 25101 450180 25121 450214
rect 25125 450180 25143 450214
rect 25725 450197 26325 450247
rect 31458 450244 32058 450294
rect 678680 450277 678704 450311
rect 681345 450253 682345 450309
rect 30245 450220 30257 450224
rect 30245 450209 30260 450220
rect 30430 450209 30445 450224
rect 21383 450146 21419 450180
rect 7389 450066 8389 450070
rect 8990 450066 9990 450070
rect 15678 450061 16678 450133
rect 17278 450061 18278 450133
rect 21383 450112 21403 450146
rect 21407 450112 21415 450146
rect 21383 450078 21419 450112
rect 7353 450016 8425 450052
rect 7353 449975 7389 450016
rect 8389 449975 8425 450016
rect 7353 449919 8425 449975
rect 7353 449903 7389 449919
rect 8389 449903 8425 449919
rect 7353 449847 8425 449903
rect 7353 449810 7389 449847
rect 8389 449810 8425 449847
rect 7353 449770 8425 449810
rect 8954 450016 10026 450052
rect 8954 449975 8990 450016
rect 9990 449975 10026 450016
rect 8954 449919 10026 449975
rect 21383 450044 21403 450078
rect 21407 450044 21415 450078
rect 21383 450010 21419 450044
rect 21481 450031 22881 450159
rect 23617 450031 25017 450159
rect 25101 450146 25147 450180
rect 25101 450112 25121 450146
rect 25125 450112 25143 450146
rect 25101 450078 25147 450112
rect 25101 450044 25121 450078
rect 25125 450044 25143 450078
rect 25725 450047 26325 450097
rect 25101 450010 25147 450044
rect 21383 449976 21403 450010
rect 21407 449976 21415 450010
rect 21383 449942 21419 449976
rect 8954 449903 8990 449919
rect 9990 449903 10026 449919
rect 15678 449906 16678 449923
rect 17278 449906 18278 449923
rect 21383 449908 21403 449942
rect 21407 449908 21415 449942
rect 8954 449847 10026 449903
rect 20250 449890 20316 449906
rect 8954 449810 8990 449847
rect 9990 449810 10026 449847
rect 8954 449770 10026 449810
rect 21383 449874 21419 449908
rect 21383 449840 21403 449874
rect 21407 449840 21415 449874
rect 21481 449868 22881 449996
rect 23617 449868 25017 449996
rect 25101 449976 25121 450010
rect 25125 449976 25143 450010
rect 25101 449942 25147 449976
rect 25101 449908 25121 449942
rect 25125 449908 25143 449942
rect 25725 449925 26325 449975
rect 25101 449874 25147 449908
rect 25101 449840 25121 449874
rect 25125 449840 25143 449874
rect 21383 449806 21419 449840
rect 21383 449772 21403 449806
rect 21407 449772 21415 449806
rect 21383 449738 21419 449772
rect 15678 449703 16678 449736
rect 17278 449703 18278 449736
rect 21383 449704 21403 449738
rect 21407 449704 21415 449738
rect 21481 449705 22881 449833
rect 23617 449705 25017 449833
rect 25101 449806 25147 449840
rect 25101 449772 25121 449806
rect 25125 449772 25143 449806
rect 25725 449775 26325 449825
rect 25101 449738 25147 449772
rect 25101 449704 25121 449738
rect 25125 449704 25143 449738
rect 21383 449670 21419 449704
rect 25101 449670 25147 449704
rect 21383 449636 21403 449670
rect 21407 449636 21415 449670
rect 7389 449559 8389 449631
rect 8990 449559 9990 449631
rect 21383 449602 21419 449636
rect 15840 449510 15870 449580
rect 15878 449546 15908 449580
rect 21383 449568 21403 449602
rect 21407 449568 21415 449602
rect 15853 449508 15870 449510
rect 21383 449534 21419 449568
rect 21481 449542 22881 449670
rect 23617 449542 25017 449670
rect 25101 449636 25121 449670
rect 25125 449636 25143 449670
rect 25725 449649 26325 449699
rect 25101 449602 25147 449636
rect 25101 449568 25121 449602
rect 25125 449568 25143 449602
rect 25101 449534 25147 449568
rect 5981 449483 6021 449493
rect 5137 449469 6021 449483
rect 21383 449500 21403 449534
rect 21407 449500 21415 449534
rect 21383 449466 21419 449500
rect 7389 449369 8389 449463
rect 7389 449359 8413 449369
rect 8990 449359 9990 449463
rect 21383 449432 21403 449466
rect 21407 449432 21415 449466
rect 21383 449398 21419 449432
rect 21383 449364 21403 449398
rect 21407 449364 21415 449398
rect 21481 449379 22881 449507
rect 23617 449379 25017 449507
rect 25101 449500 25121 449534
rect 25125 449500 25143 449534
rect 25101 449466 25147 449500
rect 25725 449499 26325 449549
rect 25101 449432 25121 449466
rect 25125 449432 25143 449466
rect 25101 449398 25147 449432
rect 25101 449364 25121 449398
rect 25125 449364 25143 449398
rect 25725 449377 26325 449427
rect 21383 449330 21419 449364
rect 25101 449330 25147 449364
rect 21383 449296 21403 449330
rect 21407 449296 21415 449330
rect 25101 449296 25121 449330
rect 25125 449296 25143 449330
rect 21383 449262 21419 449296
rect 21383 449228 21403 449262
rect 21407 449228 21415 449262
rect 21481 449229 22881 449272
rect 23617 449229 25017 449272
rect 25101 449262 25147 449296
rect 25101 449228 25121 449262
rect 25125 449228 25143 449262
rect 21383 449194 21419 449228
rect 25101 449194 25147 449228
rect 25725 449227 26325 449277
rect 21383 449160 21403 449194
rect 21407 449160 21415 449194
rect 25101 449160 25121 449194
rect 25125 449160 25143 449194
rect 27162 449170 27212 450170
rect 27312 449170 27440 450170
rect 27468 449170 27596 450170
rect 27624 449170 27752 450170
rect 27780 449170 27908 450170
rect 27936 449170 28064 450170
rect 28092 449170 28220 450170
rect 28248 449170 28376 450170
rect 28404 449170 28532 450170
rect 28560 449170 28688 450170
rect 28716 449170 28844 450170
rect 28872 449170 29000 450170
rect 29028 449170 29156 450170
rect 29184 449170 29312 450170
rect 29340 449170 29390 450170
rect 30245 450029 30445 450209
rect 30245 450018 30260 450029
rect 30245 450014 30257 450018
rect 30430 450014 30445 450029
rect 30543 450209 30558 450224
rect 678680 450209 678704 450243
rect 30543 450029 30580 450209
rect 679007 450200 679607 450250
rect 684054 450217 685054 450345
rect 686829 450303 687429 450353
rect 692515 450269 693915 450397
rect 694787 450269 696187 450397
rect 678680 450141 678704 450175
rect 678680 450073 678704 450107
rect 681345 450077 682345 450205
rect 30543 450014 30558 450029
rect 678680 450005 678704 450039
rect 680215 450024 680815 450074
rect 684054 450061 685054 450189
rect 685793 450182 685805 450186
rect 685793 450171 685808 450182
rect 685978 450171 685993 450186
rect 30245 449984 30257 449988
rect 30245 449973 30260 449984
rect 30430 449973 30445 449988
rect 30245 449793 30445 449973
rect 678680 449937 678704 449971
rect 678680 449869 678704 449903
rect 31453 449818 32053 449868
rect 680215 449848 680815 449904
rect 681345 449901 682345 450029
rect 684054 449905 685054 450033
rect 685793 449991 685993 450171
rect 685793 449980 685808 449991
rect 685793 449976 685805 449980
rect 685978 449976 685993 449991
rect 686053 450182 686065 450186
rect 686053 450171 686068 450182
rect 686238 450171 686253 450186
rect 686053 449991 686253 450171
rect 686607 450164 687607 450214
rect 697088 450171 697138 451571
rect 697238 450171 697366 451571
rect 697394 450171 697522 451571
rect 697550 450171 697678 451571
rect 697706 450171 697756 451571
rect 698030 451552 698077 451586
rect 698017 451518 698053 451552
rect 698030 451484 698077 451518
rect 698017 451450 698053 451484
rect 698030 451416 698077 451450
rect 698017 451382 698053 451416
rect 698030 451348 698077 451382
rect 698017 451314 698053 451348
rect 698030 451280 698077 451314
rect 698017 451246 698053 451280
rect 698030 451212 698077 451246
rect 698017 451178 698053 451212
rect 698030 451144 698077 451178
rect 698017 451110 698053 451144
rect 698030 451076 698077 451110
rect 698017 451042 698053 451076
rect 698030 451008 698077 451042
rect 698017 450974 698053 451008
rect 698030 450940 698077 450974
rect 698017 450906 698053 450940
rect 698030 450872 698077 450906
rect 698017 450838 698053 450872
rect 698030 450804 698077 450838
rect 698017 450770 698053 450804
rect 698030 450736 698077 450770
rect 698017 450702 698053 450736
rect 698030 450668 698077 450702
rect 698017 450634 698053 450668
rect 698030 450600 698077 450634
rect 698017 450566 698053 450600
rect 698030 450532 698077 450566
rect 698017 450498 698053 450532
rect 698030 450464 698077 450498
rect 698017 450430 698053 450464
rect 698030 450396 698077 450430
rect 698017 450362 698053 450396
rect 698030 450328 698077 450362
rect 698017 450294 698053 450328
rect 698030 450260 698077 450294
rect 698017 450226 698053 450260
rect 698030 450192 698077 450226
rect 692515 450119 693915 450162
rect 694787 450119 696187 450162
rect 698017 450158 698053 450192
rect 698030 450124 698077 450158
rect 698017 450090 698053 450124
rect 686607 450014 687607 450064
rect 698030 450056 698077 450090
rect 686053 449980 686068 449991
rect 686053 449976 686065 449980
rect 686238 449976 686253 449991
rect 685793 449946 685805 449950
rect 685793 449935 685808 449946
rect 685978 449935 685993 449950
rect 678680 449801 678704 449835
rect 30245 449782 30260 449793
rect 30245 449778 30257 449782
rect 30430 449778 30445 449793
rect 678680 449733 678704 449767
rect 681345 449731 682345 449781
rect 684054 449749 685054 449877
rect 685793 449755 685993 449935
rect 685793 449744 685808 449755
rect 685793 449740 685805 449744
rect 685978 449740 685993 449755
rect 686053 449946 686065 449950
rect 686053 449935 686068 449946
rect 686238 449935 686253 449950
rect 686053 449755 686253 449935
rect 686607 449855 687607 449905
rect 692463 449809 692511 449833
rect 696191 449809 696239 449833
rect 686053 449744 686068 449755
rect 686053 449740 686065 449744
rect 686238 449740 686253 449755
rect 31453 449648 32053 449698
rect 678680 449665 678704 449699
rect 680215 449672 680815 449728
rect 681345 449662 682345 449674
rect 678680 449597 678704 449631
rect 684054 449593 685054 449721
rect 686607 449705 687607 449755
rect 692487 449731 692511 449809
rect 696215 449755 696239 449809
rect 696191 449731 696239 449755
rect 696617 449772 696651 449773
rect 696617 449749 696626 449772
rect 696617 449731 696675 449749
rect 696651 449715 696675 449731
rect 696651 449647 696675 449681
rect 685533 449586 685545 449590
rect 685533 449575 685548 449586
rect 685718 449575 685733 449590
rect 678680 449529 678704 449563
rect 30245 449472 30845 449522
rect 680215 449502 680815 449552
rect 678680 449461 678704 449495
rect 678680 449393 678704 449427
rect 680215 449370 680815 449420
rect 681466 449411 682466 449461
rect 684054 449437 685054 449565
rect 30245 449296 30845 449352
rect 678680 449325 678704 449359
rect 678680 449257 678704 449291
rect 681466 449255 682466 449383
rect 682890 449339 683490 449389
rect 678680 449189 678704 449223
rect 680215 449194 680815 449250
rect 682890 449183 683490 449311
rect 684054 449281 685054 449409
rect 685533 449395 685733 449575
rect 685533 449384 685548 449395
rect 685533 449380 685545 449384
rect 685718 449380 685733 449395
rect 685793 449586 685805 449590
rect 685793 449575 685808 449586
rect 685978 449575 685993 449590
rect 685793 449395 685993 449575
rect 685793 449384 685808 449395
rect 685793 449380 685805 449384
rect 685978 449380 685993 449395
rect 686053 449586 686065 449590
rect 686053 449575 686068 449586
rect 686238 449575 686253 449590
rect 686053 449395 686253 449575
rect 686053 449384 686068 449395
rect 686053 449380 686065 449384
rect 686238 449380 686253 449395
rect 686313 449586 686325 449590
rect 686313 449575 686328 449586
rect 686498 449575 686513 449590
rect 686313 449395 686513 449575
rect 686313 449384 686328 449395
rect 686313 449380 686325 449384
rect 686498 449380 686513 449395
rect 686627 449586 686639 449590
rect 686627 449575 686642 449586
rect 686812 449575 686827 449590
rect 686627 449395 686827 449575
rect 686627 449384 686642 449395
rect 686627 449380 686639 449384
rect 686812 449380 686827 449395
rect 686887 449586 686899 449590
rect 686887 449575 686902 449586
rect 687072 449575 687087 449590
rect 686887 449395 687087 449575
rect 686887 449384 686902 449395
rect 686887 449380 686899 449384
rect 687072 449380 687087 449395
rect 687147 449586 687159 449590
rect 687147 449575 687162 449586
rect 687332 449575 687347 449590
rect 696651 449579 696675 449613
rect 687147 449395 687347 449575
rect 696651 449511 696675 449545
rect 696651 449443 696675 449477
rect 687147 449384 687162 449395
rect 687147 449380 687159 449384
rect 687332 449380 687347 449395
rect 696651 449375 696675 449409
rect 696651 449307 696675 449341
rect 685718 449215 685733 449230
rect 685679 449185 685733 449215
rect 21383 449126 21419 449160
rect 25101 449126 25147 449160
rect 21383 449102 21403 449126
rect 21385 449048 21403 449102
rect 21407 449082 21415 449126
rect 25101 449102 25121 449126
rect 25113 449082 25121 449102
rect 25125 449048 25143 449126
rect 30245 449120 30845 449176
rect 678680 449121 678704 449155
rect 681466 449105 682466 449155
rect 684054 449131 685054 449181
rect 685718 449170 685733 449185
rect 685793 449226 685805 449230
rect 685793 449215 685808 449226
rect 685978 449215 685993 449230
rect 685793 449185 685993 449215
rect 685793 449174 685808 449185
rect 685793 449170 685805 449174
rect 685978 449170 685993 449185
rect 686053 449226 686065 449230
rect 686053 449215 686068 449226
rect 686238 449215 686253 449230
rect 686812 449215 686827 449230
rect 686053 449185 686253 449215
rect 686807 449185 686827 449215
rect 686053 449174 686068 449185
rect 686053 449170 686065 449174
rect 686238 449170 686253 449185
rect 686812 449170 686827 449185
rect 686887 449226 686899 449230
rect 686887 449215 686902 449226
rect 687072 449215 687087 449230
rect 686887 449185 687087 449215
rect 686887 449174 686902 449185
rect 686887 449170 686899 449174
rect 687072 449170 687087 449185
rect 687147 449226 687159 449230
rect 687147 449215 687162 449226
rect 687332 449215 687347 449230
rect 687147 449185 687347 449215
rect 687147 449174 687162 449185
rect 687147 449170 687159 449174
rect 687332 449170 687347 449185
rect 685718 449129 685733 449144
rect 681794 449102 682466 449105
rect 685679 449099 685733 449129
rect 678680 449053 678704 449087
rect 685718 449084 685733 449099
rect 685793 449140 685805 449144
rect 685793 449129 685808 449140
rect 685978 449129 685993 449144
rect 685793 449099 685993 449129
rect 685793 449088 685808 449099
rect 685793 449084 685805 449088
rect 685978 449084 685993 449099
rect 686053 449140 686065 449144
rect 686053 449129 686068 449140
rect 686238 449129 686253 449144
rect 686812 449129 686827 449144
rect 686053 449099 686253 449129
rect 686807 449099 686827 449129
rect 686053 449088 686068 449099
rect 686053 449084 686065 449088
rect 686238 449084 686253 449099
rect 686812 449084 686827 449099
rect 686887 449140 686899 449144
rect 686887 449129 686902 449140
rect 687072 449129 687087 449144
rect 686887 449099 687087 449129
rect 686887 449088 686902 449099
rect 686887 449084 686899 449088
rect 687072 449084 687087 449099
rect 687147 449140 687159 449144
rect 687147 449129 687162 449140
rect 687332 449129 687347 449144
rect 687147 449099 687347 449129
rect 687147 449088 687162 449099
rect 687147 449084 687159 449088
rect 687332 449084 687347 449099
rect 30245 448950 30845 449000
rect 678680 448985 678704 449019
rect 680215 449018 680815 449074
rect 682890 449027 683490 449083
rect 21000 448800 21003 448920
rect 678680 448917 678704 448951
rect 21352 448885 21376 448909
rect 25122 448885 25146 448909
rect 21385 448861 21400 448885
rect 25098 448861 25113 448885
rect 21274 448783 21294 448851
rect 21410 448817 21430 448851
rect 25068 448817 25088 448851
rect 25204 448817 25224 448851
rect 678680 448849 678704 448883
rect 680215 448848 680815 448898
rect 21385 448807 21430 448817
rect 25102 448807 25137 448817
rect 21361 448783 21430 448807
rect 25089 448783 25137 448807
rect 25238 448783 25258 448817
rect 678680 448781 678704 448815
rect 678680 448713 678704 448747
rect 678680 448645 678704 448679
rect 679007 448672 679607 448722
rect 678680 448577 678704 448611
rect 680615 448577 680630 448592
rect 680803 448588 680815 448592
rect 680800 448577 680815 448588
rect 678680 448509 678704 448543
rect 679007 448502 679607 448552
rect 678680 448441 678704 448475
rect 678680 448373 678704 448407
rect 680615 448397 680815 448577
rect 681502 448505 681529 448995
rect 681866 448896 682466 449024
rect 682890 448871 683490 448999
rect 684004 448929 685004 448979
rect 685539 448940 685777 448972
rect 685803 448920 686119 448938
rect 681866 448740 682466 448868
rect 684004 448773 685004 448901
rect 682890 448721 683490 448771
rect 681866 448584 682466 448712
rect 682890 448605 683490 448655
rect 684004 448617 685004 448745
rect 681866 448434 682466 448484
rect 682890 448449 683490 448505
rect 684004 448461 685004 448589
rect 692427 448522 693027 448572
rect 680615 448382 680630 448397
rect 680800 448386 680815 448397
rect 680803 448382 680815 448386
rect 680502 448341 680517 448356
rect 678680 448305 678704 448339
rect 678680 448237 678704 448271
rect 678680 448169 678704 448203
rect 680480 448161 680517 448341
rect 680502 448146 680517 448161
rect 680615 448341 680630 448356
rect 680803 448352 680815 448356
rect 680800 448341 680815 448352
rect 680615 448161 680815 448341
rect 681866 448318 682466 448368
rect 682890 448293 683490 448349
rect 684004 448305 685004 448433
rect 692427 448366 693027 448494
rect 693888 448375 694194 448545
rect 694388 448375 694694 448545
rect 689309 448278 689909 448328
rect 681866 448168 682466 448218
rect 682041 448165 682385 448168
rect 680615 448146 680630 448161
rect 680800 448150 680815 448161
rect 680803 448146 680815 448150
rect 682890 448137 683490 448193
rect 684004 448149 685004 448277
rect 678680 448101 678704 448135
rect 679002 448076 679602 448126
rect 689309 448122 689909 448250
rect 692427 448210 693027 448338
rect 678680 448033 678704 448067
rect 678680 447965 678704 447999
rect 682890 447981 683490 448109
rect 684004 447993 685004 448121
rect 689309 447966 689909 448094
rect 692427 448054 693027 448110
rect 678680 447897 678704 447931
rect 679002 447900 679602 447956
rect 678680 447829 678704 447863
rect 682890 447825 683490 447953
rect 684004 447837 685004 447965
rect 692427 447898 693027 448026
rect 689309 447810 689909 447866
rect 678680 447761 678704 447795
rect 679002 447730 679602 447780
rect 679061 447727 679355 447730
rect 679380 447727 679602 447730
rect 678680 447693 678704 447727
rect 682890 447669 683490 447797
rect 684004 447687 685004 447737
rect 685803 447720 686119 447732
rect 685539 447716 686119 447720
rect 685513 447682 685537 447716
rect 685539 447682 685777 447716
rect 678680 447625 678704 447659
rect 689309 447654 689909 447782
rect 690910 447754 691110 447765
rect 692427 447742 693027 447870
rect 690910 447640 691110 447690
rect 678680 447557 678704 447591
rect 678680 447489 678704 447523
rect 682890 447513 683490 447569
rect 685718 447555 685733 447570
rect 684004 447485 685004 447535
rect 685679 447525 685733 447555
rect 685718 447510 685733 447525
rect 685793 447566 685805 447570
rect 685793 447555 685808 447566
rect 685978 447555 685993 447570
rect 685793 447525 685993 447555
rect 685793 447514 685808 447525
rect 685793 447510 685805 447514
rect 685978 447510 685993 447525
rect 686053 447566 686065 447570
rect 686053 447555 686068 447566
rect 686238 447555 686253 447570
rect 686812 447555 686827 447570
rect 686053 447525 686253 447555
rect 686807 447525 686827 447555
rect 686053 447514 686068 447525
rect 686053 447510 686065 447514
rect 686238 447510 686253 447525
rect 686812 447510 686827 447525
rect 686887 447566 686899 447570
rect 686887 447555 686902 447566
rect 687072 447555 687087 447570
rect 686887 447525 687087 447555
rect 686887 447514 686902 447525
rect 686887 447510 686899 447514
rect 687072 447510 687087 447525
rect 687147 447566 687159 447570
rect 687147 447555 687162 447566
rect 687332 447555 687347 447570
rect 687147 447525 687347 447555
rect 687147 447514 687162 447525
rect 687147 447510 687159 447514
rect 687332 447510 687347 447525
rect 689309 447498 689909 447626
rect 692427 447592 693027 447642
rect 693888 447575 694194 447745
rect 694388 447575 694694 447745
rect 678680 447421 678704 447455
rect 678680 447353 678704 447387
rect 682890 447357 683490 447485
rect 690910 447484 691110 447540
rect 685718 447469 685733 447484
rect 684004 447329 685004 447457
rect 685679 447439 685733 447469
rect 685718 447424 685733 447439
rect 685793 447480 685805 447484
rect 685793 447469 685808 447480
rect 685978 447469 685993 447484
rect 685793 447439 685993 447469
rect 685793 447428 685808 447439
rect 685793 447424 685805 447428
rect 685978 447424 685993 447439
rect 686053 447480 686065 447484
rect 686053 447469 686068 447480
rect 686238 447469 686253 447484
rect 686812 447469 686827 447484
rect 686053 447439 686253 447469
rect 686807 447439 686827 447469
rect 686053 447428 686068 447439
rect 686053 447424 686065 447428
rect 686238 447424 686253 447439
rect 686812 447424 686827 447439
rect 686887 447480 686899 447484
rect 686887 447469 686902 447480
rect 687072 447469 687087 447484
rect 686887 447439 687087 447469
rect 686887 447428 686902 447439
rect 686887 447424 686899 447428
rect 687072 447424 687087 447439
rect 687147 447480 687159 447484
rect 687147 447469 687162 447480
rect 687332 447469 687347 447484
rect 687147 447439 687347 447469
rect 692427 447462 693027 447512
rect 687147 447428 687162 447439
rect 687147 447424 687159 447428
rect 687332 447424 687347 447439
rect 689309 447348 689909 447398
rect 690910 447334 691110 447384
rect 678680 447285 678704 447319
rect 678680 447217 678704 447251
rect 682890 447201 683490 447329
rect 692427 447312 693027 447362
rect 678680 447149 678704 447183
rect 684004 447173 685004 447301
rect 685533 447270 685545 447274
rect 685533 447259 685548 447270
rect 685718 447259 685733 447274
rect 678680 447081 678704 447115
rect 679133 447101 679283 447113
rect 679452 447101 679602 447113
rect 678680 447013 678704 447047
rect 682890 447045 683490 447173
rect 679002 446988 679602 447038
rect 684004 447017 685004 447145
rect 685533 447079 685733 447259
rect 685533 447068 685548 447079
rect 685533 447064 685545 447068
rect 685718 447064 685733 447079
rect 685793 447270 685805 447274
rect 685793 447259 685808 447270
rect 685978 447259 685993 447274
rect 685793 447079 685993 447259
rect 685793 447068 685808 447079
rect 685793 447064 685805 447068
rect 685978 447064 685993 447079
rect 686053 447270 686065 447274
rect 686053 447259 686068 447270
rect 686238 447259 686253 447274
rect 686053 447079 686253 447259
rect 686053 447068 686068 447079
rect 686053 447064 686065 447068
rect 686238 447064 686253 447079
rect 686313 447270 686325 447274
rect 686313 447259 686328 447270
rect 686498 447259 686513 447274
rect 686313 447079 686513 447259
rect 686313 447068 686328 447079
rect 686313 447064 686325 447068
rect 686498 447064 686513 447079
rect 686627 447270 686639 447274
rect 686627 447259 686642 447270
rect 686812 447259 686827 447274
rect 686627 447079 686827 447259
rect 686627 447068 686642 447079
rect 686627 447064 686639 447068
rect 686812 447064 686827 447079
rect 686887 447270 686899 447274
rect 686887 447259 686902 447270
rect 687072 447259 687087 447274
rect 686887 447079 687087 447259
rect 686887 447068 686902 447079
rect 686887 447064 686899 447068
rect 687072 447064 687087 447079
rect 687147 447270 687159 447274
rect 687147 447259 687162 447270
rect 687332 447259 687347 447274
rect 687147 447079 687347 447259
rect 689309 447218 689909 447268
rect 692427 447140 693027 447190
rect 687147 447068 687162 447079
rect 687147 447064 687159 447068
rect 687332 447064 687347 447079
rect 689309 447068 689909 447118
rect 692427 446990 693027 447040
rect 678680 446945 678704 446979
rect 678680 446877 678704 446911
rect 682890 446895 683490 446945
rect 678680 446809 678704 446843
rect 679002 446812 679602 446868
rect 684004 446861 685004 446917
rect 685793 446910 685805 446914
rect 685793 446899 685808 446910
rect 685978 446899 685993 446914
rect 682890 446779 683490 446829
rect 678680 446741 678704 446775
rect 678680 446673 678704 446707
rect 679002 446642 679602 446692
rect 678680 446605 678704 446639
rect 682890 446623 683490 446751
rect 684004 446705 685004 446833
rect 685793 446719 685993 446899
rect 685793 446708 685808 446719
rect 685793 446704 685805 446708
rect 685978 446704 685993 446719
rect 686053 446910 686065 446914
rect 686053 446899 686068 446910
rect 686238 446899 686253 446914
rect 686607 446899 687607 446949
rect 690910 446934 691110 446984
rect 686053 446719 686253 446899
rect 692427 446860 693027 446910
rect 686607 446749 687607 446799
rect 690910 446778 691110 446834
rect 686053 446708 686068 446719
rect 686053 446704 686065 446708
rect 686238 446704 686253 446719
rect 692427 446704 693027 446832
rect 693888 446775 694194 446945
rect 694388 446775 694694 446945
rect 680502 446607 680517 446622
rect 678680 446537 678704 446571
rect 678680 446469 678704 446503
rect 678680 446401 678704 446435
rect 680480 446427 680517 446607
rect 680502 446412 680517 446427
rect 680615 446607 680630 446622
rect 680803 446618 680815 446622
rect 680800 446607 680815 446618
rect 680615 446427 680815 446607
rect 682890 446467 683490 446595
rect 684004 446549 685004 446677
rect 685793 446674 685805 446678
rect 685793 446663 685808 446674
rect 685978 446663 685993 446678
rect 680615 446412 680630 446427
rect 680800 446416 680815 446427
rect 680803 446412 680815 446416
rect 680615 446371 680630 446386
rect 680803 446382 680815 446386
rect 680800 446371 680815 446382
rect 678680 446333 678704 446367
rect 678680 446265 678704 446299
rect 678680 446197 678704 446231
rect 679007 446216 679607 446266
rect 680615 446191 680815 446371
rect 682890 446311 683490 446439
rect 684004 446393 685004 446521
rect 685793 446483 685993 446663
rect 685793 446472 685808 446483
rect 685793 446468 685805 446472
rect 685978 446468 685993 446483
rect 686053 446674 686065 446678
rect 686053 446663 686068 446674
rect 686238 446663 686253 446678
rect 686053 446483 686253 446663
rect 686607 446590 687607 446640
rect 690910 446628 691110 446678
rect 692427 446548 693027 446676
rect 686053 446472 686068 446483
rect 686053 446468 686065 446472
rect 686238 446468 686253 446483
rect 686607 446440 687607 446490
rect 692427 446392 693027 446448
rect 686829 446301 687429 446351
rect 684004 446243 685004 446293
rect 692427 446236 693027 446364
rect 695201 446282 695251 449282
rect 695351 446282 695479 449282
rect 695507 446282 695635 449282
rect 695663 446282 695791 449282
rect 695819 446282 695947 449282
rect 695975 446282 696103 449282
rect 696131 446282 696259 449282
rect 696287 446282 696337 449282
rect 696651 449239 696675 449273
rect 696651 449171 696675 449205
rect 696651 449103 696675 449137
rect 696651 449035 696675 449069
rect 696651 448967 696675 449001
rect 696651 448899 696675 448933
rect 696651 448831 696675 448865
rect 696651 448763 696675 448797
rect 696651 448695 696675 448729
rect 696651 448627 696675 448661
rect 697088 448641 697138 450041
rect 697238 448641 697366 450041
rect 697394 448641 697522 450041
rect 697550 448641 697678 450041
rect 697706 448641 697756 450041
rect 698017 450022 698053 450056
rect 698030 449988 698077 450022
rect 698017 449954 698053 449988
rect 698030 449920 698077 449954
rect 698017 449886 698053 449920
rect 698030 449852 698077 449886
rect 698017 449818 698053 449852
rect 698030 449784 698077 449818
rect 698017 449750 698053 449784
rect 698030 449716 698077 449750
rect 698017 449682 698053 449716
rect 698030 449648 698077 449682
rect 698017 449614 698053 449648
rect 698030 449580 698077 449614
rect 698017 449546 698053 449580
rect 698030 449512 698077 449546
rect 698017 449478 698053 449512
rect 698030 449444 698077 449478
rect 698017 449410 698053 449444
rect 698030 449376 698077 449410
rect 698017 449342 698053 449376
rect 698030 449308 698077 449342
rect 698017 449274 698053 449308
rect 698030 449240 698077 449274
rect 698017 449206 698053 449240
rect 698030 449172 698077 449206
rect 698017 449138 698053 449172
rect 698030 449104 698077 449138
rect 698017 449070 698053 449104
rect 698030 449036 698077 449070
rect 698017 449002 698053 449036
rect 698030 448968 698077 449002
rect 698017 448934 698053 448968
rect 698030 448900 698077 448934
rect 698017 448866 698053 448900
rect 698030 448832 698077 448866
rect 698017 448798 698053 448832
rect 698030 448764 698077 448798
rect 698017 448730 698053 448764
rect 698030 448696 698077 448730
rect 698017 448662 698053 448696
rect 698030 448628 698077 448662
rect 698017 448594 698053 448628
rect 696651 448559 696675 448593
rect 698030 448560 698077 448594
rect 698017 448526 698053 448560
rect 696651 448491 696675 448525
rect 698030 448492 698077 448526
rect 696651 448423 696675 448457
rect 698017 448428 698053 448492
rect 698030 448394 698077 448428
rect 696651 448355 696675 448389
rect 698017 448360 698053 448394
rect 698030 448326 698077 448360
rect 696651 448287 696675 448321
rect 698017 448292 698053 448326
rect 696651 448219 696675 448253
rect 696651 448151 696675 448185
rect 696651 448083 696675 448117
rect 696651 448015 696675 448049
rect 696651 447947 696675 447981
rect 696651 447879 696675 447913
rect 696651 447811 696675 447845
rect 696651 447743 696675 447777
rect 696651 447675 696675 447709
rect 696651 447607 696675 447641
rect 696651 447539 696675 447573
rect 696651 447471 696675 447505
rect 696651 447403 696675 447437
rect 696651 447335 696675 447369
rect 696651 447267 696675 447301
rect 696651 447199 696675 447233
rect 696651 447131 696675 447165
rect 696651 447063 696675 447097
rect 696651 446995 696675 447029
rect 696651 446927 696675 446961
rect 696651 446859 696675 446893
rect 697088 446879 697138 448279
rect 697238 446879 697366 448279
rect 697394 446879 697522 448279
rect 697550 446879 697678 448279
rect 697706 446879 697756 448279
rect 698030 448258 698077 448292
rect 698017 448224 698053 448258
rect 698030 448190 698077 448224
rect 698017 448156 698053 448190
rect 698030 448122 698077 448156
rect 698017 448088 698053 448122
rect 698030 448054 698077 448088
rect 698017 448020 698053 448054
rect 698030 447986 698077 448020
rect 698017 447952 698053 447986
rect 698030 447918 698077 447952
rect 698017 447884 698053 447918
rect 698030 447850 698077 447884
rect 698017 447816 698053 447850
rect 698030 447782 698077 447816
rect 698017 447748 698053 447782
rect 698030 447714 698077 447748
rect 698017 447680 698053 447714
rect 698030 447646 698077 447680
rect 698017 447612 698053 447646
rect 698030 447578 698077 447612
rect 698017 447544 698053 447578
rect 698030 447510 698077 447544
rect 698017 447476 698053 447510
rect 698030 447442 698077 447476
rect 698017 447408 698053 447442
rect 698030 447374 698077 447408
rect 698017 447340 698053 447374
rect 698030 447306 698077 447340
rect 698017 447272 698053 447306
rect 698030 447238 698077 447272
rect 698017 447204 698053 447238
rect 698030 447170 698077 447204
rect 698017 447136 698053 447170
rect 698030 447102 698077 447136
rect 698017 447068 698053 447102
rect 698030 447034 698077 447068
rect 698017 447000 698053 447034
rect 698030 446966 698077 447000
rect 698017 446932 698053 446966
rect 698030 446898 698077 446932
rect 698017 446864 698053 446898
rect 698030 446830 698077 446864
rect 696651 446791 696675 446825
rect 698017 446796 698053 446830
rect 698030 446762 698077 446796
rect 696651 446723 696675 446757
rect 696651 446655 696675 446689
rect 696651 446587 696675 446621
rect 696651 446519 696675 446553
rect 696651 446451 696675 446485
rect 696651 446383 696675 446417
rect 696651 446315 696675 446349
rect 696651 446247 696675 446281
rect 680615 446176 680630 446191
rect 680800 446180 680815 446191
rect 680803 446176 680815 446180
rect 678680 446129 678704 446163
rect 682890 446161 683490 446211
rect 684004 446127 685004 446177
rect 686829 446125 687429 446181
rect 678680 446061 678704 446095
rect 679007 446046 679607 446096
rect 692427 446080 693027 446208
rect 696651 446179 696675 446213
rect 696651 446111 696675 446145
rect 696651 446043 696675 446077
rect 678680 445993 678704 446027
rect 681664 446002 681812 446006
rect 681641 445994 681812 446002
rect 682113 445994 682313 446006
rect 684004 445971 685004 446027
rect 678680 445925 678704 445959
rect 686829 445955 687429 446005
rect 678680 445857 678704 445891
rect 680215 445870 680815 445920
rect 681713 445881 682313 445931
rect 682921 445899 683521 445949
rect 692427 445930 693027 445980
rect 696651 445975 696675 446009
rect 696651 445907 696675 445941
rect 678680 445789 678704 445823
rect 684004 445821 685004 445871
rect 678680 445721 678704 445755
rect 680215 445694 680815 445750
rect 681713 445705 682313 445761
rect 682921 445743 683521 445799
rect 685537 445749 686137 445799
rect 697088 445749 697138 446749
rect 697238 445749 697366 446749
rect 697394 445749 697522 446749
rect 697550 445749 697678 446749
rect 697706 445749 697756 446749
rect 698017 446728 698053 446762
rect 698030 446694 698077 446728
rect 698017 446660 698053 446694
rect 698030 446626 698077 446660
rect 698017 446592 698053 446626
rect 698030 446558 698077 446592
rect 698017 446524 698053 446558
rect 698030 446490 698077 446524
rect 698017 446456 698053 446490
rect 698030 446422 698077 446456
rect 698017 446388 698053 446422
rect 698030 446354 698077 446388
rect 698017 446320 698053 446354
rect 698030 446286 698077 446320
rect 698017 446252 698053 446286
rect 698030 446218 698077 446252
rect 698017 446184 698053 446218
rect 698030 446150 698077 446184
rect 698017 446116 698053 446150
rect 698030 446082 698077 446116
rect 698017 446048 698053 446082
rect 698030 446014 698077 446048
rect 698017 445980 698053 446014
rect 698030 445946 698077 445980
rect 698017 445912 698053 445946
rect 698030 445878 698077 445912
rect 698017 445844 698053 445878
rect 698030 445810 698077 445844
rect 698017 445776 698053 445810
rect 698030 445742 698077 445776
rect 698017 445708 698053 445742
rect 678680 445653 678704 445687
rect 698030 445674 698077 445708
rect 678680 445585 678704 445619
rect 680215 445518 680815 445574
rect 681713 445529 682313 445657
rect 682921 445593 683521 445643
rect 684070 445599 684670 445649
rect 685537 445593 686137 445649
rect 698017 445640 698053 445674
rect 698030 445606 698077 445640
rect 698017 445572 698053 445606
rect 698030 445538 698077 445572
rect 698017 445504 698053 445538
rect 684070 445443 684670 445499
rect 685537 445443 686137 445493
rect 692428 445442 693028 445492
rect 698030 445470 698077 445504
rect 698017 445436 698053 445470
rect 680215 445348 680815 445398
rect 681713 445359 682313 445409
rect 698030 445402 698077 445436
rect 698017 445368 698053 445402
rect 684070 445293 684670 445343
rect 692428 445292 693028 445342
rect 698030 445334 698077 445368
rect 698017 445300 698053 445334
rect 680215 445232 680815 445282
rect 698030 445266 698077 445300
rect 698017 445232 698053 445266
rect 692428 445162 693028 445212
rect 698030 445198 698077 445232
rect 698017 445164 698053 445198
rect 680215 445056 680815 445112
rect 692428 445006 693028 445134
rect 698030 445130 698077 445164
rect 698017 445096 698053 445130
rect 698030 445062 698077 445096
rect 698017 444983 698053 445062
rect 698084 444983 698120 451933
rect 699322 451908 700322 451964
rect 700922 451908 701922 451964
rect 707610 451953 708610 452009
rect 709211 451953 710211 452009
rect 699322 451836 700322 451892
rect 700922 451836 701922 451892
rect 707610 451881 708610 451937
rect 709211 451881 710211 451937
rect 699322 451534 700322 451606
rect 700922 451534 701922 451606
rect 707610 451579 708610 451651
rect 709211 451579 710211 451651
rect 699392 451523 699426 451534
rect 699460 451523 699494 451534
rect 699528 451523 699562 451534
rect 699596 451523 699630 451534
rect 699664 451523 699698 451534
rect 699732 451523 699766 451534
rect 699800 451523 699834 451534
rect 699868 451523 699902 451534
rect 699936 451523 699970 451534
rect 700004 451523 700038 451534
rect 700072 451523 700106 451534
rect 700140 451523 700174 451534
rect 700208 451523 700242 451534
rect 700276 451523 700310 451534
rect 700934 451523 700968 451534
rect 701002 451523 701036 451534
rect 701070 451523 701104 451534
rect 701138 451523 701172 451534
rect 701206 451523 701240 451534
rect 701274 451523 701308 451534
rect 701342 451523 701376 451534
rect 701410 451523 701444 451534
rect 701478 451523 701512 451534
rect 701546 451523 701580 451534
rect 701614 451523 701648 451534
rect 701682 451523 701716 451534
rect 701750 451523 701784 451534
rect 701818 451523 701852 451534
rect 699392 451513 699450 451523
rect 699460 451513 699518 451523
rect 699528 451513 699586 451523
rect 699596 451513 699654 451523
rect 699664 451513 699722 451523
rect 699732 451513 699790 451523
rect 699800 451513 699858 451523
rect 699868 451513 699926 451523
rect 699936 451513 699994 451523
rect 700004 451513 700062 451523
rect 700072 451513 700130 451523
rect 700140 451513 700198 451523
rect 700208 451513 700266 451523
rect 700276 451513 700334 451523
rect 700934 451513 700992 451523
rect 701002 451513 701060 451523
rect 701070 451513 701128 451523
rect 701138 451513 701196 451523
rect 701206 451513 701264 451523
rect 701274 451513 701332 451523
rect 701342 451513 701400 451523
rect 701410 451513 701468 451523
rect 701478 451513 701536 451523
rect 701546 451513 701604 451523
rect 701614 451513 701672 451523
rect 701682 451513 701740 451523
rect 701750 451513 701808 451523
rect 701818 451513 701876 451523
rect 699368 451489 700334 451513
rect 700910 451489 701876 451513
rect 699392 451474 699416 451489
rect 699460 451474 699484 451489
rect 699528 451474 699552 451489
rect 699596 451474 699620 451489
rect 699664 451474 699688 451489
rect 699732 451474 699756 451489
rect 699800 451474 699824 451489
rect 699868 451474 699892 451489
rect 699936 451474 699960 451489
rect 700004 451474 700028 451489
rect 700072 451474 700096 451489
rect 700140 451474 700164 451489
rect 700208 451474 700232 451489
rect 700276 451474 700300 451489
rect 700934 451474 700958 451489
rect 701002 451474 701026 451489
rect 701070 451474 701094 451489
rect 701138 451474 701162 451489
rect 701206 451474 701230 451489
rect 701274 451474 701298 451489
rect 701342 451474 701366 451489
rect 701410 451474 701434 451489
rect 701478 451474 701502 451489
rect 701546 451474 701570 451489
rect 701614 451474 701638 451489
rect 701682 451474 701706 451489
rect 701750 451474 701774 451489
rect 701818 451474 701842 451489
rect 699322 451319 700322 451474
rect 699322 451285 700334 451319
rect 700922 451309 701922 451474
rect 707610 451319 708610 451379
rect 709211 451319 710211 451379
rect 700910 451285 701922 451309
rect 699322 451274 700322 451285
rect 700922 451274 701922 451285
rect 699392 451261 699416 451274
rect 699460 451261 699484 451274
rect 699528 451261 699552 451274
rect 699596 451261 699620 451274
rect 699664 451261 699688 451274
rect 699732 451261 699756 451274
rect 699800 451261 699824 451274
rect 699868 451261 699892 451274
rect 699936 451261 699960 451274
rect 700004 451261 700028 451274
rect 700072 451261 700096 451274
rect 700140 451261 700164 451274
rect 700208 451261 700232 451274
rect 700276 451261 700300 451274
rect 700934 451261 700958 451274
rect 701002 451261 701026 451274
rect 701070 451261 701094 451274
rect 701138 451261 701162 451274
rect 701206 451261 701230 451274
rect 701274 451261 701298 451274
rect 701342 451261 701366 451274
rect 701410 451261 701434 451274
rect 701478 451261 701502 451274
rect 701546 451261 701570 451274
rect 701614 451261 701638 451274
rect 701682 451261 701706 451274
rect 701750 451261 701774 451274
rect 701818 451261 701842 451274
rect 699322 450916 700322 450972
rect 700922 450916 701922 450972
rect 707610 450961 708610 451017
rect 709211 450961 710211 451017
rect 699322 450844 700322 450900
rect 700922 450844 701922 450900
rect 707610 450889 708610 450945
rect 709211 450889 710211 450945
rect 699322 450542 700322 450614
rect 700922 450542 701922 450614
rect 707610 450587 708610 450659
rect 709211 450587 710211 450659
rect 699392 450531 699426 450542
rect 699460 450531 699494 450542
rect 699528 450531 699562 450542
rect 699596 450531 699630 450542
rect 699664 450531 699698 450542
rect 699732 450531 699766 450542
rect 699800 450531 699834 450542
rect 699868 450531 699902 450542
rect 699936 450531 699970 450542
rect 700004 450531 700038 450542
rect 700072 450531 700106 450542
rect 700140 450531 700174 450542
rect 700208 450531 700242 450542
rect 700276 450531 700310 450542
rect 700934 450531 700968 450542
rect 701002 450531 701036 450542
rect 701070 450531 701104 450542
rect 701138 450531 701172 450542
rect 701206 450531 701240 450542
rect 701274 450531 701308 450542
rect 701342 450531 701376 450542
rect 701410 450531 701444 450542
rect 701478 450531 701512 450542
rect 701546 450531 701580 450542
rect 701614 450531 701648 450542
rect 701682 450531 701716 450542
rect 701750 450531 701784 450542
rect 701818 450531 701852 450542
rect 699392 450521 699450 450531
rect 699460 450521 699518 450531
rect 699528 450521 699586 450531
rect 699596 450521 699654 450531
rect 699664 450521 699722 450531
rect 699732 450521 699790 450531
rect 699800 450521 699858 450531
rect 699868 450521 699926 450531
rect 699936 450521 699994 450531
rect 700004 450521 700062 450531
rect 700072 450521 700130 450531
rect 700140 450521 700198 450531
rect 700208 450521 700266 450531
rect 700276 450521 700334 450531
rect 700934 450521 700992 450531
rect 701002 450521 701060 450531
rect 701070 450521 701128 450531
rect 701138 450521 701196 450531
rect 701206 450521 701264 450531
rect 701274 450521 701332 450531
rect 701342 450521 701400 450531
rect 701410 450521 701468 450531
rect 701478 450521 701536 450531
rect 701546 450521 701604 450531
rect 701614 450521 701672 450531
rect 701682 450521 701740 450531
rect 701750 450521 701808 450531
rect 701818 450521 701876 450531
rect 699368 450497 700334 450521
rect 700910 450497 701876 450521
rect 699392 450482 699416 450497
rect 699460 450482 699484 450497
rect 699528 450482 699552 450497
rect 699596 450482 699620 450497
rect 699664 450482 699688 450497
rect 699732 450482 699756 450497
rect 699800 450482 699824 450497
rect 699868 450482 699892 450497
rect 699936 450482 699960 450497
rect 700004 450482 700028 450497
rect 700072 450482 700096 450497
rect 700140 450482 700164 450497
rect 700208 450482 700232 450497
rect 700276 450482 700300 450497
rect 700934 450482 700958 450497
rect 701002 450482 701026 450497
rect 701070 450482 701094 450497
rect 701138 450482 701162 450497
rect 701206 450482 701230 450497
rect 701274 450482 701298 450497
rect 701342 450482 701366 450497
rect 701410 450482 701434 450497
rect 701478 450482 701502 450497
rect 701546 450482 701570 450497
rect 701614 450482 701638 450497
rect 701682 450482 701706 450497
rect 701750 450482 701774 450497
rect 701818 450482 701842 450497
rect 699322 450327 700322 450482
rect 699322 450293 700334 450327
rect 700922 450317 701922 450482
rect 707610 450327 708610 450387
rect 709211 450327 710211 450387
rect 711541 450345 711629 457461
rect 711892 456200 711942 457200
rect 712062 456200 712112 457200
rect 711892 455079 711942 456079
rect 712062 455079 712112 456079
rect 711892 453958 711942 454958
rect 712062 453958 712112 454958
rect 711892 452848 711942 453848
rect 712062 452848 712112 453848
rect 711892 451727 711942 452727
rect 712062 451727 712112 452727
rect 711892 450606 711942 451606
rect 712062 450606 712112 451606
rect 712409 450371 712431 457485
rect 712469 457459 712487 457501
rect 712499 457459 712505 457467
rect 712499 457455 712511 457459
rect 712539 457455 712557 457501
rect 713640 455461 713674 457785
rect 713750 457772 714750 457822
rect 717367 457820 717413 457853
rect 717367 457819 717379 457820
rect 717401 457819 717413 457820
rect 717401 457809 717600 457819
rect 717401 457786 717413 457809
rect 713750 457562 714750 457612
rect 713750 457446 714750 457496
rect 713750 457230 714750 457358
rect 713750 457014 714750 457070
rect 713750 456798 714750 456926
rect 713750 456588 714750 456638
rect 714478 456585 714750 456588
rect 715486 455931 715536 456931
rect 715696 455931 715824 456931
rect 715912 455931 715962 456931
rect 713641 455345 713663 455461
rect 713640 455309 713674 455345
rect 713750 455314 714750 455364
rect 713750 455158 714750 455214
rect 713750 455002 714750 455130
rect 713750 454846 714750 454974
rect 713750 454690 714750 454746
rect 716425 454709 716725 454721
rect 713750 454534 714750 454662
rect 716425 454596 717425 454646
rect 713750 454378 714750 454506
rect 716425 454440 717425 454568
rect 713750 454222 714750 454350
rect 716425 454284 717425 454340
rect 713750 454072 714750 454122
rect 713750 453956 714750 454006
rect 713750 453800 714750 453928
rect 713750 453644 714750 453772
rect 713750 453488 714750 453616
rect 715354 453587 715404 454187
rect 715504 453587 715560 454187
rect 715660 453587 715716 454187
rect 715816 453587 715872 454187
rect 715972 453587 716022 454187
rect 716425 454128 717425 454256
rect 716425 453978 717425 454028
rect 716425 453862 717425 453912
rect 716425 453706 717425 453834
rect 716425 453550 717425 453606
rect 716425 453394 717425 453522
rect 713750 453332 714750 453388
rect 713750 453176 714750 453304
rect 716425 453244 717425 453294
rect 713750 453020 714750 453148
rect 713750 452870 714750 452920
rect 713750 452742 714750 452792
rect 713750 452586 714750 452642
rect 713750 452436 714750 452486
rect 713750 452320 714350 452370
rect 713750 452164 714350 452292
rect 715510 452191 715560 453191
rect 715660 452191 715788 453191
rect 715816 452191 715944 453191
rect 715972 452191 716022 453191
rect 716425 453128 717425 453178
rect 716425 452972 717425 453028
rect 716425 452822 717425 452872
rect 716425 452706 717425 452756
rect 716425 452550 717425 452678
rect 716425 452394 717425 452522
rect 716425 452238 717425 452366
rect 716425 452082 717425 452210
rect 713750 452008 714350 452064
rect 713750 451852 714350 451980
rect 716425 451932 717425 451982
rect 713750 451696 714350 451752
rect 713750 451446 714350 451496
rect 714565 451443 714765 451455
rect 713750 451330 714750 451380
rect 713750 451120 714750 451170
rect 716413 451092 716447 451150
rect 713750 451004 714750 451054
rect 713750 450794 714750 450844
rect 713750 450678 714750 450728
rect 713750 450468 714750 450518
rect 713750 450352 714750 450402
rect 700910 450293 701922 450317
rect 699322 450282 700322 450293
rect 700922 450282 701922 450293
rect 711541 450311 711633 450345
rect 699392 450269 699416 450282
rect 699460 450269 699484 450282
rect 699528 450269 699552 450282
rect 699596 450269 699620 450282
rect 699664 450269 699688 450282
rect 699732 450269 699756 450282
rect 699800 450269 699824 450282
rect 699868 450269 699892 450282
rect 699936 450269 699960 450282
rect 700004 450269 700028 450282
rect 700072 450269 700096 450282
rect 700140 450269 700164 450282
rect 700208 450269 700232 450282
rect 700276 450269 700300 450282
rect 700934 450269 700958 450282
rect 701002 450269 701026 450282
rect 701070 450269 701094 450282
rect 701138 450269 701162 450282
rect 701206 450269 701230 450282
rect 701274 450269 701298 450282
rect 701342 450269 701366 450282
rect 701410 450269 701434 450282
rect 701478 450269 701502 450282
rect 701546 450269 701570 450282
rect 701614 450269 701638 450282
rect 701682 450269 701706 450282
rect 701750 450269 701774 450282
rect 701818 450269 701842 450282
rect 699322 449924 700322 449980
rect 700922 449924 701922 449980
rect 707610 449969 708610 450025
rect 709211 449969 710211 450025
rect 699322 449852 700322 449908
rect 700922 449852 701922 449908
rect 707610 449897 708610 449953
rect 709211 449897 710211 449953
rect 699322 449550 700322 449622
rect 700922 449550 701922 449622
rect 707610 449595 708610 449667
rect 709211 449595 710211 449667
rect 699392 449539 699426 449550
rect 699460 449539 699494 449550
rect 699528 449539 699562 449550
rect 699596 449539 699630 449550
rect 699664 449539 699698 449550
rect 699732 449539 699766 449550
rect 699800 449539 699834 449550
rect 699868 449539 699902 449550
rect 699936 449539 699970 449550
rect 700004 449539 700038 449550
rect 700072 449539 700106 449550
rect 700140 449539 700174 449550
rect 700208 449539 700242 449550
rect 700276 449539 700310 449550
rect 700934 449539 700968 449550
rect 701002 449539 701036 449550
rect 701070 449539 701104 449550
rect 701138 449539 701172 449550
rect 701206 449539 701240 449550
rect 701274 449539 701308 449550
rect 701342 449539 701376 449550
rect 701410 449539 701444 449550
rect 701478 449539 701512 449550
rect 701546 449539 701580 449550
rect 701614 449539 701648 449550
rect 701682 449539 701716 449550
rect 701750 449539 701784 449550
rect 701818 449539 701852 449550
rect 699392 449529 699450 449539
rect 699460 449529 699518 449539
rect 699528 449529 699586 449539
rect 699596 449529 699654 449539
rect 699664 449529 699722 449539
rect 699732 449529 699790 449539
rect 699800 449529 699858 449539
rect 699868 449529 699926 449539
rect 699936 449529 699994 449539
rect 700004 449529 700062 449539
rect 700072 449529 700130 449539
rect 700140 449529 700198 449539
rect 700208 449529 700266 449539
rect 700276 449529 700334 449539
rect 700934 449529 700992 449539
rect 701002 449529 701060 449539
rect 701070 449529 701128 449539
rect 701138 449529 701196 449539
rect 701206 449529 701264 449539
rect 701274 449529 701332 449539
rect 701342 449529 701400 449539
rect 701410 449529 701468 449539
rect 701478 449529 701536 449539
rect 701546 449529 701604 449539
rect 701614 449529 701672 449539
rect 701682 449529 701740 449539
rect 701750 449529 701808 449539
rect 701818 449529 701876 449539
rect 699368 449505 700334 449529
rect 700910 449505 701876 449529
rect 699392 449490 699416 449505
rect 699460 449490 699484 449505
rect 699528 449490 699552 449505
rect 699596 449490 699620 449505
rect 699664 449490 699688 449505
rect 699732 449490 699756 449505
rect 699800 449490 699824 449505
rect 699868 449490 699892 449505
rect 699936 449490 699960 449505
rect 700004 449490 700028 449505
rect 700072 449490 700096 449505
rect 700140 449490 700164 449505
rect 700208 449490 700232 449505
rect 700276 449490 700300 449505
rect 700934 449490 700958 449505
rect 701002 449490 701026 449505
rect 701070 449490 701094 449505
rect 701138 449490 701162 449505
rect 701206 449490 701230 449505
rect 701274 449490 701298 449505
rect 701342 449490 701366 449505
rect 701410 449490 701434 449505
rect 701478 449490 701502 449505
rect 701546 449490 701570 449505
rect 701614 449490 701638 449505
rect 701682 449490 701706 449505
rect 701750 449490 701774 449505
rect 701818 449490 701842 449505
rect 699322 449335 700322 449490
rect 699322 449301 700334 449335
rect 700922 449325 701922 449490
rect 707610 449335 708610 449395
rect 709211 449335 710211 449395
rect 700910 449301 701922 449325
rect 699322 449290 700322 449301
rect 700922 449290 701922 449301
rect 699392 449277 699416 449290
rect 699460 449277 699484 449290
rect 699528 449277 699552 449290
rect 699596 449277 699620 449290
rect 699664 449277 699688 449290
rect 699732 449277 699756 449290
rect 699800 449277 699824 449290
rect 699868 449277 699892 449290
rect 699936 449277 699960 449290
rect 700004 449277 700028 449290
rect 700072 449277 700096 449290
rect 700140 449277 700164 449290
rect 700208 449277 700232 449290
rect 700276 449277 700300 449290
rect 700934 449277 700958 449290
rect 701002 449277 701026 449290
rect 701070 449277 701094 449290
rect 701138 449277 701162 449290
rect 701206 449277 701230 449290
rect 701274 449277 701298 449290
rect 701342 449277 701366 449290
rect 701410 449277 701434 449290
rect 701478 449277 701502 449290
rect 701546 449277 701570 449290
rect 701614 449277 701638 449290
rect 701682 449277 701706 449290
rect 701750 449277 701774 449290
rect 701818 449277 701842 449290
rect 699322 448932 700322 448988
rect 700922 448932 701922 448988
rect 707610 448977 708610 449033
rect 709211 448977 710211 449033
rect 699322 448860 700322 448916
rect 700922 448860 701922 448916
rect 707610 448905 708610 448961
rect 709211 448905 710211 448961
rect 699322 448558 700322 448630
rect 700922 448558 701922 448630
rect 707610 448603 708610 448675
rect 709211 448603 710211 448675
rect 699392 448547 699426 448558
rect 699460 448547 699494 448558
rect 699528 448547 699562 448558
rect 699596 448547 699630 448558
rect 699664 448547 699698 448558
rect 699732 448547 699766 448558
rect 699800 448547 699834 448558
rect 699868 448547 699902 448558
rect 699936 448547 699970 448558
rect 700004 448547 700038 448558
rect 700072 448547 700106 448558
rect 700140 448547 700174 448558
rect 700208 448547 700242 448558
rect 700276 448547 700310 448558
rect 700934 448547 700968 448558
rect 701002 448547 701036 448558
rect 701070 448547 701104 448558
rect 701138 448547 701172 448558
rect 701206 448547 701240 448558
rect 701274 448547 701308 448558
rect 701342 448547 701376 448558
rect 701410 448547 701444 448558
rect 701478 448547 701512 448558
rect 701546 448547 701580 448558
rect 701614 448547 701648 448558
rect 701682 448547 701716 448558
rect 701750 448547 701784 448558
rect 701818 448547 701852 448558
rect 699392 448537 699450 448547
rect 699460 448537 699518 448547
rect 699528 448537 699586 448547
rect 699596 448537 699654 448547
rect 699664 448537 699722 448547
rect 699732 448537 699790 448547
rect 699800 448537 699858 448547
rect 699868 448537 699926 448547
rect 699936 448537 699994 448547
rect 700004 448537 700062 448547
rect 700072 448537 700130 448547
rect 700140 448537 700198 448547
rect 700208 448537 700266 448547
rect 700276 448537 700334 448547
rect 700934 448537 700992 448547
rect 701002 448537 701060 448547
rect 701070 448537 701128 448547
rect 701138 448537 701196 448547
rect 701206 448537 701264 448547
rect 701274 448537 701332 448547
rect 701342 448537 701400 448547
rect 701410 448537 701468 448547
rect 701478 448537 701536 448547
rect 701546 448537 701604 448547
rect 701614 448537 701672 448547
rect 701682 448537 701740 448547
rect 701750 448537 701808 448547
rect 701818 448537 701876 448547
rect 699368 448513 700334 448537
rect 700910 448513 701876 448537
rect 699392 448498 699416 448513
rect 699460 448498 699484 448513
rect 699528 448498 699552 448513
rect 699596 448498 699620 448513
rect 699664 448498 699688 448513
rect 699732 448498 699756 448513
rect 699800 448498 699824 448513
rect 699868 448498 699892 448513
rect 699936 448498 699960 448513
rect 700004 448498 700028 448513
rect 700072 448498 700096 448513
rect 700140 448498 700164 448513
rect 700208 448498 700232 448513
rect 700276 448498 700300 448513
rect 700934 448498 700958 448513
rect 701002 448498 701026 448513
rect 701070 448498 701094 448513
rect 701138 448498 701162 448513
rect 701206 448498 701230 448513
rect 701274 448498 701298 448513
rect 701342 448498 701366 448513
rect 701410 448498 701434 448513
rect 701478 448498 701502 448513
rect 701546 448498 701570 448513
rect 701614 448498 701638 448513
rect 701682 448498 701706 448513
rect 701750 448498 701774 448513
rect 701818 448498 701842 448513
rect 699322 448343 700322 448498
rect 699322 448309 700334 448343
rect 700922 448333 701922 448498
rect 707610 448343 708610 448403
rect 709211 448343 710211 448403
rect 700910 448309 701922 448333
rect 699322 448298 700322 448309
rect 700922 448298 701922 448309
rect 699392 448285 699416 448298
rect 699460 448285 699484 448298
rect 699528 448285 699552 448298
rect 699596 448285 699620 448298
rect 699664 448285 699688 448298
rect 699732 448285 699756 448298
rect 699800 448285 699824 448298
rect 699868 448285 699892 448298
rect 699936 448285 699960 448298
rect 700004 448285 700028 448298
rect 700072 448285 700096 448298
rect 700140 448285 700164 448298
rect 700208 448285 700232 448298
rect 700276 448285 700300 448298
rect 700934 448285 700958 448298
rect 701002 448285 701026 448298
rect 701070 448285 701094 448298
rect 701138 448285 701162 448298
rect 701206 448285 701230 448298
rect 701274 448285 701298 448298
rect 701342 448285 701366 448298
rect 701410 448285 701434 448298
rect 701478 448285 701502 448298
rect 701546 448285 701570 448298
rect 701614 448285 701638 448298
rect 701682 448285 701706 448298
rect 701750 448285 701774 448298
rect 701818 448285 701842 448298
rect 699322 447940 700322 447996
rect 700922 447940 701922 447996
rect 707610 447985 708610 448041
rect 709211 447985 710211 448041
rect 699322 447868 700322 447924
rect 700922 447868 701922 447924
rect 707610 447913 708610 447969
rect 709211 447913 710211 447969
rect 699322 447566 700322 447638
rect 700922 447566 701922 447638
rect 707610 447611 708610 447683
rect 709211 447611 710211 447683
rect 699392 447555 699426 447566
rect 699460 447555 699494 447566
rect 699528 447555 699562 447566
rect 699596 447555 699630 447566
rect 699664 447555 699698 447566
rect 699732 447555 699766 447566
rect 699800 447555 699834 447566
rect 699868 447555 699902 447566
rect 699936 447555 699970 447566
rect 700004 447555 700038 447566
rect 700072 447555 700106 447566
rect 700140 447555 700174 447566
rect 700208 447555 700242 447566
rect 700276 447555 700310 447566
rect 700934 447555 700968 447566
rect 701002 447555 701036 447566
rect 701070 447555 701104 447566
rect 701138 447555 701172 447566
rect 701206 447555 701240 447566
rect 701274 447555 701308 447566
rect 701342 447555 701376 447566
rect 701410 447555 701444 447566
rect 701478 447555 701512 447566
rect 701546 447555 701580 447566
rect 701614 447555 701648 447566
rect 701682 447555 701716 447566
rect 701750 447555 701784 447566
rect 701818 447555 701852 447566
rect 699392 447545 699450 447555
rect 699460 447545 699518 447555
rect 699528 447545 699586 447555
rect 699596 447545 699654 447555
rect 699664 447545 699722 447555
rect 699732 447545 699790 447555
rect 699800 447545 699858 447555
rect 699868 447545 699926 447555
rect 699936 447545 699994 447555
rect 700004 447545 700062 447555
rect 700072 447545 700130 447555
rect 700140 447545 700198 447555
rect 700208 447545 700266 447555
rect 700276 447545 700334 447555
rect 700934 447545 700992 447555
rect 701002 447545 701060 447555
rect 701070 447545 701128 447555
rect 701138 447545 701196 447555
rect 701206 447545 701264 447555
rect 701274 447545 701332 447555
rect 701342 447545 701400 447555
rect 701410 447545 701468 447555
rect 701478 447545 701536 447555
rect 701546 447545 701604 447555
rect 701614 447545 701672 447555
rect 701682 447545 701740 447555
rect 701750 447545 701808 447555
rect 701818 447545 701876 447555
rect 699368 447521 700334 447545
rect 700910 447521 701876 447545
rect 699392 447506 699416 447521
rect 699460 447506 699484 447521
rect 699528 447506 699552 447521
rect 699596 447506 699620 447521
rect 699664 447506 699688 447521
rect 699732 447506 699756 447521
rect 699800 447506 699824 447521
rect 699868 447506 699892 447521
rect 699936 447506 699960 447521
rect 700004 447506 700028 447521
rect 700072 447506 700096 447521
rect 700140 447506 700164 447521
rect 700208 447506 700232 447521
rect 700276 447506 700300 447521
rect 700934 447506 700958 447521
rect 701002 447506 701026 447521
rect 701070 447506 701094 447521
rect 701138 447506 701162 447521
rect 701206 447506 701230 447521
rect 701274 447506 701298 447521
rect 701342 447506 701366 447521
rect 701410 447506 701434 447521
rect 701478 447506 701502 447521
rect 701546 447506 701570 447521
rect 701614 447506 701638 447521
rect 701682 447506 701706 447521
rect 701750 447506 701774 447521
rect 701818 447506 701842 447521
rect 699322 447351 700322 447506
rect 699322 447317 700334 447351
rect 700922 447341 701922 447506
rect 705107 447360 705173 447376
rect 707610 447351 708610 447411
rect 709211 447351 710211 447411
rect 700910 447317 701922 447341
rect 699322 447306 700322 447317
rect 700922 447306 701922 447317
rect 699392 447293 699416 447306
rect 699460 447293 699484 447306
rect 699528 447293 699552 447306
rect 699596 447293 699620 447306
rect 699664 447293 699688 447306
rect 699732 447293 699756 447306
rect 699800 447293 699824 447306
rect 699868 447293 699892 447306
rect 699936 447293 699960 447306
rect 700004 447293 700028 447306
rect 700072 447293 700096 447306
rect 700140 447293 700164 447306
rect 700208 447293 700232 447306
rect 700276 447293 700300 447306
rect 700934 447293 700958 447306
rect 701002 447293 701026 447306
rect 701070 447293 701094 447306
rect 701138 447293 701162 447306
rect 701206 447293 701230 447306
rect 701274 447293 701298 447306
rect 701342 447293 701366 447306
rect 701410 447293 701434 447306
rect 701478 447293 701502 447306
rect 701546 447293 701570 447306
rect 701614 447293 701638 447306
rect 701682 447293 701706 447306
rect 701750 447293 701774 447306
rect 701818 447293 701842 447306
rect 699322 446948 700322 447004
rect 700922 446948 701922 447004
rect 707610 446993 708610 447049
rect 709211 446993 710211 447049
rect 699322 446876 700322 446932
rect 700922 446876 701922 446932
rect 707610 446921 708610 446977
rect 709211 446921 710211 446977
rect 699322 446574 700322 446646
rect 700922 446574 701922 446646
rect 707610 446619 708610 446691
rect 709211 446619 710211 446691
rect 699392 446563 699426 446574
rect 699460 446563 699494 446574
rect 699528 446563 699562 446574
rect 699596 446563 699630 446574
rect 699664 446563 699698 446574
rect 699732 446563 699766 446574
rect 699800 446563 699834 446574
rect 699868 446563 699902 446574
rect 699936 446563 699970 446574
rect 700004 446563 700038 446574
rect 700072 446563 700106 446574
rect 700140 446563 700174 446574
rect 700208 446563 700242 446574
rect 700276 446563 700310 446574
rect 700934 446563 700968 446574
rect 701002 446563 701036 446574
rect 701070 446563 701104 446574
rect 701138 446563 701172 446574
rect 701206 446563 701240 446574
rect 701274 446563 701308 446574
rect 701342 446563 701376 446574
rect 701410 446563 701444 446574
rect 701478 446563 701512 446574
rect 701546 446563 701580 446574
rect 701614 446563 701648 446574
rect 701682 446563 701716 446574
rect 701750 446563 701784 446574
rect 701818 446563 701852 446574
rect 699392 446553 699450 446563
rect 699460 446553 699518 446563
rect 699528 446553 699586 446563
rect 699596 446553 699654 446563
rect 699664 446553 699722 446563
rect 699732 446553 699790 446563
rect 699800 446553 699858 446563
rect 699868 446553 699926 446563
rect 699936 446553 699994 446563
rect 700004 446553 700062 446563
rect 700072 446553 700130 446563
rect 700140 446553 700198 446563
rect 700208 446553 700266 446563
rect 700276 446553 700334 446563
rect 700934 446553 700992 446563
rect 701002 446553 701060 446563
rect 701070 446553 701128 446563
rect 701138 446553 701196 446563
rect 701206 446553 701264 446563
rect 701274 446553 701332 446563
rect 701342 446553 701400 446563
rect 701410 446553 701468 446563
rect 701478 446553 701536 446563
rect 701546 446553 701604 446563
rect 701614 446553 701672 446563
rect 701682 446553 701740 446563
rect 701750 446553 701808 446563
rect 701818 446553 701876 446563
rect 699368 446529 700334 446553
rect 700910 446529 701876 446553
rect 699392 446514 699416 446529
rect 699460 446514 699484 446529
rect 699528 446514 699552 446529
rect 699596 446514 699620 446529
rect 699664 446514 699688 446529
rect 699732 446514 699756 446529
rect 699800 446514 699824 446529
rect 699868 446514 699892 446529
rect 699936 446514 699960 446529
rect 700004 446514 700028 446529
rect 700072 446514 700096 446529
rect 700140 446514 700164 446529
rect 700208 446514 700232 446529
rect 700276 446514 700300 446529
rect 700934 446514 700958 446529
rect 701002 446514 701026 446529
rect 701070 446514 701094 446529
rect 701138 446514 701162 446529
rect 701206 446514 701230 446529
rect 701274 446514 701298 446529
rect 701342 446514 701366 446529
rect 701410 446514 701434 446529
rect 701478 446514 701502 446529
rect 701546 446514 701570 446529
rect 701614 446514 701638 446529
rect 701682 446514 701706 446529
rect 701750 446514 701774 446529
rect 701818 446514 701842 446529
rect 699322 446359 700322 446514
rect 699322 446325 700334 446359
rect 700922 446349 701922 446514
rect 707610 446359 708610 446419
rect 709211 446359 710211 446419
rect 700910 446325 701922 446349
rect 699322 446314 700322 446325
rect 700922 446314 701922 446325
rect 699392 446301 699416 446314
rect 699460 446301 699484 446314
rect 699528 446301 699552 446314
rect 699596 446301 699620 446314
rect 699664 446301 699688 446314
rect 699732 446301 699756 446314
rect 699800 446301 699824 446314
rect 699868 446301 699892 446314
rect 699936 446301 699960 446314
rect 700004 446301 700028 446314
rect 700072 446301 700096 446314
rect 700140 446301 700164 446314
rect 700208 446301 700232 446314
rect 700276 446301 700300 446314
rect 700934 446301 700958 446314
rect 701002 446301 701026 446314
rect 701070 446301 701094 446314
rect 701138 446301 701162 446314
rect 701206 446301 701230 446314
rect 701274 446301 701298 446314
rect 701342 446301 701366 446314
rect 701410 446301 701434 446314
rect 701478 446301 701502 446314
rect 701546 446301 701570 446314
rect 701614 446301 701638 446314
rect 701682 446301 701706 446314
rect 701750 446301 701774 446314
rect 701818 446301 701842 446314
rect 709211 446148 710211 446152
rect 707574 446099 707610 446134
rect 708610 446099 708646 446134
rect 707574 446098 708646 446099
rect 707574 446057 707610 446098
rect 708610 446057 708646 446098
rect 699322 445956 700322 446012
rect 700922 445956 701922 446012
rect 707574 446001 708646 446057
rect 707574 445964 707610 446001
rect 708610 445964 708646 446001
rect 707574 445959 708646 445964
rect 699322 445884 700322 445940
rect 700922 445884 701922 445940
rect 707574 445924 707610 445959
rect 708610 445924 708646 445959
rect 709175 446098 710247 446134
rect 709175 446057 709211 446098
rect 710211 446057 710247 446098
rect 709175 446001 710247 446057
rect 709175 445964 709211 446001
rect 710211 445964 710247 446001
rect 709175 445936 710247 445964
rect 709175 445924 709211 445936
rect 710211 445924 710247 445936
rect 707610 445713 708610 445785
rect 709211 445713 710211 445785
rect 699322 445623 700322 445673
rect 700922 445623 701922 445673
rect 707610 445523 708610 445617
rect 707610 445513 708644 445523
rect 709211 445513 710211 445591
rect 711541 445437 711629 450311
rect 713750 450136 714750 450264
rect 716417 450152 717417 450202
rect 711892 449049 711942 450049
rect 712062 449049 712112 450049
rect 713750 449920 714750 450048
rect 716417 449996 717417 450052
rect 716417 449846 717417 449896
rect 713750 449704 714750 449832
rect 716417 449730 717017 449780
rect 716417 449580 717017 449630
rect 713750 449488 714750 449544
rect 716417 449464 717417 449514
rect 713750 449272 714750 449400
rect 716417 449308 717417 449364
rect 713750 449056 714750 449184
rect 716417 449152 717417 449280
rect 716417 448996 717417 449052
rect 711892 447928 711942 448928
rect 712062 447928 712112 448928
rect 713750 448840 714750 448968
rect 716417 448840 717417 448968
rect 713750 448624 714750 448752
rect 716417 448684 717417 448740
rect 716417 448474 717417 448524
rect 713750 448408 714750 448464
rect 716417 448308 717417 448358
rect 713750 448192 714750 448248
rect 716417 448152 717417 448280
rect 713750 447976 714750 448104
rect 716417 447996 717417 448052
rect 711892 446807 711942 447807
rect 712062 446807 712112 447807
rect 713750 447760 714750 447888
rect 716417 447780 717417 447836
rect 713750 447544 714750 447672
rect 716417 447570 717417 447620
rect 713750 447328 714750 447456
rect 716417 447454 717417 447504
rect 716417 447298 717417 447426
rect 713750 447118 714750 447168
rect 716417 447148 717417 447198
rect 711892 445697 711942 446697
rect 712062 445697 712112 446697
rect 714686 446357 714794 446424
rect 714645 446323 714794 446357
rect 716071 446357 716074 446358
rect 716071 446356 716072 446357
rect 716073 446356 716074 446357
rect 716071 446355 716074 446356
rect 716208 446357 716211 446358
rect 716208 446356 716209 446357
rect 716210 446356 716211 446357
rect 716208 446355 716211 446356
rect 714964 446247 715998 446329
rect 716284 446247 717318 446329
rect 705107 445336 705173 445352
rect 711541 445302 711633 445437
rect 714175 445398 714225 445998
rect 714425 445398 714475 445998
rect 711579 445301 711595 445302
rect 714781 445191 714863 446226
rect 715134 445955 715828 446037
rect 714686 445123 714863 445191
rect 714645 445089 714863 445123
rect 680215 444880 680815 444936
rect 686719 444893 686739 444917
rect 686743 444893 686753 444917
rect 686719 444859 686757 444893
rect 686719 444822 686739 444859
rect 686743 444822 686753 444859
rect 692428 444850 693028 444978
rect 698017 444947 698210 444983
rect 698084 444935 698210 444947
rect 702756 444959 703645 444983
rect 702756 444935 702853 444959
rect 698084 444828 702853 444935
rect 686719 444788 686757 444822
rect 680215 444704 680815 444760
rect 686719 444751 686739 444788
rect 686743 444751 686753 444788
rect 686719 444741 686757 444751
rect 686699 444717 686767 444741
rect 686719 444704 686739 444717
rect 686743 444704 686753 444717
rect 686719 444695 686753 444704
rect 686719 444693 686743 444695
rect 692428 444694 693028 444750
rect 686685 444656 686709 444680
rect 686743 444656 686767 444680
rect 678799 444503 679399 444553
rect 680215 444534 680815 444584
rect 692428 444538 693028 444666
rect 680593 444531 680815 444534
rect 682009 444501 682069 444516
rect 682024 444465 682054 444501
rect 683708 444387 684308 444437
rect 678799 444327 679399 444383
rect 692428 444382 693028 444510
rect 714781 444308 714863 445089
rect 715063 444609 715145 445915
rect 715342 445752 715382 445792
rect 715582 445752 715622 445792
rect 715289 444777 715339 445719
rect 715382 445668 715422 445752
rect 715542 445668 715582 445752
rect 715633 444777 715683 445719
rect 715382 444672 715422 444756
rect 715542 444672 715582 444756
rect 715342 444632 715382 444672
rect 715582 444632 715622 444672
rect 715815 444609 715897 445915
rect 715134 444387 715828 444469
rect 716100 444308 716182 446226
rect 716454 445955 717148 446037
rect 716385 444609 716467 445915
rect 716660 445752 716700 445792
rect 716900 445752 716940 445792
rect 716599 444777 716649 445719
rect 716700 445668 716740 445752
rect 716860 445668 716900 445752
rect 716943 444777 716993 445719
rect 716700 444672 716740 444756
rect 716860 444672 716900 444756
rect 716660 444632 716700 444672
rect 716900 444632 716940 444672
rect 717137 444609 717219 445915
rect 716454 444387 717148 444469
rect 717419 444308 717501 446226
rect 683708 444237 684308 444287
rect 692428 444232 693028 444282
rect 678799 444157 679399 444207
rect 684565 444160 684790 444168
rect 696597 444000 696600 444120
rect 714964 444095 715998 444177
rect 716284 444095 717318 444177
rect 21000 417000 21003 417120
rect 282 416623 1316 416705
rect 1602 416623 2636 416705
rect 32810 416662 33035 416670
rect 38201 416593 38801 416643
rect 24572 416518 25172 416568
rect 33292 416513 33892 416563
rect 99 414574 181 416492
rect 452 416331 1146 416413
rect 381 414885 463 416191
rect 660 416128 700 416168
rect 900 416128 940 416168
rect 700 416044 740 416128
rect 860 416044 900 416128
rect 607 415081 657 416023
rect 951 415081 1001 416023
rect 1133 414885 1215 416191
rect 452 414763 1146 414845
rect 1418 414574 1500 416492
rect 1772 416331 2466 416413
rect 1703 414885 1785 416191
rect 1978 416128 2018 416168
rect 2218 416128 2258 416168
rect 2018 416044 2058 416128
rect 2178 416044 2218 416128
rect 1917 415081 1967 416023
rect 2261 415081 2311 416023
rect 2455 414885 2537 416191
rect 2737 415779 2819 416492
rect 24572 416362 25172 416490
rect 38201 416417 38801 416473
rect 33292 416363 33892 416413
rect 24572 416206 25172 416334
rect 35546 416299 35576 416335
rect 36785 416329 36935 416341
rect 35531 416284 35591 416299
rect 36785 416216 37385 416266
rect 38201 416247 38801 416297
rect 30833 416120 30857 416144
rect 30891 416120 30915 416144
rect 24572 416050 25172 416106
rect 30857 416105 30881 416107
rect 30857 416096 30887 416105
rect 30867 416083 30887 416096
rect 30891 416083 30907 416120
rect 30833 416059 30857 416083
rect 30867 416049 30911 416083
rect 14747 415865 19516 415972
rect 24572 415894 25172 416022
rect 30867 416012 30887 416049
rect 30891 416012 30907 416049
rect 36785 416040 37385 416096
rect 30867 415978 30911 416012
rect 30867 415941 30887 415978
rect 30891 415941 30907 415978
rect 30867 415907 30911 415941
rect 30867 415883 30887 415907
rect 30891 415883 30907 415907
rect 14747 415841 14844 415865
rect 13955 415817 14844 415841
rect 19390 415853 19516 415865
rect 19390 415841 19583 415853
rect 19390 415817 19605 415841
rect 19639 415817 19673 415841
rect 19707 415817 19741 415841
rect 19775 415817 19809 415841
rect 19843 415817 19877 415841
rect 19911 415817 19945 415841
rect 19979 415817 20013 415841
rect 20047 415817 20081 415841
rect 20115 415817 20149 415841
rect 20183 415817 20217 415841
rect 20251 415817 20285 415841
rect 20319 415817 20353 415841
rect 20387 415817 20421 415841
rect 20455 415817 20489 415841
rect 20523 415817 20557 415841
rect 20591 415817 20625 415841
rect 20659 415817 20693 415841
rect 2737 415711 2914 415779
rect 1772 414763 2466 414845
rect 2737 414574 2819 415711
rect 2848 415677 2955 415711
rect 19480 415540 19516 415817
rect 19547 415540 19583 415817
rect 24572 415738 25172 415866
rect 36785 415864 37385 415920
rect 36785 415688 37385 415744
rect 20809 415650 20833 415684
rect 20809 415582 20833 415616
rect 24572 415588 25172 415638
rect 20809 415540 20833 415548
rect 36785 415518 37385 415568
rect 3125 414802 3175 415402
rect 3375 414802 3425 415402
rect 282 414471 1316 414553
rect 1602 414471 2636 414553
rect 1389 414444 1392 414445
rect 1389 414443 1390 414444
rect 1391 414443 1392 414444
rect 1389 414442 1392 414443
rect 1526 414444 1529 414445
rect 1526 414443 1527 414444
rect 1528 414443 1529 414444
rect 2848 414443 2955 414477
rect 1526 414442 1529 414443
rect 5488 414280 5538 415103
rect 5658 414280 5708 415103
rect 6005 414280 6021 415499
rect 12427 415448 12493 415464
rect 24572 415458 25172 415508
rect 32930 415457 33530 415507
rect 35287 415391 35887 415441
rect 36785 415402 37385 415452
rect 24572 415308 25172 415358
rect 31463 415307 32063 415357
rect 32930 415301 33530 415357
rect 7389 415277 7406 415287
rect 7440 415277 7477 415287
rect 7511 415277 7551 415287
rect 7585 415277 7622 415287
rect 7656 415277 7696 415287
rect 7730 415277 7767 415287
rect 7801 415277 7841 415287
rect 7875 415277 7912 415287
rect 7946 415277 7986 415287
rect 8020 415277 8057 415287
rect 8091 415277 8131 415287
rect 8165 415277 8202 415287
rect 8236 415277 8296 415287
rect 8330 415277 8381 415287
rect 8996 415277 9044 415287
rect 9078 415277 9120 415287
rect 9154 415277 9197 415287
rect 9231 415277 9291 415287
rect 9325 415277 9362 415287
rect 9396 415277 9436 415287
rect 9470 415277 9507 415287
rect 9541 415277 9581 415287
rect 9615 415277 9652 415287
rect 9686 415277 9726 415287
rect 9760 415277 9797 415287
rect 9831 415277 9871 415287
rect 9905 415277 9942 415287
rect 9976 415277 9990 415287
rect 7389 415209 8389 415277
rect 8990 415183 9990 415277
rect 36785 415226 37385 415282
rect 15678 415127 16678 415177
rect 17278 415127 18278 415177
rect 31463 415151 32063 415207
rect 32930 415151 33530 415201
rect 34079 415157 34679 415207
rect 7389 414840 8389 414864
rect 15678 414860 16678 414916
rect 17278 414860 18278 414916
rect 8990 414840 9990 414841
rect 7389 414743 8389 414799
rect 8990 414743 9990 414799
rect 15678 414788 16678 414844
rect 17278 414788 18278 414844
rect 8990 414701 9990 414702
rect 15678 414286 16678 414426
rect 17278 414286 18278 414426
rect 19844 414280 19894 415051
rect 20462 414280 20512 415051
rect 31463 415001 32063 415051
rect 34079 415001 34679 415057
rect 35287 415039 35887 415095
rect 36785 415050 37385 415106
rect 32596 414929 33596 414979
rect 24573 414820 25173 414870
rect 34079 414851 34679 414901
rect 35287 414869 35887 414919
rect 36785 414880 37385 414930
rect 30171 414795 30771 414845
rect 32596 414773 33596 414829
rect 37993 414704 38593 414754
rect 30171 414619 30771 414675
rect 32596 414623 33596 414673
rect 34110 414589 34710 414639
rect 21263 414280 21313 414518
rect 22349 414280 22399 414518
rect 32596 414507 33596 414557
rect 30171 414449 30771 414499
rect 36785 414429 36985 414609
rect 37993 414534 38593 414584
rect 24573 414352 25173 414408
rect 29993 414310 30993 414360
rect 31347 414280 31547 414317
rect 31607 414280 31807 414317
rect 36785 414280 36985 414373
rect 37083 414280 37120 414373
rect 696597 412200 696600 412320
rect 692376 411983 692396 412017
rect 692463 411993 692532 412017
rect 696191 411993 696239 412017
rect 692487 411983 692532 411993
rect 696204 411983 696239 411993
rect 696340 411983 696360 412017
rect 692487 411915 692502 411939
rect 696200 411915 696215 411939
rect 692454 411891 692478 411915
rect 696224 411891 696248 411915
rect 686755 411800 687355 411850
rect 692487 411748 692505 411752
rect 692479 411718 692505 411748
rect 692487 411698 692505 411718
rect 686755 411624 687355 411680
rect 692485 411674 692505 411698
rect 692509 411674 692517 411718
rect 696215 411698 696223 411748
rect 696203 411674 696223 411698
rect 696227 411674 696245 411752
rect 692485 411640 692521 411674
rect 696203 411640 696249 411674
rect 686755 411448 687355 411504
rect 686755 411278 687355 411328
rect 685547 411102 686147 411152
rect 687155 411007 687170 411022
rect 687343 411018 687355 411022
rect 687340 411007 687355 411018
rect 685547 410932 686147 410982
rect 687155 410827 687355 411007
rect 687155 410812 687170 410827
rect 687340 410816 687355 410827
rect 687343 410812 687355 410816
rect 687042 410771 687057 410786
rect 687020 410591 687057 410771
rect 687155 410771 687170 410786
rect 687343 410782 687355 410786
rect 687340 410771 687355 410782
rect 687155 410591 687355 410771
rect 688210 410630 688260 411630
rect 688360 410740 688488 411630
rect 688516 410740 688644 411630
rect 688672 410740 688800 411630
rect 688828 410740 688956 411630
rect 688984 410740 689112 411630
rect 689140 410740 689268 411630
rect 689296 410740 689424 411630
rect 689452 410740 689580 411630
rect 689608 410740 689736 411630
rect 689764 410740 689892 411630
rect 689920 410740 690048 411630
rect 690076 410740 690204 411630
rect 690232 410740 690360 411630
rect 690388 410630 690438 411630
rect 692485 411606 692505 411640
rect 692509 411606 692517 411640
rect 696203 411606 696223 411640
rect 696227 411606 696245 411640
rect 691275 411523 691875 411573
rect 692485 411572 692521 411606
rect 696203 411572 696249 411606
rect 692485 411538 692505 411572
rect 692509 411538 692517 411572
rect 692485 411504 692521 411538
rect 692583 411528 693983 411571
rect 694719 411528 696119 411571
rect 696203 411538 696223 411572
rect 696227 411538 696245 411572
rect 696203 411504 696249 411538
rect 692485 411470 692505 411504
rect 692509 411470 692517 411504
rect 692485 411436 692521 411470
rect 691275 411373 691875 411423
rect 692485 411402 692505 411436
rect 692509 411402 692517 411436
rect 692485 411368 692521 411402
rect 692485 411334 692505 411368
rect 692509 411334 692517 411368
rect 692583 411365 693983 411493
rect 694719 411365 696119 411493
rect 696203 411470 696223 411504
rect 696227 411470 696245 411504
rect 696203 411436 696249 411470
rect 707624 411441 707658 411475
rect 707695 411441 707729 411475
rect 707769 411441 707803 411475
rect 707840 411441 707874 411475
rect 707914 411441 707948 411475
rect 707985 411441 708019 411475
rect 708059 411441 708093 411475
rect 708130 411441 708164 411475
rect 708204 411441 708238 411475
rect 708275 411441 708309 411475
rect 708369 411441 708403 411475
rect 708446 411441 708480 411475
rect 708520 411441 708554 411465
rect 708588 411441 708610 411465
rect 709211 411441 709234 411465
rect 709270 411441 709304 411475
rect 709364 411441 709398 411475
rect 709435 411441 709469 411475
rect 709509 411441 709543 411475
rect 709580 411441 709614 411475
rect 709654 411441 709688 411475
rect 709725 411441 709759 411475
rect 709799 411441 709833 411475
rect 709870 411441 709904 411475
rect 709944 411441 709978 411475
rect 710015 411441 710049 411475
rect 710089 411441 710123 411475
rect 710160 411441 710194 411475
rect 696203 411402 696223 411436
rect 696227 411402 696245 411436
rect 707610 411431 707624 411441
rect 707658 411431 707695 411441
rect 707729 411431 707769 411441
rect 707803 411431 707840 411441
rect 707874 411431 707914 411441
rect 707948 411431 707985 411441
rect 708019 411431 708059 411441
rect 708093 411431 708130 411441
rect 708164 411431 708204 411441
rect 708238 411431 708275 411441
rect 708309 411431 708369 411441
rect 708403 411431 708446 411441
rect 708480 411431 708520 411441
rect 708554 411431 708588 411441
rect 708610 411431 708634 411441
rect 709211 411431 709270 411441
rect 709304 411431 709364 411441
rect 709398 411431 709435 411441
rect 709469 411431 709509 411441
rect 709543 411431 709580 411441
rect 709614 411431 709654 411441
rect 709688 411431 709725 411441
rect 709759 411431 709799 411441
rect 709833 411431 709870 411441
rect 709904 411431 709944 411441
rect 709978 411431 710015 411441
rect 710049 411431 710089 411441
rect 710123 411431 710160 411441
rect 710194 411431 710211 411441
rect 696203 411368 696249 411402
rect 696203 411334 696223 411368
rect 696227 411334 696245 411368
rect 707610 411337 708610 411431
rect 709211 411337 710211 411431
rect 691275 411251 691875 411301
rect 692485 411300 692521 411334
rect 692485 411266 692505 411300
rect 692509 411266 692517 411300
rect 692485 411232 692521 411266
rect 692485 411198 692505 411232
rect 692509 411198 692517 411232
rect 692583 411202 693983 411330
rect 694719 411202 696119 411330
rect 696203 411300 696249 411334
rect 711579 411317 712463 411331
rect 711579 411307 711619 411317
rect 696203 411266 696223 411300
rect 696227 411266 696245 411300
rect 701730 411290 701747 411292
rect 696203 411232 696249 411266
rect 696203 411198 696223 411232
rect 696227 411198 696245 411232
rect 701692 411220 701722 411254
rect 701730 411220 701760 411290
rect 707610 411241 708610 411301
rect 709211 411241 710211 411301
rect 692485 411164 692521 411198
rect 691275 411101 691875 411151
rect 692485 411130 692505 411164
rect 692509 411130 692517 411164
rect 692485 411096 692521 411130
rect 692485 411062 692505 411096
rect 692509 411062 692517 411096
rect 692485 411028 692521 411062
rect 692583 411039 693983 411167
rect 694719 411039 696119 411167
rect 696203 411164 696249 411198
rect 696203 411130 696223 411164
rect 696227 411130 696245 411164
rect 696203 411096 696249 411130
rect 696203 411062 696223 411096
rect 696227 411062 696245 411096
rect 699322 411064 700322 411097
rect 700922 411064 701922 411097
rect 696203 411028 696249 411062
rect 707610 411044 708610 411048
rect 709211 411044 710211 411048
rect 691275 410975 691875 411025
rect 692485 410994 692505 411028
rect 692509 410994 692517 411028
rect 692485 410960 692521 410994
rect 692485 410926 692505 410960
rect 692509 410926 692517 410960
rect 692485 410892 692521 410926
rect 691275 410825 691875 410875
rect 692485 410858 692505 410892
rect 692509 410858 692517 410892
rect 692583 410876 693983 411004
rect 694719 410876 696119 411004
rect 696203 410994 696223 411028
rect 696227 410994 696245 411028
rect 707574 410994 708646 411030
rect 696203 410960 696249 410994
rect 696203 410926 696223 410960
rect 696227 410926 696245 410960
rect 707574 410953 707610 410994
rect 708610 410953 708646 410994
rect 696203 410892 696249 410926
rect 697284 410894 697350 410910
rect 707574 410897 708646 410953
rect 696203 410858 696223 410892
rect 696227 410858 696245 410892
rect 699322 410877 700322 410894
rect 700922 410877 701922 410894
rect 707574 410881 707610 410897
rect 708610 410881 708646 410897
rect 692485 410824 692521 410858
rect 692485 410790 692505 410824
rect 692509 410790 692517 410824
rect 692485 410756 692521 410790
rect 691275 410703 691875 410753
rect 692485 410740 692505 410756
rect 692509 410740 692517 410756
rect 692583 410740 693983 410841
rect 694719 410740 696119 410841
rect 696203 410824 696249 410858
rect 707574 410825 708646 410881
rect 696203 410790 696223 410824
rect 696227 410790 696245 410824
rect 696203 410756 696249 410790
rect 696203 410740 696223 410756
rect 696227 410740 696245 410756
rect 699322 410740 700322 410811
rect 700922 410740 701922 410811
rect 707574 410788 707610 410825
rect 708610 410788 708646 410825
rect 707574 410748 708646 410788
rect 709175 410994 710247 411030
rect 709175 410953 709211 410994
rect 710211 410953 710247 410994
rect 709175 410897 710247 410953
rect 709175 410881 709211 410897
rect 710211 410881 710247 410897
rect 709175 410825 710247 410881
rect 709175 410788 709211 410825
rect 710211 410788 710247 410825
rect 709175 410748 710247 410788
rect 685542 410506 686142 410556
rect 691275 410553 691875 410603
rect 685542 410330 686142 410386
rect 692583 410237 693983 410280
rect 694719 410237 696119 410280
rect 699322 410278 700322 410418
rect 700922 410278 701922 410418
rect 685542 410160 686142 410210
rect 692583 410101 693983 410144
rect 694719 410101 696119 410144
rect 680215 409678 680815 409728
rect 680215 409502 680815 409558
rect 685551 409516 686551 409566
rect 689154 409480 689204 409897
rect 689304 409480 689360 409897
rect 689460 409480 689516 409897
rect 689616 409480 689672 409897
rect 689772 409480 689828 409897
rect 689928 409480 689978 409897
rect 699322 409860 700322 409916
rect 700922 409860 701922 409916
rect 707610 409905 708610 409961
rect 709211 409905 710211 409961
rect 699322 409788 700322 409844
rect 700922 409788 701922 409844
rect 707610 409833 708610 409889
rect 709211 409833 710211 409889
rect 711579 409525 711605 411307
rect 715956 410297 716006 411297
rect 716106 410740 716234 411297
rect 716262 410297 716312 411297
rect 711579 409480 711595 409495
rect 712409 409480 712431 409485
rect 713640 409480 713641 409785
rect 713750 409772 714750 409822
rect 713750 409562 714750 409612
rect 713750 409480 714750 409496
rect 2850 403304 3850 403320
rect 2850 403188 3850 403238
rect 2850 402978 3850 403028
rect 3959 403015 3960 403320
rect 5169 403315 5191 403320
rect 6005 403305 6021 403320
rect 1288 401503 1338 402503
rect 1438 401503 1566 402060
rect 1594 401503 1644 402503
rect 5995 401493 6021 403275
rect 7389 402911 8389 402967
rect 8990 402911 9990 402967
rect 15678 402956 16678 403012
rect 17278 402956 18278 403012
rect 7389 402839 8389 402895
rect 8990 402839 9990 402895
rect 15678 402884 16678 402940
rect 17278 402884 18278 402940
rect 27622 402903 27672 403320
rect 27772 402903 27828 403320
rect 27928 402903 27984 403320
rect 28084 402903 28140 403320
rect 28240 402903 28296 403320
rect 28396 402903 28446 403320
rect 31049 403234 32049 403284
rect 36785 403242 37385 403298
rect 36785 403072 37385 403122
rect 21481 402656 22881 402699
rect 23617 402656 25017 402699
rect 31458 402590 32058 402640
rect 15678 402382 16678 402522
rect 17278 402382 18278 402522
rect 21481 402520 22881 402563
rect 23617 402520 25017 402563
rect 31458 402414 32058 402470
rect 25725 402197 26325 402247
rect 31458 402244 32058 402294
rect 7353 402016 8425 402052
rect 7353 401975 7389 402016
rect 8389 401975 8425 402016
rect 7353 401919 8425 401975
rect 7353 401903 7389 401919
rect 8389 401903 8425 401919
rect 7353 401847 8425 401903
rect 7353 401810 7389 401847
rect 8389 401810 8425 401847
rect 7353 401770 8425 401810
rect 8954 402016 10026 402052
rect 8954 401975 8990 402016
rect 9990 401975 10026 402016
rect 8954 401919 10026 401975
rect 21383 402044 21403 402060
rect 21407 402044 21415 402060
rect 21383 402010 21419 402044
rect 21481 402031 22881 402060
rect 23617 402031 25017 402060
rect 25101 402044 25121 402060
rect 25125 402044 25143 402060
rect 25725 402047 26325 402097
rect 25101 402010 25147 402044
rect 21383 401976 21403 402010
rect 21407 401976 21415 402010
rect 21383 401942 21419 401976
rect 8954 401903 8990 401919
rect 9990 401903 10026 401919
rect 15678 401906 16678 401923
rect 17278 401906 18278 401923
rect 21383 401908 21403 401942
rect 21407 401908 21415 401942
rect 8954 401847 10026 401903
rect 20250 401890 20316 401906
rect 8954 401810 8990 401847
rect 9990 401810 10026 401847
rect 8954 401770 10026 401810
rect 21383 401874 21419 401908
rect 21383 401840 21403 401874
rect 21407 401840 21415 401874
rect 21481 401868 22881 401996
rect 23617 401868 25017 401996
rect 25101 401976 25121 402010
rect 25125 401976 25143 402010
rect 25101 401942 25147 401976
rect 25101 401908 25121 401942
rect 25125 401908 25143 401942
rect 25725 401925 26325 401975
rect 25101 401874 25147 401908
rect 25101 401840 25121 401874
rect 25125 401840 25143 401874
rect 21383 401806 21419 401840
rect 21383 401772 21403 401806
rect 21407 401772 21415 401806
rect 21383 401738 21419 401772
rect 15678 401703 16678 401736
rect 17278 401703 18278 401736
rect 21383 401704 21403 401738
rect 21407 401704 21415 401738
rect 21481 401705 22881 401833
rect 23617 401705 25017 401833
rect 25101 401806 25147 401840
rect 25101 401772 25121 401806
rect 25125 401772 25143 401806
rect 25725 401775 26325 401825
rect 25101 401738 25147 401772
rect 25101 401704 25121 401738
rect 25125 401704 25143 401738
rect 21383 401670 21419 401704
rect 25101 401670 25147 401704
rect 21383 401636 21403 401670
rect 21407 401636 21415 401670
rect 7389 401559 8389 401631
rect 8990 401559 9990 401631
rect 21383 401602 21419 401636
rect 15840 401510 15870 401580
rect 15878 401546 15908 401580
rect 21383 401568 21403 401602
rect 21407 401568 21415 401602
rect 15853 401508 15870 401510
rect 21383 401534 21419 401568
rect 21481 401542 22881 401670
rect 23617 401542 25017 401670
rect 25101 401636 25121 401670
rect 25125 401636 25143 401670
rect 25725 401649 26325 401699
rect 25101 401602 25147 401636
rect 25101 401568 25121 401602
rect 25125 401568 25143 401602
rect 25101 401534 25147 401568
rect 5981 401483 6021 401493
rect 5137 401469 6021 401483
rect 21383 401500 21403 401534
rect 21407 401500 21415 401534
rect 21383 401466 21419 401500
rect 7389 401369 8389 401463
rect 7389 401359 8413 401369
rect 8990 401359 9990 401463
rect 21383 401432 21403 401466
rect 21407 401432 21415 401466
rect 21383 401398 21419 401432
rect 21383 401364 21403 401398
rect 21407 401364 21415 401398
rect 21481 401379 22881 401507
rect 23617 401379 25017 401507
rect 25101 401500 25121 401534
rect 25125 401500 25143 401534
rect 25101 401466 25147 401500
rect 25725 401499 26325 401549
rect 25101 401432 25121 401466
rect 25125 401432 25143 401466
rect 25101 401398 25147 401432
rect 25101 401364 25121 401398
rect 25125 401364 25143 401398
rect 25725 401377 26325 401427
rect 21383 401330 21419 401364
rect 25101 401330 25147 401364
rect 21383 401296 21403 401330
rect 21407 401296 21415 401330
rect 25101 401296 25121 401330
rect 25125 401296 25143 401330
rect 21383 401262 21419 401296
rect 21383 401228 21403 401262
rect 21407 401228 21415 401262
rect 21481 401229 22881 401272
rect 23617 401229 25017 401272
rect 25101 401262 25147 401296
rect 25101 401228 25121 401262
rect 25125 401228 25143 401262
rect 21383 401194 21419 401228
rect 25101 401194 25147 401228
rect 25725 401227 26325 401277
rect 21383 401160 21403 401194
rect 21407 401160 21415 401194
rect 25101 401160 25121 401194
rect 25125 401160 25143 401194
rect 27162 401170 27212 402170
rect 27312 401170 27440 402060
rect 27468 401170 27596 402060
rect 27624 401170 27752 402060
rect 27780 401170 27908 402060
rect 27936 401170 28064 402060
rect 28092 401170 28220 402060
rect 28248 401170 28376 402060
rect 28404 401170 28532 402060
rect 28560 401170 28688 402060
rect 28716 401170 28844 402060
rect 28872 401170 29000 402060
rect 29028 401170 29156 402060
rect 29184 401170 29312 402060
rect 29340 401170 29390 402170
rect 30245 402029 30445 402209
rect 30245 402018 30260 402029
rect 30245 402014 30257 402018
rect 30430 402014 30445 402029
rect 30543 402029 30580 402209
rect 30543 402014 30558 402029
rect 30245 401984 30257 401988
rect 30245 401973 30260 401984
rect 30430 401973 30445 401988
rect 30245 401793 30445 401973
rect 31453 401818 32053 401868
rect 30245 401782 30260 401793
rect 30245 401778 30257 401782
rect 30430 401778 30445 401793
rect 31453 401648 32053 401698
rect 30245 401472 30845 401522
rect 30245 401296 30845 401352
rect 21383 401126 21419 401160
rect 25101 401126 25147 401160
rect 21383 401102 21403 401126
rect 21385 401048 21403 401102
rect 21407 401082 21415 401126
rect 25101 401102 25121 401126
rect 25113 401082 25121 401102
rect 25125 401048 25143 401126
rect 30245 401120 30845 401176
rect 30245 400950 30845 401000
rect 21000 400800 21003 400920
rect 21352 400885 21376 400909
rect 25122 400885 25146 400909
rect 21385 400861 21400 400885
rect 25098 400861 25113 400885
rect 21274 400783 21294 400851
rect 21410 400817 21430 400851
rect 25068 400817 25088 400851
rect 25204 400817 25224 400851
rect 21385 400807 21430 400817
rect 25102 400807 25137 400817
rect 21361 400783 21430 400807
rect 25089 400783 25137 400807
rect 25238 400783 25258 400817
rect 680480 398427 680517 398520
rect 680615 398427 680815 398520
rect 685793 398483 685993 398520
rect 686053 398483 686253 398520
rect 686607 398440 687607 398490
rect 692427 398392 693027 398448
rect 679007 398216 679607 398266
rect 680615 398191 680815 398371
rect 686829 398301 687429 398351
rect 684004 398243 685004 398293
rect 695201 398282 695251 398520
rect 696287 398282 696337 398520
rect 682890 398161 683490 398211
rect 684004 398127 685004 398177
rect 686829 398125 687429 398181
rect 679007 398046 679607 398096
rect 684004 397971 685004 398027
rect 686829 397955 687429 398005
rect 680215 397870 680815 397920
rect 681713 397881 682313 397931
rect 682921 397899 683521 397949
rect 692427 397930 693027 397980
rect 684004 397821 685004 397871
rect 680215 397694 680815 397750
rect 681713 397705 682313 397761
rect 682921 397743 683521 397799
rect 685537 397749 686137 397799
rect 697088 397749 697138 398520
rect 697706 397749 697756 398520
rect 699322 398374 700322 398514
rect 700922 398374 701922 398514
rect 707610 398098 708610 398099
rect 699322 397956 700322 398012
rect 700922 397956 701922 398012
rect 707610 398001 708610 398057
rect 709211 398001 710211 398057
rect 707610 397959 708610 397960
rect 699322 397884 700322 397940
rect 700922 397884 701922 397940
rect 709211 397936 710211 397960
rect 682921 397593 683521 397643
rect 684070 397599 684670 397649
rect 685537 397593 686137 397649
rect 699322 397623 700322 397673
rect 700922 397623 701922 397673
rect 680215 397518 680815 397574
rect 707610 397523 708610 397617
rect 709211 397523 710211 397591
rect 707610 397513 707624 397523
rect 707658 397513 707695 397523
rect 707729 397513 707769 397523
rect 707803 397513 707840 397523
rect 707874 397513 707914 397523
rect 707948 397513 707985 397523
rect 708019 397513 708059 397523
rect 708093 397513 708130 397523
rect 708164 397513 708204 397523
rect 708238 397513 708275 397523
rect 708309 397513 708369 397523
rect 708403 397513 708446 397523
rect 708480 397513 708522 397523
rect 708556 397513 708604 397523
rect 709219 397513 709270 397523
rect 709304 397513 709364 397523
rect 709398 397513 709435 397523
rect 709469 397513 709509 397523
rect 709543 397513 709580 397523
rect 709614 397513 709654 397523
rect 709688 397513 709725 397523
rect 709759 397513 709799 397523
rect 709833 397513 709870 397523
rect 709904 397513 709944 397523
rect 709978 397513 710015 397523
rect 710049 397513 710089 397523
rect 710123 397513 710160 397523
rect 710194 397513 710211 397523
rect 684070 397443 684670 397499
rect 685537 397443 686137 397493
rect 692428 397442 693028 397492
rect 680215 397348 680815 397398
rect 681713 397359 682313 397409
rect 684070 397293 684670 397343
rect 692428 397292 693028 397342
rect 705107 397336 705173 397352
rect 711579 397301 711595 398520
rect 711892 397697 711942 398520
rect 712062 397697 712112 398520
rect 716071 398357 716074 398358
rect 714645 398323 714752 398357
rect 716071 398356 716072 398357
rect 716073 398356 716074 398357
rect 716071 398355 716074 398356
rect 716208 398357 716211 398358
rect 716208 398356 716209 398357
rect 716210 398356 716211 398357
rect 716208 398355 716211 398356
rect 714964 398247 715998 398329
rect 716284 398247 717318 398329
rect 714175 397398 714225 397998
rect 714425 397398 714475 397998
rect 680215 397232 680815 397282
rect 698017 397232 698053 397260
rect 692428 397162 693028 397212
rect 698030 397198 698077 397232
rect 698017 397164 698053 397198
rect 680215 397056 680815 397112
rect 692428 397006 693028 397134
rect 698030 397130 698077 397164
rect 698017 397096 698053 397130
rect 698030 397062 698077 397096
rect 698017 396983 698053 397062
rect 698084 396983 698120 397260
rect 714781 397191 714863 398226
rect 715134 397955 715828 398037
rect 714686 397123 714863 397191
rect 714645 397089 714863 397123
rect 680215 396880 680815 396936
rect 686719 396893 686739 396917
rect 686743 396893 686753 396917
rect 686719 396859 686757 396893
rect 686719 396822 686739 396859
rect 686743 396822 686753 396859
rect 692428 396850 693028 396978
rect 698017 396947 698210 396983
rect 698084 396935 698210 396947
rect 702756 396959 703645 396983
rect 702756 396935 702853 396959
rect 698084 396828 702853 396935
rect 686719 396788 686757 396822
rect 680215 396704 680815 396760
rect 686719 396751 686739 396788
rect 686743 396751 686753 396788
rect 686719 396741 686757 396751
rect 686699 396717 686767 396741
rect 686719 396704 686739 396717
rect 686743 396704 686753 396717
rect 686719 396695 686753 396704
rect 686719 396693 686743 396695
rect 692428 396694 693028 396750
rect 686685 396656 686709 396680
rect 686743 396656 686767 396680
rect 678799 396503 679399 396553
rect 680215 396534 680815 396584
rect 692428 396538 693028 396666
rect 680593 396531 680815 396534
rect 682009 396501 682069 396516
rect 682024 396465 682054 396501
rect 683708 396387 684308 396437
rect 678799 396327 679399 396383
rect 692428 396382 693028 396510
rect 714781 396308 714863 397089
rect 715063 396609 715145 397915
rect 715289 396777 715339 397719
rect 715633 396777 715683 397719
rect 715382 396672 715422 396756
rect 715542 396672 715582 396756
rect 715342 396632 715382 396672
rect 715582 396632 715622 396672
rect 715815 396609 715897 397915
rect 715134 396387 715828 396469
rect 716100 396308 716182 398226
rect 716454 397955 717148 398037
rect 716385 396609 716467 397915
rect 716599 396777 716649 397719
rect 716943 396777 716993 397719
rect 716700 396672 716740 396756
rect 716860 396672 716900 396756
rect 716660 396632 716700 396672
rect 716900 396632 716940 396672
rect 717137 396609 717219 397915
rect 716454 396387 717148 396469
rect 717419 396308 717501 398226
rect 683708 396237 684308 396287
rect 692428 396232 693028 396282
rect 678799 396157 679399 396207
rect 684565 396160 684790 396168
rect 696597 396000 696600 396120
rect 714964 396095 715998 396177
rect 716284 396095 717318 396177
rect 21000 369000 21003 369120
rect 282 368623 1316 368705
rect 1602 368623 2636 368705
rect 32810 368662 33035 368670
rect 38201 368593 38801 368643
rect 24572 368518 25172 368568
rect 33292 368513 33892 368563
rect 99 366574 181 368492
rect 452 368331 1146 368413
rect 381 366885 463 368191
rect 660 368128 700 368168
rect 900 368128 940 368168
rect 700 368044 740 368128
rect 860 368044 900 368128
rect 607 367081 657 368023
rect 951 367081 1001 368023
rect 1133 366885 1215 368191
rect 452 366763 1146 366845
rect 1418 366574 1500 368492
rect 1772 368331 2466 368413
rect 1703 366885 1785 368191
rect 1978 368128 2018 368168
rect 2218 368128 2258 368168
rect 2018 368044 2058 368128
rect 2178 368044 2218 368128
rect 1917 367081 1967 368023
rect 2261 367081 2311 368023
rect 2455 366885 2537 368191
rect 2737 367779 2819 368492
rect 24572 368362 25172 368490
rect 38201 368417 38801 368473
rect 33292 368363 33892 368413
rect 24572 368206 25172 368334
rect 35546 368299 35576 368335
rect 36785 368329 36935 368341
rect 35531 368284 35591 368299
rect 36785 368216 37385 368266
rect 38201 368247 38801 368297
rect 30833 368120 30857 368144
rect 30891 368120 30915 368144
rect 24572 368050 25172 368106
rect 30857 368105 30881 368107
rect 30857 368096 30887 368105
rect 30867 368083 30887 368096
rect 30891 368083 30907 368120
rect 30833 368059 30857 368083
rect 30867 368049 30911 368083
rect 14747 367865 19516 367972
rect 24572 367894 25172 368022
rect 30867 368012 30887 368049
rect 30891 368012 30907 368049
rect 36785 368040 37385 368096
rect 30867 367978 30911 368012
rect 30867 367941 30887 367978
rect 30891 367941 30907 367978
rect 30867 367907 30911 367941
rect 30867 367883 30887 367907
rect 30891 367883 30907 367907
rect 14747 367841 14844 367865
rect 13955 367817 14844 367841
rect 19390 367853 19516 367865
rect 19390 367841 19583 367853
rect 19390 367817 19605 367841
rect 19639 367817 19673 367841
rect 19707 367817 19741 367841
rect 19775 367817 19809 367841
rect 19843 367817 19877 367841
rect 19911 367817 19945 367841
rect 19979 367817 20013 367841
rect 20047 367817 20081 367841
rect 20115 367817 20149 367841
rect 20183 367817 20217 367841
rect 20251 367817 20285 367841
rect 20319 367817 20353 367841
rect 20387 367817 20421 367841
rect 20455 367817 20489 367841
rect 20523 367817 20557 367841
rect 20591 367817 20625 367841
rect 20659 367817 20693 367841
rect 2737 367711 2914 367779
rect 1772 366763 2466 366845
rect 2737 366574 2819 367711
rect 2848 367677 2955 367711
rect 19480 367540 19516 367817
rect 19547 367540 19583 367817
rect 24572 367738 25172 367866
rect 36785 367864 37385 367920
rect 36785 367688 37385 367744
rect 20809 367650 20833 367684
rect 20809 367582 20833 367616
rect 24572 367588 25172 367638
rect 20809 367540 20833 367548
rect 36785 367518 37385 367568
rect 3125 366802 3175 367402
rect 3375 366802 3425 367402
rect 282 366471 1316 366553
rect 1602 366471 2636 366553
rect 1389 366444 1392 366445
rect 1389 366443 1390 366444
rect 1391 366443 1392 366444
rect 1389 366442 1392 366443
rect 1526 366444 1529 366445
rect 1526 366443 1527 366444
rect 1528 366443 1529 366444
rect 2848 366443 2955 366477
rect 1526 366442 1529 366443
rect 5488 366280 5538 367103
rect 5658 366280 5708 367103
rect 6005 366280 6021 367499
rect 12427 367448 12493 367464
rect 24572 367458 25172 367508
rect 32930 367457 33530 367507
rect 35287 367391 35887 367441
rect 36785 367402 37385 367452
rect 24572 367308 25172 367358
rect 31463 367307 32063 367357
rect 32930 367301 33530 367357
rect 7389 367277 7406 367287
rect 7440 367277 7477 367287
rect 7511 367277 7551 367287
rect 7585 367277 7622 367287
rect 7656 367277 7696 367287
rect 7730 367277 7767 367287
rect 7801 367277 7841 367287
rect 7875 367277 7912 367287
rect 7946 367277 7986 367287
rect 8020 367277 8057 367287
rect 8091 367277 8131 367287
rect 8165 367277 8202 367287
rect 8236 367277 8296 367287
rect 8330 367277 8381 367287
rect 8996 367277 9044 367287
rect 9078 367277 9120 367287
rect 9154 367277 9197 367287
rect 9231 367277 9291 367287
rect 9325 367277 9362 367287
rect 9396 367277 9436 367287
rect 9470 367277 9507 367287
rect 9541 367277 9581 367287
rect 9615 367277 9652 367287
rect 9686 367277 9726 367287
rect 9760 367277 9797 367287
rect 9831 367277 9871 367287
rect 9905 367277 9942 367287
rect 9976 367277 9990 367287
rect 7389 367209 8389 367277
rect 8990 367183 9990 367277
rect 36785 367226 37385 367282
rect 15678 367127 16678 367177
rect 17278 367127 18278 367177
rect 31463 367151 32063 367207
rect 32930 367151 33530 367201
rect 34079 367157 34679 367207
rect 7389 366840 8389 366864
rect 15678 366860 16678 366916
rect 17278 366860 18278 366916
rect 8990 366840 9990 366841
rect 7389 366743 8389 366799
rect 8990 366743 9990 366799
rect 15678 366788 16678 366844
rect 17278 366788 18278 366844
rect 8990 366701 9990 366702
rect 15678 366286 16678 366426
rect 17278 366286 18278 366426
rect 19844 366280 19894 367051
rect 20462 366280 20512 367051
rect 31463 367001 32063 367051
rect 34079 367001 34679 367057
rect 35287 367039 35887 367095
rect 36785 367050 37385 367106
rect 32596 366929 33596 366979
rect 24573 366820 25173 366870
rect 34079 366851 34679 366901
rect 35287 366869 35887 366919
rect 36785 366880 37385 366930
rect 30171 366795 30771 366845
rect 32596 366773 33596 366829
rect 37993 366704 38593 366754
rect 30171 366619 30771 366675
rect 32596 366623 33596 366673
rect 34110 366589 34710 366639
rect 21263 366280 21313 366518
rect 22349 366280 22399 366518
rect 32596 366507 33596 366557
rect 30171 366449 30771 366499
rect 36785 366429 36985 366609
rect 37993 366534 38593 366584
rect 24573 366352 25173 366408
rect 29993 366310 30993 366360
rect 31347 366280 31547 366317
rect 31607 366280 31807 366317
rect 36785 366280 36985 366373
rect 37083 366280 37120 366373
rect 696597 364200 696600 364320
rect 692376 363983 692396 364017
rect 692463 363993 692532 364017
rect 696191 363993 696239 364017
rect 692487 363983 692532 363993
rect 696204 363983 696239 363993
rect 696340 363983 696360 364017
rect 692487 363915 692502 363939
rect 696200 363915 696215 363939
rect 692454 363891 692478 363915
rect 696224 363891 696248 363915
rect 686755 363800 687355 363850
rect 692487 363748 692505 363752
rect 692479 363718 692505 363748
rect 692487 363698 692505 363718
rect 686755 363624 687355 363680
rect 692485 363674 692505 363698
rect 692509 363674 692517 363718
rect 696215 363698 696223 363748
rect 696203 363674 696223 363698
rect 696227 363674 696245 363752
rect 692485 363640 692521 363674
rect 696203 363640 696249 363674
rect 686755 363448 687355 363504
rect 686755 363278 687355 363328
rect 685547 363102 686147 363152
rect 687155 363007 687170 363022
rect 687343 363018 687355 363022
rect 687340 363007 687355 363018
rect 685547 362932 686147 362982
rect 687155 362827 687355 363007
rect 687155 362812 687170 362827
rect 687340 362816 687355 362827
rect 687343 362812 687355 362816
rect 687042 362771 687057 362786
rect 687020 362591 687057 362771
rect 687042 362576 687057 362591
rect 687155 362771 687170 362786
rect 687343 362782 687355 362786
rect 687340 362771 687355 362782
rect 687155 362591 687355 362771
rect 688210 362630 688260 363630
rect 688360 362630 688488 363630
rect 688516 362630 688644 363630
rect 688672 362630 688800 363630
rect 688828 362630 688956 363630
rect 688984 362630 689112 363630
rect 689140 362630 689268 363630
rect 689296 362630 689424 363630
rect 689452 362630 689580 363630
rect 689608 362630 689736 363630
rect 689764 362630 689892 363630
rect 689920 362630 690048 363630
rect 690076 362630 690204 363630
rect 690232 362630 690360 363630
rect 690388 362630 690438 363630
rect 692485 363606 692505 363640
rect 692509 363606 692517 363640
rect 696203 363606 696223 363640
rect 696227 363606 696245 363640
rect 691275 363523 691875 363573
rect 692485 363572 692521 363606
rect 696203 363572 696249 363606
rect 692485 363538 692505 363572
rect 692509 363538 692517 363572
rect 692485 363504 692521 363538
rect 692583 363528 693983 363571
rect 694719 363528 696119 363571
rect 696203 363538 696223 363572
rect 696227 363538 696245 363572
rect 696203 363504 696249 363538
rect 692485 363470 692505 363504
rect 692509 363470 692517 363504
rect 692485 363436 692521 363470
rect 691275 363373 691875 363423
rect 692485 363402 692505 363436
rect 692509 363402 692517 363436
rect 692485 363368 692521 363402
rect 692485 363334 692505 363368
rect 692509 363334 692517 363368
rect 692583 363365 693983 363493
rect 694719 363365 696119 363493
rect 696203 363470 696223 363504
rect 696227 363470 696245 363504
rect 696203 363436 696249 363470
rect 707624 363441 707658 363475
rect 707695 363441 707729 363475
rect 707769 363441 707803 363475
rect 707840 363441 707874 363475
rect 707914 363441 707948 363475
rect 707985 363441 708019 363475
rect 708059 363441 708093 363475
rect 708130 363441 708164 363475
rect 708204 363441 708238 363475
rect 708275 363441 708309 363475
rect 708369 363441 708403 363475
rect 708446 363441 708480 363475
rect 708520 363441 708554 363465
rect 708588 363441 708610 363465
rect 709211 363441 709234 363465
rect 709270 363441 709304 363475
rect 709364 363441 709398 363475
rect 709435 363441 709469 363475
rect 709509 363441 709543 363475
rect 709580 363441 709614 363475
rect 709654 363441 709688 363475
rect 709725 363441 709759 363475
rect 709799 363441 709833 363475
rect 709870 363441 709904 363475
rect 709944 363441 709978 363475
rect 710015 363441 710049 363475
rect 710089 363441 710123 363475
rect 710160 363441 710194 363475
rect 696203 363402 696223 363436
rect 696227 363402 696245 363436
rect 707610 363431 707624 363441
rect 707658 363431 707695 363441
rect 707729 363431 707769 363441
rect 707803 363431 707840 363441
rect 707874 363431 707914 363441
rect 707948 363431 707985 363441
rect 708019 363431 708059 363441
rect 708093 363431 708130 363441
rect 708164 363431 708204 363441
rect 708238 363431 708275 363441
rect 708309 363431 708369 363441
rect 708403 363431 708446 363441
rect 708480 363431 708520 363441
rect 708554 363431 708588 363441
rect 708610 363431 708634 363441
rect 709211 363431 709270 363441
rect 709304 363431 709364 363441
rect 709398 363431 709435 363441
rect 709469 363431 709509 363441
rect 709543 363431 709580 363441
rect 709614 363431 709654 363441
rect 709688 363431 709725 363441
rect 709759 363431 709799 363441
rect 709833 363431 709870 363441
rect 709904 363431 709944 363441
rect 709978 363431 710015 363441
rect 710049 363431 710089 363441
rect 710123 363431 710160 363441
rect 710194 363431 710211 363441
rect 696203 363368 696249 363402
rect 696203 363334 696223 363368
rect 696227 363334 696245 363368
rect 707610 363337 708610 363431
rect 709211 363337 710211 363431
rect 691275 363251 691875 363301
rect 692485 363300 692521 363334
rect 692485 363266 692505 363300
rect 692509 363266 692517 363300
rect 692485 363232 692521 363266
rect 692485 363198 692505 363232
rect 692509 363198 692517 363232
rect 692583 363202 693983 363330
rect 694719 363202 696119 363330
rect 696203 363300 696249 363334
rect 711579 363317 712463 363331
rect 711579 363307 711619 363317
rect 696203 363266 696223 363300
rect 696227 363266 696245 363300
rect 701730 363290 701747 363292
rect 696203 363232 696249 363266
rect 696203 363198 696223 363232
rect 696227 363198 696245 363232
rect 701692 363220 701722 363254
rect 701730 363220 701760 363290
rect 707610 363241 708610 363301
rect 709211 363241 710211 363301
rect 692485 363164 692521 363198
rect 691275 363101 691875 363151
rect 692485 363130 692505 363164
rect 692509 363130 692517 363164
rect 692485 363096 692521 363130
rect 692485 363062 692505 363096
rect 692509 363062 692517 363096
rect 692485 363028 692521 363062
rect 692583 363039 693983 363167
rect 694719 363039 696119 363167
rect 696203 363164 696249 363198
rect 696203 363130 696223 363164
rect 696227 363130 696245 363164
rect 696203 363096 696249 363130
rect 696203 363062 696223 363096
rect 696227 363062 696245 363096
rect 699322 363064 700322 363097
rect 700922 363064 701922 363097
rect 696203 363028 696249 363062
rect 707610 363044 708610 363048
rect 709211 363044 710211 363048
rect 691275 362975 691875 363025
rect 692485 362994 692505 363028
rect 692509 362994 692517 363028
rect 692485 362960 692521 362994
rect 692485 362926 692505 362960
rect 692509 362926 692517 362960
rect 692485 362892 692521 362926
rect 691275 362825 691875 362875
rect 692485 362858 692505 362892
rect 692509 362858 692517 362892
rect 692583 362876 693983 363004
rect 694719 362876 696119 363004
rect 696203 362994 696223 363028
rect 696227 362994 696245 363028
rect 707574 362994 708646 363030
rect 696203 362960 696249 362994
rect 696203 362926 696223 362960
rect 696227 362926 696245 362960
rect 707574 362953 707610 362994
rect 708610 362953 708646 362994
rect 696203 362892 696249 362926
rect 697284 362894 697350 362910
rect 707574 362897 708646 362953
rect 696203 362858 696223 362892
rect 696227 362858 696245 362892
rect 699322 362877 700322 362894
rect 700922 362877 701922 362894
rect 707574 362881 707610 362897
rect 708610 362881 708646 362897
rect 692485 362824 692521 362858
rect 692485 362790 692505 362824
rect 692509 362790 692517 362824
rect 692485 362756 692521 362790
rect 691275 362703 691875 362753
rect 692485 362722 692505 362756
rect 692509 362722 692517 362756
rect 692485 362688 692521 362722
rect 692583 362713 693983 362841
rect 694719 362713 696119 362841
rect 696203 362824 696249 362858
rect 707574 362825 708646 362881
rect 696203 362790 696223 362824
rect 696227 362790 696245 362824
rect 696203 362756 696249 362790
rect 696203 362722 696223 362756
rect 696227 362722 696245 362756
rect 699322 362739 700322 362811
rect 700922 362739 701922 362811
rect 707574 362788 707610 362825
rect 708610 362788 708646 362825
rect 707574 362748 708646 362788
rect 709175 362994 710247 363030
rect 709175 362953 709211 362994
rect 710211 362953 710247 362994
rect 709175 362897 710247 362953
rect 709175 362881 709211 362897
rect 710211 362881 710247 362897
rect 709175 362825 710247 362881
rect 709175 362788 709211 362825
rect 710211 362788 710247 362825
rect 709175 362748 710247 362788
rect 696203 362688 696249 362722
rect 692485 362654 692505 362688
rect 692509 362654 692517 362688
rect 692485 362620 692521 362654
rect 687155 362576 687170 362591
rect 687340 362580 687355 362591
rect 687343 362576 687355 362580
rect 685542 362506 686142 362556
rect 691275 362553 691875 362603
rect 692485 362586 692505 362620
rect 692509 362586 692517 362620
rect 692485 362552 692521 362586
rect 692485 362518 692505 362552
rect 692509 362518 692517 362552
rect 692583 362550 693983 362678
rect 694719 362550 696119 362678
rect 696203 362654 696223 362688
rect 696227 362654 696245 362688
rect 696203 362620 696249 362654
rect 696203 362586 696223 362620
rect 696227 362586 696245 362620
rect 696203 362552 696249 362586
rect 696203 362518 696223 362552
rect 696227 362518 696245 362552
rect 692485 362484 692521 362518
rect 692485 362450 692505 362484
rect 692509 362450 692517 362484
rect 692485 362416 692521 362450
rect 679817 362330 679841 362354
rect 685542 362330 686142 362386
rect 692485 362382 692505 362416
rect 692509 362382 692517 362416
rect 692583 362387 693983 362515
rect 694719 362387 696119 362515
rect 696203 362484 696249 362518
rect 696203 362450 696223 362484
rect 696227 362450 696245 362484
rect 699322 362478 700322 362550
rect 700922 362478 701922 362550
rect 707610 362523 708610 362595
rect 709211 362523 710211 362595
rect 699392 362467 699426 362478
rect 699460 362467 699494 362478
rect 699528 362467 699562 362478
rect 699596 362467 699630 362478
rect 699664 362467 699698 362478
rect 699732 362467 699766 362478
rect 699800 362467 699834 362478
rect 699868 362467 699902 362478
rect 699936 362467 699970 362478
rect 700004 362467 700038 362478
rect 700072 362467 700106 362478
rect 700140 362467 700174 362478
rect 700208 362467 700242 362478
rect 700276 362467 700310 362478
rect 700934 362467 700968 362478
rect 701002 362467 701036 362478
rect 701070 362467 701104 362478
rect 701138 362467 701172 362478
rect 701206 362467 701240 362478
rect 701274 362467 701308 362478
rect 701342 362467 701376 362478
rect 701410 362467 701444 362478
rect 701478 362467 701512 362478
rect 701546 362467 701580 362478
rect 701614 362467 701648 362478
rect 701682 362467 701716 362478
rect 701750 362467 701784 362478
rect 701818 362467 701852 362478
rect 699392 362457 699450 362467
rect 699460 362457 699518 362467
rect 699528 362457 699586 362467
rect 699596 362457 699654 362467
rect 699664 362457 699722 362467
rect 699732 362457 699790 362467
rect 699800 362457 699858 362467
rect 699868 362457 699926 362467
rect 699936 362457 699994 362467
rect 700004 362457 700062 362467
rect 700072 362457 700130 362467
rect 700140 362457 700198 362467
rect 700208 362457 700266 362467
rect 700276 362457 700334 362467
rect 700934 362457 700992 362467
rect 701002 362457 701060 362467
rect 701070 362457 701128 362467
rect 701138 362457 701196 362467
rect 701206 362457 701264 362467
rect 701274 362457 701332 362467
rect 701342 362457 701400 362467
rect 701410 362457 701468 362467
rect 701478 362457 701536 362467
rect 701546 362457 701604 362467
rect 701614 362457 701672 362467
rect 701682 362457 701740 362467
rect 701750 362457 701808 362467
rect 701818 362457 701876 362467
rect 696203 362416 696249 362450
rect 699368 362433 700334 362457
rect 700910 362433 701876 362457
rect 699392 362418 699416 362433
rect 699460 362418 699484 362433
rect 699528 362418 699552 362433
rect 699596 362418 699620 362433
rect 699664 362418 699688 362433
rect 699732 362418 699756 362433
rect 699800 362418 699824 362433
rect 699868 362418 699892 362433
rect 699936 362418 699960 362433
rect 700004 362418 700028 362433
rect 700072 362418 700096 362433
rect 700140 362418 700164 362433
rect 700208 362418 700232 362433
rect 700276 362418 700300 362433
rect 700934 362418 700958 362433
rect 701002 362418 701026 362433
rect 701070 362418 701094 362433
rect 701138 362418 701162 362433
rect 701206 362418 701230 362433
rect 701274 362418 701298 362433
rect 701342 362418 701366 362433
rect 701410 362418 701434 362433
rect 701478 362418 701502 362433
rect 701546 362418 701570 362433
rect 701614 362418 701638 362433
rect 701682 362418 701706 362433
rect 701750 362418 701774 362433
rect 701818 362418 701842 362433
rect 696203 362382 696223 362416
rect 696227 362382 696245 362416
rect 692485 362348 692521 362382
rect 696203 362348 696249 362382
rect 679549 362307 679573 362330
rect 679793 362306 679808 362330
rect 692485 362314 692505 362348
rect 692509 362314 692517 362348
rect 696203 362314 696223 362348
rect 696227 362314 696245 362348
rect 692485 362280 692521 362314
rect 696203 362280 696249 362314
rect 679549 362237 679573 362271
rect 692485 362246 692505 362280
rect 692509 362246 692517 362280
rect 692485 362212 692521 362246
rect 692583 362237 693983 362280
rect 694719 362237 696119 362280
rect 696203 362246 696223 362280
rect 696227 362246 696245 362280
rect 699322 362263 700322 362418
rect 696203 362212 696249 362246
rect 699322 362229 700334 362263
rect 700922 362253 701922 362418
rect 700910 362229 701922 362253
rect 699322 362218 700322 362229
rect 700922 362218 701922 362229
rect 707574 362263 708646 362299
rect 707574 362226 707610 362263
rect 708610 362226 708646 362263
rect 679549 362167 679573 362201
rect 685542 362160 686142 362210
rect 685601 362157 685895 362160
rect 685920 362157 686142 362160
rect 692485 362178 692505 362212
rect 692509 362178 692517 362212
rect 696203 362178 696223 362212
rect 696227 362178 696245 362212
rect 699392 362205 699416 362218
rect 699460 362205 699484 362218
rect 699528 362205 699552 362218
rect 699596 362205 699620 362218
rect 699664 362205 699688 362218
rect 699732 362205 699756 362218
rect 699800 362205 699824 362218
rect 699868 362205 699892 362218
rect 699936 362205 699960 362218
rect 700004 362205 700028 362218
rect 700072 362205 700096 362218
rect 700140 362205 700164 362218
rect 700208 362205 700232 362218
rect 700276 362205 700300 362218
rect 700934 362205 700958 362218
rect 701002 362205 701026 362218
rect 701070 362205 701094 362218
rect 701138 362205 701162 362218
rect 701206 362205 701230 362218
rect 701274 362205 701298 362218
rect 701342 362205 701366 362218
rect 701410 362205 701434 362218
rect 701478 362205 701502 362218
rect 701546 362205 701570 362218
rect 701614 362205 701638 362218
rect 701682 362205 701706 362218
rect 701750 362205 701774 362218
rect 701818 362205 701842 362218
rect 707574 362186 708646 362226
rect 709175 362263 710247 362299
rect 709175 362226 709211 362263
rect 710211 362226 710247 362263
rect 709175 362186 710247 362226
rect 692485 362144 692521 362178
rect 696203 362144 696249 362178
rect 679549 362097 679573 362131
rect 692485 362110 692505 362144
rect 692509 362110 692517 362144
rect 692485 362076 692521 362110
rect 692583 362101 693983 362144
rect 694719 362101 696119 362144
rect 696203 362110 696223 362144
rect 696227 362110 696245 362144
rect 696203 362076 696249 362110
rect 679549 362027 679573 362061
rect 692485 362042 692505 362076
rect 692509 362042 692517 362076
rect 692485 362008 692521 362042
rect 679549 361957 679573 361991
rect 692485 361974 692505 362008
rect 692509 361974 692517 362008
rect 679793 361933 679808 361957
rect 692485 361940 692521 361974
rect 679817 361909 679841 361933
rect 692485 361906 692505 361940
rect 692509 361906 692517 361940
rect 692583 361938 693983 362066
rect 694719 361938 696119 362066
rect 696203 362042 696223 362076
rect 696227 362042 696245 362076
rect 696203 362008 696249 362042
rect 696203 361974 696223 362008
rect 696227 361974 696245 362008
rect 696203 361940 696249 361974
rect 696203 361906 696223 361940
rect 696227 361906 696245 361940
rect 687685 361838 687709 361862
rect 687661 361814 687675 361838
rect 687669 361797 687675 361814
rect 679515 361762 679539 361785
rect 679613 361762 679637 361785
rect 679491 361737 679515 361761
rect 679637 361737 679661 361761
rect 680215 361678 680815 361728
rect 680215 361502 680815 361558
rect 685551 361516 686551 361566
rect 680215 361326 680815 361382
rect 685551 361360 686551 361488
rect 689154 361439 689204 361897
rect 689151 361355 689204 361439
rect 680215 361156 680815 361206
rect 685551 361204 686551 361332
rect 685551 361048 686551 361176
rect 686865 361116 687465 361166
rect 679007 360980 679607 361030
rect 680615 360885 680630 360900
rect 680803 360896 680815 360900
rect 680800 360885 680815 360896
rect 685551 360892 686551 360948
rect 686865 360940 687465 361068
rect 679007 360810 679607 360860
rect 680615 360705 680815 360885
rect 683328 360793 683928 360843
rect 682573 360717 683173 360767
rect 680615 360690 680630 360705
rect 680800 360694 680815 360705
rect 680803 360690 680815 360694
rect 680502 360649 680517 360664
rect 680480 360469 680517 360649
rect 680502 360454 680517 360469
rect 680615 360649 680630 360664
rect 680803 360660 680815 360664
rect 680800 360649 680815 360660
rect 680615 360469 680815 360649
rect 682573 360541 683173 360669
rect 683328 360617 683928 360745
rect 685551 360736 686551 360864
rect 686865 360764 687465 360820
rect 685551 360580 686551 360708
rect 686865 360588 687465 360716
rect 680615 360454 680630 360469
rect 680800 360458 680815 360469
rect 680803 360454 680815 360458
rect 683328 360441 683928 360497
rect 679002 360384 679602 360434
rect 685551 360424 686551 360552
rect 682573 360365 683173 360421
rect 686865 360412 687465 360468
rect 679002 360208 679602 360264
rect 682573 360189 683173 360317
rect 683328 360265 683928 360321
rect 685551 360274 686551 360324
rect 686865 360236 687465 360364
rect 685551 360158 686551 360208
rect 678680 360123 678704 360157
rect 678680 360055 678704 360089
rect 679002 360038 679602 360088
rect 679061 360035 679355 360038
rect 679380 360035 679602 360038
rect 678680 359987 678704 360021
rect 682573 360013 683173 360141
rect 683328 360089 683928 360145
rect 678680 359919 678704 359953
rect 678680 359851 678704 359885
rect 682573 359837 683173 359965
rect 683328 359913 683928 360041
rect 685551 359982 686551 360110
rect 686865 360060 687465 360116
rect 678680 359783 678704 359817
rect 685551 359806 686551 359934
rect 686865 359884 687465 360012
rect 678680 359715 678704 359749
rect 678680 359647 678704 359681
rect 682573 359661 683173 359789
rect 683328 359737 683928 359793
rect 685551 359630 686551 359758
rect 686865 359708 687465 359836
rect 678680 359579 678704 359613
rect 683328 359567 683928 359617
rect 678680 359511 678704 359545
rect 682573 359491 683173 359541
rect 684519 359498 685119 359548
rect 678680 359443 678704 359477
rect 685551 359454 686551 359582
rect 686865 359532 687465 359660
rect 679133 359409 679283 359421
rect 679452 359409 679602 359421
rect 678680 359375 678704 359409
rect 678680 359307 678704 359341
rect 679002 359296 679602 359346
rect 684519 359342 685119 359398
rect 685551 359278 686551 359406
rect 686865 359356 687465 359484
rect 678680 359239 678704 359273
rect 678680 359171 678704 359205
rect 684519 359192 685119 359242
rect 678680 359103 678704 359137
rect 679002 359120 679602 359176
rect 681745 359081 682345 359131
rect 682509 359069 683109 359119
rect 678680 359035 678704 359069
rect 683739 359027 684339 359077
rect 684519 359062 685119 359112
rect 685551 359102 686551 359230
rect 686865 359180 687465 359308
rect 678680 358967 678704 359001
rect 679002 358950 679602 359000
rect 678680 358899 678704 358933
rect 680502 358915 680517 358930
rect 678680 358831 678704 358865
rect 678680 358763 678704 358797
rect 680480 358735 680517 358915
rect 678680 358695 678704 358729
rect 680502 358720 680517 358735
rect 680615 358915 680630 358930
rect 680803 358926 680815 358930
rect 680800 358915 680815 358926
rect 681745 358925 682345 358981
rect 680615 358735 680815 358915
rect 681745 358769 682345 358897
rect 682509 358893 683109 359021
rect 684519 358906 685119 359034
rect 685551 358926 686551 359054
rect 686865 359004 687465 359060
rect 683739 358837 684339 358893
rect 686865 358828 687465 358956
rect 680615 358720 680630 358735
rect 680800 358724 680815 358735
rect 680803 358720 680815 358724
rect 680615 358679 680630 358694
rect 680803 358690 680815 358694
rect 680800 358679 680815 358690
rect 678680 358627 678704 358661
rect 678680 358559 678704 358593
rect 678680 358491 678704 358525
rect 679007 358524 679607 358574
rect 680615 358499 680815 358679
rect 681745 358613 682345 358741
rect 682509 358717 683109 358773
rect 684519 358750 685119 358806
rect 685551 358750 686551 358806
rect 682509 358541 683109 358669
rect 684519 358594 685119 358722
rect 685551 358594 686551 358722
rect 686865 358652 687465 358780
rect 680615 358484 680630 358499
rect 680800 358488 680815 358499
rect 680803 358484 680815 358488
rect 681745 358463 682345 358513
rect 683739 358477 684339 358513
rect 678680 358423 678704 358457
rect 684519 358444 685119 358494
rect 685551 358438 686551 358566
rect 686865 358476 687465 358604
rect 678680 358355 678704 358389
rect 679007 358354 679607 358404
rect 682509 358371 683109 358421
rect 678680 358287 678704 358321
rect 684519 358314 685119 358364
rect 678680 358219 678704 358253
rect 678680 358151 678704 358185
rect 680215 358178 680815 358228
rect 681745 358209 682345 358259
rect 678680 358083 678704 358117
rect 678680 358015 678704 358049
rect 680215 358002 680815 358058
rect 681745 358053 682345 358181
rect 682509 358030 683109 358080
rect 678680 357947 678704 357981
rect 678680 357879 678704 357913
rect 681745 357897 682345 357953
rect 678680 357811 678704 357845
rect 680215 357826 680815 357882
rect 678680 357743 678704 357777
rect 681745 357741 682345 357869
rect 682509 357854 683109 357910
rect 678680 357675 678704 357709
rect 680215 357656 680815 357706
rect 682509 357684 683109 357734
rect 683248 357680 683298 358268
rect 683398 357680 683448 358268
rect 684519 358158 685119 358286
rect 685551 358282 686551 358410
rect 686865 358300 687465 358428
rect 684519 358002 685119 358130
rect 685551 358126 686551 358254
rect 686865 358124 687465 358252
rect 685551 357970 686551 358098
rect 686865 357954 687465 358004
rect 684519 357852 685119 357902
rect 685551 357814 686551 357870
rect 686865 357838 687465 357888
rect 683248 357668 683448 357680
rect 685551 357658 686551 357786
rect 686865 357662 687465 357790
rect 678680 357607 678704 357641
rect 681745 357591 682345 357641
rect 683571 357605 683581 357646
rect 678680 357539 678704 357573
rect 680215 357524 680815 357574
rect 682509 357555 683509 357605
rect 678680 357471 678704 357505
rect 685551 357502 686551 357630
rect 686865 357486 687465 357542
rect 678680 357403 678704 357437
rect 678680 357335 678704 357369
rect 680215 357348 680815 357404
rect 681745 357389 682345 357439
rect 682509 357385 683509 357435
rect 683278 357382 683398 357385
rect 683571 357382 683581 357385
rect 685551 357346 686551 357474
rect 678680 357267 678704 357301
rect 678680 357199 678704 357233
rect 680215 357172 680815 357228
rect 681745 357213 682345 357341
rect 682509 357247 683109 357297
rect 678680 357131 678704 357165
rect 678680 357063 678704 357097
rect 678654 357013 678680 357039
rect 680215 357002 680815 357052
rect 681745 357037 682345 357093
rect 682509 357071 683109 357127
rect 678680 356929 678704 356963
rect 678680 356861 678704 356895
rect 678680 356793 678704 356827
rect 679007 356826 679607 356876
rect 681745 356867 682345 356917
rect 682509 356901 683109 356951
rect 678680 356725 678704 356759
rect 680615 356731 680630 356746
rect 680803 356742 680815 356746
rect 680800 356731 680815 356742
rect 678680 356657 678704 356691
rect 679007 356656 679607 356706
rect 678680 356589 678704 356623
rect 678680 356521 678704 356555
rect 680615 356551 680815 356731
rect 681345 356651 682345 356701
rect 682508 356631 683108 356681
rect 680615 356536 680630 356551
rect 680800 356540 680815 356551
rect 680803 356536 680815 356540
rect 680502 356495 680517 356510
rect 678680 356453 678704 356487
rect 678680 356385 678704 356419
rect 678680 356317 678704 356351
rect 680480 356315 680517 356495
rect 680502 356300 680517 356315
rect 680615 356495 680630 356510
rect 680803 356506 680815 356510
rect 680800 356495 680815 356506
rect 680615 356315 680815 356495
rect 681345 356475 682345 356531
rect 682508 356455 683108 356511
rect 680615 356300 680630 356315
rect 680800 356304 680815 356315
rect 680803 356300 680815 356304
rect 681345 356299 682345 356427
rect 682508 356285 683108 356335
rect 683228 356322 683278 357322
rect 683398 356322 683448 357322
rect 685551 357190 686551 357318
rect 686865 357310 687465 357438
rect 685551 357034 686551 357162
rect 686865 357140 687465 357190
rect 686865 357024 687465 357074
rect 685551 356884 686551 356934
rect 686865 356848 687465 356976
rect 685551 356768 686551 356818
rect 686865 356672 687465 356800
rect 684404 356609 685004 356659
rect 685551 356612 686551 356668
rect 685551 356456 686551 356512
rect 686865 356496 687465 356624
rect 685551 356300 686551 356356
rect 686865 356320 687465 356376
rect 678680 356249 678704 356283
rect 679002 356230 679602 356280
rect 678680 356181 678704 356215
rect 678680 356113 678704 356147
rect 681345 356129 682345 356179
rect 684404 356175 685004 356225
rect 685551 356150 686551 356200
rect 686865 356150 687465 356200
rect 678680 356045 678704 356079
rect 679002 356054 679602 356110
rect 681390 356070 681424 356080
rect 681458 356070 681492 356080
rect 681526 356070 681560 356080
rect 681594 356070 681628 356080
rect 681662 356070 681696 356080
rect 681730 356070 681764 356080
rect 681798 356070 681832 356080
rect 681866 356070 681900 356080
rect 681934 356070 681968 356080
rect 682002 356070 682036 356080
rect 682077 356070 682111 356080
rect 682145 356070 682179 356080
rect 682213 356070 682247 356080
rect 682281 356070 682315 356080
rect 681345 356034 682345 356046
rect 678680 355977 678704 356011
rect 678680 355909 678704 355943
rect 679002 355884 679602 355934
rect 681345 355927 682345 355977
rect 684004 355973 685004 356023
rect 685551 356014 686551 356064
rect 686865 356034 687465 356084
rect 679061 355881 679355 355884
rect 679380 355881 679602 355884
rect 678680 355841 678704 355875
rect 678680 355773 678704 355807
rect 681345 355751 682345 355879
rect 684004 355817 685004 355873
rect 685551 355858 686551 355914
rect 686865 355858 687465 355914
rect 686686 355812 686714 355840
rect 678680 355705 678704 355739
rect 678680 355637 678704 355671
rect 678680 355569 678704 355603
rect 681345 355575 682345 355703
rect 684004 355661 685004 355789
rect 685551 355708 686551 355758
rect 686865 355688 687465 355738
rect 678680 355501 678704 355535
rect 684004 355505 685004 355633
rect 687573 355554 687585 361277
rect 689154 361107 689204 361355
rect 689151 361023 689204 361107
rect 689154 360897 689204 361023
rect 689304 360897 689360 361897
rect 689460 360897 689516 361897
rect 689616 360897 689672 361897
rect 689772 360897 689828 361897
rect 689928 360897 689978 361897
rect 692485 361872 692521 361906
rect 692485 361838 692505 361872
rect 692509 361838 692517 361872
rect 690952 361509 691122 361815
rect 692485 361804 692521 361838
rect 692485 361770 692505 361804
rect 692509 361770 692517 361804
rect 692583 361775 693983 361903
rect 694719 361775 696119 361903
rect 696203 361872 696249 361906
rect 696203 361838 696223 361872
rect 696227 361838 696245 361872
rect 699322 361860 700322 361916
rect 700922 361860 701922 361916
rect 707610 361905 708610 361961
rect 709211 361905 710211 361961
rect 696203 361804 696249 361838
rect 696203 361770 696223 361804
rect 696227 361770 696245 361804
rect 699322 361788 700322 361844
rect 700922 361788 701922 361844
rect 707610 361833 708610 361889
rect 709211 361833 710211 361889
rect 692485 361736 692521 361770
rect 692485 361702 692505 361736
rect 692509 361702 692517 361736
rect 692485 361668 692521 361702
rect 692485 361634 692505 361668
rect 692509 361634 692517 361668
rect 692485 361600 692521 361634
rect 692583 361612 693983 361740
rect 694719 361612 696119 361740
rect 696203 361736 696249 361770
rect 696203 361702 696223 361736
rect 696227 361702 696245 361736
rect 696203 361668 696249 361702
rect 696203 361634 696223 361668
rect 696227 361634 696245 361668
rect 696203 361600 696249 361634
rect 692485 361566 692505 361600
rect 692509 361566 692517 361600
rect 692485 361532 692521 361566
rect 692485 361498 692505 361532
rect 692509 361498 692517 361532
rect 692485 361464 692521 361498
rect 692485 361430 692505 361464
rect 692509 361430 692517 361464
rect 692583 361449 693983 361577
rect 694719 361449 696119 361577
rect 696203 361566 696223 361600
rect 696227 361566 696245 361600
rect 696203 361532 696249 361566
rect 696203 361498 696223 361532
rect 696227 361498 696245 361532
rect 696203 361464 696249 361498
rect 699322 361486 700322 361558
rect 700922 361486 701922 361558
rect 707610 361531 708610 361603
rect 709211 361531 710211 361603
rect 711579 361553 711605 363307
rect 715956 362297 716006 363297
rect 716106 362297 716234 363297
rect 716262 362297 716312 363297
rect 699392 361475 699426 361486
rect 699460 361475 699494 361486
rect 699528 361475 699562 361486
rect 699596 361475 699630 361486
rect 699664 361475 699698 361486
rect 699732 361475 699766 361486
rect 699800 361475 699834 361486
rect 699868 361475 699902 361486
rect 699936 361475 699970 361486
rect 700004 361475 700038 361486
rect 700072 361475 700106 361486
rect 700140 361475 700174 361486
rect 700208 361475 700242 361486
rect 700276 361475 700310 361486
rect 700934 361475 700968 361486
rect 701002 361475 701036 361486
rect 701070 361475 701104 361486
rect 701138 361475 701172 361486
rect 701206 361475 701240 361486
rect 701274 361475 701308 361486
rect 701342 361475 701376 361486
rect 701410 361475 701444 361486
rect 701478 361475 701512 361486
rect 701546 361475 701580 361486
rect 701614 361475 701648 361486
rect 701682 361475 701716 361486
rect 701750 361475 701784 361486
rect 701818 361475 701852 361486
rect 711511 361485 711663 361553
rect 712447 361501 712557 361511
rect 711579 361482 711663 361485
rect 699392 361465 699450 361475
rect 699460 361465 699518 361475
rect 699528 361465 699586 361475
rect 699596 361465 699654 361475
rect 699664 361465 699722 361475
rect 699732 361465 699790 361475
rect 699800 361465 699858 361475
rect 699868 361465 699926 361475
rect 699936 361465 699994 361475
rect 700004 361465 700062 361475
rect 700072 361465 700130 361475
rect 700140 361465 700198 361475
rect 700208 361465 700266 361475
rect 700276 361465 700334 361475
rect 700934 361465 700992 361475
rect 701002 361465 701060 361475
rect 701070 361465 701128 361475
rect 701138 361465 701196 361475
rect 701206 361465 701264 361475
rect 701274 361465 701332 361475
rect 701342 361465 701400 361475
rect 701410 361465 701468 361475
rect 701478 361465 701536 361475
rect 701546 361465 701604 361475
rect 701614 361465 701672 361475
rect 701682 361465 701740 361475
rect 701750 361465 701808 361475
rect 701818 361465 701876 361475
rect 696203 361430 696223 361464
rect 696227 361430 696245 361464
rect 699368 361441 700334 361465
rect 700910 361441 701876 361465
rect 711541 361461 711633 361482
rect 692485 361396 692521 361430
rect 692485 361362 692505 361396
rect 692509 361362 692517 361396
rect 692485 361328 692521 361362
rect 692485 361294 692505 361328
rect 692509 361294 692517 361328
rect 692485 361260 692521 361294
rect 692583 361286 693983 361414
rect 694719 361286 696119 361414
rect 696203 361396 696249 361430
rect 699392 361426 699416 361441
rect 699460 361426 699484 361441
rect 699528 361426 699552 361441
rect 699596 361426 699620 361441
rect 699664 361426 699688 361441
rect 699732 361426 699756 361441
rect 699800 361426 699824 361441
rect 699868 361426 699892 361441
rect 699936 361426 699960 361441
rect 700004 361426 700028 361441
rect 700072 361426 700096 361441
rect 700140 361426 700164 361441
rect 700208 361426 700232 361441
rect 700276 361426 700300 361441
rect 700934 361426 700958 361441
rect 701002 361426 701026 361441
rect 701070 361426 701094 361441
rect 701138 361426 701162 361441
rect 701206 361426 701230 361441
rect 701274 361426 701298 361441
rect 701342 361426 701366 361441
rect 701410 361426 701434 361441
rect 701478 361426 701502 361441
rect 701546 361426 701570 361441
rect 701614 361426 701638 361441
rect 701682 361426 701706 361441
rect 701750 361426 701774 361441
rect 701818 361426 701842 361441
rect 696203 361362 696223 361396
rect 696227 361362 696245 361396
rect 696203 361328 696249 361362
rect 696203 361294 696223 361328
rect 696227 361294 696245 361328
rect 696203 361260 696249 361294
rect 699322 361271 700322 361426
rect 692485 361226 692505 361260
rect 692509 361226 692517 361260
rect 692485 361192 692521 361226
rect 692485 361158 692505 361192
rect 692509 361158 692517 361192
rect 692485 361124 692521 361158
rect 692485 361090 692505 361124
rect 692509 361090 692517 361124
rect 692583 361123 693983 361251
rect 694719 361123 696119 361251
rect 696203 361226 696223 361260
rect 696227 361226 696245 361260
rect 699322 361237 700334 361271
rect 700922 361261 701922 361426
rect 707610 361271 708610 361331
rect 709211 361271 710211 361331
rect 700910 361237 701922 361261
rect 699322 361226 700322 361237
rect 700922 361226 701922 361237
rect 696203 361192 696249 361226
rect 699392 361213 699416 361226
rect 699460 361213 699484 361226
rect 699528 361213 699552 361226
rect 699596 361213 699620 361226
rect 699664 361213 699688 361226
rect 699732 361213 699756 361226
rect 699800 361213 699824 361226
rect 699868 361213 699892 361226
rect 699936 361213 699960 361226
rect 700004 361213 700028 361226
rect 700072 361213 700096 361226
rect 700140 361213 700164 361226
rect 700208 361213 700232 361226
rect 700276 361213 700300 361226
rect 700934 361213 700958 361226
rect 701002 361213 701026 361226
rect 701070 361213 701094 361226
rect 701138 361213 701162 361226
rect 701206 361213 701230 361226
rect 701274 361213 701298 361226
rect 701342 361213 701366 361226
rect 701410 361213 701434 361226
rect 701478 361213 701502 361226
rect 701546 361213 701570 361226
rect 701614 361213 701638 361226
rect 701682 361213 701706 361226
rect 701750 361213 701774 361226
rect 701818 361213 701842 361226
rect 696203 361158 696223 361192
rect 696227 361158 696245 361192
rect 696203 361124 696249 361158
rect 696203 361090 696223 361124
rect 696227 361090 696245 361124
rect 692485 361056 692521 361090
rect 696203 361056 696249 361090
rect 692485 361022 692505 361056
rect 692509 361022 692517 361056
rect 696203 361022 696223 361056
rect 696227 361022 696245 361056
rect 692485 360988 692521 361022
rect 692485 360954 692505 360988
rect 692509 360954 692517 360988
rect 692583 360966 693983 361016
rect 694719 360966 696119 361016
rect 696203 360988 696249 361022
rect 696203 360954 696223 360988
rect 696227 360954 696245 360988
rect 692485 360920 692521 360954
rect 696203 360920 696249 360954
rect 692485 360896 692505 360920
rect 692487 360852 692505 360896
rect 692509 360886 692517 360920
rect 696203 360896 696223 360920
rect 696215 360886 696223 360896
rect 696227 360852 696245 360920
rect 697284 360870 697350 360886
rect 699322 360868 700322 360924
rect 700922 360868 701922 360924
rect 707610 360913 708610 360969
rect 709211 360913 710211 360969
rect 692174 360787 692186 360811
rect 692288 360787 692312 360811
rect 696390 360787 696414 360811
rect 696516 360787 696528 360811
rect 699322 360796 700322 360852
rect 700922 360796 701922 360852
rect 707610 360841 708610 360897
rect 709211 360841 710211 360897
rect 692264 360763 692288 360777
rect 696414 360763 696438 360777
rect 692288 360729 692312 360753
rect 696390 360729 696414 360753
rect 688940 360475 688990 360675
rect 689110 360475 689238 360675
rect 689286 360475 689342 360675
rect 689462 360475 689590 360675
rect 689638 360559 689688 360675
rect 692736 360597 695966 360699
rect 689638 360475 689691 360559
rect 699322 360494 700322 360566
rect 700922 360494 701922 360566
rect 707610 360539 708610 360611
rect 709211 360539 710211 360611
rect 699392 360483 699426 360494
rect 699460 360483 699494 360494
rect 699528 360483 699562 360494
rect 699596 360483 699630 360494
rect 699664 360483 699698 360494
rect 699732 360483 699766 360494
rect 699800 360483 699834 360494
rect 699868 360483 699902 360494
rect 699936 360483 699970 360494
rect 700004 360483 700038 360494
rect 700072 360483 700106 360494
rect 700140 360483 700174 360494
rect 700208 360483 700242 360494
rect 700276 360483 700310 360494
rect 700934 360483 700968 360494
rect 701002 360483 701036 360494
rect 701070 360483 701104 360494
rect 701138 360483 701172 360494
rect 701206 360483 701240 360494
rect 701274 360483 701308 360494
rect 701342 360483 701376 360494
rect 701410 360483 701444 360494
rect 701478 360483 701512 360494
rect 701546 360483 701580 360494
rect 701614 360483 701648 360494
rect 701682 360483 701716 360494
rect 701750 360483 701784 360494
rect 701818 360483 701852 360494
rect 689649 360471 689683 360475
rect 699392 360473 699450 360483
rect 699460 360473 699518 360483
rect 699528 360473 699586 360483
rect 699596 360473 699654 360483
rect 699664 360473 699722 360483
rect 699732 360473 699790 360483
rect 699800 360473 699858 360483
rect 699868 360473 699926 360483
rect 699936 360473 699994 360483
rect 700004 360473 700062 360483
rect 700072 360473 700130 360483
rect 700140 360473 700198 360483
rect 700208 360473 700266 360483
rect 700276 360473 700334 360483
rect 700934 360473 700992 360483
rect 701002 360473 701060 360483
rect 701070 360473 701128 360483
rect 701138 360473 701196 360483
rect 701206 360473 701264 360483
rect 701274 360473 701332 360483
rect 701342 360473 701400 360483
rect 701410 360473 701468 360483
rect 701478 360473 701536 360483
rect 701546 360473 701604 360483
rect 701614 360473 701672 360483
rect 701682 360473 701740 360483
rect 701750 360473 701808 360483
rect 701818 360473 701876 360483
rect 692451 360444 692475 360468
rect 692509 360444 692533 360468
rect 696169 360444 696193 360468
rect 696227 360444 696251 360468
rect 699368 360449 700334 360473
rect 700910 360449 701876 360473
rect 692485 360410 692499 360444
rect 696203 360410 696217 360444
rect 699392 360434 699416 360449
rect 699460 360434 699484 360449
rect 699528 360434 699552 360449
rect 699596 360434 699620 360449
rect 699664 360434 699688 360449
rect 699732 360434 699756 360449
rect 699800 360434 699824 360449
rect 699868 360434 699892 360449
rect 699936 360434 699960 360449
rect 700004 360434 700028 360449
rect 700072 360434 700096 360449
rect 700140 360434 700164 360449
rect 700208 360434 700232 360449
rect 700276 360434 700300 360449
rect 700934 360434 700958 360449
rect 701002 360434 701026 360449
rect 701070 360434 701094 360449
rect 701138 360434 701162 360449
rect 701206 360434 701230 360449
rect 701274 360434 701298 360449
rect 701342 360434 701366 360449
rect 701410 360434 701434 360449
rect 701478 360434 701502 360449
rect 701546 360434 701570 360449
rect 701614 360434 701638 360449
rect 701682 360434 701706 360449
rect 701750 360434 701774 360449
rect 701818 360434 701842 360449
rect 692451 360386 692475 360410
rect 692509 360386 692533 360410
rect 696169 360386 696193 360410
rect 696227 360386 696251 360410
rect 690664 360318 691664 360368
rect 692515 360280 693915 360330
rect 694787 360280 696187 360330
rect 699322 360279 700322 360434
rect 699322 360245 700334 360279
rect 700922 360269 701922 360434
rect 703539 360286 703699 360290
rect 707610 360279 708610 360339
rect 709211 360279 710211 360339
rect 700910 360245 701922 360269
rect 690242 360219 690326 360222
rect 690242 360214 690442 360219
rect 690238 360180 690442 360214
rect 690242 360169 690442 360180
rect 690664 360162 691664 360218
rect 687686 360128 687720 360162
rect 687686 360104 687710 360128
rect 689649 360127 689683 360131
rect 688940 359927 688990 360127
rect 689110 359927 689238 360127
rect 689286 359927 689342 360127
rect 689462 359927 689590 360127
rect 689638 360043 689691 360127
rect 689638 359927 689688 360043
rect 690242 359993 690442 360121
rect 692515 360117 693915 360245
rect 694787 360117 696187 360245
rect 699322 360234 700322 360245
rect 700922 360234 701922 360245
rect 699392 360221 699416 360234
rect 699460 360221 699484 360234
rect 699528 360221 699552 360234
rect 699596 360221 699620 360234
rect 699664 360221 699688 360234
rect 699732 360221 699756 360234
rect 699800 360221 699824 360234
rect 699868 360221 699892 360234
rect 699936 360221 699960 360234
rect 700004 360221 700028 360234
rect 700072 360221 700096 360234
rect 700140 360221 700164 360234
rect 700208 360221 700232 360234
rect 700276 360221 700300 360234
rect 700934 360221 700958 360234
rect 701002 360221 701026 360234
rect 701070 360221 701094 360234
rect 701138 360221 701162 360234
rect 701206 360221 701230 360234
rect 701274 360221 701298 360234
rect 701342 360221 701366 360234
rect 701410 360221 701434 360234
rect 701478 360221 701502 360234
rect 701546 360221 701570 360234
rect 701614 360221 701638 360234
rect 701682 360221 701706 360234
rect 701750 360221 701774 360234
rect 701818 360221 701842 360234
rect 703541 360140 703701 360144
rect 690664 360006 691664 360062
rect 692515 359954 693915 360082
rect 694787 359954 696187 360082
rect 690242 359817 690442 359873
rect 690664 359850 691664 359906
rect 692515 359791 693915 359919
rect 694787 359791 696187 359919
rect 699322 359876 700322 359932
rect 700922 359876 701922 359932
rect 707610 359921 708610 359977
rect 709211 359921 710211 359977
rect 699322 359804 700322 359860
rect 700922 359804 701922 359860
rect 707610 359849 708610 359905
rect 709211 359849 710211 359905
rect 689154 359579 689204 359705
rect 687686 359501 687720 359535
rect 687798 359515 687822 359539
rect 687774 359491 687798 359504
rect 689151 359495 689204 359579
rect 687798 359456 687822 359480
rect 689154 359247 689204 359495
rect 689151 359163 689204 359247
rect 689154 358705 689204 359163
rect 689304 358705 689360 359705
rect 689460 358705 689516 359705
rect 689616 358705 689672 359705
rect 689772 358705 689828 359705
rect 689928 358705 689978 359705
rect 690242 359641 690442 359769
rect 690664 359700 691664 359750
rect 690790 359697 690874 359700
rect 691123 359697 691207 359700
rect 692515 359628 693915 359756
rect 694787 359628 696187 359756
rect 704735 359731 705041 359833
rect 704719 359715 705057 359731
rect 690242 359465 690442 359521
rect 692515 359465 693915 359593
rect 694787 359465 696187 359593
rect 699322 359502 700322 359574
rect 700922 359502 701922 359574
rect 707610 359547 708610 359619
rect 709211 359547 710211 359619
rect 699392 359491 699426 359502
rect 699460 359491 699494 359502
rect 699528 359491 699562 359502
rect 699596 359491 699630 359502
rect 699664 359491 699698 359502
rect 699732 359491 699766 359502
rect 699800 359491 699834 359502
rect 699868 359491 699902 359502
rect 699936 359491 699970 359502
rect 700004 359491 700038 359502
rect 700072 359491 700106 359502
rect 700140 359491 700174 359502
rect 700208 359491 700242 359502
rect 700276 359491 700310 359502
rect 700934 359491 700968 359502
rect 701002 359491 701036 359502
rect 701070 359491 701104 359502
rect 701138 359491 701172 359502
rect 701206 359491 701240 359502
rect 701274 359491 701308 359502
rect 701342 359491 701376 359502
rect 701410 359491 701444 359502
rect 701478 359491 701512 359502
rect 701546 359491 701580 359502
rect 701614 359491 701648 359502
rect 701682 359491 701716 359502
rect 701750 359491 701784 359502
rect 701818 359491 701852 359502
rect 699392 359481 699450 359491
rect 699460 359481 699518 359491
rect 699528 359481 699586 359491
rect 699596 359481 699654 359491
rect 699664 359481 699722 359491
rect 699732 359481 699790 359491
rect 699800 359481 699858 359491
rect 699868 359481 699926 359491
rect 699936 359481 699994 359491
rect 700004 359481 700062 359491
rect 700072 359481 700130 359491
rect 700140 359481 700198 359491
rect 700208 359481 700266 359491
rect 700276 359481 700334 359491
rect 700934 359481 700992 359491
rect 701002 359481 701060 359491
rect 701070 359481 701128 359491
rect 701138 359481 701196 359491
rect 701206 359481 701264 359491
rect 701274 359481 701332 359491
rect 701342 359481 701400 359491
rect 701410 359481 701468 359491
rect 701478 359481 701536 359491
rect 701546 359481 701604 359491
rect 701614 359481 701672 359491
rect 701682 359481 701740 359491
rect 701750 359481 701808 359491
rect 701818 359481 701876 359491
rect 699368 359457 700334 359481
rect 700910 359457 701876 359481
rect 699392 359442 699416 359457
rect 699460 359442 699484 359457
rect 699528 359442 699552 359457
rect 699596 359442 699620 359457
rect 699664 359442 699688 359457
rect 699732 359442 699756 359457
rect 699800 359442 699824 359457
rect 699868 359442 699892 359457
rect 699936 359442 699960 359457
rect 700004 359442 700028 359457
rect 700072 359442 700096 359457
rect 700140 359442 700164 359457
rect 700208 359442 700232 359457
rect 700276 359442 700300 359457
rect 700934 359442 700958 359457
rect 701002 359442 701026 359457
rect 701070 359442 701094 359457
rect 701138 359442 701162 359457
rect 701206 359442 701230 359457
rect 701274 359442 701298 359457
rect 701342 359442 701366 359457
rect 701410 359442 701434 359457
rect 701478 359442 701502 359457
rect 701546 359442 701570 359457
rect 701614 359442 701638 359457
rect 701682 359442 701706 359457
rect 701750 359442 701774 359457
rect 701818 359442 701842 359457
rect 690242 359289 690442 359417
rect 692515 359302 693915 359430
rect 694787 359302 696187 359430
rect 690790 359286 690874 359289
rect 691123 359286 691207 359289
rect 699322 359287 700322 359442
rect 690664 359236 691664 359286
rect 699322 359253 700334 359287
rect 700922 359277 701922 359442
rect 707610 359287 708610 359347
rect 709211 359287 710211 359347
rect 700910 359253 701922 359277
rect 699322 359242 700322 359253
rect 700922 359242 701922 359253
rect 699392 359229 699416 359242
rect 699460 359229 699484 359242
rect 699528 359229 699552 359242
rect 699596 359229 699620 359242
rect 699664 359229 699688 359242
rect 699732 359229 699756 359242
rect 699800 359229 699824 359242
rect 699868 359229 699892 359242
rect 699936 359229 699960 359242
rect 700004 359229 700028 359242
rect 700072 359229 700096 359242
rect 700140 359229 700164 359242
rect 700208 359229 700232 359242
rect 700276 359229 700300 359242
rect 700934 359229 700958 359242
rect 701002 359229 701026 359242
rect 701070 359229 701094 359242
rect 701138 359229 701162 359242
rect 701206 359229 701230 359242
rect 701274 359229 701298 359242
rect 701342 359229 701366 359242
rect 701410 359229 701434 359242
rect 701478 359229 701502 359242
rect 701546 359229 701570 359242
rect 701614 359229 701638 359242
rect 701682 359229 701706 359242
rect 701750 359229 701774 359242
rect 701818 359229 701842 359242
rect 690242 359113 690442 359169
rect 692515 359152 693915 359195
rect 694787 359152 696187 359195
rect 690664 359080 691664 359136
rect 690242 358937 690442 359065
rect 692515 359016 693915 359059
rect 694787 359016 696187 359059
rect 690664 358924 691664 358980
rect 692515 358853 693915 358981
rect 694787 358853 696187 358981
rect 703541 358944 703701 358948
rect 699322 358884 700322 358940
rect 700922 358884 701922 358940
rect 707610 358929 708610 358985
rect 709211 358929 710211 358985
rect 690242 358806 690442 358817
rect 690238 358772 690442 358806
rect 690242 358767 690442 358772
rect 690664 358768 691664 358824
rect 690242 358764 690326 358767
rect 692515 358690 693915 358818
rect 694787 358690 696187 358818
rect 699322 358812 700322 358868
rect 700922 358812 701922 358868
rect 707610 358857 708610 358913
rect 709211 358857 710211 358913
rect 703541 358798 703701 358802
rect 690664 358618 691664 358668
rect 692515 358527 693915 358655
rect 694787 358527 696187 358655
rect 699322 358510 700322 358582
rect 700922 358510 701922 358582
rect 707610 358555 708610 358627
rect 709211 358555 710211 358627
rect 699392 358499 699426 358510
rect 699460 358499 699494 358510
rect 699528 358499 699562 358510
rect 699596 358499 699630 358510
rect 699664 358499 699698 358510
rect 699732 358499 699766 358510
rect 699800 358499 699834 358510
rect 699868 358499 699902 358510
rect 699936 358499 699970 358510
rect 700004 358499 700038 358510
rect 700072 358499 700106 358510
rect 700140 358499 700174 358510
rect 700208 358499 700242 358510
rect 700276 358499 700310 358510
rect 700934 358499 700968 358510
rect 701002 358499 701036 358510
rect 701070 358499 701104 358510
rect 701138 358499 701172 358510
rect 701206 358499 701240 358510
rect 701274 358499 701308 358510
rect 701342 358499 701376 358510
rect 701410 358499 701444 358510
rect 701478 358499 701512 358510
rect 701546 358499 701580 358510
rect 701614 358499 701648 358510
rect 701682 358499 701716 358510
rect 701750 358499 701784 358510
rect 701818 358499 701852 358510
rect 692515 358364 693915 358492
rect 694787 358364 696187 358492
rect 699392 358489 699450 358499
rect 699460 358489 699518 358499
rect 699528 358489 699586 358499
rect 699596 358489 699654 358499
rect 699664 358489 699722 358499
rect 699732 358489 699790 358499
rect 699800 358489 699858 358499
rect 699868 358489 699926 358499
rect 699936 358489 699994 358499
rect 700004 358489 700062 358499
rect 700072 358489 700130 358499
rect 700140 358489 700198 358499
rect 700208 358489 700266 358499
rect 700276 358489 700334 358499
rect 700934 358489 700992 358499
rect 701002 358489 701060 358499
rect 701070 358489 701128 358499
rect 701138 358489 701196 358499
rect 701206 358489 701264 358499
rect 701274 358489 701332 358499
rect 701342 358489 701400 358499
rect 701410 358489 701468 358499
rect 701478 358489 701536 358499
rect 701546 358489 701604 358499
rect 701614 358489 701672 358499
rect 701682 358489 701740 358499
rect 701750 358489 701808 358499
rect 701818 358489 701876 358499
rect 699368 358465 700334 358489
rect 700910 358465 701876 358489
rect 699392 358450 699416 358465
rect 699460 358450 699484 358465
rect 699528 358450 699552 358465
rect 699596 358450 699620 358465
rect 699664 358450 699688 358465
rect 699732 358450 699756 358465
rect 699800 358450 699824 358465
rect 699868 358450 699892 358465
rect 699936 358450 699960 358465
rect 700004 358450 700028 358465
rect 700072 358450 700096 358465
rect 700140 358450 700164 358465
rect 700208 358450 700232 358465
rect 700276 358450 700300 358465
rect 700934 358450 700958 358465
rect 701002 358450 701026 358465
rect 701070 358450 701094 358465
rect 701138 358450 701162 358465
rect 701206 358450 701230 358465
rect 701274 358450 701298 358465
rect 701342 358450 701366 358465
rect 701410 358450 701434 358465
rect 701478 358450 701502 358465
rect 701546 358450 701570 358465
rect 701614 358450 701638 358465
rect 701682 358450 701706 358465
rect 701750 358450 701774 358465
rect 701818 358450 701842 358465
rect 692515 358201 693915 358329
rect 694787 358201 696187 358329
rect 699322 358295 700322 358450
rect 699322 358261 700334 358295
rect 700922 358285 701922 358450
rect 707610 358295 708610 358355
rect 709211 358295 710211 358355
rect 700910 358261 701922 358285
rect 699322 358250 700322 358261
rect 700922 358250 701922 358261
rect 699392 358237 699416 358250
rect 699460 358237 699484 358250
rect 699528 358237 699552 358250
rect 699596 358237 699620 358250
rect 699664 358237 699688 358250
rect 699732 358237 699756 358250
rect 699800 358237 699824 358250
rect 699868 358237 699892 358250
rect 699936 358237 699960 358250
rect 700004 358237 700028 358250
rect 700072 358237 700096 358250
rect 700140 358237 700164 358250
rect 700208 358237 700232 358250
rect 700276 358237 700300 358250
rect 700934 358237 700958 358250
rect 701002 358237 701026 358250
rect 701070 358237 701094 358250
rect 701138 358237 701162 358250
rect 701206 358237 701230 358250
rect 701274 358237 701298 358250
rect 701342 358237 701366 358250
rect 701410 358237 701434 358250
rect 701478 358237 701502 358250
rect 701546 358237 701570 358250
rect 701614 358237 701638 358250
rect 701682 358237 701706 358250
rect 701750 358237 701774 358250
rect 701818 358237 701842 358250
rect 692515 358038 693915 358166
rect 694787 358038 696187 358166
rect 692047 357468 696655 358004
rect 699322 357892 700322 357948
rect 700922 357892 701922 357948
rect 707610 357937 708610 357993
rect 709211 357937 710211 357993
rect 699322 357820 700322 357876
rect 700922 357820 701922 357876
rect 707610 357865 708610 357921
rect 709211 357865 710211 357921
rect 697314 357582 697620 357752
rect 699322 357518 700322 357590
rect 700922 357518 701922 357590
rect 707610 357563 708610 357635
rect 709211 357563 710211 357635
rect 704719 357527 705057 357543
rect 699392 357507 699426 357518
rect 699460 357507 699494 357518
rect 699528 357507 699562 357518
rect 699596 357507 699630 357518
rect 699664 357507 699698 357518
rect 699732 357507 699766 357518
rect 699800 357507 699834 357518
rect 699868 357507 699902 357518
rect 699936 357507 699970 357518
rect 700004 357507 700038 357518
rect 700072 357507 700106 357518
rect 700140 357507 700174 357518
rect 700208 357507 700242 357518
rect 700276 357507 700310 357518
rect 700934 357507 700968 357518
rect 701002 357507 701036 357518
rect 701070 357507 701104 357518
rect 701138 357507 701172 357518
rect 701206 357507 701240 357518
rect 701274 357507 701308 357518
rect 701342 357507 701376 357518
rect 701410 357507 701444 357518
rect 701478 357507 701512 357518
rect 701546 357507 701580 357518
rect 701614 357507 701648 357518
rect 701682 357507 701716 357518
rect 701750 357507 701784 357518
rect 701818 357507 701852 357518
rect 699392 357497 699450 357507
rect 699460 357497 699518 357507
rect 699528 357497 699586 357507
rect 699596 357497 699654 357507
rect 699664 357497 699722 357507
rect 699732 357497 699790 357507
rect 699800 357497 699858 357507
rect 699868 357497 699926 357507
rect 699936 357497 699994 357507
rect 700004 357497 700062 357507
rect 700072 357497 700130 357507
rect 700140 357497 700198 357507
rect 700208 357497 700266 357507
rect 700276 357497 700334 357507
rect 700934 357497 700992 357507
rect 701002 357497 701060 357507
rect 701070 357497 701128 357507
rect 701138 357497 701196 357507
rect 701206 357497 701264 357507
rect 701274 357497 701332 357507
rect 701342 357497 701400 357507
rect 701410 357497 701468 357507
rect 701478 357497 701536 357507
rect 701546 357497 701604 357507
rect 701614 357497 701672 357507
rect 701682 357497 701740 357507
rect 701750 357497 701808 357507
rect 701818 357497 701876 357507
rect 699368 357473 700334 357497
rect 700910 357473 701876 357497
rect 699392 357458 699416 357473
rect 699460 357458 699484 357473
rect 699528 357458 699552 357473
rect 699596 357458 699620 357473
rect 699664 357458 699688 357473
rect 699732 357458 699756 357473
rect 699800 357458 699824 357473
rect 699868 357458 699892 357473
rect 699936 357458 699960 357473
rect 700004 357458 700028 357473
rect 700072 357458 700096 357473
rect 700140 357458 700164 357473
rect 700208 357458 700232 357473
rect 700276 357458 700300 357473
rect 700934 357458 700958 357473
rect 701002 357458 701026 357473
rect 701070 357458 701094 357473
rect 701138 357458 701162 357473
rect 701206 357458 701230 357473
rect 701274 357458 701298 357473
rect 701342 357458 701366 357473
rect 701410 357458 701434 357473
rect 701478 357458 701502 357473
rect 701546 357458 701570 357473
rect 701614 357458 701638 357473
rect 701682 357458 701706 357473
rect 701750 357458 701774 357473
rect 701818 357458 701842 357473
rect 699322 357303 700322 357458
rect 692463 357268 692511 357292
rect 696191 357268 696239 357292
rect 692487 357214 692511 357268
rect 696215 357214 696239 357268
rect 699322 357269 700334 357303
rect 700922 357293 701922 357458
rect 704735 357425 705041 357527
rect 707610 357303 708610 357363
rect 709211 357303 710211 357363
rect 700910 357269 701922 357293
rect 699322 357258 700322 357269
rect 700922 357258 701922 357269
rect 699392 357245 699416 357258
rect 699460 357245 699484 357258
rect 699528 357245 699552 357258
rect 699596 357245 699620 357258
rect 699664 357245 699688 357258
rect 699732 357245 699756 357258
rect 699800 357245 699824 357258
rect 699868 357245 699892 357258
rect 699936 357245 699960 357258
rect 700004 357245 700028 357258
rect 700072 357245 700096 357258
rect 700140 357245 700164 357258
rect 700208 357245 700232 357258
rect 700276 357245 700300 357258
rect 700934 357245 700958 357258
rect 701002 357245 701026 357258
rect 701070 357245 701094 357258
rect 701138 357245 701162 357258
rect 701206 357245 701230 357258
rect 701274 357245 701298 357258
rect 701342 357245 701366 357258
rect 701410 357245 701434 357258
rect 701478 357245 701502 357258
rect 701546 357245 701570 357258
rect 701614 357245 701638 357258
rect 701682 357245 701706 357258
rect 701750 357245 701774 357258
rect 701818 357245 701842 357258
rect 692463 357190 692511 357214
rect 696191 357190 696239 357214
rect 687686 357119 687720 357153
rect 687798 357141 687822 357165
rect 687686 357095 687710 357119
rect 687774 357117 687798 357129
rect 687798 357081 687822 357105
rect 692450 357037 692474 357061
rect 692508 357037 692532 357061
rect 696170 357037 696194 357061
rect 696228 357037 696252 357061
rect 692484 357013 692498 357037
rect 696204 357013 696218 357037
rect 692484 356935 692487 356959
rect 696215 356935 696218 356959
rect 692508 356911 692532 356935
rect 696170 356911 696194 356935
rect 699322 356900 700322 356956
rect 700922 356900 701922 356956
rect 707610 356945 708610 357001
rect 709211 356945 710211 357001
rect 692515 356805 693915 356848
rect 694787 356805 696187 356848
rect 699322 356828 700322 356884
rect 700922 356828 701922 356884
rect 707610 356873 708610 356929
rect 709211 356873 710211 356929
rect 692515 356642 693915 356770
rect 694787 356642 696187 356770
rect 688883 356473 688918 356502
rect 692515 356479 693915 356607
rect 694787 356479 696187 356607
rect 699322 356526 700322 356598
rect 700922 356526 701922 356598
rect 707610 356571 708610 356643
rect 709211 356571 710211 356643
rect 699392 356515 699426 356526
rect 699460 356515 699494 356526
rect 699528 356515 699562 356526
rect 699596 356515 699630 356526
rect 699664 356515 699698 356526
rect 699732 356515 699766 356526
rect 699800 356515 699834 356526
rect 699868 356515 699902 356526
rect 699936 356515 699970 356526
rect 700004 356515 700038 356526
rect 700072 356515 700106 356526
rect 700140 356515 700174 356526
rect 700208 356515 700242 356526
rect 700276 356515 700310 356526
rect 700934 356515 700968 356526
rect 701002 356515 701036 356526
rect 701070 356515 701104 356526
rect 701138 356515 701172 356526
rect 701206 356515 701240 356526
rect 701274 356515 701308 356526
rect 701342 356515 701376 356526
rect 701410 356515 701444 356526
rect 701478 356515 701512 356526
rect 701546 356515 701580 356526
rect 701614 356515 701648 356526
rect 701682 356515 701716 356526
rect 701750 356515 701784 356526
rect 701818 356515 701852 356526
rect 699392 356505 699450 356515
rect 699460 356505 699518 356515
rect 699528 356505 699586 356515
rect 699596 356505 699654 356515
rect 699664 356505 699722 356515
rect 699732 356505 699790 356515
rect 699800 356505 699858 356515
rect 699868 356505 699926 356515
rect 699936 356505 699994 356515
rect 700004 356505 700062 356515
rect 700072 356505 700130 356515
rect 700140 356505 700198 356515
rect 700208 356505 700266 356515
rect 700276 356505 700334 356515
rect 700934 356505 700992 356515
rect 701002 356505 701060 356515
rect 701070 356505 701128 356515
rect 701138 356505 701196 356515
rect 701206 356505 701264 356515
rect 701274 356505 701332 356515
rect 701342 356505 701400 356515
rect 701410 356505 701468 356515
rect 701478 356505 701536 356515
rect 701546 356505 701604 356515
rect 701614 356505 701672 356515
rect 701682 356505 701740 356515
rect 701750 356505 701808 356515
rect 701818 356505 701876 356515
rect 699368 356481 700334 356505
rect 700910 356481 701876 356505
rect 688883 356468 688884 356473
rect 688917 356468 688918 356473
rect 688917 356439 688951 356468
rect 699392 356466 699416 356481
rect 699460 356466 699484 356481
rect 699528 356466 699552 356481
rect 699596 356466 699620 356481
rect 699664 356466 699688 356481
rect 699732 356466 699756 356481
rect 699800 356466 699824 356481
rect 699868 356466 699892 356481
rect 699936 356466 699960 356481
rect 700004 356466 700028 356481
rect 700072 356466 700096 356481
rect 700140 356466 700164 356481
rect 700208 356466 700232 356481
rect 700276 356466 700300 356481
rect 700934 356466 700958 356481
rect 701002 356466 701026 356481
rect 701070 356466 701094 356481
rect 701138 356466 701162 356481
rect 701206 356466 701230 356481
rect 701274 356466 701298 356481
rect 701342 356466 701366 356481
rect 701410 356466 701434 356481
rect 701478 356466 701502 356481
rect 701546 356466 701570 356481
rect 701614 356466 701638 356481
rect 701682 356466 701706 356481
rect 701750 356466 701774 356481
rect 701818 356466 701842 356481
rect 688917 356370 688951 356404
rect 688917 356301 688951 356335
rect 692515 356316 693915 356444
rect 694787 356316 696187 356444
rect 699322 356311 700322 356466
rect 688917 356232 688951 356266
rect 688917 356163 688951 356197
rect 692515 356153 693915 356281
rect 694787 356153 696187 356281
rect 699322 356277 700334 356311
rect 700922 356301 701922 356466
rect 707610 356311 708610 356371
rect 709211 356311 710211 356371
rect 700910 356277 701922 356301
rect 699322 356266 700322 356277
rect 700922 356266 701922 356277
rect 699392 356253 699416 356266
rect 699460 356253 699484 356266
rect 699528 356253 699552 356266
rect 699596 356253 699620 356266
rect 699664 356253 699688 356266
rect 699732 356253 699756 356266
rect 699800 356253 699824 356266
rect 699868 356253 699892 356266
rect 699936 356253 699960 356266
rect 700004 356253 700028 356266
rect 700072 356253 700096 356266
rect 700140 356253 700164 356266
rect 700208 356253 700232 356266
rect 700276 356253 700300 356266
rect 700934 356253 700958 356266
rect 701002 356253 701026 356266
rect 701070 356253 701094 356266
rect 701138 356253 701162 356266
rect 701206 356253 701230 356266
rect 701274 356253 701298 356266
rect 701342 356253 701366 356266
rect 701410 356253 701434 356266
rect 701478 356253 701502 356266
rect 701546 356253 701570 356266
rect 701614 356253 701638 356266
rect 701682 356253 701706 356266
rect 701750 356253 701774 356266
rect 701818 356253 701842 356266
rect 688917 356094 688951 356128
rect 688917 356025 688951 356059
rect 692515 355996 693915 356046
rect 694787 355996 696187 356046
rect 688917 355956 688951 355990
rect 698017 355933 698120 355969
rect 688917 355887 688951 355921
rect 692463 355885 692511 355909
rect 696191 355885 696239 355909
rect 688917 355818 688951 355852
rect 692487 355831 692511 355885
rect 696215 355831 696239 355885
rect 698017 355858 698053 355933
rect 692463 355807 692511 355831
rect 696191 355807 696239 355831
rect 698030 355824 698077 355858
rect 698017 355790 698053 355824
rect 688917 355749 688951 355783
rect 698030 355756 698077 355790
rect 698017 355722 698053 355756
rect 688917 355680 688951 355714
rect 698030 355688 698077 355722
rect 698017 355654 698053 355688
rect 688917 355611 688951 355645
rect 692463 355629 692521 355653
rect 696191 355629 696249 355653
rect 692487 355619 692521 355629
rect 696215 355619 696249 355629
rect 698030 355620 698077 355654
rect 698017 355586 698053 355620
rect 686879 355544 687585 355554
rect 686882 355528 687585 355544
rect 688917 355542 688951 355576
rect 692487 355547 692521 355581
rect 696215 355547 696249 355581
rect 678680 355433 678704 355467
rect 681345 355399 682345 355455
rect 678680 355365 678704 355399
rect 684004 355349 685004 355477
rect 688917 355473 688951 355507
rect 692487 355475 692521 355509
rect 696215 355475 696249 355509
rect 688917 355404 688951 355438
rect 692487 355427 692521 355437
rect 696215 355427 696249 355437
rect 692463 355403 692521 355427
rect 696191 355403 696249 355427
rect 688917 355335 688951 355369
rect 2850 355304 3850 355320
rect 2850 355188 3850 355238
rect 2850 354978 3850 355028
rect 3959 355015 3960 355320
rect 5169 355315 5191 355320
rect 6005 355305 6021 355320
rect 1288 353503 1338 354503
rect 1438 353503 1566 354060
rect 1594 353503 1644 354503
rect 5995 353493 6021 355275
rect 7389 354911 8389 354967
rect 8990 354911 9990 354967
rect 15678 354956 16678 355012
rect 17278 354956 18278 355012
rect 7389 354839 8389 354895
rect 8990 354839 9990 354895
rect 15678 354884 16678 354940
rect 17278 354884 18278 354940
rect 27622 354903 27672 355320
rect 27772 354903 27828 355320
rect 27928 354903 27984 355320
rect 28084 354903 28140 355320
rect 28240 354903 28296 355320
rect 28396 354903 28446 355320
rect 31049 355234 32049 355284
rect 36785 355242 37385 355298
rect 678680 355297 678704 355331
rect 678680 355229 678704 355263
rect 679133 355255 679283 355267
rect 679452 355255 679602 355267
rect 681345 355229 682345 355279
rect 678680 355161 678704 355195
rect 684004 355193 685004 355321
rect 688917 355266 688951 355300
rect 679002 355142 679602 355192
rect 36785 355072 37385 355122
rect 678680 355093 678704 355127
rect 681441 355064 681457 355130
rect 682225 355064 682241 355130
rect 678680 355025 678704 355059
rect 684004 355037 685004 355165
rect 685537 355161 686137 355211
rect 688917 355197 688951 355231
rect 692463 355214 692521 355248
rect 696191 355214 696249 355248
rect 688917 355128 688951 355162
rect 678680 354957 678704 354991
rect 679002 354966 679602 355022
rect 678680 354889 678704 354923
rect 681441 354902 681457 354968
rect 683625 354902 683641 354968
rect 684004 354881 685004 355009
rect 685537 355005 686137 355061
rect 688917 355059 688951 355093
rect 692515 355084 693915 355127
rect 694787 355084 696187 355127
rect 688917 354990 688951 355024
rect 688917 354921 688951 354955
rect 692515 354921 693915 355049
rect 694787 354921 696187 355049
rect 685537 354855 686137 354905
rect 678680 354821 678704 354855
rect 679002 354796 679602 354846
rect 678680 354753 678704 354787
rect 680502 354761 680517 354776
rect 21481 354656 22881 354699
rect 23617 354656 25017 354699
rect 678680 354685 678704 354719
rect 31458 354590 32058 354640
rect 678680 354617 678704 354651
rect 15678 354382 16678 354522
rect 17278 354382 18278 354522
rect 21481 354520 22881 354563
rect 23617 354520 25017 354563
rect 678680 354549 678704 354583
rect 680480 354581 680517 354761
rect 680502 354566 680517 354581
rect 680615 354761 680630 354776
rect 680803 354772 680815 354776
rect 680800 354761 680815 354772
rect 680615 354581 680815 354761
rect 681441 354740 681457 354806
rect 683625 354740 683641 354806
rect 684004 354725 685004 354853
rect 688917 354852 688951 354886
rect 688917 354783 688951 354817
rect 692515 354758 693915 354886
rect 694787 354758 696187 354886
rect 688917 354714 688951 354748
rect 686829 354649 687429 354699
rect 688917 354645 688951 354679
rect 680615 354566 680630 354581
rect 680800 354570 680815 354581
rect 681441 354578 681457 354644
rect 682225 354578 682241 354644
rect 684004 354575 685004 354625
rect 688917 354576 688951 354610
rect 692515 354595 693915 354723
rect 694787 354595 696187 354723
rect 680803 354566 680815 354570
rect 680615 354525 680630 354540
rect 680803 354536 680815 354540
rect 680800 354525 680815 354536
rect 678680 354481 678704 354515
rect 31458 354414 32058 354470
rect 678680 354413 678704 354447
rect 678680 354345 678704 354379
rect 679007 354370 679607 354420
rect 680615 354345 680815 354525
rect 681345 354429 682345 354479
rect 686829 354473 687429 354529
rect 688917 354507 688951 354541
rect 688917 354438 688951 354472
rect 692515 354432 693915 354560
rect 694787 354432 696187 354560
rect 684054 354373 685054 354423
rect 688917 354393 688951 354403
rect 688893 354369 688951 354393
rect 680615 354330 680630 354345
rect 680800 354334 680815 354345
rect 680803 354330 680815 354334
rect 25725 354197 26325 354247
rect 31458 354244 32058 354294
rect 678680 354277 678704 354311
rect 681345 354253 682345 354309
rect 678680 354209 678704 354243
rect 7353 354016 8425 354052
rect 7353 353975 7389 354016
rect 8389 353975 8425 354016
rect 7353 353919 8425 353975
rect 7353 353903 7389 353919
rect 8389 353903 8425 353919
rect 7353 353847 8425 353903
rect 7353 353810 7389 353847
rect 8389 353810 8425 353847
rect 7353 353770 8425 353810
rect 8954 354016 10026 354052
rect 8954 353975 8990 354016
rect 9990 353975 10026 354016
rect 8954 353919 10026 353975
rect 21383 354044 21403 354060
rect 21407 354044 21415 354060
rect 21383 354010 21419 354044
rect 21481 354031 22881 354060
rect 23617 354031 25017 354060
rect 25101 354044 25121 354060
rect 25125 354044 25143 354060
rect 25725 354047 26325 354097
rect 25101 354010 25147 354044
rect 21383 353976 21403 354010
rect 21407 353976 21415 354010
rect 21383 353942 21419 353976
rect 8954 353903 8990 353919
rect 9990 353903 10026 353919
rect 15678 353906 16678 353923
rect 17278 353906 18278 353923
rect 21383 353908 21403 353942
rect 21407 353908 21415 353942
rect 8954 353847 10026 353903
rect 20250 353890 20316 353906
rect 8954 353810 8990 353847
rect 9990 353810 10026 353847
rect 8954 353770 10026 353810
rect 21383 353874 21419 353908
rect 21383 353840 21403 353874
rect 21407 353840 21415 353874
rect 21481 353868 22881 353996
rect 23617 353868 25017 353996
rect 25101 353976 25121 354010
rect 25125 353976 25143 354010
rect 25101 353942 25147 353976
rect 25101 353908 25121 353942
rect 25125 353908 25143 353942
rect 25725 353925 26325 353975
rect 25101 353874 25147 353908
rect 25101 353840 25121 353874
rect 25125 353840 25143 353874
rect 21383 353806 21419 353840
rect 21383 353772 21403 353806
rect 21407 353772 21415 353806
rect 21383 353738 21419 353772
rect 15678 353703 16678 353736
rect 17278 353703 18278 353736
rect 21383 353704 21403 353738
rect 21407 353704 21415 353738
rect 21481 353705 22881 353833
rect 23617 353705 25017 353833
rect 25101 353806 25147 353840
rect 25101 353772 25121 353806
rect 25125 353772 25143 353806
rect 25725 353775 26325 353825
rect 25101 353738 25147 353772
rect 25101 353704 25121 353738
rect 25125 353704 25143 353738
rect 21383 353670 21419 353704
rect 25101 353670 25147 353704
rect 21383 353636 21403 353670
rect 21407 353636 21415 353670
rect 7389 353559 8389 353631
rect 8990 353559 9990 353631
rect 21383 353602 21419 353636
rect 15840 353510 15870 353580
rect 15878 353546 15908 353580
rect 21383 353568 21403 353602
rect 21407 353568 21415 353602
rect 15853 353508 15870 353510
rect 21383 353534 21419 353568
rect 21481 353542 22881 353670
rect 23617 353542 25017 353670
rect 25101 353636 25121 353670
rect 25125 353636 25143 353670
rect 25725 353649 26325 353699
rect 25101 353602 25147 353636
rect 25101 353568 25121 353602
rect 25125 353568 25143 353602
rect 25101 353534 25147 353568
rect 5981 353483 6021 353493
rect 5137 353469 6021 353483
rect 21383 353500 21403 353534
rect 21407 353500 21415 353534
rect 21383 353466 21419 353500
rect 7389 353369 8389 353463
rect 7389 353359 8413 353369
rect 8990 353359 9990 353463
rect 21383 353432 21403 353466
rect 21407 353432 21415 353466
rect 21383 353398 21419 353432
rect 21383 353364 21403 353398
rect 21407 353364 21415 353398
rect 21481 353379 22881 353507
rect 23617 353379 25017 353507
rect 25101 353500 25121 353534
rect 25125 353500 25143 353534
rect 25101 353466 25147 353500
rect 25725 353499 26325 353549
rect 25101 353432 25121 353466
rect 25125 353432 25143 353466
rect 25101 353398 25147 353432
rect 25101 353364 25121 353398
rect 25125 353364 25143 353398
rect 25725 353377 26325 353427
rect 21383 353330 21419 353364
rect 25101 353330 25147 353364
rect 21383 353296 21403 353330
rect 21407 353296 21415 353330
rect 25101 353296 25121 353330
rect 25125 353296 25143 353330
rect 21383 353262 21419 353296
rect 21383 353228 21403 353262
rect 21407 353228 21415 353262
rect 21481 353229 22881 353272
rect 23617 353229 25017 353272
rect 25101 353262 25147 353296
rect 25101 353228 25121 353262
rect 25125 353228 25143 353262
rect 21383 353194 21419 353228
rect 25101 353194 25147 353228
rect 25725 353227 26325 353277
rect 21383 353160 21403 353194
rect 21407 353160 21415 353194
rect 25101 353160 25121 353194
rect 25125 353160 25143 353194
rect 27162 353170 27212 354170
rect 27312 353170 27440 354060
rect 27468 353170 27596 354060
rect 27624 353170 27752 354060
rect 27780 353170 27908 354060
rect 27936 353170 28064 354060
rect 28092 353170 28220 354060
rect 28248 353170 28376 354060
rect 28404 353170 28532 354060
rect 28560 353170 28688 354060
rect 28716 353170 28844 354060
rect 28872 353170 29000 354060
rect 29028 353170 29156 354060
rect 29184 353170 29312 354060
rect 29340 353170 29390 354170
rect 30245 354029 30445 354209
rect 30245 354018 30260 354029
rect 30245 354014 30257 354018
rect 30430 354014 30445 354029
rect 30543 354029 30580 354209
rect 679007 354200 679607 354250
rect 684054 354217 685054 354345
rect 686829 354303 687429 354353
rect 692515 354269 693915 354397
rect 694787 354269 696187 354397
rect 678680 354141 678704 354175
rect 678680 354073 678704 354107
rect 681345 354077 682345 354205
rect 30543 354014 30558 354029
rect 678680 354005 678704 354039
rect 680215 354024 680815 354074
rect 684054 354061 685054 354189
rect 685793 354182 685805 354186
rect 685793 354171 685808 354182
rect 685978 354171 685993 354186
rect 30245 353984 30257 353988
rect 30245 353973 30260 353984
rect 30430 353973 30445 353988
rect 30245 353793 30445 353973
rect 678680 353937 678704 353971
rect 678680 353869 678704 353903
rect 31453 353818 32053 353868
rect 680215 353848 680815 353904
rect 681345 353901 682345 354029
rect 684054 353905 685054 354033
rect 685793 353991 685993 354171
rect 685793 353980 685808 353991
rect 685793 353976 685805 353980
rect 685978 353976 685993 353991
rect 686053 354182 686065 354186
rect 686053 354171 686068 354182
rect 686238 354171 686253 354186
rect 686053 353991 686253 354171
rect 686607 354164 687607 354214
rect 697088 354171 697138 355571
rect 697238 354171 697366 355571
rect 697394 354171 697522 355571
rect 697550 354171 697678 355571
rect 697706 354171 697756 355571
rect 698030 355552 698077 355586
rect 698017 355518 698053 355552
rect 698030 355484 698077 355518
rect 698017 355450 698053 355484
rect 698030 355416 698077 355450
rect 698017 355382 698053 355416
rect 698030 355348 698077 355382
rect 698017 355314 698053 355348
rect 698030 355280 698077 355314
rect 698017 355246 698053 355280
rect 698030 355212 698077 355246
rect 698017 355178 698053 355212
rect 698030 355144 698077 355178
rect 698017 355110 698053 355144
rect 698030 355076 698077 355110
rect 698017 355042 698053 355076
rect 698030 355008 698077 355042
rect 698017 354974 698053 355008
rect 698030 354940 698077 354974
rect 698017 354906 698053 354940
rect 698030 354872 698077 354906
rect 698017 354838 698053 354872
rect 698030 354804 698077 354838
rect 698017 354770 698053 354804
rect 698030 354736 698077 354770
rect 698017 354702 698053 354736
rect 698030 354668 698077 354702
rect 698017 354634 698053 354668
rect 698030 354600 698077 354634
rect 698017 354566 698053 354600
rect 698030 354532 698077 354566
rect 698017 354498 698053 354532
rect 698030 354464 698077 354498
rect 698017 354430 698053 354464
rect 698030 354396 698077 354430
rect 698017 354362 698053 354396
rect 698030 354328 698077 354362
rect 698017 354294 698053 354328
rect 698030 354260 698077 354294
rect 698017 354226 698053 354260
rect 698030 354192 698077 354226
rect 692515 354119 693915 354162
rect 694787 354119 696187 354162
rect 698017 354158 698053 354192
rect 698030 354124 698077 354158
rect 698017 354090 698053 354124
rect 686607 354014 687607 354064
rect 698030 354056 698077 354090
rect 686053 353980 686068 353991
rect 686053 353976 686065 353980
rect 686238 353976 686253 353991
rect 685793 353946 685805 353950
rect 685793 353935 685808 353946
rect 685978 353935 685993 353950
rect 678680 353801 678704 353835
rect 30245 353782 30260 353793
rect 30245 353778 30257 353782
rect 30430 353778 30445 353793
rect 678680 353733 678704 353767
rect 681345 353731 682345 353781
rect 684054 353749 685054 353877
rect 685793 353755 685993 353935
rect 685793 353744 685808 353755
rect 685793 353740 685805 353744
rect 685978 353740 685993 353755
rect 686053 353946 686065 353950
rect 686053 353935 686068 353946
rect 686238 353935 686253 353950
rect 686053 353755 686253 353935
rect 686607 353855 687607 353905
rect 692463 353809 692511 353833
rect 696191 353809 696239 353833
rect 686053 353744 686068 353755
rect 686053 353740 686065 353744
rect 686238 353740 686253 353755
rect 31453 353648 32053 353698
rect 678680 353665 678704 353699
rect 680215 353672 680815 353728
rect 681345 353662 682345 353674
rect 678680 353597 678704 353631
rect 684054 353593 685054 353721
rect 686607 353705 687607 353755
rect 692487 353731 692511 353809
rect 696215 353755 696239 353809
rect 696191 353731 696239 353755
rect 696617 353772 696651 353773
rect 696617 353749 696626 353772
rect 696617 353731 696675 353749
rect 696651 353715 696675 353731
rect 696651 353647 696675 353681
rect 685533 353586 685545 353590
rect 685533 353575 685548 353586
rect 685718 353575 685733 353590
rect 678680 353529 678704 353563
rect 30245 353472 30845 353522
rect 680215 353502 680815 353552
rect 678680 353461 678704 353495
rect 678680 353393 678704 353427
rect 680215 353370 680815 353420
rect 681466 353411 682466 353461
rect 684054 353437 685054 353565
rect 30245 353296 30845 353352
rect 678680 353325 678704 353359
rect 678680 353257 678704 353291
rect 681466 353255 682466 353383
rect 682890 353339 683490 353389
rect 678680 353189 678704 353223
rect 680215 353194 680815 353250
rect 682890 353183 683490 353311
rect 684054 353281 685054 353409
rect 685533 353395 685733 353575
rect 685533 353384 685548 353395
rect 685533 353380 685545 353384
rect 685718 353380 685733 353395
rect 685793 353586 685805 353590
rect 685793 353575 685808 353586
rect 685978 353575 685993 353590
rect 685793 353395 685993 353575
rect 685793 353384 685808 353395
rect 685793 353380 685805 353384
rect 685978 353380 685993 353395
rect 686053 353586 686065 353590
rect 686053 353575 686068 353586
rect 686238 353575 686253 353590
rect 686053 353395 686253 353575
rect 686053 353384 686068 353395
rect 686053 353380 686065 353384
rect 686238 353380 686253 353395
rect 686313 353586 686325 353590
rect 686313 353575 686328 353586
rect 686498 353575 686513 353590
rect 686313 353395 686513 353575
rect 686313 353384 686328 353395
rect 686313 353380 686325 353384
rect 686498 353380 686513 353395
rect 686627 353586 686639 353590
rect 686627 353575 686642 353586
rect 686812 353575 686827 353590
rect 686627 353395 686827 353575
rect 686627 353384 686642 353395
rect 686627 353380 686639 353384
rect 686812 353380 686827 353395
rect 686887 353586 686899 353590
rect 686887 353575 686902 353586
rect 687072 353575 687087 353590
rect 686887 353395 687087 353575
rect 686887 353384 686902 353395
rect 686887 353380 686899 353384
rect 687072 353380 687087 353395
rect 687147 353586 687159 353590
rect 687147 353575 687162 353586
rect 687332 353575 687347 353590
rect 696651 353579 696675 353613
rect 687147 353395 687347 353575
rect 696651 353511 696675 353545
rect 696651 353443 696675 353477
rect 687147 353384 687162 353395
rect 687147 353380 687159 353384
rect 687332 353380 687347 353395
rect 696651 353375 696675 353409
rect 696651 353307 696675 353341
rect 685718 353215 685733 353230
rect 685679 353185 685733 353215
rect 21383 353126 21419 353160
rect 25101 353126 25147 353160
rect 21383 353102 21403 353126
rect 21385 353048 21403 353102
rect 21407 353082 21415 353126
rect 25101 353102 25121 353126
rect 25113 353082 25121 353102
rect 25125 353048 25143 353126
rect 30245 353120 30845 353176
rect 678680 353121 678704 353155
rect 681466 353105 682466 353155
rect 684054 353131 685054 353181
rect 685718 353170 685733 353185
rect 685793 353226 685805 353230
rect 685793 353215 685808 353226
rect 685978 353215 685993 353230
rect 685793 353185 685993 353215
rect 685793 353174 685808 353185
rect 685793 353170 685805 353174
rect 685978 353170 685993 353185
rect 686053 353226 686065 353230
rect 686053 353215 686068 353226
rect 686238 353215 686253 353230
rect 686812 353215 686827 353230
rect 686053 353185 686253 353215
rect 686807 353185 686827 353215
rect 686053 353174 686068 353185
rect 686053 353170 686065 353174
rect 686238 353170 686253 353185
rect 686812 353170 686827 353185
rect 686887 353226 686899 353230
rect 686887 353215 686902 353226
rect 687072 353215 687087 353230
rect 686887 353185 687087 353215
rect 686887 353174 686902 353185
rect 686887 353170 686899 353174
rect 687072 353170 687087 353185
rect 687147 353226 687159 353230
rect 687147 353215 687162 353226
rect 687332 353215 687347 353230
rect 687147 353185 687347 353215
rect 687147 353174 687162 353185
rect 687147 353170 687159 353174
rect 687332 353170 687347 353185
rect 685718 353129 685733 353144
rect 681794 353102 682466 353105
rect 685679 353099 685733 353129
rect 678680 353053 678704 353087
rect 685718 353084 685733 353099
rect 685793 353140 685805 353144
rect 685793 353129 685808 353140
rect 685978 353129 685993 353144
rect 685793 353099 685993 353129
rect 685793 353088 685808 353099
rect 685793 353084 685805 353088
rect 685978 353084 685993 353099
rect 686053 353140 686065 353144
rect 686053 353129 686068 353140
rect 686238 353129 686253 353144
rect 686812 353129 686827 353144
rect 686053 353099 686253 353129
rect 686807 353099 686827 353129
rect 686053 353088 686068 353099
rect 686053 353084 686065 353088
rect 686238 353084 686253 353099
rect 686812 353084 686827 353099
rect 686887 353140 686899 353144
rect 686887 353129 686902 353140
rect 687072 353129 687087 353144
rect 686887 353099 687087 353129
rect 686887 353088 686902 353099
rect 686887 353084 686899 353088
rect 687072 353084 687087 353099
rect 687147 353140 687159 353144
rect 687147 353129 687162 353140
rect 687332 353129 687347 353144
rect 687147 353099 687347 353129
rect 687147 353088 687162 353099
rect 687147 353084 687159 353088
rect 687332 353084 687347 353099
rect 30245 352950 30845 353000
rect 678680 352985 678704 353019
rect 680215 353018 680815 353074
rect 682890 353027 683490 353083
rect 21000 352800 21003 352920
rect 678680 352917 678704 352951
rect 21352 352885 21376 352909
rect 25122 352885 25146 352909
rect 21385 352861 21400 352885
rect 25098 352861 25113 352885
rect 21274 352783 21294 352851
rect 21410 352817 21430 352851
rect 25068 352817 25088 352851
rect 25204 352817 25224 352851
rect 678680 352849 678704 352883
rect 680215 352848 680815 352898
rect 21385 352807 21430 352817
rect 25102 352807 25137 352817
rect 21361 352783 21430 352807
rect 25089 352783 25137 352807
rect 25238 352783 25258 352817
rect 678680 352781 678704 352815
rect 678680 352713 678704 352747
rect 678680 352645 678704 352679
rect 679007 352672 679607 352722
rect 678680 352577 678704 352611
rect 680615 352577 680630 352592
rect 680803 352588 680815 352592
rect 680800 352577 680815 352588
rect 678680 352509 678704 352543
rect 679007 352502 679607 352552
rect 678680 352441 678704 352475
rect 678680 352373 678704 352407
rect 680615 352397 680815 352577
rect 681502 352505 681529 352995
rect 681866 352896 682466 353024
rect 682890 352871 683490 352999
rect 684004 352929 685004 352979
rect 685539 352940 685777 352972
rect 685803 352920 686119 352938
rect 681866 352740 682466 352868
rect 684004 352773 685004 352901
rect 682890 352721 683490 352771
rect 681866 352584 682466 352712
rect 682890 352605 683490 352655
rect 684004 352617 685004 352745
rect 681866 352434 682466 352484
rect 682890 352449 683490 352505
rect 684004 352461 685004 352589
rect 692427 352522 693027 352572
rect 680615 352382 680630 352397
rect 680800 352386 680815 352397
rect 680803 352382 680815 352386
rect 680502 352341 680517 352356
rect 678680 352305 678704 352339
rect 678680 352237 678704 352271
rect 678680 352169 678704 352203
rect 680480 352161 680517 352341
rect 680502 352146 680517 352161
rect 680615 352341 680630 352356
rect 680803 352352 680815 352356
rect 680800 352341 680815 352352
rect 680615 352161 680815 352341
rect 681866 352318 682466 352368
rect 682890 352293 683490 352349
rect 684004 352305 685004 352433
rect 692427 352366 693027 352494
rect 693888 352375 694194 352545
rect 694388 352375 694694 352545
rect 689309 352278 689909 352328
rect 681866 352168 682466 352218
rect 682041 352165 682385 352168
rect 680615 352146 680630 352161
rect 680800 352150 680815 352161
rect 680803 352146 680815 352150
rect 682890 352137 683490 352193
rect 684004 352149 685004 352277
rect 678680 352101 678704 352135
rect 679002 352076 679602 352126
rect 689309 352122 689909 352250
rect 692427 352210 693027 352338
rect 678680 352033 678704 352067
rect 678680 351965 678704 351999
rect 682890 351981 683490 352109
rect 684004 351993 685004 352121
rect 689309 351966 689909 352094
rect 692427 352054 693027 352110
rect 678680 351897 678704 351931
rect 679002 351900 679602 351956
rect 678680 351829 678704 351863
rect 682890 351825 683490 351953
rect 684004 351837 685004 351965
rect 692427 351898 693027 352026
rect 689309 351810 689909 351866
rect 678680 351761 678704 351795
rect 679002 351730 679602 351780
rect 679061 351727 679355 351730
rect 679380 351727 679602 351730
rect 678680 351693 678704 351727
rect 682890 351669 683490 351797
rect 684004 351687 685004 351737
rect 685803 351720 686119 351732
rect 685539 351716 686119 351720
rect 685513 351682 685537 351716
rect 685539 351682 685777 351716
rect 678680 351625 678704 351659
rect 689309 351654 689909 351782
rect 690910 351754 691110 351765
rect 692427 351742 693027 351870
rect 690910 351640 691110 351690
rect 678680 351557 678704 351591
rect 678680 351489 678704 351523
rect 682890 351513 683490 351569
rect 685718 351555 685733 351570
rect 684004 351485 685004 351535
rect 685679 351525 685733 351555
rect 685718 351510 685733 351525
rect 685793 351566 685805 351570
rect 685793 351555 685808 351566
rect 685978 351555 685993 351570
rect 685793 351525 685993 351555
rect 685793 351514 685808 351525
rect 685793 351510 685805 351514
rect 685978 351510 685993 351525
rect 686053 351566 686065 351570
rect 686053 351555 686068 351566
rect 686238 351555 686253 351570
rect 686812 351555 686827 351570
rect 686053 351525 686253 351555
rect 686807 351525 686827 351555
rect 686053 351514 686068 351525
rect 686053 351510 686065 351514
rect 686238 351510 686253 351525
rect 686812 351510 686827 351525
rect 686887 351566 686899 351570
rect 686887 351555 686902 351566
rect 687072 351555 687087 351570
rect 686887 351525 687087 351555
rect 686887 351514 686902 351525
rect 686887 351510 686899 351514
rect 687072 351510 687087 351525
rect 687147 351566 687159 351570
rect 687147 351555 687162 351566
rect 687332 351555 687347 351570
rect 687147 351525 687347 351555
rect 687147 351514 687162 351525
rect 687147 351510 687159 351514
rect 687332 351510 687347 351525
rect 689309 351498 689909 351626
rect 692427 351592 693027 351642
rect 693888 351575 694194 351745
rect 694388 351575 694694 351745
rect 678680 351421 678704 351455
rect 678680 351353 678704 351387
rect 682890 351357 683490 351485
rect 690910 351484 691110 351540
rect 685718 351469 685733 351484
rect 684004 351329 685004 351457
rect 685679 351439 685733 351469
rect 685718 351424 685733 351439
rect 685793 351480 685805 351484
rect 685793 351469 685808 351480
rect 685978 351469 685993 351484
rect 685793 351439 685993 351469
rect 685793 351428 685808 351439
rect 685793 351424 685805 351428
rect 685978 351424 685993 351439
rect 686053 351480 686065 351484
rect 686053 351469 686068 351480
rect 686238 351469 686253 351484
rect 686812 351469 686827 351484
rect 686053 351439 686253 351469
rect 686807 351439 686827 351469
rect 686053 351428 686068 351439
rect 686053 351424 686065 351428
rect 686238 351424 686253 351439
rect 686812 351424 686827 351439
rect 686887 351480 686899 351484
rect 686887 351469 686902 351480
rect 687072 351469 687087 351484
rect 686887 351439 687087 351469
rect 686887 351428 686902 351439
rect 686887 351424 686899 351428
rect 687072 351424 687087 351439
rect 687147 351480 687159 351484
rect 687147 351469 687162 351480
rect 687332 351469 687347 351484
rect 687147 351439 687347 351469
rect 692427 351462 693027 351512
rect 687147 351428 687162 351439
rect 687147 351424 687159 351428
rect 687332 351424 687347 351439
rect 689309 351348 689909 351398
rect 690910 351334 691110 351384
rect 678680 351285 678704 351319
rect 678680 351217 678704 351251
rect 682890 351201 683490 351329
rect 692427 351312 693027 351362
rect 678680 351149 678704 351183
rect 684004 351173 685004 351301
rect 685533 351270 685545 351274
rect 685533 351259 685548 351270
rect 685718 351259 685733 351274
rect 678680 351081 678704 351115
rect 679133 351101 679283 351113
rect 679452 351101 679602 351113
rect 678680 351013 678704 351047
rect 682890 351045 683490 351173
rect 679002 350988 679602 351038
rect 684004 351017 685004 351145
rect 685533 351079 685733 351259
rect 685533 351068 685548 351079
rect 685533 351064 685545 351068
rect 685718 351064 685733 351079
rect 685793 351270 685805 351274
rect 685793 351259 685808 351270
rect 685978 351259 685993 351274
rect 685793 351079 685993 351259
rect 685793 351068 685808 351079
rect 685793 351064 685805 351068
rect 685978 351064 685993 351079
rect 686053 351270 686065 351274
rect 686053 351259 686068 351270
rect 686238 351259 686253 351274
rect 686053 351079 686253 351259
rect 686053 351068 686068 351079
rect 686053 351064 686065 351068
rect 686238 351064 686253 351079
rect 686313 351270 686325 351274
rect 686313 351259 686328 351270
rect 686498 351259 686513 351274
rect 686313 351079 686513 351259
rect 686313 351068 686328 351079
rect 686313 351064 686325 351068
rect 686498 351064 686513 351079
rect 686627 351270 686639 351274
rect 686627 351259 686642 351270
rect 686812 351259 686827 351274
rect 686627 351079 686827 351259
rect 686627 351068 686642 351079
rect 686627 351064 686639 351068
rect 686812 351064 686827 351079
rect 686887 351270 686899 351274
rect 686887 351259 686902 351270
rect 687072 351259 687087 351274
rect 686887 351079 687087 351259
rect 686887 351068 686902 351079
rect 686887 351064 686899 351068
rect 687072 351064 687087 351079
rect 687147 351270 687159 351274
rect 687147 351259 687162 351270
rect 687332 351259 687347 351274
rect 687147 351079 687347 351259
rect 689309 351218 689909 351268
rect 692427 351140 693027 351190
rect 687147 351068 687162 351079
rect 687147 351064 687159 351068
rect 687332 351064 687347 351079
rect 689309 351068 689909 351118
rect 692427 350990 693027 351040
rect 678680 350945 678704 350979
rect 678680 350877 678704 350911
rect 682890 350895 683490 350945
rect 678680 350809 678704 350843
rect 679002 350812 679602 350868
rect 684004 350861 685004 350917
rect 685793 350910 685805 350914
rect 685793 350899 685808 350910
rect 685978 350899 685993 350914
rect 682890 350779 683490 350829
rect 678680 350741 678704 350775
rect 678680 350673 678704 350707
rect 679002 350642 679602 350692
rect 678680 350605 678704 350639
rect 682890 350623 683490 350751
rect 684004 350705 685004 350833
rect 685793 350719 685993 350899
rect 685793 350708 685808 350719
rect 685793 350704 685805 350708
rect 685978 350704 685993 350719
rect 686053 350910 686065 350914
rect 686053 350899 686068 350910
rect 686238 350899 686253 350914
rect 686607 350899 687607 350949
rect 690910 350934 691110 350984
rect 686053 350719 686253 350899
rect 692427 350860 693027 350910
rect 686607 350749 687607 350799
rect 690910 350778 691110 350834
rect 686053 350708 686068 350719
rect 686053 350704 686065 350708
rect 686238 350704 686253 350719
rect 692427 350704 693027 350832
rect 693888 350775 694194 350945
rect 694388 350775 694694 350945
rect 680502 350607 680517 350622
rect 678680 350537 678704 350571
rect 678680 350469 678704 350503
rect 678680 350401 678704 350435
rect 680480 350427 680517 350607
rect 680502 350412 680517 350427
rect 680615 350607 680630 350622
rect 680803 350618 680815 350622
rect 680800 350607 680815 350618
rect 680615 350427 680815 350607
rect 682890 350467 683490 350595
rect 684004 350549 685004 350677
rect 685793 350674 685805 350678
rect 685793 350663 685808 350674
rect 685978 350663 685993 350678
rect 680615 350412 680630 350427
rect 680800 350416 680815 350427
rect 680803 350412 680815 350416
rect 680615 350371 680630 350386
rect 680803 350382 680815 350386
rect 680800 350371 680815 350382
rect 678680 350333 678704 350367
rect 678680 350265 678704 350299
rect 678680 350197 678704 350231
rect 679007 350216 679607 350266
rect 680615 350191 680815 350371
rect 682890 350311 683490 350439
rect 684004 350393 685004 350521
rect 685793 350483 685993 350663
rect 685793 350472 685808 350483
rect 685793 350468 685805 350472
rect 685978 350468 685993 350483
rect 686053 350674 686065 350678
rect 686053 350663 686068 350674
rect 686238 350663 686253 350678
rect 686053 350483 686253 350663
rect 686607 350590 687607 350640
rect 690910 350628 691110 350678
rect 692427 350548 693027 350676
rect 686053 350472 686068 350483
rect 686053 350468 686065 350472
rect 686238 350468 686253 350483
rect 686607 350440 687607 350490
rect 692427 350392 693027 350448
rect 686829 350301 687429 350351
rect 684004 350243 685004 350293
rect 692427 350236 693027 350364
rect 695201 350282 695251 353282
rect 695351 350282 695479 353282
rect 695507 350282 695635 353282
rect 695663 350282 695791 353282
rect 695819 350282 695947 353282
rect 695975 350282 696103 353282
rect 696131 350282 696259 353282
rect 696287 350282 696337 353282
rect 696651 353239 696675 353273
rect 696651 353171 696675 353205
rect 696651 353103 696675 353137
rect 696651 353035 696675 353069
rect 696651 352967 696675 353001
rect 696651 352899 696675 352933
rect 696651 352831 696675 352865
rect 696651 352763 696675 352797
rect 696651 352695 696675 352729
rect 696651 352627 696675 352661
rect 697088 352641 697138 354041
rect 697238 352641 697366 354041
rect 697394 352641 697522 354041
rect 697550 352641 697678 354041
rect 697706 352641 697756 354041
rect 698017 354022 698053 354056
rect 698030 353988 698077 354022
rect 698017 353954 698053 353988
rect 698030 353920 698077 353954
rect 698017 353886 698053 353920
rect 698030 353852 698077 353886
rect 698017 353818 698053 353852
rect 698030 353784 698077 353818
rect 698017 353750 698053 353784
rect 698030 353716 698077 353750
rect 698017 353682 698053 353716
rect 698030 353648 698077 353682
rect 698017 353614 698053 353648
rect 698030 353580 698077 353614
rect 698017 353546 698053 353580
rect 698030 353512 698077 353546
rect 698017 353478 698053 353512
rect 698030 353444 698077 353478
rect 698017 353410 698053 353444
rect 698030 353376 698077 353410
rect 698017 353342 698053 353376
rect 698030 353308 698077 353342
rect 698017 353274 698053 353308
rect 698030 353240 698077 353274
rect 698017 353206 698053 353240
rect 698030 353172 698077 353206
rect 698017 353138 698053 353172
rect 698030 353104 698077 353138
rect 698017 353070 698053 353104
rect 698030 353036 698077 353070
rect 698017 353002 698053 353036
rect 698030 352968 698077 353002
rect 698017 352934 698053 352968
rect 698030 352900 698077 352934
rect 698017 352866 698053 352900
rect 698030 352832 698077 352866
rect 698017 352798 698053 352832
rect 698030 352764 698077 352798
rect 698017 352730 698053 352764
rect 698030 352696 698077 352730
rect 698017 352662 698053 352696
rect 698030 352628 698077 352662
rect 698017 352594 698053 352628
rect 696651 352559 696675 352593
rect 698030 352560 698077 352594
rect 698017 352526 698053 352560
rect 696651 352491 696675 352525
rect 698030 352492 698077 352526
rect 696651 352423 696675 352457
rect 698017 352428 698053 352492
rect 698030 352394 698077 352428
rect 696651 352355 696675 352389
rect 698017 352360 698053 352394
rect 698030 352326 698077 352360
rect 696651 352287 696675 352321
rect 698017 352292 698053 352326
rect 696651 352219 696675 352253
rect 696651 352151 696675 352185
rect 696651 352083 696675 352117
rect 696651 352015 696675 352049
rect 696651 351947 696675 351981
rect 696651 351879 696675 351913
rect 696651 351811 696675 351845
rect 696651 351743 696675 351777
rect 696651 351675 696675 351709
rect 696651 351607 696675 351641
rect 696651 351539 696675 351573
rect 696651 351471 696675 351505
rect 696651 351403 696675 351437
rect 696651 351335 696675 351369
rect 696651 351267 696675 351301
rect 696651 351199 696675 351233
rect 696651 351131 696675 351165
rect 696651 351063 696675 351097
rect 696651 350995 696675 351029
rect 696651 350927 696675 350961
rect 696651 350859 696675 350893
rect 697088 350879 697138 352279
rect 697238 350879 697366 352279
rect 697394 350879 697522 352279
rect 697550 350879 697678 352279
rect 697706 350879 697756 352279
rect 698030 352258 698077 352292
rect 698017 352224 698053 352258
rect 698030 352190 698077 352224
rect 698017 352156 698053 352190
rect 698030 352122 698077 352156
rect 698017 352088 698053 352122
rect 698030 352054 698077 352088
rect 698017 352020 698053 352054
rect 698030 351986 698077 352020
rect 698017 351952 698053 351986
rect 698030 351918 698077 351952
rect 698017 351884 698053 351918
rect 698030 351850 698077 351884
rect 698017 351816 698053 351850
rect 698030 351782 698077 351816
rect 698017 351748 698053 351782
rect 698030 351714 698077 351748
rect 698017 351680 698053 351714
rect 698030 351646 698077 351680
rect 698017 351612 698053 351646
rect 698030 351578 698077 351612
rect 698017 351544 698053 351578
rect 698030 351510 698077 351544
rect 698017 351476 698053 351510
rect 698030 351442 698077 351476
rect 698017 351408 698053 351442
rect 698030 351374 698077 351408
rect 698017 351340 698053 351374
rect 698030 351306 698077 351340
rect 698017 351272 698053 351306
rect 698030 351238 698077 351272
rect 698017 351204 698053 351238
rect 698030 351170 698077 351204
rect 698017 351136 698053 351170
rect 698030 351102 698077 351136
rect 698017 351068 698053 351102
rect 698030 351034 698077 351068
rect 698017 351000 698053 351034
rect 698030 350966 698077 351000
rect 698017 350932 698053 350966
rect 698030 350898 698077 350932
rect 698017 350864 698053 350898
rect 698030 350830 698077 350864
rect 696651 350791 696675 350825
rect 698017 350796 698053 350830
rect 698030 350762 698077 350796
rect 696651 350723 696675 350757
rect 696651 350655 696675 350689
rect 696651 350587 696675 350621
rect 696651 350519 696675 350553
rect 696651 350451 696675 350485
rect 696651 350383 696675 350417
rect 696651 350315 696675 350349
rect 696651 350247 696675 350281
rect 680615 350176 680630 350191
rect 680800 350180 680815 350191
rect 680803 350176 680815 350180
rect 678680 350129 678704 350163
rect 682890 350161 683490 350211
rect 684004 350127 685004 350177
rect 686829 350125 687429 350181
rect 678680 350061 678704 350095
rect 679007 350046 679607 350096
rect 692427 350080 693027 350208
rect 696651 350179 696675 350213
rect 696651 350111 696675 350145
rect 696651 350043 696675 350077
rect 678680 349993 678704 350027
rect 681664 350002 681812 350006
rect 681641 349994 681812 350002
rect 682113 349994 682313 350006
rect 684004 349971 685004 350027
rect 678680 349925 678704 349959
rect 686829 349955 687429 350005
rect 678680 349857 678704 349891
rect 680215 349870 680815 349920
rect 681713 349881 682313 349931
rect 682921 349899 683521 349949
rect 692427 349930 693027 349980
rect 696651 349975 696675 350009
rect 696651 349907 696675 349941
rect 678680 349789 678704 349823
rect 684004 349821 685004 349871
rect 678680 349721 678704 349755
rect 680215 349694 680815 349750
rect 681713 349705 682313 349761
rect 682921 349743 683521 349799
rect 685537 349749 686137 349799
rect 697088 349749 697138 350749
rect 697238 349749 697366 350749
rect 697394 349749 697522 350749
rect 697550 349749 697678 350749
rect 697706 349749 697756 350749
rect 698017 350728 698053 350762
rect 698030 350694 698077 350728
rect 698017 350660 698053 350694
rect 698030 350626 698077 350660
rect 698017 350592 698053 350626
rect 698030 350558 698077 350592
rect 698017 350524 698053 350558
rect 698030 350490 698077 350524
rect 698017 350456 698053 350490
rect 698030 350422 698077 350456
rect 698017 350388 698053 350422
rect 698030 350354 698077 350388
rect 698017 350320 698053 350354
rect 698030 350286 698077 350320
rect 698017 350252 698053 350286
rect 698030 350218 698077 350252
rect 698017 350184 698053 350218
rect 698030 350150 698077 350184
rect 698017 350116 698053 350150
rect 698030 350082 698077 350116
rect 698017 350048 698053 350082
rect 698030 350014 698077 350048
rect 698017 349980 698053 350014
rect 698030 349946 698077 349980
rect 698017 349912 698053 349946
rect 698030 349878 698077 349912
rect 698017 349844 698053 349878
rect 698030 349810 698077 349844
rect 698017 349776 698053 349810
rect 698030 349742 698077 349776
rect 698017 349708 698053 349742
rect 678680 349653 678704 349687
rect 698030 349674 698077 349708
rect 678680 349585 678704 349619
rect 680215 349518 680815 349574
rect 681713 349529 682313 349657
rect 682921 349593 683521 349643
rect 684070 349599 684670 349649
rect 685537 349593 686137 349649
rect 698017 349640 698053 349674
rect 698030 349606 698077 349640
rect 698017 349572 698053 349606
rect 698030 349538 698077 349572
rect 698017 349504 698053 349538
rect 684070 349443 684670 349499
rect 685537 349443 686137 349493
rect 692428 349442 693028 349492
rect 698030 349470 698077 349504
rect 698017 349436 698053 349470
rect 680215 349348 680815 349398
rect 681713 349359 682313 349409
rect 698030 349402 698077 349436
rect 698017 349368 698053 349402
rect 684070 349293 684670 349343
rect 692428 349292 693028 349342
rect 698030 349334 698077 349368
rect 698017 349300 698053 349334
rect 680215 349232 680815 349282
rect 698030 349266 698077 349300
rect 698017 349232 698053 349266
rect 692428 349162 693028 349212
rect 698030 349198 698077 349232
rect 698017 349164 698053 349198
rect 680215 349056 680815 349112
rect 692428 349006 693028 349134
rect 698030 349130 698077 349164
rect 698017 349096 698053 349130
rect 698030 349062 698077 349096
rect 698017 348983 698053 349062
rect 698084 348983 698120 355933
rect 699322 355908 700322 355964
rect 700922 355908 701922 355964
rect 707610 355953 708610 356009
rect 709211 355953 710211 356009
rect 699322 355836 700322 355892
rect 700922 355836 701922 355892
rect 707610 355881 708610 355937
rect 709211 355881 710211 355937
rect 699322 355534 700322 355606
rect 700922 355534 701922 355606
rect 707610 355579 708610 355651
rect 709211 355579 710211 355651
rect 699392 355523 699426 355534
rect 699460 355523 699494 355534
rect 699528 355523 699562 355534
rect 699596 355523 699630 355534
rect 699664 355523 699698 355534
rect 699732 355523 699766 355534
rect 699800 355523 699834 355534
rect 699868 355523 699902 355534
rect 699936 355523 699970 355534
rect 700004 355523 700038 355534
rect 700072 355523 700106 355534
rect 700140 355523 700174 355534
rect 700208 355523 700242 355534
rect 700276 355523 700310 355534
rect 700934 355523 700968 355534
rect 701002 355523 701036 355534
rect 701070 355523 701104 355534
rect 701138 355523 701172 355534
rect 701206 355523 701240 355534
rect 701274 355523 701308 355534
rect 701342 355523 701376 355534
rect 701410 355523 701444 355534
rect 701478 355523 701512 355534
rect 701546 355523 701580 355534
rect 701614 355523 701648 355534
rect 701682 355523 701716 355534
rect 701750 355523 701784 355534
rect 701818 355523 701852 355534
rect 699392 355513 699450 355523
rect 699460 355513 699518 355523
rect 699528 355513 699586 355523
rect 699596 355513 699654 355523
rect 699664 355513 699722 355523
rect 699732 355513 699790 355523
rect 699800 355513 699858 355523
rect 699868 355513 699926 355523
rect 699936 355513 699994 355523
rect 700004 355513 700062 355523
rect 700072 355513 700130 355523
rect 700140 355513 700198 355523
rect 700208 355513 700266 355523
rect 700276 355513 700334 355523
rect 700934 355513 700992 355523
rect 701002 355513 701060 355523
rect 701070 355513 701128 355523
rect 701138 355513 701196 355523
rect 701206 355513 701264 355523
rect 701274 355513 701332 355523
rect 701342 355513 701400 355523
rect 701410 355513 701468 355523
rect 701478 355513 701536 355523
rect 701546 355513 701604 355523
rect 701614 355513 701672 355523
rect 701682 355513 701740 355523
rect 701750 355513 701808 355523
rect 701818 355513 701876 355523
rect 699368 355489 700334 355513
rect 700910 355489 701876 355513
rect 699392 355474 699416 355489
rect 699460 355474 699484 355489
rect 699528 355474 699552 355489
rect 699596 355474 699620 355489
rect 699664 355474 699688 355489
rect 699732 355474 699756 355489
rect 699800 355474 699824 355489
rect 699868 355474 699892 355489
rect 699936 355474 699960 355489
rect 700004 355474 700028 355489
rect 700072 355474 700096 355489
rect 700140 355474 700164 355489
rect 700208 355474 700232 355489
rect 700276 355474 700300 355489
rect 700934 355474 700958 355489
rect 701002 355474 701026 355489
rect 701070 355474 701094 355489
rect 701138 355474 701162 355489
rect 701206 355474 701230 355489
rect 701274 355474 701298 355489
rect 701342 355474 701366 355489
rect 701410 355474 701434 355489
rect 701478 355474 701502 355489
rect 701546 355474 701570 355489
rect 701614 355474 701638 355489
rect 701682 355474 701706 355489
rect 701750 355474 701774 355489
rect 701818 355474 701842 355489
rect 699322 355319 700322 355474
rect 699322 355285 700334 355319
rect 700922 355309 701922 355474
rect 707610 355319 708610 355379
rect 709211 355319 710211 355379
rect 700910 355285 701922 355309
rect 699322 355274 700322 355285
rect 700922 355274 701922 355285
rect 699392 355261 699416 355274
rect 699460 355261 699484 355274
rect 699528 355261 699552 355274
rect 699596 355261 699620 355274
rect 699664 355261 699688 355274
rect 699732 355261 699756 355274
rect 699800 355261 699824 355274
rect 699868 355261 699892 355274
rect 699936 355261 699960 355274
rect 700004 355261 700028 355274
rect 700072 355261 700096 355274
rect 700140 355261 700164 355274
rect 700208 355261 700232 355274
rect 700276 355261 700300 355274
rect 700934 355261 700958 355274
rect 701002 355261 701026 355274
rect 701070 355261 701094 355274
rect 701138 355261 701162 355274
rect 701206 355261 701230 355274
rect 701274 355261 701298 355274
rect 701342 355261 701366 355274
rect 701410 355261 701434 355274
rect 701478 355261 701502 355274
rect 701546 355261 701570 355274
rect 701614 355261 701638 355274
rect 701682 355261 701706 355274
rect 701750 355261 701774 355274
rect 701818 355261 701842 355274
rect 699322 354916 700322 354972
rect 700922 354916 701922 354972
rect 707610 354961 708610 355017
rect 709211 354961 710211 355017
rect 699322 354844 700322 354900
rect 700922 354844 701922 354900
rect 707610 354889 708610 354945
rect 709211 354889 710211 354945
rect 699322 354542 700322 354614
rect 700922 354542 701922 354614
rect 707610 354587 708610 354659
rect 709211 354587 710211 354659
rect 699392 354531 699426 354542
rect 699460 354531 699494 354542
rect 699528 354531 699562 354542
rect 699596 354531 699630 354542
rect 699664 354531 699698 354542
rect 699732 354531 699766 354542
rect 699800 354531 699834 354542
rect 699868 354531 699902 354542
rect 699936 354531 699970 354542
rect 700004 354531 700038 354542
rect 700072 354531 700106 354542
rect 700140 354531 700174 354542
rect 700208 354531 700242 354542
rect 700276 354531 700310 354542
rect 700934 354531 700968 354542
rect 701002 354531 701036 354542
rect 701070 354531 701104 354542
rect 701138 354531 701172 354542
rect 701206 354531 701240 354542
rect 701274 354531 701308 354542
rect 701342 354531 701376 354542
rect 701410 354531 701444 354542
rect 701478 354531 701512 354542
rect 701546 354531 701580 354542
rect 701614 354531 701648 354542
rect 701682 354531 701716 354542
rect 701750 354531 701784 354542
rect 701818 354531 701852 354542
rect 699392 354521 699450 354531
rect 699460 354521 699518 354531
rect 699528 354521 699586 354531
rect 699596 354521 699654 354531
rect 699664 354521 699722 354531
rect 699732 354521 699790 354531
rect 699800 354521 699858 354531
rect 699868 354521 699926 354531
rect 699936 354521 699994 354531
rect 700004 354521 700062 354531
rect 700072 354521 700130 354531
rect 700140 354521 700198 354531
rect 700208 354521 700266 354531
rect 700276 354521 700334 354531
rect 700934 354521 700992 354531
rect 701002 354521 701060 354531
rect 701070 354521 701128 354531
rect 701138 354521 701196 354531
rect 701206 354521 701264 354531
rect 701274 354521 701332 354531
rect 701342 354521 701400 354531
rect 701410 354521 701468 354531
rect 701478 354521 701536 354531
rect 701546 354521 701604 354531
rect 701614 354521 701672 354531
rect 701682 354521 701740 354531
rect 701750 354521 701808 354531
rect 701818 354521 701876 354531
rect 699368 354497 700334 354521
rect 700910 354497 701876 354521
rect 699392 354482 699416 354497
rect 699460 354482 699484 354497
rect 699528 354482 699552 354497
rect 699596 354482 699620 354497
rect 699664 354482 699688 354497
rect 699732 354482 699756 354497
rect 699800 354482 699824 354497
rect 699868 354482 699892 354497
rect 699936 354482 699960 354497
rect 700004 354482 700028 354497
rect 700072 354482 700096 354497
rect 700140 354482 700164 354497
rect 700208 354482 700232 354497
rect 700276 354482 700300 354497
rect 700934 354482 700958 354497
rect 701002 354482 701026 354497
rect 701070 354482 701094 354497
rect 701138 354482 701162 354497
rect 701206 354482 701230 354497
rect 701274 354482 701298 354497
rect 701342 354482 701366 354497
rect 701410 354482 701434 354497
rect 701478 354482 701502 354497
rect 701546 354482 701570 354497
rect 701614 354482 701638 354497
rect 701682 354482 701706 354497
rect 701750 354482 701774 354497
rect 701818 354482 701842 354497
rect 699322 354327 700322 354482
rect 699322 354293 700334 354327
rect 700922 354317 701922 354482
rect 707610 354327 708610 354387
rect 709211 354327 710211 354387
rect 711541 354345 711629 361461
rect 711892 360200 711942 361200
rect 712062 360200 712112 361200
rect 711892 359079 711942 360079
rect 712062 359079 712112 360079
rect 711892 357958 711942 358958
rect 712062 357958 712112 358958
rect 711892 356848 711942 357848
rect 712062 356848 712112 357848
rect 711892 355727 711942 356727
rect 712062 355727 712112 356727
rect 711892 354606 711942 355606
rect 712062 354606 712112 355606
rect 712409 354371 712431 361485
rect 712469 361459 712487 361501
rect 712499 361459 712505 361467
rect 712499 361455 712511 361459
rect 712539 361455 712557 361501
rect 713640 359461 713674 361785
rect 713750 361772 714750 361822
rect 717367 361820 717413 361853
rect 717367 361819 717379 361820
rect 717401 361819 717413 361820
rect 717401 361809 717600 361819
rect 717401 361786 717413 361809
rect 713750 361562 714750 361612
rect 713750 361446 714750 361496
rect 713750 361230 714750 361358
rect 713750 361014 714750 361070
rect 713750 360798 714750 360926
rect 713750 360588 714750 360638
rect 714478 360585 714750 360588
rect 715486 359931 715536 360931
rect 715696 359931 715824 360931
rect 715912 359931 715962 360931
rect 713641 359345 713663 359461
rect 713640 359309 713674 359345
rect 713750 359314 714750 359364
rect 713750 359158 714750 359214
rect 713750 359002 714750 359130
rect 713750 358846 714750 358974
rect 713750 358690 714750 358746
rect 716425 358709 716725 358721
rect 713750 358534 714750 358662
rect 716425 358596 717425 358646
rect 713750 358378 714750 358506
rect 716425 358440 717425 358568
rect 713750 358222 714750 358350
rect 716425 358284 717425 358340
rect 713750 358072 714750 358122
rect 713750 357956 714750 358006
rect 713750 357800 714750 357928
rect 713750 357644 714750 357772
rect 713750 357488 714750 357616
rect 715354 357587 715404 358187
rect 715504 357587 715560 358187
rect 715660 357587 715716 358187
rect 715816 357587 715872 358187
rect 715972 357587 716022 358187
rect 716425 358128 717425 358256
rect 716425 357978 717425 358028
rect 716425 357862 717425 357912
rect 716425 357706 717425 357834
rect 716425 357550 717425 357606
rect 716425 357394 717425 357522
rect 713750 357332 714750 357388
rect 713750 357176 714750 357304
rect 716425 357244 717425 357294
rect 713750 357020 714750 357148
rect 713750 356870 714750 356920
rect 713750 356742 714750 356792
rect 713750 356586 714750 356642
rect 713750 356436 714750 356486
rect 713750 356320 714350 356370
rect 713750 356164 714350 356292
rect 715510 356191 715560 357191
rect 715660 356191 715788 357191
rect 715816 356191 715944 357191
rect 715972 356191 716022 357191
rect 716425 357128 717425 357178
rect 716425 356972 717425 357028
rect 716425 356822 717425 356872
rect 716425 356706 717425 356756
rect 716425 356550 717425 356678
rect 716425 356394 717425 356522
rect 716425 356238 717425 356366
rect 716425 356082 717425 356210
rect 713750 356008 714350 356064
rect 713750 355852 714350 355980
rect 716425 355932 717425 355982
rect 713750 355696 714350 355752
rect 713750 355446 714350 355496
rect 714565 355443 714765 355455
rect 713750 355330 714750 355380
rect 713750 355120 714750 355170
rect 716413 355092 716447 355150
rect 713750 355004 714750 355054
rect 713750 354794 714750 354844
rect 713750 354678 714750 354728
rect 713750 354468 714750 354518
rect 713750 354352 714750 354402
rect 700910 354293 701922 354317
rect 699322 354282 700322 354293
rect 700922 354282 701922 354293
rect 711541 354311 711633 354345
rect 699392 354269 699416 354282
rect 699460 354269 699484 354282
rect 699528 354269 699552 354282
rect 699596 354269 699620 354282
rect 699664 354269 699688 354282
rect 699732 354269 699756 354282
rect 699800 354269 699824 354282
rect 699868 354269 699892 354282
rect 699936 354269 699960 354282
rect 700004 354269 700028 354282
rect 700072 354269 700096 354282
rect 700140 354269 700164 354282
rect 700208 354269 700232 354282
rect 700276 354269 700300 354282
rect 700934 354269 700958 354282
rect 701002 354269 701026 354282
rect 701070 354269 701094 354282
rect 701138 354269 701162 354282
rect 701206 354269 701230 354282
rect 701274 354269 701298 354282
rect 701342 354269 701366 354282
rect 701410 354269 701434 354282
rect 701478 354269 701502 354282
rect 701546 354269 701570 354282
rect 701614 354269 701638 354282
rect 701682 354269 701706 354282
rect 701750 354269 701774 354282
rect 701818 354269 701842 354282
rect 699322 353924 700322 353980
rect 700922 353924 701922 353980
rect 707610 353969 708610 354025
rect 709211 353969 710211 354025
rect 699322 353852 700322 353908
rect 700922 353852 701922 353908
rect 707610 353897 708610 353953
rect 709211 353897 710211 353953
rect 699322 353550 700322 353622
rect 700922 353550 701922 353622
rect 707610 353595 708610 353667
rect 709211 353595 710211 353667
rect 699392 353539 699426 353550
rect 699460 353539 699494 353550
rect 699528 353539 699562 353550
rect 699596 353539 699630 353550
rect 699664 353539 699698 353550
rect 699732 353539 699766 353550
rect 699800 353539 699834 353550
rect 699868 353539 699902 353550
rect 699936 353539 699970 353550
rect 700004 353539 700038 353550
rect 700072 353539 700106 353550
rect 700140 353539 700174 353550
rect 700208 353539 700242 353550
rect 700276 353539 700310 353550
rect 700934 353539 700968 353550
rect 701002 353539 701036 353550
rect 701070 353539 701104 353550
rect 701138 353539 701172 353550
rect 701206 353539 701240 353550
rect 701274 353539 701308 353550
rect 701342 353539 701376 353550
rect 701410 353539 701444 353550
rect 701478 353539 701512 353550
rect 701546 353539 701580 353550
rect 701614 353539 701648 353550
rect 701682 353539 701716 353550
rect 701750 353539 701784 353550
rect 701818 353539 701852 353550
rect 699392 353529 699450 353539
rect 699460 353529 699518 353539
rect 699528 353529 699586 353539
rect 699596 353529 699654 353539
rect 699664 353529 699722 353539
rect 699732 353529 699790 353539
rect 699800 353529 699858 353539
rect 699868 353529 699926 353539
rect 699936 353529 699994 353539
rect 700004 353529 700062 353539
rect 700072 353529 700130 353539
rect 700140 353529 700198 353539
rect 700208 353529 700266 353539
rect 700276 353529 700334 353539
rect 700934 353529 700992 353539
rect 701002 353529 701060 353539
rect 701070 353529 701128 353539
rect 701138 353529 701196 353539
rect 701206 353529 701264 353539
rect 701274 353529 701332 353539
rect 701342 353529 701400 353539
rect 701410 353529 701468 353539
rect 701478 353529 701536 353539
rect 701546 353529 701604 353539
rect 701614 353529 701672 353539
rect 701682 353529 701740 353539
rect 701750 353529 701808 353539
rect 701818 353529 701876 353539
rect 699368 353505 700334 353529
rect 700910 353505 701876 353529
rect 699392 353490 699416 353505
rect 699460 353490 699484 353505
rect 699528 353490 699552 353505
rect 699596 353490 699620 353505
rect 699664 353490 699688 353505
rect 699732 353490 699756 353505
rect 699800 353490 699824 353505
rect 699868 353490 699892 353505
rect 699936 353490 699960 353505
rect 700004 353490 700028 353505
rect 700072 353490 700096 353505
rect 700140 353490 700164 353505
rect 700208 353490 700232 353505
rect 700276 353490 700300 353505
rect 700934 353490 700958 353505
rect 701002 353490 701026 353505
rect 701070 353490 701094 353505
rect 701138 353490 701162 353505
rect 701206 353490 701230 353505
rect 701274 353490 701298 353505
rect 701342 353490 701366 353505
rect 701410 353490 701434 353505
rect 701478 353490 701502 353505
rect 701546 353490 701570 353505
rect 701614 353490 701638 353505
rect 701682 353490 701706 353505
rect 701750 353490 701774 353505
rect 701818 353490 701842 353505
rect 699322 353335 700322 353490
rect 699322 353301 700334 353335
rect 700922 353325 701922 353490
rect 707610 353335 708610 353395
rect 709211 353335 710211 353395
rect 700910 353301 701922 353325
rect 699322 353290 700322 353301
rect 700922 353290 701922 353301
rect 699392 353277 699416 353290
rect 699460 353277 699484 353290
rect 699528 353277 699552 353290
rect 699596 353277 699620 353290
rect 699664 353277 699688 353290
rect 699732 353277 699756 353290
rect 699800 353277 699824 353290
rect 699868 353277 699892 353290
rect 699936 353277 699960 353290
rect 700004 353277 700028 353290
rect 700072 353277 700096 353290
rect 700140 353277 700164 353290
rect 700208 353277 700232 353290
rect 700276 353277 700300 353290
rect 700934 353277 700958 353290
rect 701002 353277 701026 353290
rect 701070 353277 701094 353290
rect 701138 353277 701162 353290
rect 701206 353277 701230 353290
rect 701274 353277 701298 353290
rect 701342 353277 701366 353290
rect 701410 353277 701434 353290
rect 701478 353277 701502 353290
rect 701546 353277 701570 353290
rect 701614 353277 701638 353290
rect 701682 353277 701706 353290
rect 701750 353277 701774 353290
rect 701818 353277 701842 353290
rect 699322 352932 700322 352988
rect 700922 352932 701922 352988
rect 707610 352977 708610 353033
rect 709211 352977 710211 353033
rect 699322 352860 700322 352916
rect 700922 352860 701922 352916
rect 707610 352905 708610 352961
rect 709211 352905 710211 352961
rect 699322 352558 700322 352630
rect 700922 352558 701922 352630
rect 707610 352603 708610 352675
rect 709211 352603 710211 352675
rect 699392 352547 699426 352558
rect 699460 352547 699494 352558
rect 699528 352547 699562 352558
rect 699596 352547 699630 352558
rect 699664 352547 699698 352558
rect 699732 352547 699766 352558
rect 699800 352547 699834 352558
rect 699868 352547 699902 352558
rect 699936 352547 699970 352558
rect 700004 352547 700038 352558
rect 700072 352547 700106 352558
rect 700140 352547 700174 352558
rect 700208 352547 700242 352558
rect 700276 352547 700310 352558
rect 700934 352547 700968 352558
rect 701002 352547 701036 352558
rect 701070 352547 701104 352558
rect 701138 352547 701172 352558
rect 701206 352547 701240 352558
rect 701274 352547 701308 352558
rect 701342 352547 701376 352558
rect 701410 352547 701444 352558
rect 701478 352547 701512 352558
rect 701546 352547 701580 352558
rect 701614 352547 701648 352558
rect 701682 352547 701716 352558
rect 701750 352547 701784 352558
rect 701818 352547 701852 352558
rect 699392 352537 699450 352547
rect 699460 352537 699518 352547
rect 699528 352537 699586 352547
rect 699596 352537 699654 352547
rect 699664 352537 699722 352547
rect 699732 352537 699790 352547
rect 699800 352537 699858 352547
rect 699868 352537 699926 352547
rect 699936 352537 699994 352547
rect 700004 352537 700062 352547
rect 700072 352537 700130 352547
rect 700140 352537 700198 352547
rect 700208 352537 700266 352547
rect 700276 352537 700334 352547
rect 700934 352537 700992 352547
rect 701002 352537 701060 352547
rect 701070 352537 701128 352547
rect 701138 352537 701196 352547
rect 701206 352537 701264 352547
rect 701274 352537 701332 352547
rect 701342 352537 701400 352547
rect 701410 352537 701468 352547
rect 701478 352537 701536 352547
rect 701546 352537 701604 352547
rect 701614 352537 701672 352547
rect 701682 352537 701740 352547
rect 701750 352537 701808 352547
rect 701818 352537 701876 352547
rect 699368 352513 700334 352537
rect 700910 352513 701876 352537
rect 699392 352498 699416 352513
rect 699460 352498 699484 352513
rect 699528 352498 699552 352513
rect 699596 352498 699620 352513
rect 699664 352498 699688 352513
rect 699732 352498 699756 352513
rect 699800 352498 699824 352513
rect 699868 352498 699892 352513
rect 699936 352498 699960 352513
rect 700004 352498 700028 352513
rect 700072 352498 700096 352513
rect 700140 352498 700164 352513
rect 700208 352498 700232 352513
rect 700276 352498 700300 352513
rect 700934 352498 700958 352513
rect 701002 352498 701026 352513
rect 701070 352498 701094 352513
rect 701138 352498 701162 352513
rect 701206 352498 701230 352513
rect 701274 352498 701298 352513
rect 701342 352498 701366 352513
rect 701410 352498 701434 352513
rect 701478 352498 701502 352513
rect 701546 352498 701570 352513
rect 701614 352498 701638 352513
rect 701682 352498 701706 352513
rect 701750 352498 701774 352513
rect 701818 352498 701842 352513
rect 699322 352343 700322 352498
rect 699322 352309 700334 352343
rect 700922 352333 701922 352498
rect 707610 352343 708610 352403
rect 709211 352343 710211 352403
rect 700910 352309 701922 352333
rect 699322 352298 700322 352309
rect 700922 352298 701922 352309
rect 699392 352285 699416 352298
rect 699460 352285 699484 352298
rect 699528 352285 699552 352298
rect 699596 352285 699620 352298
rect 699664 352285 699688 352298
rect 699732 352285 699756 352298
rect 699800 352285 699824 352298
rect 699868 352285 699892 352298
rect 699936 352285 699960 352298
rect 700004 352285 700028 352298
rect 700072 352285 700096 352298
rect 700140 352285 700164 352298
rect 700208 352285 700232 352298
rect 700276 352285 700300 352298
rect 700934 352285 700958 352298
rect 701002 352285 701026 352298
rect 701070 352285 701094 352298
rect 701138 352285 701162 352298
rect 701206 352285 701230 352298
rect 701274 352285 701298 352298
rect 701342 352285 701366 352298
rect 701410 352285 701434 352298
rect 701478 352285 701502 352298
rect 701546 352285 701570 352298
rect 701614 352285 701638 352298
rect 701682 352285 701706 352298
rect 701750 352285 701774 352298
rect 701818 352285 701842 352298
rect 699322 351940 700322 351996
rect 700922 351940 701922 351996
rect 707610 351985 708610 352041
rect 709211 351985 710211 352041
rect 699322 351868 700322 351924
rect 700922 351868 701922 351924
rect 707610 351913 708610 351969
rect 709211 351913 710211 351969
rect 699322 351566 700322 351638
rect 700922 351566 701922 351638
rect 707610 351611 708610 351683
rect 709211 351611 710211 351683
rect 699392 351555 699426 351566
rect 699460 351555 699494 351566
rect 699528 351555 699562 351566
rect 699596 351555 699630 351566
rect 699664 351555 699698 351566
rect 699732 351555 699766 351566
rect 699800 351555 699834 351566
rect 699868 351555 699902 351566
rect 699936 351555 699970 351566
rect 700004 351555 700038 351566
rect 700072 351555 700106 351566
rect 700140 351555 700174 351566
rect 700208 351555 700242 351566
rect 700276 351555 700310 351566
rect 700934 351555 700968 351566
rect 701002 351555 701036 351566
rect 701070 351555 701104 351566
rect 701138 351555 701172 351566
rect 701206 351555 701240 351566
rect 701274 351555 701308 351566
rect 701342 351555 701376 351566
rect 701410 351555 701444 351566
rect 701478 351555 701512 351566
rect 701546 351555 701580 351566
rect 701614 351555 701648 351566
rect 701682 351555 701716 351566
rect 701750 351555 701784 351566
rect 701818 351555 701852 351566
rect 699392 351545 699450 351555
rect 699460 351545 699518 351555
rect 699528 351545 699586 351555
rect 699596 351545 699654 351555
rect 699664 351545 699722 351555
rect 699732 351545 699790 351555
rect 699800 351545 699858 351555
rect 699868 351545 699926 351555
rect 699936 351545 699994 351555
rect 700004 351545 700062 351555
rect 700072 351545 700130 351555
rect 700140 351545 700198 351555
rect 700208 351545 700266 351555
rect 700276 351545 700334 351555
rect 700934 351545 700992 351555
rect 701002 351545 701060 351555
rect 701070 351545 701128 351555
rect 701138 351545 701196 351555
rect 701206 351545 701264 351555
rect 701274 351545 701332 351555
rect 701342 351545 701400 351555
rect 701410 351545 701468 351555
rect 701478 351545 701536 351555
rect 701546 351545 701604 351555
rect 701614 351545 701672 351555
rect 701682 351545 701740 351555
rect 701750 351545 701808 351555
rect 701818 351545 701876 351555
rect 699368 351521 700334 351545
rect 700910 351521 701876 351545
rect 699392 351506 699416 351521
rect 699460 351506 699484 351521
rect 699528 351506 699552 351521
rect 699596 351506 699620 351521
rect 699664 351506 699688 351521
rect 699732 351506 699756 351521
rect 699800 351506 699824 351521
rect 699868 351506 699892 351521
rect 699936 351506 699960 351521
rect 700004 351506 700028 351521
rect 700072 351506 700096 351521
rect 700140 351506 700164 351521
rect 700208 351506 700232 351521
rect 700276 351506 700300 351521
rect 700934 351506 700958 351521
rect 701002 351506 701026 351521
rect 701070 351506 701094 351521
rect 701138 351506 701162 351521
rect 701206 351506 701230 351521
rect 701274 351506 701298 351521
rect 701342 351506 701366 351521
rect 701410 351506 701434 351521
rect 701478 351506 701502 351521
rect 701546 351506 701570 351521
rect 701614 351506 701638 351521
rect 701682 351506 701706 351521
rect 701750 351506 701774 351521
rect 701818 351506 701842 351521
rect 699322 351351 700322 351506
rect 699322 351317 700334 351351
rect 700922 351341 701922 351506
rect 705107 351360 705173 351376
rect 707610 351351 708610 351411
rect 709211 351351 710211 351411
rect 700910 351317 701922 351341
rect 699322 351306 700322 351317
rect 700922 351306 701922 351317
rect 699392 351293 699416 351306
rect 699460 351293 699484 351306
rect 699528 351293 699552 351306
rect 699596 351293 699620 351306
rect 699664 351293 699688 351306
rect 699732 351293 699756 351306
rect 699800 351293 699824 351306
rect 699868 351293 699892 351306
rect 699936 351293 699960 351306
rect 700004 351293 700028 351306
rect 700072 351293 700096 351306
rect 700140 351293 700164 351306
rect 700208 351293 700232 351306
rect 700276 351293 700300 351306
rect 700934 351293 700958 351306
rect 701002 351293 701026 351306
rect 701070 351293 701094 351306
rect 701138 351293 701162 351306
rect 701206 351293 701230 351306
rect 701274 351293 701298 351306
rect 701342 351293 701366 351306
rect 701410 351293 701434 351306
rect 701478 351293 701502 351306
rect 701546 351293 701570 351306
rect 701614 351293 701638 351306
rect 701682 351293 701706 351306
rect 701750 351293 701774 351306
rect 701818 351293 701842 351306
rect 699322 350948 700322 351004
rect 700922 350948 701922 351004
rect 707610 350993 708610 351049
rect 709211 350993 710211 351049
rect 699322 350876 700322 350932
rect 700922 350876 701922 350932
rect 707610 350921 708610 350977
rect 709211 350921 710211 350977
rect 699322 350574 700322 350646
rect 700922 350574 701922 350646
rect 707610 350619 708610 350691
rect 709211 350619 710211 350691
rect 699392 350563 699426 350574
rect 699460 350563 699494 350574
rect 699528 350563 699562 350574
rect 699596 350563 699630 350574
rect 699664 350563 699698 350574
rect 699732 350563 699766 350574
rect 699800 350563 699834 350574
rect 699868 350563 699902 350574
rect 699936 350563 699970 350574
rect 700004 350563 700038 350574
rect 700072 350563 700106 350574
rect 700140 350563 700174 350574
rect 700208 350563 700242 350574
rect 700276 350563 700310 350574
rect 700934 350563 700968 350574
rect 701002 350563 701036 350574
rect 701070 350563 701104 350574
rect 701138 350563 701172 350574
rect 701206 350563 701240 350574
rect 701274 350563 701308 350574
rect 701342 350563 701376 350574
rect 701410 350563 701444 350574
rect 701478 350563 701512 350574
rect 701546 350563 701580 350574
rect 701614 350563 701648 350574
rect 701682 350563 701716 350574
rect 701750 350563 701784 350574
rect 701818 350563 701852 350574
rect 699392 350553 699450 350563
rect 699460 350553 699518 350563
rect 699528 350553 699586 350563
rect 699596 350553 699654 350563
rect 699664 350553 699722 350563
rect 699732 350553 699790 350563
rect 699800 350553 699858 350563
rect 699868 350553 699926 350563
rect 699936 350553 699994 350563
rect 700004 350553 700062 350563
rect 700072 350553 700130 350563
rect 700140 350553 700198 350563
rect 700208 350553 700266 350563
rect 700276 350553 700334 350563
rect 700934 350553 700992 350563
rect 701002 350553 701060 350563
rect 701070 350553 701128 350563
rect 701138 350553 701196 350563
rect 701206 350553 701264 350563
rect 701274 350553 701332 350563
rect 701342 350553 701400 350563
rect 701410 350553 701468 350563
rect 701478 350553 701536 350563
rect 701546 350553 701604 350563
rect 701614 350553 701672 350563
rect 701682 350553 701740 350563
rect 701750 350553 701808 350563
rect 701818 350553 701876 350563
rect 699368 350529 700334 350553
rect 700910 350529 701876 350553
rect 699392 350514 699416 350529
rect 699460 350514 699484 350529
rect 699528 350514 699552 350529
rect 699596 350514 699620 350529
rect 699664 350514 699688 350529
rect 699732 350514 699756 350529
rect 699800 350514 699824 350529
rect 699868 350514 699892 350529
rect 699936 350514 699960 350529
rect 700004 350514 700028 350529
rect 700072 350514 700096 350529
rect 700140 350514 700164 350529
rect 700208 350514 700232 350529
rect 700276 350514 700300 350529
rect 700934 350514 700958 350529
rect 701002 350514 701026 350529
rect 701070 350514 701094 350529
rect 701138 350514 701162 350529
rect 701206 350514 701230 350529
rect 701274 350514 701298 350529
rect 701342 350514 701366 350529
rect 701410 350514 701434 350529
rect 701478 350514 701502 350529
rect 701546 350514 701570 350529
rect 701614 350514 701638 350529
rect 701682 350514 701706 350529
rect 701750 350514 701774 350529
rect 701818 350514 701842 350529
rect 699322 350359 700322 350514
rect 699322 350325 700334 350359
rect 700922 350349 701922 350514
rect 707610 350359 708610 350419
rect 709211 350359 710211 350419
rect 700910 350325 701922 350349
rect 699322 350314 700322 350325
rect 700922 350314 701922 350325
rect 699392 350301 699416 350314
rect 699460 350301 699484 350314
rect 699528 350301 699552 350314
rect 699596 350301 699620 350314
rect 699664 350301 699688 350314
rect 699732 350301 699756 350314
rect 699800 350301 699824 350314
rect 699868 350301 699892 350314
rect 699936 350301 699960 350314
rect 700004 350301 700028 350314
rect 700072 350301 700096 350314
rect 700140 350301 700164 350314
rect 700208 350301 700232 350314
rect 700276 350301 700300 350314
rect 700934 350301 700958 350314
rect 701002 350301 701026 350314
rect 701070 350301 701094 350314
rect 701138 350301 701162 350314
rect 701206 350301 701230 350314
rect 701274 350301 701298 350314
rect 701342 350301 701366 350314
rect 701410 350301 701434 350314
rect 701478 350301 701502 350314
rect 701546 350301 701570 350314
rect 701614 350301 701638 350314
rect 701682 350301 701706 350314
rect 701750 350301 701774 350314
rect 701818 350301 701842 350314
rect 709211 350148 710211 350152
rect 707574 350099 707610 350134
rect 708610 350099 708646 350134
rect 707574 350098 708646 350099
rect 707574 350057 707610 350098
rect 708610 350057 708646 350098
rect 699322 349956 700322 350012
rect 700922 349956 701922 350012
rect 707574 350001 708646 350057
rect 707574 349964 707610 350001
rect 708610 349964 708646 350001
rect 707574 349959 708646 349964
rect 699322 349884 700322 349940
rect 700922 349884 701922 349940
rect 707574 349924 707610 349959
rect 708610 349924 708646 349959
rect 709175 350098 710247 350134
rect 709175 350057 709211 350098
rect 710211 350057 710247 350098
rect 709175 350001 710247 350057
rect 709175 349964 709211 350001
rect 710211 349964 710247 350001
rect 709175 349936 710247 349964
rect 709175 349924 709211 349936
rect 710211 349924 710247 349936
rect 707610 349713 708610 349785
rect 709211 349713 710211 349785
rect 699322 349623 700322 349673
rect 700922 349623 701922 349673
rect 707610 349523 708610 349617
rect 707610 349513 708644 349523
rect 709211 349513 710211 349591
rect 711541 349437 711629 354311
rect 713750 354136 714750 354264
rect 716417 354152 717417 354202
rect 711892 353049 711942 354049
rect 712062 353049 712112 354049
rect 713750 353920 714750 354048
rect 716417 353996 717417 354052
rect 716417 353846 717417 353896
rect 713750 353704 714750 353832
rect 716417 353730 717017 353780
rect 716417 353580 717017 353630
rect 713750 353488 714750 353544
rect 716417 353464 717417 353514
rect 713750 353272 714750 353400
rect 716417 353308 717417 353364
rect 713750 353056 714750 353184
rect 716417 353152 717417 353280
rect 716417 352996 717417 353052
rect 711892 351928 711942 352928
rect 712062 351928 712112 352928
rect 713750 352840 714750 352968
rect 716417 352840 717417 352968
rect 713750 352624 714750 352752
rect 716417 352684 717417 352740
rect 716417 352474 717417 352524
rect 713750 352408 714750 352464
rect 716417 352308 717417 352358
rect 713750 352192 714750 352248
rect 716417 352152 717417 352280
rect 713750 351976 714750 352104
rect 716417 351996 717417 352052
rect 711892 350807 711942 351807
rect 712062 350807 712112 351807
rect 713750 351760 714750 351888
rect 716417 351780 717417 351836
rect 713750 351544 714750 351672
rect 716417 351570 717417 351620
rect 713750 351328 714750 351456
rect 716417 351454 717417 351504
rect 716417 351298 717417 351426
rect 713750 351118 714750 351168
rect 716417 351148 717417 351198
rect 711892 349697 711942 350697
rect 712062 349697 712112 350697
rect 714686 350357 714794 350424
rect 714645 350323 714794 350357
rect 716071 350357 716074 350358
rect 716071 350356 716072 350357
rect 716073 350356 716074 350357
rect 716071 350355 716074 350356
rect 716208 350357 716211 350358
rect 716208 350356 716209 350357
rect 716210 350356 716211 350357
rect 716208 350355 716211 350356
rect 714964 350247 715998 350329
rect 716284 350247 717318 350329
rect 705107 349336 705173 349352
rect 711541 349302 711633 349437
rect 714175 349398 714225 349998
rect 714425 349398 714475 349998
rect 711579 349301 711595 349302
rect 714781 349191 714863 350226
rect 715134 349955 715828 350037
rect 714686 349123 714863 349191
rect 714645 349089 714863 349123
rect 680215 348880 680815 348936
rect 686719 348893 686739 348917
rect 686743 348893 686753 348917
rect 686719 348859 686757 348893
rect 686719 348822 686739 348859
rect 686743 348822 686753 348859
rect 692428 348850 693028 348978
rect 698017 348947 698210 348983
rect 698084 348935 698210 348947
rect 702756 348959 703645 348983
rect 702756 348935 702853 348959
rect 698084 348828 702853 348935
rect 686719 348788 686757 348822
rect 680215 348704 680815 348760
rect 686719 348751 686739 348788
rect 686743 348751 686753 348788
rect 686719 348741 686757 348751
rect 686699 348717 686767 348741
rect 686719 348704 686739 348717
rect 686743 348704 686753 348717
rect 686719 348695 686753 348704
rect 686719 348693 686743 348695
rect 692428 348694 693028 348750
rect 686685 348656 686709 348680
rect 686743 348656 686767 348680
rect 678799 348503 679399 348553
rect 680215 348534 680815 348584
rect 692428 348538 693028 348666
rect 680593 348531 680815 348534
rect 682009 348501 682069 348516
rect 682024 348465 682054 348501
rect 683708 348387 684308 348437
rect 678799 348327 679399 348383
rect 692428 348382 693028 348510
rect 714781 348308 714863 349089
rect 715063 348609 715145 349915
rect 715342 349752 715382 349792
rect 715582 349752 715622 349792
rect 715289 348777 715339 349719
rect 715382 349668 715422 349752
rect 715542 349668 715582 349752
rect 715633 348777 715683 349719
rect 715382 348672 715422 348756
rect 715542 348672 715582 348756
rect 715342 348632 715382 348672
rect 715582 348632 715622 348672
rect 715815 348609 715897 349915
rect 715134 348387 715828 348469
rect 716100 348308 716182 350226
rect 716454 349955 717148 350037
rect 716385 348609 716467 349915
rect 716660 349752 716700 349792
rect 716900 349752 716940 349792
rect 716599 348777 716649 349719
rect 716700 349668 716740 349752
rect 716860 349668 716900 349752
rect 716943 348777 716993 349719
rect 716700 348672 716740 348756
rect 716860 348672 716900 348756
rect 716660 348632 716700 348672
rect 716900 348632 716940 348672
rect 717137 348609 717219 349915
rect 716454 348387 717148 348469
rect 717419 348308 717501 350226
rect 683708 348237 684308 348287
rect 692428 348232 693028 348282
rect 678799 348157 679399 348207
rect 684565 348160 684790 348168
rect 696597 348000 696600 348120
rect 714964 348095 715998 348177
rect 716284 348095 717318 348177
rect 21000 321000 21003 321120
rect 282 320623 1316 320705
rect 1602 320623 2636 320705
rect 32810 320662 33035 320670
rect 38201 320593 38801 320643
rect 24572 320518 25172 320568
rect 33292 320513 33892 320563
rect 99 318574 181 320492
rect 452 320331 1146 320413
rect 381 318885 463 320191
rect 660 320128 700 320168
rect 900 320128 940 320168
rect 700 320044 740 320128
rect 860 320044 900 320128
rect 607 319081 657 320023
rect 700 319048 740 319132
rect 860 319048 900 319132
rect 951 319081 1001 320023
rect 660 319008 700 319048
rect 900 319008 940 319048
rect 1133 318885 1215 320191
rect 452 318763 1146 318845
rect 1418 318574 1500 320492
rect 1772 320331 2466 320413
rect 1703 318885 1785 320191
rect 1978 320128 2018 320168
rect 2218 320128 2258 320168
rect 2018 320044 2058 320128
rect 2178 320044 2218 320128
rect 1917 319081 1967 320023
rect 2018 319048 2058 319132
rect 2178 319048 2218 319132
rect 2261 319081 2311 320023
rect 1978 319008 2018 319048
rect 2218 319008 2258 319048
rect 2455 318885 2537 320191
rect 2737 319779 2819 320492
rect 24572 320362 25172 320490
rect 38201 320417 38801 320473
rect 33292 320363 33892 320413
rect 24572 320206 25172 320334
rect 35546 320299 35576 320335
rect 36785 320329 36935 320341
rect 35531 320284 35591 320299
rect 36785 320216 37385 320266
rect 38201 320247 38801 320297
rect 30833 320120 30857 320144
rect 30891 320120 30915 320144
rect 24572 320050 25172 320106
rect 30857 320105 30881 320107
rect 30857 320096 30887 320105
rect 30867 320083 30887 320096
rect 30891 320083 30907 320120
rect 30833 320059 30857 320083
rect 30867 320049 30911 320083
rect 14747 319865 19516 319972
rect 24572 319894 25172 320022
rect 30867 320012 30887 320049
rect 30891 320012 30907 320049
rect 36785 320040 37385 320096
rect 30867 319978 30911 320012
rect 30867 319941 30887 319978
rect 30891 319941 30907 319978
rect 30867 319907 30911 319941
rect 30867 319883 30887 319907
rect 30891 319883 30907 319907
rect 14747 319841 14844 319865
rect 13955 319817 14844 319841
rect 19390 319853 19516 319865
rect 19390 319841 19583 319853
rect 19390 319817 19605 319841
rect 19639 319817 19673 319841
rect 19707 319817 19741 319841
rect 19775 319817 19809 319841
rect 19843 319817 19877 319841
rect 19911 319817 19945 319841
rect 19979 319817 20013 319841
rect 20047 319817 20081 319841
rect 20115 319817 20149 319841
rect 20183 319817 20217 319841
rect 20251 319817 20285 319841
rect 20319 319817 20353 319841
rect 20387 319817 20421 319841
rect 20455 319817 20489 319841
rect 20523 319817 20557 319841
rect 20591 319817 20625 319841
rect 20659 319817 20693 319841
rect 2737 319711 2914 319779
rect 1772 318763 2466 318845
rect 2737 318574 2819 319711
rect 2848 319677 2955 319711
rect 6005 319498 6021 319499
rect 3125 318802 3175 319402
rect 3375 318802 3425 319402
rect 5967 319363 6059 319498
rect 12427 319448 12493 319464
rect 282 318471 1316 318553
rect 1602 318471 2636 318553
rect 2806 318477 2914 318545
rect 1389 318444 1392 318445
rect 1389 318443 1390 318444
rect 1391 318443 1392 318444
rect 1389 318442 1392 318443
rect 1526 318444 1529 318445
rect 1526 318443 1527 318444
rect 1528 318443 1529 318444
rect 2848 318443 2955 318477
rect 1526 318442 1529 318443
rect 5488 318103 5538 319103
rect 5658 318103 5708 319103
rect 183 317602 1183 317652
rect 2850 317632 3850 317682
rect 183 317446 1183 317574
rect 2850 317416 3850 317544
rect 183 317296 1183 317346
rect 183 317180 1183 317230
rect 2850 317200 3850 317328
rect 183 316964 1183 317020
rect 2850 316984 3850 317112
rect 5488 316993 5538 317993
rect 5658 316993 5708 317993
rect 183 316748 1183 316804
rect 2850 316768 3850 316896
rect 183 316592 1183 316720
rect 2850 316552 3850 316608
rect 183 316442 1183 316492
rect 2850 316336 3850 316392
rect 183 316276 1183 316326
rect 2850 316120 3850 316248
rect 183 316060 1183 316116
rect 183 315904 1183 316032
rect 2850 315904 3850 316032
rect 5488 315872 5538 316872
rect 5658 315872 5708 316872
rect 183 315748 1183 315804
rect 183 315592 1183 315720
rect 2850 315688 3850 315816
rect 183 315436 1183 315492
rect 2850 315472 3850 315600
rect 183 315286 1183 315336
rect 2850 315256 3850 315312
rect 583 315170 1183 315220
rect 583 315020 1183 315070
rect 2850 315040 3850 315168
rect 183 314904 1183 314954
rect 2850 314824 3850 314952
rect 183 314748 1183 314804
rect 5488 314751 5538 315751
rect 5658 314751 5708 315751
rect 183 314598 1183 314648
rect 2850 314608 3850 314736
rect 5971 314489 6059 319363
rect 7406 319287 7440 319321
rect 7477 319287 7511 319321
rect 7551 319287 7585 319321
rect 7622 319287 7656 319321
rect 7696 319287 7730 319321
rect 7767 319287 7801 319321
rect 7841 319287 7875 319321
rect 7912 319287 7946 319321
rect 7986 319287 8020 319321
rect 8057 319287 8091 319321
rect 8131 319287 8165 319321
rect 8202 319287 8236 319321
rect 8296 319287 8330 319321
rect 8381 319311 8423 319321
rect 8381 319287 8389 319311
rect 8415 319287 8423 319311
rect 8956 319311 8996 319321
rect 8956 319287 8962 319311
rect 8990 319287 8996 319311
rect 9044 319287 9078 319321
rect 9120 319287 9154 319321
rect 9197 319287 9231 319321
rect 9291 319287 9325 319321
rect 9362 319287 9396 319321
rect 9436 319287 9470 319321
rect 9507 319287 9541 319321
rect 9581 319287 9615 319321
rect 9652 319287 9686 319321
rect 9726 319287 9760 319321
rect 9797 319287 9831 319321
rect 9871 319287 9905 319321
rect 9942 319287 9976 319321
rect 7389 319277 7406 319287
rect 7440 319277 7477 319287
rect 7511 319277 7551 319287
rect 7585 319277 7622 319287
rect 7656 319277 7696 319287
rect 7730 319277 7767 319287
rect 7801 319277 7841 319287
rect 7875 319277 7912 319287
rect 7946 319277 7986 319287
rect 8020 319277 8057 319287
rect 8091 319277 8131 319287
rect 8165 319277 8202 319287
rect 8236 319277 8296 319287
rect 8330 319277 8381 319287
rect 8389 319277 8423 319287
rect 8990 319277 9044 319287
rect 9078 319277 9120 319287
rect 9154 319277 9197 319287
rect 9231 319277 9291 319287
rect 9325 319277 9362 319287
rect 9396 319277 9436 319287
rect 9470 319277 9507 319287
rect 9541 319277 9581 319287
rect 9615 319277 9652 319287
rect 9686 319277 9726 319287
rect 9760 319277 9797 319287
rect 9831 319277 9871 319287
rect 9905 319277 9942 319287
rect 9976 319277 9990 319287
rect 7389 319209 8389 319277
rect 8990 319183 9990 319277
rect 7389 319087 8389 319147
rect 8990 319087 9990 319147
rect 15678 319127 16678 319177
rect 17278 319127 18278 319177
rect 7353 318864 7389 318876
rect 8389 318864 8425 318876
rect 7353 318840 8425 318864
rect 7353 318799 7389 318840
rect 8389 318799 8425 318840
rect 7353 318743 8425 318799
rect 7353 318706 7389 318743
rect 8389 318706 8425 318743
rect 7353 318666 8425 318706
rect 8954 318841 8990 318876
rect 9990 318841 10026 318876
rect 15678 318860 16678 318916
rect 17278 318860 18278 318916
rect 8954 318840 10026 318841
rect 8954 318799 8990 318840
rect 9990 318799 10026 318840
rect 8954 318743 10026 318799
rect 15678 318788 16678 318844
rect 17278 318788 18278 318844
rect 8954 318706 8990 318743
rect 9990 318706 10026 318743
rect 8954 318701 10026 318706
rect 8954 318666 8990 318701
rect 9990 318666 10026 318701
rect 7389 318441 8389 318513
rect 8990 318441 9990 318513
rect 15678 318486 16678 318558
rect 17278 318486 18278 318558
rect 15748 318475 15782 318486
rect 15816 318475 15850 318486
rect 15884 318475 15918 318486
rect 15952 318475 15986 318486
rect 16020 318475 16054 318486
rect 16088 318475 16122 318486
rect 16156 318475 16190 318486
rect 16224 318475 16258 318486
rect 16292 318475 16326 318486
rect 16360 318475 16394 318486
rect 16428 318475 16462 318486
rect 16496 318475 16530 318486
rect 16564 318475 16598 318486
rect 16632 318475 16666 318486
rect 17290 318475 17324 318486
rect 17358 318475 17392 318486
rect 17426 318475 17460 318486
rect 17494 318475 17528 318486
rect 17562 318475 17596 318486
rect 17630 318475 17664 318486
rect 17698 318475 17732 318486
rect 17766 318475 17800 318486
rect 17834 318475 17868 318486
rect 17902 318475 17936 318486
rect 17970 318475 18004 318486
rect 18038 318475 18072 318486
rect 18106 318475 18140 318486
rect 18174 318475 18208 318486
rect 15748 318465 15806 318475
rect 15816 318465 15874 318475
rect 15884 318465 15942 318475
rect 15952 318465 16010 318475
rect 16020 318465 16078 318475
rect 16088 318465 16146 318475
rect 16156 318465 16214 318475
rect 16224 318465 16282 318475
rect 16292 318465 16350 318475
rect 16360 318465 16418 318475
rect 16428 318465 16486 318475
rect 16496 318465 16554 318475
rect 16564 318465 16622 318475
rect 16632 318465 16690 318475
rect 17290 318465 17348 318475
rect 17358 318465 17416 318475
rect 17426 318465 17484 318475
rect 17494 318465 17552 318475
rect 17562 318465 17620 318475
rect 17630 318465 17688 318475
rect 17698 318465 17756 318475
rect 17766 318465 17824 318475
rect 17834 318465 17892 318475
rect 17902 318465 17960 318475
rect 17970 318465 18028 318475
rect 18038 318465 18096 318475
rect 18106 318465 18164 318475
rect 18174 318465 18232 318475
rect 15724 318441 16690 318465
rect 17266 318441 18232 318465
rect 15748 318426 15772 318441
rect 15816 318426 15840 318441
rect 15884 318426 15908 318441
rect 15952 318426 15976 318441
rect 16020 318426 16044 318441
rect 16088 318426 16112 318441
rect 16156 318426 16180 318441
rect 16224 318426 16248 318441
rect 16292 318426 16316 318441
rect 16360 318426 16384 318441
rect 16428 318426 16452 318441
rect 16496 318426 16520 318441
rect 16564 318426 16588 318441
rect 16632 318426 16656 318441
rect 17290 318426 17314 318441
rect 17358 318426 17382 318441
rect 17426 318426 17450 318441
rect 17494 318426 17518 318441
rect 17562 318426 17586 318441
rect 17630 318426 17654 318441
rect 17698 318426 17722 318441
rect 17766 318426 17790 318441
rect 17834 318426 17858 318441
rect 17902 318426 17926 318441
rect 17970 318426 17994 318441
rect 18038 318426 18062 318441
rect 18106 318426 18130 318441
rect 18174 318426 18198 318441
rect 15678 318271 16678 318426
rect 7389 318181 8389 318241
rect 8990 318181 9990 318241
rect 15678 318237 16690 318271
rect 17278 318261 18278 318426
rect 17266 318237 18278 318261
rect 15678 318226 16678 318237
rect 17278 318226 18278 318237
rect 15748 318213 15772 318226
rect 15816 318213 15840 318226
rect 15884 318213 15908 318226
rect 15952 318213 15976 318226
rect 16020 318213 16044 318226
rect 16088 318213 16112 318226
rect 16156 318213 16180 318226
rect 16224 318213 16248 318226
rect 16292 318213 16316 318226
rect 16360 318213 16384 318226
rect 16428 318213 16452 318226
rect 16496 318213 16520 318226
rect 16564 318213 16588 318226
rect 16632 318213 16656 318226
rect 17290 318213 17314 318226
rect 17358 318213 17382 318226
rect 17426 318213 17450 318226
rect 17494 318213 17518 318226
rect 17562 318213 17586 318226
rect 17630 318213 17654 318226
rect 17698 318213 17722 318226
rect 17766 318213 17790 318226
rect 17834 318213 17858 318226
rect 17902 318213 17926 318226
rect 17970 318213 17994 318226
rect 18038 318213 18062 318226
rect 18106 318213 18130 318226
rect 18174 318213 18198 318226
rect 7389 317823 8389 317879
rect 8990 317823 9990 317879
rect 15678 317868 16678 317924
rect 17278 317868 18278 317924
rect 7389 317751 8389 317807
rect 8990 317751 9990 317807
rect 15678 317796 16678 317852
rect 17278 317796 18278 317852
rect 7389 317449 8389 317521
rect 8990 317449 9990 317521
rect 15678 317494 16678 317566
rect 17278 317494 18278 317566
rect 15748 317483 15782 317494
rect 15816 317483 15850 317494
rect 15884 317483 15918 317494
rect 15952 317483 15986 317494
rect 16020 317483 16054 317494
rect 16088 317483 16122 317494
rect 16156 317483 16190 317494
rect 16224 317483 16258 317494
rect 16292 317483 16326 317494
rect 16360 317483 16394 317494
rect 16428 317483 16462 317494
rect 16496 317483 16530 317494
rect 16564 317483 16598 317494
rect 16632 317483 16666 317494
rect 17290 317483 17324 317494
rect 17358 317483 17392 317494
rect 17426 317483 17460 317494
rect 17494 317483 17528 317494
rect 17562 317483 17596 317494
rect 17630 317483 17664 317494
rect 17698 317483 17732 317494
rect 17766 317483 17800 317494
rect 17834 317483 17868 317494
rect 17902 317483 17936 317494
rect 17970 317483 18004 317494
rect 18038 317483 18072 317494
rect 18106 317483 18140 317494
rect 18174 317483 18208 317494
rect 15748 317473 15806 317483
rect 15816 317473 15874 317483
rect 15884 317473 15942 317483
rect 15952 317473 16010 317483
rect 16020 317473 16078 317483
rect 16088 317473 16146 317483
rect 16156 317473 16214 317483
rect 16224 317473 16282 317483
rect 16292 317473 16350 317483
rect 16360 317473 16418 317483
rect 16428 317473 16486 317483
rect 16496 317473 16554 317483
rect 16564 317473 16622 317483
rect 16632 317473 16690 317483
rect 17290 317473 17348 317483
rect 17358 317473 17416 317483
rect 17426 317473 17484 317483
rect 17494 317473 17552 317483
rect 17562 317473 17620 317483
rect 17630 317473 17688 317483
rect 17698 317473 17756 317483
rect 17766 317473 17824 317483
rect 17834 317473 17892 317483
rect 17902 317473 17960 317483
rect 17970 317473 18028 317483
rect 18038 317473 18096 317483
rect 18106 317473 18164 317483
rect 18174 317473 18232 317483
rect 15724 317449 16690 317473
rect 17266 317449 18232 317473
rect 12427 317424 12493 317440
rect 15748 317434 15772 317449
rect 15816 317434 15840 317449
rect 15884 317434 15908 317449
rect 15952 317434 15976 317449
rect 16020 317434 16044 317449
rect 16088 317434 16112 317449
rect 16156 317434 16180 317449
rect 16224 317434 16248 317449
rect 16292 317434 16316 317449
rect 16360 317434 16384 317449
rect 16428 317434 16452 317449
rect 16496 317434 16520 317449
rect 16564 317434 16588 317449
rect 16632 317434 16656 317449
rect 17290 317434 17314 317449
rect 17358 317434 17382 317449
rect 17426 317434 17450 317449
rect 17494 317434 17518 317449
rect 17562 317434 17586 317449
rect 17630 317434 17654 317449
rect 17698 317434 17722 317449
rect 17766 317434 17790 317449
rect 17834 317434 17858 317449
rect 17902 317434 17926 317449
rect 17970 317434 17994 317449
rect 18038 317434 18062 317449
rect 18106 317434 18130 317449
rect 18174 317434 18198 317449
rect 15678 317279 16678 317434
rect 7389 317189 8389 317249
rect 8990 317189 9990 317249
rect 15678 317245 16690 317279
rect 17278 317269 18278 317434
rect 17266 317245 18278 317269
rect 15678 317234 16678 317245
rect 17278 317234 18278 317245
rect 15748 317221 15772 317234
rect 15816 317221 15840 317234
rect 15884 317221 15908 317234
rect 15952 317221 15976 317234
rect 16020 317221 16044 317234
rect 16088 317221 16112 317234
rect 16156 317221 16180 317234
rect 16224 317221 16248 317234
rect 16292 317221 16316 317234
rect 16360 317221 16384 317234
rect 16428 317221 16452 317234
rect 16496 317221 16520 317234
rect 16564 317221 16588 317234
rect 16632 317221 16656 317234
rect 17290 317221 17314 317234
rect 17358 317221 17382 317234
rect 17426 317221 17450 317234
rect 17494 317221 17518 317234
rect 17562 317221 17586 317234
rect 17630 317221 17654 317234
rect 17698 317221 17722 317234
rect 17766 317221 17790 317234
rect 17834 317221 17858 317234
rect 17902 317221 17926 317234
rect 17970 317221 17994 317234
rect 18038 317221 18062 317234
rect 18106 317221 18130 317234
rect 18174 317221 18198 317234
rect 7389 316831 8389 316887
rect 8990 316831 9990 316887
rect 15678 316876 16678 316932
rect 17278 316876 18278 316932
rect 7389 316759 8389 316815
rect 8990 316759 9990 316815
rect 15678 316804 16678 316860
rect 17278 316804 18278 316860
rect 7389 316457 8389 316529
rect 8990 316457 9990 316529
rect 15678 316502 16678 316574
rect 17278 316502 18278 316574
rect 15748 316491 15782 316502
rect 15816 316491 15850 316502
rect 15884 316491 15918 316502
rect 15952 316491 15986 316502
rect 16020 316491 16054 316502
rect 16088 316491 16122 316502
rect 16156 316491 16190 316502
rect 16224 316491 16258 316502
rect 16292 316491 16326 316502
rect 16360 316491 16394 316502
rect 16428 316491 16462 316502
rect 16496 316491 16530 316502
rect 16564 316491 16598 316502
rect 16632 316491 16666 316502
rect 17290 316491 17324 316502
rect 17358 316491 17392 316502
rect 17426 316491 17460 316502
rect 17494 316491 17528 316502
rect 17562 316491 17596 316502
rect 17630 316491 17664 316502
rect 17698 316491 17732 316502
rect 17766 316491 17800 316502
rect 17834 316491 17868 316502
rect 17902 316491 17936 316502
rect 17970 316491 18004 316502
rect 18038 316491 18072 316502
rect 18106 316491 18140 316502
rect 18174 316491 18208 316502
rect 15748 316481 15806 316491
rect 15816 316481 15874 316491
rect 15884 316481 15942 316491
rect 15952 316481 16010 316491
rect 16020 316481 16078 316491
rect 16088 316481 16146 316491
rect 16156 316481 16214 316491
rect 16224 316481 16282 316491
rect 16292 316481 16350 316491
rect 16360 316481 16418 316491
rect 16428 316481 16486 316491
rect 16496 316481 16554 316491
rect 16564 316481 16622 316491
rect 16632 316481 16690 316491
rect 17290 316481 17348 316491
rect 17358 316481 17416 316491
rect 17426 316481 17484 316491
rect 17494 316481 17552 316491
rect 17562 316481 17620 316491
rect 17630 316481 17688 316491
rect 17698 316481 17756 316491
rect 17766 316481 17824 316491
rect 17834 316481 17892 316491
rect 17902 316481 17960 316491
rect 17970 316481 18028 316491
rect 18038 316481 18096 316491
rect 18106 316481 18164 316491
rect 18174 316481 18232 316491
rect 15724 316457 16690 316481
rect 17266 316457 18232 316481
rect 15748 316442 15772 316457
rect 15816 316442 15840 316457
rect 15884 316442 15908 316457
rect 15952 316442 15976 316457
rect 16020 316442 16044 316457
rect 16088 316442 16112 316457
rect 16156 316442 16180 316457
rect 16224 316442 16248 316457
rect 16292 316442 16316 316457
rect 16360 316442 16384 316457
rect 16428 316442 16452 316457
rect 16496 316442 16520 316457
rect 16564 316442 16588 316457
rect 16632 316442 16656 316457
rect 17290 316442 17314 316457
rect 17358 316442 17382 316457
rect 17426 316442 17450 316457
rect 17494 316442 17518 316457
rect 17562 316442 17586 316457
rect 17630 316442 17654 316457
rect 17698 316442 17722 316457
rect 17766 316442 17790 316457
rect 17834 316442 17858 316457
rect 17902 316442 17926 316457
rect 17970 316442 17994 316457
rect 18038 316442 18062 316457
rect 18106 316442 18130 316457
rect 18174 316442 18198 316457
rect 15678 316287 16678 316442
rect 7389 316197 8389 316257
rect 8990 316197 9990 316257
rect 15678 316253 16690 316287
rect 17278 316277 18278 316442
rect 17266 316253 18278 316277
rect 15678 316242 16678 316253
rect 17278 316242 18278 316253
rect 15748 316229 15772 316242
rect 15816 316229 15840 316242
rect 15884 316229 15908 316242
rect 15952 316229 15976 316242
rect 16020 316229 16044 316242
rect 16088 316229 16112 316242
rect 16156 316229 16180 316242
rect 16224 316229 16248 316242
rect 16292 316229 16316 316242
rect 16360 316229 16384 316242
rect 16428 316229 16452 316242
rect 16496 316229 16520 316242
rect 16564 316229 16588 316242
rect 16632 316229 16656 316242
rect 17290 316229 17314 316242
rect 17358 316229 17382 316242
rect 17426 316229 17450 316242
rect 17494 316229 17518 316242
rect 17562 316229 17586 316242
rect 17630 316229 17654 316242
rect 17698 316229 17722 316242
rect 17766 316229 17790 316242
rect 17834 316229 17858 316242
rect 17902 316229 17926 316242
rect 17970 316229 17994 316242
rect 18038 316229 18062 316242
rect 18106 316229 18130 316242
rect 18174 316229 18198 316242
rect 7389 315839 8389 315895
rect 8990 315839 9990 315895
rect 15678 315884 16678 315940
rect 17278 315884 18278 315940
rect 7389 315767 8389 315823
rect 8990 315767 9990 315823
rect 15678 315812 16678 315868
rect 17278 315812 18278 315868
rect 7389 315465 8389 315537
rect 8990 315465 9990 315537
rect 15678 315510 16678 315582
rect 17278 315510 18278 315582
rect 15748 315499 15782 315510
rect 15816 315499 15850 315510
rect 15884 315499 15918 315510
rect 15952 315499 15986 315510
rect 16020 315499 16054 315510
rect 16088 315499 16122 315510
rect 16156 315499 16190 315510
rect 16224 315499 16258 315510
rect 16292 315499 16326 315510
rect 16360 315499 16394 315510
rect 16428 315499 16462 315510
rect 16496 315499 16530 315510
rect 16564 315499 16598 315510
rect 16632 315499 16666 315510
rect 17290 315499 17324 315510
rect 17358 315499 17392 315510
rect 17426 315499 17460 315510
rect 17494 315499 17528 315510
rect 17562 315499 17596 315510
rect 17630 315499 17664 315510
rect 17698 315499 17732 315510
rect 17766 315499 17800 315510
rect 17834 315499 17868 315510
rect 17902 315499 17936 315510
rect 17970 315499 18004 315510
rect 18038 315499 18072 315510
rect 18106 315499 18140 315510
rect 18174 315499 18208 315510
rect 15748 315489 15806 315499
rect 15816 315489 15874 315499
rect 15884 315489 15942 315499
rect 15952 315489 16010 315499
rect 16020 315489 16078 315499
rect 16088 315489 16146 315499
rect 16156 315489 16214 315499
rect 16224 315489 16282 315499
rect 16292 315489 16350 315499
rect 16360 315489 16418 315499
rect 16428 315489 16486 315499
rect 16496 315489 16554 315499
rect 16564 315489 16622 315499
rect 16632 315489 16690 315499
rect 17290 315489 17348 315499
rect 17358 315489 17416 315499
rect 17426 315489 17484 315499
rect 17494 315489 17552 315499
rect 17562 315489 17620 315499
rect 17630 315489 17688 315499
rect 17698 315489 17756 315499
rect 17766 315489 17824 315499
rect 17834 315489 17892 315499
rect 17902 315489 17960 315499
rect 17970 315489 18028 315499
rect 18038 315489 18096 315499
rect 18106 315489 18164 315499
rect 18174 315489 18232 315499
rect 15724 315465 16690 315489
rect 17266 315465 18232 315489
rect 15748 315450 15772 315465
rect 15816 315450 15840 315465
rect 15884 315450 15908 315465
rect 15952 315450 15976 315465
rect 16020 315450 16044 315465
rect 16088 315450 16112 315465
rect 16156 315450 16180 315465
rect 16224 315450 16248 315465
rect 16292 315450 16316 315465
rect 16360 315450 16384 315465
rect 16428 315450 16452 315465
rect 16496 315450 16520 315465
rect 16564 315450 16588 315465
rect 16632 315450 16656 315465
rect 17290 315450 17314 315465
rect 17358 315450 17382 315465
rect 17426 315450 17450 315465
rect 17494 315450 17518 315465
rect 17562 315450 17586 315465
rect 17630 315450 17654 315465
rect 17698 315450 17722 315465
rect 17766 315450 17790 315465
rect 17834 315450 17858 315465
rect 17902 315450 17926 315465
rect 17970 315450 17994 315465
rect 18038 315450 18062 315465
rect 18106 315450 18130 315465
rect 18174 315450 18198 315465
rect 15678 315295 16678 315450
rect 7389 315205 8389 315265
rect 8990 315205 9990 315265
rect 15678 315261 16690 315295
rect 17278 315285 18278 315450
rect 17266 315261 18278 315285
rect 15678 315250 16678 315261
rect 17278 315250 18278 315261
rect 15748 315237 15772 315250
rect 15816 315237 15840 315250
rect 15884 315237 15908 315250
rect 15952 315237 15976 315250
rect 16020 315237 16044 315250
rect 16088 315237 16112 315250
rect 16156 315237 16180 315250
rect 16224 315237 16248 315250
rect 16292 315237 16316 315250
rect 16360 315237 16384 315250
rect 16428 315237 16452 315250
rect 16496 315237 16520 315250
rect 16564 315237 16588 315250
rect 16632 315237 16656 315250
rect 17290 315237 17314 315250
rect 17358 315237 17382 315250
rect 17426 315237 17450 315250
rect 17494 315237 17518 315250
rect 17562 315237 17586 315250
rect 17630 315237 17654 315250
rect 17698 315237 17722 315250
rect 17766 315237 17790 315250
rect 17834 315237 17858 315250
rect 17902 315237 17926 315250
rect 17970 315237 17994 315250
rect 18038 315237 18062 315250
rect 18106 315237 18130 315250
rect 18174 315237 18198 315250
rect 7389 314847 8389 314903
rect 8990 314847 9990 314903
rect 15678 314892 16678 314948
rect 17278 314892 18278 314948
rect 7389 314775 8389 314831
rect 8990 314775 9990 314831
rect 15678 314820 16678 314876
rect 17278 314820 18278 314876
rect 5967 314455 6059 314489
rect 7389 314473 8389 314545
rect 8990 314473 9990 314545
rect 15678 314518 16678 314590
rect 17278 314518 18278 314590
rect 15748 314507 15782 314518
rect 15816 314507 15850 314518
rect 15884 314507 15918 314518
rect 15952 314507 15986 314518
rect 16020 314507 16054 314518
rect 16088 314507 16122 314518
rect 16156 314507 16190 314518
rect 16224 314507 16258 314518
rect 16292 314507 16326 314518
rect 16360 314507 16394 314518
rect 16428 314507 16462 314518
rect 16496 314507 16530 314518
rect 16564 314507 16598 314518
rect 16632 314507 16666 314518
rect 17290 314507 17324 314518
rect 17358 314507 17392 314518
rect 17426 314507 17460 314518
rect 17494 314507 17528 314518
rect 17562 314507 17596 314518
rect 17630 314507 17664 314518
rect 17698 314507 17732 314518
rect 17766 314507 17800 314518
rect 17834 314507 17868 314518
rect 17902 314507 17936 314518
rect 17970 314507 18004 314518
rect 18038 314507 18072 314518
rect 18106 314507 18140 314518
rect 18174 314507 18208 314518
rect 15748 314497 15806 314507
rect 15816 314497 15874 314507
rect 15884 314497 15942 314507
rect 15952 314497 16010 314507
rect 16020 314497 16078 314507
rect 16088 314497 16146 314507
rect 16156 314497 16214 314507
rect 16224 314497 16282 314507
rect 16292 314497 16350 314507
rect 16360 314497 16418 314507
rect 16428 314497 16486 314507
rect 16496 314497 16554 314507
rect 16564 314497 16622 314507
rect 16632 314497 16690 314507
rect 17290 314497 17348 314507
rect 17358 314497 17416 314507
rect 17426 314497 17484 314507
rect 17494 314497 17552 314507
rect 17562 314497 17620 314507
rect 17630 314497 17688 314507
rect 17698 314497 17756 314507
rect 17766 314497 17824 314507
rect 17834 314497 17892 314507
rect 17902 314497 17960 314507
rect 17970 314497 18028 314507
rect 18038 314497 18096 314507
rect 18106 314497 18164 314507
rect 18174 314497 18232 314507
rect 15724 314473 16690 314497
rect 17266 314473 18232 314497
rect 15748 314458 15772 314473
rect 15816 314458 15840 314473
rect 15884 314458 15908 314473
rect 15952 314458 15976 314473
rect 16020 314458 16044 314473
rect 16088 314458 16112 314473
rect 16156 314458 16180 314473
rect 16224 314458 16248 314473
rect 16292 314458 16316 314473
rect 16360 314458 16384 314473
rect 16428 314458 16452 314473
rect 16496 314458 16520 314473
rect 16564 314458 16588 314473
rect 16632 314458 16656 314473
rect 17290 314458 17314 314473
rect 17358 314458 17382 314473
rect 17426 314458 17450 314473
rect 17494 314458 17518 314473
rect 17562 314458 17586 314473
rect 17630 314458 17654 314473
rect 17698 314458 17722 314473
rect 17766 314458 17790 314473
rect 17834 314458 17858 314473
rect 17902 314458 17926 314473
rect 17970 314458 17994 314473
rect 18038 314458 18062 314473
rect 18106 314458 18130 314473
rect 18174 314458 18198 314473
rect 2850 314398 3850 314448
rect 2850 314282 3850 314332
rect 2850 314072 3850 314122
rect 2850 313956 3850 314006
rect 2850 313746 3850 313796
rect 1153 313660 1187 313718
rect 2850 313630 3850 313680
rect 2850 313420 3850 313470
rect 2850 313417 3107 313420
rect 3250 313304 3850 313354
rect 3250 313048 3850 313104
rect 3250 312892 3850 313020
rect 175 312818 1175 312868
rect 175 312662 1175 312790
rect 3250 312736 3850 312792
rect 175 312506 1175 312634
rect 175 312350 1175 312478
rect 175 312194 1175 312322
rect 175 312044 1175 312094
rect 175 311928 1175 311978
rect 175 311772 1175 311828
rect 175 311622 1175 311672
rect 1578 311609 1628 312609
rect 1728 311609 1856 312609
rect 1884 311609 2012 312609
rect 2040 311609 2090 312609
rect 3250 312580 3850 312708
rect 3250 312430 3850 312480
rect 2850 312314 3850 312364
rect 2850 312158 3850 312214
rect 2850 312008 3850 312058
rect 2850 311880 3850 311930
rect 2850 311724 3850 311852
rect 2850 311568 3850 311696
rect 175 311506 1175 311556
rect 175 311350 1175 311478
rect 2850 311412 3850 311468
rect 2850 311256 3850 311384
rect 175 311194 1175 311250
rect 175 311038 1175 311166
rect 175 310888 1175 310938
rect 175 310772 1175 310822
rect 175 310616 1175 310744
rect 1578 310613 1628 311213
rect 1728 310613 1784 311213
rect 1884 310613 1940 311213
rect 2040 310613 2096 311213
rect 2196 310613 2246 311213
rect 2850 311100 3850 311228
rect 2850 310944 3850 311072
rect 2850 310794 3850 310844
rect 2850 310678 3850 310728
rect 2850 310522 3850 310650
rect 175 310460 1175 310516
rect 175 310304 1175 310432
rect 2850 310366 3850 310494
rect 2850 310210 3850 310338
rect 175 310154 1175 310204
rect 803 310151 1175 310154
rect 2850 310054 3850 310110
rect 2850 309898 3850 310026
rect 2850 309742 3850 309870
rect 2850 309586 3850 309642
rect 2850 309436 3850 309486
rect 3926 309455 3960 309491
rect 3967 309339 3989 309455
rect 1638 307869 1688 308869
rect 1848 307869 1976 308869
rect 2064 307869 2114 308869
rect 2850 308275 3050 308287
rect 2850 308162 3850 308212
rect 2850 307946 3850 308074
rect 2850 307730 3850 307786
rect 2850 307514 3850 307642
rect 2850 307304 3850 307354
rect 2850 307188 3850 307238
rect 2850 306978 3850 307028
rect 3926 307015 3960 309339
rect 5169 307315 5191 314429
rect 5488 313194 5538 314194
rect 5658 313194 5708 314194
rect 5488 312073 5538 313073
rect 5658 312073 5708 313073
rect 5488 310952 5538 311952
rect 5658 310952 5708 311952
rect 5488 309842 5538 310842
rect 5658 309842 5708 310842
rect 5488 308721 5538 309721
rect 5658 308721 5708 309721
rect 5488 307600 5538 308600
rect 5658 307600 5708 308600
rect 5971 307386 6059 314455
rect 15678 314303 16678 314458
rect 7389 314213 8389 314273
rect 8990 314213 9990 314273
rect 15678 314269 16690 314303
rect 17278 314293 18278 314458
rect 17266 314269 18278 314293
rect 15678 314258 16678 314269
rect 17278 314258 18278 314269
rect 15748 314245 15772 314258
rect 15816 314245 15840 314258
rect 15884 314245 15908 314258
rect 15952 314245 15976 314258
rect 16020 314245 16044 314258
rect 16088 314245 16112 314258
rect 16156 314245 16180 314258
rect 16224 314245 16248 314258
rect 16292 314245 16316 314258
rect 16360 314245 16384 314258
rect 16428 314245 16452 314258
rect 16496 314245 16520 314258
rect 16564 314245 16588 314258
rect 16632 314245 16656 314258
rect 17290 314245 17314 314258
rect 17358 314245 17382 314258
rect 17426 314245 17450 314258
rect 17494 314245 17518 314258
rect 17562 314245 17586 314258
rect 17630 314245 17654 314258
rect 17698 314245 17722 314258
rect 17766 314245 17790 314258
rect 17834 314245 17858 314258
rect 17902 314245 17926 314258
rect 17970 314245 17994 314258
rect 18038 314245 18062 314258
rect 18106 314245 18130 314258
rect 18174 314245 18198 314258
rect 7389 313855 8389 313911
rect 8990 313855 9990 313911
rect 15678 313900 16678 313956
rect 17278 313900 18278 313956
rect 7389 313783 8389 313839
rect 8990 313783 9990 313839
rect 15678 313828 16678 313884
rect 17278 313828 18278 313884
rect 7389 313481 8389 313553
rect 8990 313481 9990 313553
rect 15678 313526 16678 313598
rect 17278 313526 18278 313598
rect 15748 313515 15782 313526
rect 15816 313515 15850 313526
rect 15884 313515 15918 313526
rect 15952 313515 15986 313526
rect 16020 313515 16054 313526
rect 16088 313515 16122 313526
rect 16156 313515 16190 313526
rect 16224 313515 16258 313526
rect 16292 313515 16326 313526
rect 16360 313515 16394 313526
rect 16428 313515 16462 313526
rect 16496 313515 16530 313526
rect 16564 313515 16598 313526
rect 16632 313515 16666 313526
rect 17290 313515 17324 313526
rect 17358 313515 17392 313526
rect 17426 313515 17460 313526
rect 17494 313515 17528 313526
rect 17562 313515 17596 313526
rect 17630 313515 17664 313526
rect 17698 313515 17732 313526
rect 17766 313515 17800 313526
rect 17834 313515 17868 313526
rect 17902 313515 17936 313526
rect 17970 313515 18004 313526
rect 18038 313515 18072 313526
rect 18106 313515 18140 313526
rect 18174 313515 18208 313526
rect 15748 313505 15806 313515
rect 15816 313505 15874 313515
rect 15884 313505 15942 313515
rect 15952 313505 16010 313515
rect 16020 313505 16078 313515
rect 16088 313505 16146 313515
rect 16156 313505 16214 313515
rect 16224 313505 16282 313515
rect 16292 313505 16350 313515
rect 16360 313505 16418 313515
rect 16428 313505 16486 313515
rect 16496 313505 16554 313515
rect 16564 313505 16622 313515
rect 16632 313505 16690 313515
rect 17290 313505 17348 313515
rect 17358 313505 17416 313515
rect 17426 313505 17484 313515
rect 17494 313505 17552 313515
rect 17562 313505 17620 313515
rect 17630 313505 17688 313515
rect 17698 313505 17756 313515
rect 17766 313505 17824 313515
rect 17834 313505 17892 313515
rect 17902 313505 17960 313515
rect 17970 313505 18028 313515
rect 18038 313505 18096 313515
rect 18106 313505 18164 313515
rect 18174 313505 18232 313515
rect 15724 313481 16690 313505
rect 17266 313481 18232 313505
rect 15748 313466 15772 313481
rect 15816 313466 15840 313481
rect 15884 313466 15908 313481
rect 15952 313466 15976 313481
rect 16020 313466 16044 313481
rect 16088 313466 16112 313481
rect 16156 313466 16180 313481
rect 16224 313466 16248 313481
rect 16292 313466 16316 313481
rect 16360 313466 16384 313481
rect 16428 313466 16452 313481
rect 16496 313466 16520 313481
rect 16564 313466 16588 313481
rect 16632 313466 16656 313481
rect 17290 313466 17314 313481
rect 17358 313466 17382 313481
rect 17426 313466 17450 313481
rect 17494 313466 17518 313481
rect 17562 313466 17586 313481
rect 17630 313466 17654 313481
rect 17698 313466 17722 313481
rect 17766 313466 17790 313481
rect 17834 313466 17858 313481
rect 17902 313466 17926 313481
rect 17970 313466 17994 313481
rect 18038 313466 18062 313481
rect 18106 313466 18130 313481
rect 18174 313466 18198 313481
rect 15678 313311 16678 313466
rect 7389 313221 8389 313281
rect 8990 313221 9990 313281
rect 15678 313277 16690 313311
rect 17278 313301 18278 313466
rect 17266 313277 18278 313301
rect 15678 313266 16678 313277
rect 17278 313266 18278 313277
rect 15748 313253 15772 313266
rect 15816 313253 15840 313266
rect 15884 313253 15908 313266
rect 15952 313253 15976 313266
rect 16020 313253 16044 313266
rect 16088 313253 16112 313266
rect 16156 313253 16180 313266
rect 16224 313253 16248 313266
rect 16292 313253 16316 313266
rect 16360 313253 16384 313266
rect 16428 313253 16452 313266
rect 16496 313253 16520 313266
rect 16564 313253 16588 313266
rect 16632 313253 16656 313266
rect 17290 313253 17314 313266
rect 17358 313253 17382 313266
rect 17426 313253 17450 313266
rect 17494 313253 17518 313266
rect 17562 313253 17586 313266
rect 17630 313253 17654 313266
rect 17698 313253 17722 313266
rect 17766 313253 17790 313266
rect 17834 313253 17858 313266
rect 17902 313253 17926 313266
rect 17970 313253 17994 313266
rect 18038 313253 18062 313266
rect 18106 313253 18130 313266
rect 18174 313253 18198 313266
rect 7389 312863 8389 312919
rect 8990 312863 9990 312919
rect 15678 312908 16678 312964
rect 17278 312908 18278 312964
rect 7389 312791 8389 312847
rect 8990 312791 9990 312847
rect 15678 312836 16678 312892
rect 17278 312836 18278 312892
rect 19480 312867 19516 319817
rect 19547 312867 19583 319817
rect 24572 319738 25172 319866
rect 36785 319864 37385 319920
rect 36785 319688 37385 319744
rect 20809 319650 20833 319684
rect 20809 319582 20833 319616
rect 24572 319588 25172 319638
rect 20809 319514 20833 319548
rect 36785 319518 37385 319568
rect 20809 319446 20833 319480
rect 24572 319458 25172 319508
rect 32930 319457 33530 319507
rect 20809 319378 20833 319412
rect 35287 319391 35887 319441
rect 36785 319402 37385 319452
rect 20809 319310 20833 319344
rect 24572 319308 25172 319358
rect 31463 319307 32063 319357
rect 32930 319301 33530 319357
rect 20809 319242 20833 319276
rect 35287 319215 35887 319343
rect 36785 319226 37385 319282
rect 20809 319174 20833 319208
rect 31463 319151 32063 319207
rect 32930 319151 33530 319201
rect 34079 319157 34679 319207
rect 20809 319106 20833 319140
rect 19844 318051 19894 319051
rect 19994 318051 20122 319051
rect 20150 318051 20278 319051
rect 20306 318051 20434 319051
rect 20462 318051 20512 319051
rect 20809 319038 20833 319072
rect 20809 318970 20833 319004
rect 20973 319000 21007 319024
rect 21041 319000 21075 319024
rect 21109 319000 21143 319024
rect 21177 319000 21211 319024
rect 21245 319000 21279 319024
rect 21313 319000 21347 319024
rect 21381 319000 21415 319024
rect 21449 319000 21483 319024
rect 21517 319000 21551 319024
rect 21585 319000 21619 319024
rect 21653 319000 21687 319024
rect 21721 319000 21755 319024
rect 21789 319000 21823 319024
rect 21857 319000 21891 319024
rect 21925 319000 21959 319024
rect 21993 319000 22027 319024
rect 22061 319000 22095 319024
rect 22129 319000 22163 319024
rect 22197 319000 22210 319024
rect 31463 319001 32063 319051
rect 34079 319001 34679 319057
rect 35287 319039 35887 319095
rect 36785 319050 37385 319106
rect 20809 318902 20833 318936
rect 32596 318929 33596 318979
rect 20809 318834 20833 318868
rect 24573 318820 25173 318870
rect 34079 318851 34679 318901
rect 35287 318869 35887 318919
rect 36785 318880 37385 318930
rect 35287 318866 35559 318869
rect 35716 318866 35887 318869
rect 20809 318766 20833 318800
rect 30171 318795 30771 318845
rect 20809 318698 20833 318732
rect 24573 318664 25173 318792
rect 32596 318773 33596 318829
rect 37993 318704 38593 318754
rect 19844 316521 19894 317921
rect 19994 316521 20122 317921
rect 20150 316521 20278 317921
rect 20306 316521 20434 317921
rect 20462 316521 20512 317921
rect 20809 316219 20833 316253
rect 19844 314759 19894 316159
rect 19994 314759 20122 316159
rect 20150 314759 20278 316159
rect 20306 314759 20434 316159
rect 20462 314759 20512 316159
rect 20809 316151 20833 316185
rect 20809 316083 20833 316117
rect 20809 316015 20833 316049
rect 20809 315947 20833 315981
rect 20809 315879 20833 315913
rect 20809 315811 20833 315845
rect 20809 315743 20833 315777
rect 20809 315675 20833 315709
rect 20809 315607 20833 315641
rect 20809 315539 20833 315573
rect 21263 315518 21313 318518
rect 21413 315518 21541 318518
rect 21569 315518 21697 318518
rect 21725 315518 21853 318518
rect 21881 315518 22009 318518
rect 22037 315518 22165 318518
rect 22193 315518 22321 318518
rect 22349 315518 22399 318518
rect 24573 318508 25173 318636
rect 30171 318619 30771 318675
rect 32596 318623 33596 318673
rect 34110 318589 34710 318639
rect 36785 318620 36797 318624
rect 36785 318609 36800 318620
rect 36970 318609 36985 318624
rect 26348 318530 26372 318564
rect 32596 318507 33596 318557
rect 26348 318461 26372 318495
rect 30171 318449 30771 318499
rect 24573 318352 25173 318408
rect 24573 318196 25173 318324
rect 29993 318310 30993 318360
rect 32596 318351 33596 318479
rect 34110 318433 34710 318561
rect 36785 318429 36985 318609
rect 37993 318534 38593 318584
rect 36785 318418 36800 318429
rect 36785 318414 36797 318418
rect 36970 318414 36985 318429
rect 31347 318317 31362 318332
rect 31535 318328 31547 318332
rect 31532 318317 31547 318328
rect 24573 318040 25173 318168
rect 26490 318122 26690 318172
rect 29993 318160 30993 318210
rect 31347 318137 31547 318317
rect 31347 318122 31362 318137
rect 31532 318126 31547 318137
rect 31535 318122 31547 318126
rect 31607 318317 31622 318332
rect 31795 318328 31807 318332
rect 31792 318317 31807 318328
rect 31607 318137 31807 318317
rect 32596 318195 33596 318323
rect 34110 318277 34710 318405
rect 36785 318384 36797 318388
rect 36785 318373 36800 318384
rect 36970 318373 36985 318388
rect 31607 318122 31622 318137
rect 31792 318126 31807 318137
rect 31795 318122 31807 318126
rect 31347 318081 31362 318096
rect 31535 318092 31547 318096
rect 31532 318081 31547 318092
rect 22906 317855 23212 318025
rect 23406 317855 23712 318025
rect 26490 317966 26690 318022
rect 29993 318001 30993 318051
rect 24573 317890 25173 317940
rect 31347 317901 31547 318081
rect 26490 317816 26690 317866
rect 29993 317851 30993 317901
rect 31347 317886 31362 317901
rect 31532 317890 31547 317901
rect 31535 317886 31547 317890
rect 31607 318081 31622 318096
rect 31795 318092 31807 318096
rect 31792 318081 31807 318092
rect 31607 317901 31807 318081
rect 32596 318039 33596 318167
rect 34110 318121 34710 318249
rect 36785 318193 36985 318373
rect 36785 318182 36800 318193
rect 36785 318178 36797 318182
rect 36970 318178 36985 318193
rect 37083 318373 37098 318388
rect 37083 318193 37120 318373
rect 37083 318178 37098 318193
rect 37998 318108 38598 318158
rect 34110 317971 34710 318021
rect 31607 317886 31622 317901
rect 31792 317890 31807 317901
rect 31795 317886 31807 317890
rect 32596 317883 33596 317939
rect 37998 317932 38598 317988
rect 34110 317855 34710 317905
rect 24573 317760 25173 317810
rect 27691 317682 28291 317732
rect 30253 317721 30268 317736
rect 30441 317732 30453 317736
rect 30438 317721 30453 317732
rect 24573 317610 25173 317660
rect 27691 317532 28291 317582
rect 30253 317541 30453 317721
rect 30253 317526 30268 317541
rect 30438 317530 30453 317541
rect 30441 317526 30453 317530
rect 30513 317721 30528 317736
rect 30701 317732 30713 317736
rect 30698 317721 30713 317732
rect 30513 317541 30713 317721
rect 30513 317526 30528 317541
rect 30698 317530 30713 317541
rect 30701 317526 30713 317530
rect 30773 317721 30788 317736
rect 30961 317732 30973 317736
rect 30958 317721 30973 317732
rect 30773 317541 30973 317721
rect 30773 317526 30788 317541
rect 30958 317530 30973 317541
rect 30961 317526 30973 317530
rect 31087 317721 31102 317736
rect 31275 317732 31287 317736
rect 31272 317721 31287 317732
rect 31087 317541 31287 317721
rect 31087 317526 31102 317541
rect 31272 317530 31287 317541
rect 31275 317526 31287 317530
rect 31347 317721 31362 317736
rect 31535 317732 31547 317736
rect 31532 317721 31547 317732
rect 31347 317541 31547 317721
rect 31347 317526 31362 317541
rect 31532 317530 31547 317541
rect 31535 317526 31547 317530
rect 31607 317721 31622 317736
rect 31795 317732 31807 317736
rect 31792 317721 31807 317732
rect 31607 317541 31807 317721
rect 31607 317526 31622 317541
rect 31792 317530 31807 317541
rect 31795 317526 31807 317530
rect 31867 317721 31882 317736
rect 32055 317732 32067 317736
rect 32052 317721 32067 317732
rect 32596 317727 33596 317855
rect 31867 317541 32067 317721
rect 34110 317699 34710 317827
rect 37998 317762 38598 317812
rect 37998 317759 38220 317762
rect 38245 317759 38539 317762
rect 32596 317571 33596 317699
rect 34110 317543 34710 317671
rect 31867 317526 31882 317541
rect 32052 317530 32067 317541
rect 32055 317526 32067 317530
rect 22619 317446 22647 317474
rect 24573 317438 25173 317488
rect 26490 317416 26690 317466
rect 27691 317402 28291 317452
rect 32596 317415 33596 317543
rect 34110 317387 34710 317515
rect 24573 317288 25173 317338
rect 26490 317260 26690 317316
rect 27691 317246 28291 317374
rect 30253 317361 30268 317376
rect 30441 317372 30453 317376
rect 30438 317361 30453 317372
rect 30253 317331 30453 317361
rect 30253 317316 30268 317331
rect 30438 317320 30453 317331
rect 30441 317316 30453 317320
rect 30513 317361 30528 317376
rect 30701 317372 30713 317376
rect 30698 317361 30713 317372
rect 30513 317331 30713 317361
rect 30513 317316 30528 317331
rect 30698 317320 30713 317331
rect 30701 317316 30713 317320
rect 30773 317361 30788 317376
rect 31347 317361 31362 317376
rect 31535 317372 31547 317376
rect 31532 317361 31547 317372
rect 30773 317331 30793 317361
rect 31347 317331 31547 317361
rect 30773 317316 30788 317331
rect 31347 317316 31362 317331
rect 31532 317320 31547 317331
rect 31535 317316 31547 317320
rect 31607 317361 31622 317376
rect 31795 317372 31807 317376
rect 31792 317361 31807 317372
rect 31607 317331 31807 317361
rect 31607 317316 31622 317331
rect 31792 317320 31807 317331
rect 31795 317316 31807 317320
rect 31867 317361 31882 317376
rect 31867 317331 31921 317361
rect 31867 317316 31882 317331
rect 30253 317275 30268 317290
rect 30441 317286 30453 317290
rect 30438 317275 30453 317286
rect 30253 317245 30453 317275
rect 30253 317230 30268 317245
rect 30438 317234 30453 317245
rect 30441 317230 30453 317234
rect 30513 317275 30528 317290
rect 30701 317286 30713 317290
rect 30698 317275 30713 317286
rect 30513 317245 30713 317275
rect 30513 317230 30528 317245
rect 30698 317234 30713 317245
rect 30701 317230 30713 317234
rect 30773 317275 30788 317290
rect 31347 317275 31362 317290
rect 31535 317286 31547 317290
rect 31532 317275 31547 317286
rect 30773 317245 30793 317275
rect 31347 317245 31547 317275
rect 30773 317230 30788 317245
rect 31347 317230 31362 317245
rect 31532 317234 31547 317245
rect 31535 317230 31547 317234
rect 31607 317275 31622 317290
rect 31795 317286 31807 317290
rect 31792 317275 31807 317286
rect 31607 317245 31807 317275
rect 31607 317230 31622 317245
rect 31792 317234 31807 317245
rect 31795 317230 31807 317234
rect 31867 317275 31882 317290
rect 31867 317245 31921 317275
rect 32596 317265 33596 317315
rect 31867 317230 31882 317245
rect 34110 317231 34710 317287
rect 22906 317055 23212 317225
rect 23406 317055 23712 317225
rect 24573 317158 25173 317208
rect 24573 317002 25173 317130
rect 26490 317107 26690 317160
rect 27691 317090 28291 317218
rect 31823 317084 32061 317118
rect 31481 317080 32061 317084
rect 31481 317068 31797 317080
rect 32596 317063 33596 317113
rect 34110 317075 34710 317203
rect 37998 317133 38148 317145
rect 38317 317133 38467 317145
rect 24573 316846 25173 316974
rect 27691 316934 28291 316990
rect 32596 316907 33596 317035
rect 34110 316919 34710 317047
rect 37998 317020 38598 317070
rect 27691 316778 28291 316906
rect 25286 316758 25310 316762
rect 32596 316751 33596 316879
rect 34110 316763 34710 316891
rect 37998 316844 38598 316900
rect 24573 316690 25173 316746
rect 25286 316687 25310 316721
rect 24573 316534 25173 316662
rect 25286 316615 25310 316649
rect 27691 316622 28291 316750
rect 32596 316595 33596 316723
rect 35287 316695 35487 316707
rect 37998 316674 38598 316724
rect 34110 316607 34710 316663
rect 36785 316650 36797 316654
rect 36785 316639 36800 316650
rect 36970 316639 36985 316654
rect 35134 316582 35734 316632
rect 25286 316543 25310 316577
rect 22906 316255 23212 316425
rect 23406 316255 23712 316425
rect 24573 316378 25173 316506
rect 25286 316471 25310 316505
rect 27691 316472 28291 316522
rect 32596 316439 33596 316567
rect 34110 316451 34710 316507
rect 35134 316432 35734 316482
rect 36785 316459 36985 316639
rect 36785 316448 36800 316459
rect 36785 316444 36797 316448
rect 36970 316444 36985 316459
rect 37083 316639 37098 316654
rect 37083 316459 37120 316639
rect 37083 316444 37098 316459
rect 36785 316414 36797 316418
rect 32596 316283 33596 316411
rect 36785 316403 36800 316414
rect 36970 316403 36985 316418
rect 34110 316295 34710 316351
rect 35134 316316 35734 316366
rect 24573 316228 25173 316278
rect 32596 316127 33596 316255
rect 34110 316145 34710 316195
rect 35134 316160 35734 316288
rect 32596 315971 33596 316099
rect 34110 316029 34710 316079
rect 35134 316004 35734 316132
rect 31481 315862 31797 315880
rect 34110 315873 34710 316001
rect 31823 315828 32061 315860
rect 32596 315821 33596 315871
rect 35134 315848 35734 315976
rect 36071 315805 36098 316295
rect 36785 316223 36985 316403
rect 37993 316248 38593 316298
rect 36785 316212 36800 316223
rect 36785 316208 36797 316212
rect 36970 316208 36985 316223
rect 37993 316078 38593 316128
rect 36785 315902 37385 315952
rect 34110 315717 34710 315773
rect 30253 315701 30268 315716
rect 30441 315712 30453 315716
rect 30438 315701 30453 315712
rect 30253 315671 30453 315701
rect 30253 315656 30268 315671
rect 30438 315660 30453 315671
rect 30441 315656 30453 315660
rect 30513 315701 30528 315716
rect 30701 315712 30713 315716
rect 30698 315701 30713 315712
rect 30513 315671 30713 315701
rect 30513 315656 30528 315671
rect 30698 315660 30713 315671
rect 30701 315656 30713 315660
rect 30773 315701 30788 315716
rect 31347 315701 31362 315716
rect 31535 315712 31547 315716
rect 31532 315701 31547 315712
rect 30773 315671 30793 315701
rect 31347 315671 31547 315701
rect 30773 315656 30788 315671
rect 31347 315656 31362 315671
rect 31532 315660 31547 315671
rect 31535 315656 31547 315660
rect 31607 315701 31622 315716
rect 31795 315712 31807 315716
rect 31792 315701 31807 315712
rect 31607 315671 31807 315701
rect 31607 315656 31622 315671
rect 31792 315660 31807 315671
rect 31795 315656 31807 315660
rect 31867 315701 31882 315716
rect 31867 315671 31921 315701
rect 35134 315698 35734 315770
rect 36785 315726 37385 315782
rect 31867 315656 31882 315671
rect 30253 315615 30268 315630
rect 30441 315626 30453 315630
rect 30438 315615 30453 315626
rect 30253 315585 30453 315615
rect 30253 315570 30268 315585
rect 30438 315574 30453 315585
rect 30441 315570 30453 315574
rect 30513 315615 30528 315630
rect 30701 315626 30713 315630
rect 30698 315615 30713 315626
rect 30513 315585 30713 315615
rect 30513 315570 30528 315585
rect 30698 315574 30713 315585
rect 30701 315570 30713 315574
rect 30773 315615 30788 315630
rect 31347 315615 31362 315630
rect 31535 315626 31547 315630
rect 31532 315615 31547 315626
rect 30773 315585 30793 315615
rect 31347 315585 31547 315615
rect 30773 315570 30788 315585
rect 31347 315570 31362 315585
rect 31532 315574 31547 315585
rect 31535 315570 31547 315574
rect 31607 315615 31622 315630
rect 31795 315626 31807 315630
rect 31792 315615 31807 315626
rect 31607 315585 31807 315615
rect 31607 315570 31622 315585
rect 31792 315574 31807 315585
rect 31795 315570 31807 315574
rect 31867 315615 31882 315630
rect 32546 315619 33546 315669
rect 31867 315585 31921 315615
rect 31867 315570 31882 315585
rect 20809 315471 20833 315505
rect 32546 315463 33546 315591
rect 34110 315561 34710 315689
rect 35134 315645 36134 315695
rect 35134 315489 36134 315617
rect 36785 315550 37385 315606
rect 20809 315403 20833 315437
rect 30253 315405 30268 315420
rect 30441 315416 30453 315420
rect 30438 315405 30453 315416
rect 20809 315335 20833 315369
rect 20809 315267 20833 315301
rect 20809 315199 20833 315233
rect 30253 315225 30453 315405
rect 30253 315210 30268 315225
rect 30438 315214 30453 315225
rect 30441 315210 30453 315214
rect 30513 315405 30528 315420
rect 30701 315416 30713 315420
rect 30698 315405 30713 315416
rect 30513 315225 30713 315405
rect 30513 315210 30528 315225
rect 30698 315214 30713 315225
rect 30701 315210 30713 315214
rect 30773 315405 30788 315420
rect 30961 315416 30973 315420
rect 30958 315405 30973 315416
rect 30773 315225 30973 315405
rect 30773 315210 30788 315225
rect 30958 315214 30973 315225
rect 30961 315210 30973 315214
rect 31087 315405 31102 315420
rect 31275 315416 31287 315420
rect 31272 315405 31287 315416
rect 31087 315225 31287 315405
rect 31087 315210 31102 315225
rect 31272 315214 31287 315225
rect 31275 315210 31287 315214
rect 31347 315405 31362 315420
rect 31535 315416 31547 315420
rect 31532 315405 31547 315416
rect 31347 315225 31547 315405
rect 31347 315210 31362 315225
rect 31532 315214 31547 315225
rect 31535 315210 31547 315214
rect 31607 315405 31622 315420
rect 31795 315416 31807 315420
rect 31792 315405 31807 315416
rect 31607 315225 31807 315405
rect 31607 315210 31622 315225
rect 31792 315214 31807 315225
rect 31795 315210 31807 315214
rect 31867 315405 31882 315420
rect 32055 315416 32067 315420
rect 32052 315405 32067 315416
rect 31867 315225 32067 315405
rect 32546 315307 33546 315435
rect 34110 315411 34710 315461
rect 35134 315339 36134 315389
rect 36785 315380 37385 315430
rect 31867 315210 31882 315225
rect 32052 315214 32067 315225
rect 32055 315210 32067 315214
rect 20809 315131 20833 315165
rect 32546 315151 33546 315279
rect 36785 315248 37385 315298
rect 35285 315162 35319 315172
rect 35353 315162 35387 315172
rect 35421 315162 35455 315172
rect 35489 315162 35523 315172
rect 35564 315162 35598 315172
rect 35632 315162 35666 315172
rect 35700 315162 35734 315172
rect 35768 315162 35802 315172
rect 35836 315162 35870 315172
rect 35904 315162 35938 315172
rect 35972 315162 36006 315172
rect 36040 315162 36074 315172
rect 36108 315162 36142 315172
rect 36176 315162 36210 315172
rect 35255 315126 36255 315138
rect 20809 315063 20833 315097
rect 20940 315085 20983 315103
rect 20940 315069 20949 315085
rect 20974 315069 20983 315085
rect 25113 315069 25349 315093
rect 25383 315069 25417 315093
rect 20974 315051 21008 315069
rect 20809 314995 20833 315029
rect 20974 315028 21003 315051
rect 21361 315045 21409 315069
rect 20949 315027 20983 315028
rect 21385 314991 21409 315045
rect 25113 314991 25137 315069
rect 29993 315045 30993 315095
rect 31347 315045 31362 315060
rect 31535 315056 31547 315060
rect 31532 315045 31547 315056
rect 21361 314967 21409 314991
rect 25089 314967 25137 314991
rect 20809 314927 20833 314961
rect 20809 314859 20833 314893
rect 20809 314791 20833 314825
rect 20809 314723 20833 314757
rect 20809 314655 20833 314689
rect 21413 314638 22813 314681
rect 23685 314638 25085 314681
rect 19844 313229 19894 314629
rect 19994 313229 20122 314629
rect 20150 313229 20278 314629
rect 20306 313229 20434 314629
rect 20462 313229 20512 314629
rect 20809 314587 20833 314621
rect 20809 314519 20833 314553
rect 20809 314451 20833 314485
rect 21413 314475 22813 314603
rect 23685 314475 25085 314603
rect 20809 314383 20833 314417
rect 20809 314315 20833 314349
rect 21413 314312 22813 314440
rect 23685 314312 25085 314440
rect 20809 314247 20833 314281
rect 20809 314179 20833 314213
rect 21413 314149 22813 314277
rect 23685 314149 25085 314277
rect 20809 314111 20833 314145
rect 20809 314043 20833 314077
rect 20809 313975 20833 314009
rect 21413 313986 22813 314114
rect 23685 313986 25085 314114
rect 20809 313907 20833 313941
rect 20809 313839 20833 313873
rect 21413 313823 22813 313951
rect 23685 313823 25085 313951
rect 20809 313771 20833 313805
rect 20809 313703 20833 313737
rect 21413 313673 22813 313716
rect 23685 313673 25085 313716
rect 20809 313635 20833 313669
rect 20809 313567 20833 313601
rect 21361 313552 21419 313586
rect 25089 313552 25147 313586
rect 20809 313499 20833 313533
rect 20809 313431 20833 313465
rect 20809 313363 20833 313397
rect 21361 313373 21419 313397
rect 25089 313373 25147 313397
rect 21385 313363 21419 313373
rect 25113 313363 25147 313373
rect 20809 313295 20833 313329
rect 21385 313291 21419 313325
rect 25113 313291 25147 313325
rect 20809 313227 20833 313261
rect 21385 313219 21419 313253
rect 25113 313219 25147 313253
rect 20809 313159 20833 313193
rect 21385 313171 21419 313181
rect 25113 313171 25147 313181
rect 21361 313147 21419 313171
rect 25089 313147 25147 313171
rect 20809 313091 20833 313125
rect 20809 313023 20833 313057
rect 20809 312955 20833 312989
rect 21361 312969 21409 312993
rect 25089 312969 25137 312993
rect 20809 312887 20833 312921
rect 21385 312915 21409 312969
rect 25113 312915 25137 312969
rect 21361 312891 21409 312915
rect 25089 312891 25137 312915
rect 19480 312831 19583 312867
rect 21413 312754 22813 312804
rect 23685 312754 25085 312804
rect 7389 312489 8389 312561
rect 8990 312489 9990 312561
rect 15678 312534 16678 312606
rect 17278 312534 18278 312606
rect 21413 312591 22813 312719
rect 23685 312591 25085 312719
rect 15748 312523 15782 312534
rect 15816 312523 15850 312534
rect 15884 312523 15918 312534
rect 15952 312523 15986 312534
rect 16020 312523 16054 312534
rect 16088 312523 16122 312534
rect 16156 312523 16190 312534
rect 16224 312523 16258 312534
rect 16292 312523 16326 312534
rect 16360 312523 16394 312534
rect 16428 312523 16462 312534
rect 16496 312523 16530 312534
rect 16564 312523 16598 312534
rect 16632 312523 16666 312534
rect 17290 312523 17324 312534
rect 17358 312523 17392 312534
rect 17426 312523 17460 312534
rect 17494 312523 17528 312534
rect 17562 312523 17596 312534
rect 17630 312523 17664 312534
rect 17698 312523 17732 312534
rect 17766 312523 17800 312534
rect 17834 312523 17868 312534
rect 17902 312523 17936 312534
rect 17970 312523 18004 312534
rect 18038 312523 18072 312534
rect 18106 312523 18140 312534
rect 18174 312523 18208 312534
rect 15748 312513 15806 312523
rect 15816 312513 15874 312523
rect 15884 312513 15942 312523
rect 15952 312513 16010 312523
rect 16020 312513 16078 312523
rect 16088 312513 16146 312523
rect 16156 312513 16214 312523
rect 16224 312513 16282 312523
rect 16292 312513 16350 312523
rect 16360 312513 16418 312523
rect 16428 312513 16486 312523
rect 16496 312513 16554 312523
rect 16564 312513 16622 312523
rect 16632 312513 16690 312523
rect 17290 312513 17348 312523
rect 17358 312513 17416 312523
rect 17426 312513 17484 312523
rect 17494 312513 17552 312523
rect 17562 312513 17620 312523
rect 17630 312513 17688 312523
rect 17698 312513 17756 312523
rect 17766 312513 17824 312523
rect 17834 312513 17892 312523
rect 17902 312513 17960 312523
rect 17970 312513 18028 312523
rect 18038 312513 18096 312523
rect 18106 312513 18164 312523
rect 18174 312513 18232 312523
rect 15724 312489 16690 312513
rect 17266 312489 18232 312513
rect 15748 312474 15772 312489
rect 15816 312474 15840 312489
rect 15884 312474 15908 312489
rect 15952 312474 15976 312489
rect 16020 312474 16044 312489
rect 16088 312474 16112 312489
rect 16156 312474 16180 312489
rect 16224 312474 16248 312489
rect 16292 312474 16316 312489
rect 16360 312474 16384 312489
rect 16428 312474 16452 312489
rect 16496 312474 16520 312489
rect 16564 312474 16588 312489
rect 16632 312474 16656 312489
rect 17290 312474 17314 312489
rect 17358 312474 17382 312489
rect 17426 312474 17450 312489
rect 17494 312474 17518 312489
rect 17562 312474 17586 312489
rect 17630 312474 17654 312489
rect 17698 312474 17722 312489
rect 17766 312474 17790 312489
rect 17834 312474 17858 312489
rect 17902 312474 17926 312489
rect 17970 312474 17994 312489
rect 18038 312474 18062 312489
rect 18106 312474 18130 312489
rect 18174 312474 18198 312489
rect 15678 312319 16678 312474
rect 7389 312229 8389 312289
rect 8990 312229 9990 312289
rect 15678 312285 16690 312319
rect 17278 312309 18278 312474
rect 21413 312428 22813 312556
rect 23685 312428 25085 312556
rect 17266 312285 18278 312309
rect 15678 312274 16678 312285
rect 17278 312274 18278 312285
rect 15748 312261 15772 312274
rect 15816 312261 15840 312274
rect 15884 312261 15908 312274
rect 15952 312261 15976 312274
rect 16020 312261 16044 312274
rect 16088 312261 16112 312274
rect 16156 312261 16180 312274
rect 16224 312261 16248 312274
rect 16292 312261 16316 312274
rect 16360 312261 16384 312274
rect 16428 312261 16452 312274
rect 16496 312261 16520 312274
rect 16564 312261 16588 312274
rect 16632 312261 16656 312274
rect 17290 312261 17314 312274
rect 17358 312261 17382 312274
rect 17426 312261 17450 312274
rect 17494 312261 17518 312274
rect 17562 312261 17586 312274
rect 17630 312261 17654 312274
rect 17698 312261 17722 312274
rect 17766 312261 17790 312274
rect 17834 312261 17858 312274
rect 17902 312261 17926 312274
rect 17970 312261 17994 312274
rect 18038 312261 18062 312274
rect 18106 312261 18130 312274
rect 18174 312261 18198 312274
rect 21413 312265 22813 312393
rect 23685 312265 25085 312393
rect 21413 312102 22813 312230
rect 23685 312102 25085 312230
rect 7389 311871 8389 311927
rect 8990 311871 9990 311927
rect 15678 311916 16678 311972
rect 17278 311916 18278 311972
rect 21413 311952 22813 311995
rect 23685 311952 25085 311995
rect 7389 311799 8389 311855
rect 8990 311799 9990 311855
rect 15678 311844 16678 311900
rect 17278 311844 18278 311900
rect 21406 311865 21430 311889
rect 25068 311865 25092 311889
rect 21382 311841 21385 311865
rect 25113 311841 25116 311865
rect 21382 311763 21396 311787
rect 25102 311763 25116 311787
rect 21348 311739 21372 311763
rect 21406 311739 21430 311763
rect 25068 311739 25092 311763
rect 25126 311739 25150 311763
rect 25524 311703 25548 315001
rect 29993 314895 30993 314945
rect 31347 314865 31547 315045
rect 31347 314850 31362 314865
rect 31532 314854 31547 314865
rect 31535 314850 31547 314854
rect 31607 315045 31622 315060
rect 31795 315056 31807 315060
rect 31792 315045 31807 315056
rect 31607 314865 31807 315045
rect 32546 314995 33546 315123
rect 36785 315072 37385 315128
rect 35255 315019 36255 315069
rect 31607 314850 31622 314865
rect 31792 314854 31807 314865
rect 31795 314850 31807 314854
rect 32546 314839 33546 314967
rect 35255 314843 36255 314971
rect 36785 314896 37385 314952
rect 31347 314809 31362 314824
rect 31535 314820 31547 314824
rect 31532 314809 31547 314820
rect 29993 314736 30993 314786
rect 29993 314586 30993 314636
rect 31347 314629 31547 314809
rect 31347 314614 31362 314629
rect 31532 314618 31547 314629
rect 31535 314614 31547 314618
rect 31607 314809 31622 314824
rect 31795 314820 31807 314824
rect 31792 314809 31807 314820
rect 31607 314629 31807 314809
rect 32546 314683 33546 314811
rect 35255 314667 36255 314795
rect 36785 314726 37385 314776
rect 31607 314614 31622 314629
rect 31792 314618 31807 314629
rect 31795 314614 31807 314618
rect 32546 314527 33546 314655
rect 37993 314550 38593 314600
rect 28647 314450 28671 314477
rect 30171 314447 30771 314497
rect 35255 314491 36255 314547
rect 36785 314466 36797 314470
rect 36785 314455 36800 314466
rect 36970 314455 36985 314470
rect 28683 314397 28717 314431
rect 32546 314377 33546 314427
rect 28683 314328 28717 314362
rect 28683 314259 28717 314293
rect 30171 314271 30771 314327
rect 35255 314321 36255 314371
rect 36785 314275 36985 314455
rect 37993 314380 38593 314430
rect 36785 314264 36800 314275
rect 36785 314260 36797 314264
rect 36970 314260 36985 314275
rect 36785 314230 36797 314234
rect 28683 314190 28717 314224
rect 32596 314175 33596 314225
rect 35359 314156 35375 314222
rect 36143 314156 36159 314222
rect 36785 314219 36800 314230
rect 36970 314219 36985 314234
rect 28683 314121 28717 314155
rect 30171 314101 30771 314151
rect 28683 314052 28717 314086
rect 32596 314019 33596 314147
rect 28683 313983 28717 314017
rect 33959 313994 33975 314060
rect 36143 313994 36159 314060
rect 36785 314039 36985 314219
rect 36785 314028 36800 314039
rect 36785 314024 36797 314028
rect 36970 314024 36985 314039
rect 37083 314219 37098 314234
rect 37083 314039 37120 314219
rect 37083 314024 37098 314039
rect 28683 313914 28717 313948
rect 31463 313895 32063 313945
rect 28683 313845 28717 313879
rect 32596 313863 33596 313991
rect 37998 313954 38598 314004
rect 28683 313776 28717 313810
rect 28683 313707 28717 313741
rect 31463 313739 32063 313795
rect 32596 313707 33596 313835
rect 33959 313832 33975 313898
rect 36143 313832 36159 313898
rect 37998 313778 38598 313834
rect 28683 313638 28717 313672
rect 28683 313569 28717 313603
rect 31463 313589 32063 313639
rect 32596 313551 33596 313679
rect 35359 313670 35375 313736
rect 36143 313670 36159 313736
rect 37998 313608 38598 313658
rect 37998 313605 38220 313608
rect 38245 313605 38539 313608
rect 28683 313500 28717 313534
rect 28683 313431 28717 313465
rect 28683 313362 28717 313396
rect 32596 313395 33596 313523
rect 35255 313521 36255 313571
rect 28683 313293 28717 313327
rect 28683 313224 28717 313258
rect 30015 313256 30718 313272
rect 30015 313246 30721 313256
rect 28683 313155 28717 313189
rect 28683 313086 28717 313120
rect 28683 313017 28717 313051
rect 28683 312948 28717 312982
rect 28683 312879 28717 312913
rect 28683 312810 28717 312844
rect 28683 312741 28717 312775
rect 28683 312672 28717 312706
rect 28683 312603 28717 312637
rect 28683 312534 28717 312568
rect 28683 312465 28717 312499
rect 28683 312396 28717 312430
rect 28682 312361 28683 312366
rect 28682 312332 28717 312361
rect 28647 312303 28671 312332
rect 28647 312234 28671 312268
rect 28647 312165 28671 312199
rect 28647 312096 28671 312130
rect 28647 312027 28671 312061
rect 28647 311958 28671 311992
rect 28647 311889 28671 311923
rect 28647 311820 28671 311854
rect 28647 311751 28671 311785
rect 28647 311682 28671 311716
rect 29778 311695 29802 311719
rect 29802 311671 29826 311683
rect 29880 311681 29914 311715
rect 25524 311635 25548 311669
rect 7389 311497 8389 311569
rect 8990 311497 9990 311569
rect 15678 311542 16678 311614
rect 17278 311542 18278 311614
rect 28647 311613 28671 311647
rect 29778 311635 29802 311659
rect 21361 311586 21409 311610
rect 25089 311586 25137 311610
rect 15748 311531 15782 311542
rect 15816 311531 15850 311542
rect 15884 311531 15918 311542
rect 15952 311531 15986 311542
rect 16020 311531 16054 311542
rect 16088 311531 16122 311542
rect 16156 311531 16190 311542
rect 16224 311531 16258 311542
rect 16292 311531 16326 311542
rect 16360 311531 16394 311542
rect 16428 311531 16462 311542
rect 16496 311531 16530 311542
rect 16564 311531 16598 311542
rect 16632 311531 16666 311542
rect 17290 311531 17324 311542
rect 17358 311531 17392 311542
rect 17426 311531 17460 311542
rect 17494 311531 17528 311542
rect 17562 311531 17596 311542
rect 17630 311531 17664 311542
rect 17698 311531 17732 311542
rect 17766 311531 17800 311542
rect 17834 311531 17868 311542
rect 17902 311531 17936 311542
rect 17970 311531 18004 311542
rect 18038 311531 18072 311542
rect 18106 311531 18140 311542
rect 18174 311531 18208 311542
rect 21385 311532 21409 311586
rect 25113 311532 25137 311586
rect 28647 311544 28671 311578
rect 15748 311521 15806 311531
rect 15816 311521 15874 311531
rect 15884 311521 15942 311531
rect 15952 311521 16010 311531
rect 16020 311521 16078 311531
rect 16088 311521 16146 311531
rect 16156 311521 16214 311531
rect 16224 311521 16282 311531
rect 16292 311521 16350 311531
rect 16360 311521 16418 311531
rect 16428 311521 16486 311531
rect 16496 311521 16554 311531
rect 16564 311521 16622 311531
rect 16632 311521 16690 311531
rect 17290 311521 17348 311531
rect 17358 311521 17416 311531
rect 17426 311521 17484 311531
rect 17494 311521 17552 311531
rect 17562 311521 17620 311531
rect 17630 311521 17688 311531
rect 17698 311521 17756 311531
rect 17766 311521 17824 311531
rect 17834 311521 17892 311531
rect 17902 311521 17960 311531
rect 17970 311521 18028 311531
rect 18038 311521 18096 311531
rect 18106 311521 18164 311531
rect 18174 311521 18232 311531
rect 15724 311497 16690 311521
rect 17266 311497 18232 311521
rect 21361 311508 21409 311532
rect 25089 311508 25137 311532
rect 15748 311482 15772 311497
rect 15816 311482 15840 311497
rect 15884 311482 15908 311497
rect 15952 311482 15976 311497
rect 16020 311482 16044 311497
rect 16088 311482 16112 311497
rect 16156 311482 16180 311497
rect 16224 311482 16248 311497
rect 16292 311482 16316 311497
rect 16360 311482 16384 311497
rect 16428 311482 16452 311497
rect 16496 311482 16520 311497
rect 16564 311482 16588 311497
rect 16632 311482 16656 311497
rect 17290 311482 17314 311497
rect 17358 311482 17382 311497
rect 17426 311482 17450 311497
rect 17494 311482 17518 311497
rect 17562 311482 17586 311497
rect 17630 311482 17654 311497
rect 17698 311482 17722 311497
rect 17766 311482 17790 311497
rect 17834 311482 17858 311497
rect 17902 311482 17926 311497
rect 17970 311482 17994 311497
rect 18038 311482 18062 311497
rect 18106 311482 18130 311497
rect 18174 311482 18198 311497
rect 7389 311237 8389 311297
rect 8990 311237 9990 311297
rect 12559 311273 12865 311375
rect 15678 311327 16678 311482
rect 15678 311293 16690 311327
rect 17278 311317 18278 311482
rect 28647 311475 28671 311509
rect 28647 311406 28671 311440
rect 28647 311337 28671 311371
rect 17266 311293 18278 311317
rect 15678 311282 16678 311293
rect 17278 311282 18278 311293
rect 12543 311257 12881 311273
rect 15748 311269 15772 311282
rect 15816 311269 15840 311282
rect 15884 311269 15908 311282
rect 15952 311269 15976 311282
rect 16020 311269 16044 311282
rect 16088 311269 16112 311282
rect 16156 311269 16180 311282
rect 16224 311269 16248 311282
rect 16292 311269 16316 311282
rect 16360 311269 16384 311282
rect 16428 311269 16452 311282
rect 16496 311269 16520 311282
rect 16564 311269 16588 311282
rect 16632 311269 16656 311282
rect 17290 311269 17314 311282
rect 17358 311269 17382 311282
rect 17426 311269 17450 311282
rect 17494 311269 17518 311282
rect 17562 311269 17586 311282
rect 17630 311269 17654 311282
rect 17698 311269 17722 311282
rect 17766 311269 17790 311282
rect 17834 311269 17858 311282
rect 17902 311269 17926 311282
rect 17970 311269 17994 311282
rect 18038 311269 18062 311282
rect 18106 311269 18130 311282
rect 18174 311269 18198 311282
rect 19980 311048 20286 311218
rect 7389 310879 8389 310935
rect 8990 310879 9990 310935
rect 15678 310924 16678 310980
rect 17278 310924 18278 310980
rect 7389 310807 8389 310863
rect 8990 310807 9990 310863
rect 15678 310852 16678 310908
rect 17278 310852 18278 310908
rect 20945 310796 25553 311332
rect 28647 311268 28671 311302
rect 28647 311199 28671 311233
rect 28647 311154 28671 311164
rect 21413 310706 22813 310796
rect 23685 310706 25085 310796
rect 7389 310505 8389 310577
rect 8990 310505 9990 310577
rect 15678 310550 16678 310622
rect 17278 310550 18278 310622
rect 15748 310539 15782 310550
rect 15816 310539 15850 310550
rect 15884 310539 15918 310550
rect 15952 310539 15986 310550
rect 16020 310539 16054 310550
rect 16088 310539 16122 310550
rect 16156 310539 16190 310550
rect 16224 310539 16258 310550
rect 16292 310539 16326 310550
rect 16360 310539 16394 310550
rect 16428 310539 16462 310550
rect 16496 310539 16530 310550
rect 16564 310539 16598 310550
rect 16632 310539 16666 310550
rect 17290 310539 17324 310550
rect 17358 310539 17392 310550
rect 17426 310539 17460 310550
rect 17494 310539 17528 310550
rect 17562 310539 17596 310550
rect 17630 310539 17664 310550
rect 17698 310539 17732 310550
rect 17766 310539 17800 310550
rect 17834 310539 17868 310550
rect 17902 310539 17936 310550
rect 17970 310539 18004 310550
rect 18038 310539 18072 310550
rect 18106 310539 18140 310550
rect 18174 310539 18208 310550
rect 21413 310543 22813 310671
rect 23685 310543 25085 310671
rect 15748 310529 15806 310539
rect 15816 310529 15874 310539
rect 15884 310529 15942 310539
rect 15952 310529 16010 310539
rect 16020 310529 16078 310539
rect 16088 310529 16146 310539
rect 16156 310529 16214 310539
rect 16224 310529 16282 310539
rect 16292 310529 16350 310539
rect 16360 310529 16418 310539
rect 16428 310529 16486 310539
rect 16496 310529 16554 310539
rect 16564 310529 16622 310539
rect 16632 310529 16690 310539
rect 17290 310529 17348 310539
rect 17358 310529 17416 310539
rect 17426 310529 17484 310539
rect 17494 310529 17552 310539
rect 17562 310529 17620 310539
rect 17630 310529 17688 310539
rect 17698 310529 17756 310539
rect 17766 310529 17824 310539
rect 17834 310529 17892 310539
rect 17902 310529 17960 310539
rect 17970 310529 18028 310539
rect 18038 310529 18096 310539
rect 18106 310529 18164 310539
rect 18174 310529 18232 310539
rect 15724 310505 16690 310529
rect 17266 310505 18232 310529
rect 15748 310490 15772 310505
rect 15816 310490 15840 310505
rect 15884 310490 15908 310505
rect 15952 310490 15976 310505
rect 16020 310490 16044 310505
rect 16088 310490 16112 310505
rect 16156 310490 16180 310505
rect 16224 310490 16248 310505
rect 16292 310490 16316 310505
rect 16360 310490 16384 310505
rect 16428 310490 16452 310505
rect 16496 310490 16520 310505
rect 16564 310490 16588 310505
rect 16632 310490 16656 310505
rect 17290 310490 17314 310505
rect 17358 310490 17382 310505
rect 17426 310490 17450 310505
rect 17494 310490 17518 310505
rect 17562 310490 17586 310505
rect 17630 310490 17654 310505
rect 17698 310490 17722 310505
rect 17766 310490 17790 310505
rect 17834 310490 17858 310505
rect 17902 310490 17926 310505
rect 17970 310490 17994 310505
rect 18038 310490 18062 310505
rect 18106 310490 18130 310505
rect 18174 310490 18198 310505
rect 15678 310335 16678 310490
rect 7389 310245 8389 310305
rect 8990 310245 9990 310305
rect 15678 310301 16690 310335
rect 17278 310325 18278 310490
rect 21413 310380 22813 310508
rect 23685 310380 25085 310508
rect 17266 310301 18278 310325
rect 15678 310290 16678 310301
rect 17278 310290 18278 310301
rect 15748 310277 15772 310290
rect 15816 310277 15840 310290
rect 15884 310277 15908 310290
rect 15952 310277 15976 310290
rect 16020 310277 16044 310290
rect 16088 310277 16112 310290
rect 16156 310277 16180 310290
rect 16224 310277 16248 310290
rect 16292 310277 16316 310290
rect 16360 310277 16384 310290
rect 16428 310277 16452 310290
rect 16496 310277 16520 310290
rect 16564 310277 16588 310290
rect 16632 310277 16656 310290
rect 17290 310277 17314 310290
rect 17358 310277 17382 310290
rect 17426 310277 17450 310290
rect 17494 310277 17518 310290
rect 17562 310277 17586 310290
rect 17630 310277 17654 310290
rect 17698 310277 17722 310290
rect 17766 310277 17790 310290
rect 17834 310277 17858 310290
rect 17902 310277 17926 310290
rect 17970 310277 17994 310290
rect 18038 310277 18062 310290
rect 18106 310277 18130 310290
rect 18174 310277 18198 310290
rect 21413 310217 22813 310345
rect 23685 310217 25085 310345
rect 21413 310054 22813 310182
rect 23685 310054 25085 310182
rect 25936 310132 26936 310182
rect 27274 310033 27358 310036
rect 13899 309998 14059 310002
rect 7389 309887 8389 309943
rect 8990 309887 9990 309943
rect 15678 309932 16678 309988
rect 17278 309932 18278 309988
rect 7389 309815 8389 309871
rect 8990 309815 9990 309871
rect 15678 309860 16678 309916
rect 17278 309860 18278 309916
rect 21413 309891 22813 310019
rect 23685 309891 25085 310019
rect 25936 309976 26936 310032
rect 27158 309983 27358 310033
rect 13899 309852 14059 309856
rect 25936 309820 26936 309876
rect 27158 309807 27358 309935
rect 21413 309741 22813 309784
rect 23685 309741 25085 309784
rect 25936 309664 26936 309720
rect 7389 309513 8389 309585
rect 8990 309513 9990 309585
rect 15678 309558 16678 309630
rect 17278 309558 18278 309630
rect 21413 309605 22813 309648
rect 23685 309605 25085 309648
rect 27158 309631 27358 309687
rect 15748 309547 15782 309558
rect 15816 309547 15850 309558
rect 15884 309547 15918 309558
rect 15952 309547 15986 309558
rect 16020 309547 16054 309558
rect 16088 309547 16122 309558
rect 16156 309547 16190 309558
rect 16224 309547 16258 309558
rect 16292 309547 16326 309558
rect 16360 309547 16394 309558
rect 16428 309547 16462 309558
rect 16496 309547 16530 309558
rect 16564 309547 16598 309558
rect 16632 309547 16666 309558
rect 17290 309547 17324 309558
rect 17358 309547 17392 309558
rect 17426 309547 17460 309558
rect 17494 309547 17528 309558
rect 17562 309547 17596 309558
rect 17630 309547 17664 309558
rect 17698 309547 17732 309558
rect 17766 309547 17800 309558
rect 17834 309547 17868 309558
rect 17902 309547 17936 309558
rect 17970 309547 18004 309558
rect 18038 309547 18072 309558
rect 18106 309547 18140 309558
rect 18174 309547 18208 309558
rect 15748 309537 15806 309547
rect 15816 309537 15874 309547
rect 15884 309537 15942 309547
rect 15952 309537 16010 309547
rect 16020 309537 16078 309547
rect 16088 309537 16146 309547
rect 16156 309537 16214 309547
rect 16224 309537 16282 309547
rect 16292 309537 16350 309547
rect 16360 309537 16418 309547
rect 16428 309537 16486 309547
rect 16496 309537 16554 309547
rect 16564 309537 16622 309547
rect 16632 309537 16690 309547
rect 17290 309537 17348 309547
rect 17358 309537 17416 309547
rect 17426 309537 17484 309547
rect 17494 309537 17552 309547
rect 17562 309537 17620 309547
rect 17630 309537 17688 309547
rect 17698 309537 17756 309547
rect 17766 309537 17824 309547
rect 17834 309537 17892 309547
rect 17902 309537 17960 309547
rect 17970 309537 18028 309547
rect 18038 309537 18096 309547
rect 18106 309537 18164 309547
rect 18174 309537 18232 309547
rect 15724 309513 16690 309537
rect 17266 309513 18232 309537
rect 15748 309498 15772 309513
rect 15816 309498 15840 309513
rect 15884 309498 15908 309513
rect 15952 309498 15976 309513
rect 16020 309498 16044 309513
rect 16088 309498 16112 309513
rect 16156 309498 16180 309513
rect 16224 309498 16248 309513
rect 16292 309498 16316 309513
rect 16360 309498 16384 309513
rect 16428 309498 16452 309513
rect 16496 309498 16520 309513
rect 16564 309498 16588 309513
rect 16632 309498 16656 309513
rect 17290 309498 17314 309513
rect 17358 309498 17382 309513
rect 17426 309498 17450 309513
rect 17494 309498 17518 309513
rect 17562 309498 17586 309513
rect 17630 309498 17654 309513
rect 17698 309498 17722 309513
rect 17766 309498 17790 309513
rect 17834 309498 17858 309513
rect 17902 309498 17926 309513
rect 17970 309498 17994 309513
rect 18038 309498 18062 309513
rect 18106 309498 18130 309513
rect 18174 309498 18198 309513
rect 15678 309343 16678 309498
rect 7389 309253 8389 309313
rect 8990 309253 9990 309313
rect 15678 309309 16690 309343
rect 17278 309333 18278 309498
rect 21413 309442 22813 309570
rect 23685 309442 25085 309570
rect 25936 309514 26936 309564
rect 26393 309511 26477 309514
rect 26726 309511 26810 309514
rect 27158 309455 27358 309583
rect 17266 309309 18278 309333
rect 15678 309298 16678 309309
rect 17278 309298 18278 309309
rect 15748 309285 15772 309298
rect 15816 309285 15840 309298
rect 15884 309285 15908 309298
rect 15952 309285 15976 309298
rect 16020 309285 16044 309298
rect 16088 309285 16112 309298
rect 16156 309285 16180 309298
rect 16224 309285 16248 309298
rect 16292 309285 16316 309298
rect 16360 309285 16384 309298
rect 16428 309285 16452 309298
rect 16496 309285 16520 309298
rect 16564 309285 16588 309298
rect 16632 309285 16656 309298
rect 17290 309285 17314 309298
rect 17358 309285 17382 309298
rect 17426 309285 17450 309298
rect 17494 309285 17518 309298
rect 17562 309285 17586 309298
rect 17630 309285 17654 309298
rect 17698 309285 17722 309298
rect 17766 309285 17790 309298
rect 17834 309285 17858 309298
rect 17902 309285 17926 309298
rect 17970 309285 17994 309298
rect 18038 309285 18062 309298
rect 18106 309285 18130 309298
rect 18174 309285 18198 309298
rect 21413 309279 22813 309407
rect 23685 309279 25085 309407
rect 27158 309279 27358 309335
rect 21413 309116 22813 309244
rect 23685 309116 25085 309244
rect 27158 309103 27358 309231
rect 26393 309100 26477 309103
rect 26726 309100 26810 309103
rect 12543 309069 12881 309085
rect 12559 308967 12865 309069
rect 7389 308895 8389 308951
rect 8990 308895 9990 308951
rect 15678 308940 16678 308996
rect 17278 308940 18278 308996
rect 21413 308953 22813 309081
rect 23685 308953 25085 309081
rect 25936 309050 26936 309100
rect 27622 309095 27672 310095
rect 27772 309095 27828 310095
rect 27928 309095 27984 310095
rect 28084 309095 28140 310095
rect 28240 309095 28296 310095
rect 28396 309637 28446 310095
rect 28396 309553 28449 309637
rect 28396 309305 28446 309553
rect 29778 309320 29802 309344
rect 28396 309221 28449 309305
rect 29802 309296 29826 309309
rect 29880 309299 29914 309333
rect 29778 309261 29802 309285
rect 29890 309275 29914 309299
rect 28396 309095 28446 309221
rect 7389 308823 8389 308879
rect 8990 308823 9990 308879
rect 15678 308868 16678 308924
rect 17278 308868 18278 308924
rect 21413 308790 22813 308918
rect 23685 308790 25085 308918
rect 25936 308894 26936 308950
rect 27158 308927 27358 308983
rect 13899 308656 14059 308660
rect 7389 308521 8389 308593
rect 8990 308521 9990 308593
rect 15678 308566 16678 308638
rect 17278 308566 18278 308638
rect 21413 308627 22813 308755
rect 23685 308627 25085 308755
rect 25936 308738 26936 308794
rect 27158 308751 27358 308879
rect 27912 308757 27962 308873
rect 27909 308673 27962 308757
rect 28082 308673 28210 308873
rect 28258 308673 28314 308873
rect 28434 308673 28562 308873
rect 28610 308673 28660 308873
rect 27917 308669 27951 308673
rect 29880 308672 29914 308706
rect 25936 308582 26936 308638
rect 27158 308581 27358 308631
rect 27274 308578 27358 308581
rect 15748 308555 15782 308566
rect 15816 308555 15850 308566
rect 15884 308555 15918 308566
rect 15952 308555 15986 308566
rect 16020 308555 16054 308566
rect 16088 308555 16122 308566
rect 16156 308555 16190 308566
rect 16224 308555 16258 308566
rect 16292 308555 16326 308566
rect 16360 308555 16394 308566
rect 16428 308555 16462 308566
rect 16496 308555 16530 308566
rect 16564 308555 16598 308566
rect 16632 308555 16666 308566
rect 17290 308555 17324 308566
rect 17358 308555 17392 308566
rect 17426 308555 17460 308566
rect 17494 308555 17528 308566
rect 17562 308555 17596 308566
rect 17630 308555 17664 308566
rect 17698 308555 17732 308566
rect 17766 308555 17800 308566
rect 17834 308555 17868 308566
rect 17902 308555 17936 308566
rect 17970 308555 18004 308566
rect 18038 308555 18072 308566
rect 18106 308555 18140 308566
rect 18174 308555 18208 308566
rect 15748 308545 15806 308555
rect 15816 308545 15874 308555
rect 15884 308545 15942 308555
rect 15952 308545 16010 308555
rect 16020 308545 16078 308555
rect 16088 308545 16146 308555
rect 16156 308545 16214 308555
rect 16224 308545 16282 308555
rect 16292 308545 16350 308555
rect 16360 308545 16418 308555
rect 16428 308545 16486 308555
rect 16496 308545 16554 308555
rect 16564 308545 16622 308555
rect 16632 308545 16690 308555
rect 17290 308545 17348 308555
rect 17358 308545 17416 308555
rect 17426 308545 17484 308555
rect 17494 308545 17552 308555
rect 17562 308545 17620 308555
rect 17630 308545 17688 308555
rect 17698 308545 17756 308555
rect 17766 308545 17824 308555
rect 17834 308545 17892 308555
rect 17902 308545 17960 308555
rect 17970 308545 18028 308555
rect 18038 308545 18096 308555
rect 18106 308545 18164 308555
rect 18174 308545 18232 308555
rect 15724 308521 16690 308545
rect 17266 308521 18232 308545
rect 13901 308510 14061 308514
rect 15748 308506 15772 308521
rect 15816 308506 15840 308521
rect 15884 308506 15908 308521
rect 15952 308506 15976 308521
rect 16020 308506 16044 308521
rect 16088 308506 16112 308521
rect 16156 308506 16180 308521
rect 16224 308506 16248 308521
rect 16292 308506 16316 308521
rect 16360 308506 16384 308521
rect 16428 308506 16452 308521
rect 16496 308506 16520 308521
rect 16564 308506 16588 308521
rect 16632 308506 16656 308521
rect 17290 308506 17314 308521
rect 17358 308506 17382 308521
rect 17426 308506 17450 308521
rect 17494 308506 17518 308521
rect 17562 308506 17586 308521
rect 17630 308506 17654 308521
rect 17698 308506 17722 308521
rect 17766 308506 17790 308521
rect 17834 308506 17858 308521
rect 17902 308506 17926 308521
rect 17970 308506 17994 308521
rect 18038 308506 18062 308521
rect 18106 308506 18130 308521
rect 18174 308506 18198 308521
rect 15678 308351 16678 308506
rect 7389 308261 8389 308321
rect 8990 308261 9990 308321
rect 15678 308317 16690 308351
rect 17278 308341 18278 308506
rect 21413 308470 22813 308520
rect 23685 308470 25085 308520
rect 25936 308432 26936 308482
rect 21349 308390 21373 308414
rect 21407 308390 21431 308414
rect 25067 308390 25091 308414
rect 25125 308390 25149 308414
rect 21383 308356 21397 308390
rect 25101 308356 25115 308390
rect 17266 308317 18278 308341
rect 21349 308332 21373 308356
rect 21407 308332 21431 308356
rect 25067 308332 25091 308356
rect 25125 308332 25149 308356
rect 27917 308325 27951 308329
rect 15678 308306 16678 308317
rect 17278 308306 18278 308317
rect 15748 308293 15772 308306
rect 15816 308293 15840 308306
rect 15884 308293 15908 308306
rect 15952 308293 15976 308306
rect 16020 308293 16044 308306
rect 16088 308293 16112 308306
rect 16156 308293 16180 308306
rect 16224 308293 16248 308306
rect 16292 308293 16316 308306
rect 16360 308293 16384 308306
rect 16428 308293 16452 308306
rect 16496 308293 16520 308306
rect 16564 308293 16588 308306
rect 16632 308293 16656 308306
rect 17290 308293 17314 308306
rect 17358 308293 17382 308306
rect 17426 308293 17450 308306
rect 17494 308293 17518 308306
rect 17562 308293 17586 308306
rect 17630 308293 17654 308306
rect 17698 308293 17722 308306
rect 17766 308293 17790 308306
rect 17834 308293 17858 308306
rect 17902 308293 17926 308306
rect 17970 308293 17994 308306
rect 18038 308293 18062 308306
rect 18106 308293 18130 308306
rect 18174 308293 18198 308306
rect 27909 308241 27962 308325
rect 21634 308101 24864 308203
rect 27912 308125 27962 308241
rect 28082 308125 28210 308325
rect 28258 308125 28314 308325
rect 28434 308125 28562 308325
rect 28610 308125 28660 308325
rect 21186 308047 21210 308071
rect 25288 308047 25312 308071
rect 21162 308023 21186 308037
rect 25312 308023 25336 308037
rect 7389 307903 8389 307959
rect 8990 307903 9990 307959
rect 15678 307948 16678 308004
rect 17278 307948 18278 308004
rect 21072 307989 21084 308013
rect 21186 307989 21210 308013
rect 25288 307989 25312 308013
rect 25414 307989 25426 308013
rect 21385 307944 21403 307948
rect 7389 307831 8389 307887
rect 8990 307831 9990 307887
rect 15678 307876 16678 307932
rect 17278 307876 18278 307932
rect 20250 307914 20316 307930
rect 21377 307914 21403 307944
rect 21385 307904 21403 307914
rect 21383 307880 21403 307904
rect 21407 307880 21415 307914
rect 25113 307904 25121 307944
rect 25101 307880 25121 307904
rect 25125 307880 25143 307948
rect 21383 307846 21419 307880
rect 25101 307846 25147 307880
rect 21383 307812 21403 307846
rect 21407 307812 21415 307846
rect 21383 307778 21419 307812
rect 21481 307784 22881 307834
rect 23617 307784 25017 307834
rect 25101 307812 25121 307846
rect 25125 307812 25143 307846
rect 25101 307778 25147 307812
rect 21383 307744 21403 307778
rect 21407 307744 21415 307778
rect 21383 307710 21419 307744
rect 21383 307676 21403 307710
rect 21407 307676 21415 307710
rect 7389 307529 8389 307601
rect 8990 307529 9990 307601
rect 15678 307574 16678 307646
rect 17278 307574 18278 307646
rect 21383 307642 21419 307676
rect 21383 307608 21403 307642
rect 21407 307608 21415 307642
rect 21481 307621 22881 307749
rect 23617 307621 25017 307749
rect 25101 307744 25121 307778
rect 25125 307744 25143 307778
rect 25101 307710 25147 307744
rect 25101 307676 25121 307710
rect 25125 307676 25143 307710
rect 25101 307642 25147 307676
rect 25101 307608 25121 307642
rect 25125 307608 25143 307642
rect 21383 307574 21419 307608
rect 15748 307563 15782 307574
rect 15816 307563 15850 307574
rect 15884 307563 15918 307574
rect 15952 307563 15986 307574
rect 16020 307563 16054 307574
rect 16088 307563 16122 307574
rect 16156 307563 16190 307574
rect 16224 307563 16258 307574
rect 16292 307563 16326 307574
rect 16360 307563 16394 307574
rect 16428 307563 16462 307574
rect 16496 307563 16530 307574
rect 16564 307563 16598 307574
rect 16632 307563 16666 307574
rect 17290 307563 17324 307574
rect 17358 307563 17392 307574
rect 17426 307563 17460 307574
rect 17494 307563 17528 307574
rect 17562 307563 17596 307574
rect 17630 307563 17664 307574
rect 17698 307563 17732 307574
rect 17766 307563 17800 307574
rect 17834 307563 17868 307574
rect 17902 307563 17936 307574
rect 17970 307563 18004 307574
rect 18038 307563 18072 307574
rect 18106 307563 18140 307574
rect 18174 307563 18208 307574
rect 15748 307553 15806 307563
rect 15816 307553 15874 307563
rect 15884 307553 15942 307563
rect 15952 307553 16010 307563
rect 16020 307553 16078 307563
rect 16088 307553 16146 307563
rect 16156 307553 16214 307563
rect 16224 307553 16282 307563
rect 16292 307553 16350 307563
rect 16360 307553 16418 307563
rect 16428 307553 16486 307563
rect 16496 307553 16554 307563
rect 16564 307553 16622 307563
rect 16632 307553 16690 307563
rect 17290 307553 17348 307563
rect 17358 307553 17416 307563
rect 17426 307553 17484 307563
rect 17494 307553 17552 307563
rect 17562 307553 17620 307563
rect 17630 307553 17688 307563
rect 17698 307553 17756 307563
rect 17766 307553 17824 307563
rect 17834 307553 17892 307563
rect 17902 307553 17960 307563
rect 17970 307553 18028 307563
rect 18038 307553 18096 307563
rect 18106 307553 18164 307563
rect 18174 307553 18232 307563
rect 15724 307529 16690 307553
rect 17266 307529 18232 307553
rect 21383 307540 21403 307574
rect 21407 307540 21415 307574
rect 15748 307514 15772 307529
rect 15816 307514 15840 307529
rect 15884 307514 15908 307529
rect 15952 307514 15976 307529
rect 16020 307514 16044 307529
rect 16088 307514 16112 307529
rect 16156 307514 16180 307529
rect 16224 307514 16248 307529
rect 16292 307514 16316 307529
rect 16360 307514 16384 307529
rect 16428 307514 16452 307529
rect 16496 307514 16520 307529
rect 16564 307514 16588 307529
rect 16632 307514 16656 307529
rect 17290 307514 17314 307529
rect 17358 307514 17382 307529
rect 17426 307514 17450 307529
rect 17494 307514 17518 307529
rect 17562 307514 17586 307529
rect 17630 307514 17654 307529
rect 17698 307514 17722 307529
rect 17766 307514 17790 307529
rect 17834 307514 17858 307529
rect 17902 307514 17926 307529
rect 17970 307514 17994 307529
rect 18038 307514 18062 307529
rect 18106 307514 18130 307529
rect 18174 307514 18198 307529
rect 5937 307318 6089 307386
rect 15678 307359 16678 307514
rect 6005 307315 6089 307318
rect 5967 307305 6059 307315
rect 6005 307275 6021 307305
rect 1288 305503 1338 306503
rect 1438 305503 1566 306503
rect 1594 305503 1644 306503
rect 5995 305493 6021 307275
rect 7389 307269 8389 307329
rect 8990 307269 9990 307329
rect 15678 307325 16690 307359
rect 17278 307349 18278 307514
rect 17266 307325 18278 307349
rect 15678 307314 16678 307325
rect 17278 307314 18278 307325
rect 21383 307506 21419 307540
rect 21383 307472 21403 307506
rect 21407 307472 21415 307506
rect 21383 307438 21419 307472
rect 21481 307458 22881 307586
rect 23617 307458 25017 307586
rect 25101 307574 25147 307608
rect 25101 307540 25121 307574
rect 25125 307540 25143 307574
rect 25101 307506 25147 307540
rect 25101 307472 25121 307506
rect 25125 307472 25143 307506
rect 25101 307438 25147 307472
rect 21383 307404 21403 307438
rect 21407 307404 21415 307438
rect 21383 307370 21419 307404
rect 21383 307336 21403 307370
rect 21407 307336 21415 307370
rect 15748 307301 15772 307314
rect 15816 307301 15840 307314
rect 15884 307301 15908 307314
rect 15952 307301 15976 307314
rect 16020 307301 16044 307314
rect 16088 307301 16112 307314
rect 16156 307301 16180 307314
rect 16224 307301 16248 307314
rect 16292 307301 16316 307314
rect 16360 307301 16384 307314
rect 16428 307301 16452 307314
rect 16496 307301 16520 307314
rect 16564 307301 16588 307314
rect 16632 307301 16656 307314
rect 17290 307301 17314 307314
rect 17358 307301 17382 307314
rect 17426 307301 17450 307314
rect 17494 307301 17518 307314
rect 17562 307301 17586 307314
rect 17630 307301 17654 307314
rect 17698 307301 17722 307314
rect 17766 307301 17790 307314
rect 17834 307301 17858 307314
rect 17902 307301 17926 307314
rect 17970 307301 17994 307314
rect 18038 307301 18062 307314
rect 18106 307301 18130 307314
rect 18174 307301 18198 307314
rect 21383 307302 21419 307336
rect 21383 307268 21403 307302
rect 21407 307268 21415 307302
rect 21481 307295 22881 307423
rect 23617 307295 25017 307423
rect 25101 307404 25121 307438
rect 25125 307404 25143 307438
rect 25101 307370 25147 307404
rect 25101 307336 25121 307370
rect 25125 307336 25143 307370
rect 25101 307302 25147 307336
rect 25101 307268 25121 307302
rect 25125 307268 25143 307302
rect 21383 307234 21419 307268
rect 21383 307200 21403 307234
rect 21407 307200 21415 307234
rect 21383 307166 21419 307200
rect 21383 307132 21403 307166
rect 21407 307132 21415 307166
rect 21481 307132 22881 307260
rect 23617 307132 25017 307260
rect 25101 307234 25147 307268
rect 25101 307200 25121 307234
rect 25125 307200 25143 307234
rect 25101 307166 25147 307200
rect 25101 307132 25121 307166
rect 25125 307132 25143 307166
rect 21383 307098 21419 307132
rect 25101 307098 25147 307132
rect 21383 307064 21403 307098
rect 21407 307064 21415 307098
rect 21383 307030 21419 307064
rect 7389 306911 8389 306967
rect 8990 306911 9990 306967
rect 15678 306956 16678 307012
rect 17278 306956 18278 307012
rect 21383 306996 21403 307030
rect 21407 306996 21415 307030
rect 21383 306962 21419 306996
rect 21481 306969 22881 307097
rect 23617 306969 25017 307097
rect 25101 307064 25121 307098
rect 25125 307064 25143 307098
rect 25101 307030 25147 307064
rect 25101 306996 25121 307030
rect 25125 306996 25143 307030
rect 25101 306962 25147 306996
rect 26478 306985 26648 307291
rect 7389 306839 8389 306895
rect 8990 306839 9990 306895
rect 15678 306884 16678 306940
rect 17278 306884 18278 306940
rect 21383 306928 21403 306962
rect 21407 306928 21415 306962
rect 21383 306894 21419 306928
rect 21383 306860 21403 306894
rect 21407 306860 21415 306894
rect 21383 306826 21419 306860
rect 21383 306792 21403 306826
rect 21407 306792 21415 306826
rect 21481 306806 22881 306934
rect 23617 306806 25017 306934
rect 25101 306928 25121 306962
rect 25125 306928 25143 306962
rect 25101 306894 25147 306928
rect 27622 306903 27672 307903
rect 27772 306903 27828 307903
rect 27928 306903 27984 307903
rect 28084 306903 28140 307903
rect 28240 306903 28296 307903
rect 28396 307777 28446 307903
rect 28396 307693 28449 307777
rect 28396 307445 28446 307693
rect 30015 307523 30027 313246
rect 32596 313239 33596 313367
rect 35255 313345 36255 313401
rect 30135 313062 30735 313112
rect 31049 313042 32049 313092
rect 32596 313083 33596 313211
rect 35255 313169 36255 313297
rect 35255 312993 36255 313121
rect 30135 312886 30735 312942
rect 31049 312886 32049 312942
rect 32596 312927 33596 312983
rect 37998 312979 38148 312991
rect 38317 312979 38467 312991
rect 30135 312716 30735 312766
rect 31049 312736 32049 312786
rect 32596 312777 33596 312827
rect 35255 312823 36255 312873
rect 37998 312866 38598 312916
rect 35255 312754 36255 312766
rect 37998 312690 38598 312746
rect 30135 312600 30735 312650
rect 31049 312600 32049 312650
rect 32596 312575 33196 312625
rect 35255 312621 36255 312671
rect 30135 312424 30735 312480
rect 31049 312444 32049 312500
rect 30135 312248 30735 312376
rect 31049 312288 32049 312344
rect 30135 312072 30735 312200
rect 31049 312132 32049 312188
rect 32596 312141 33196 312191
rect 30135 311896 30735 312024
rect 31049 311982 32049 312032
rect 31049 311866 32049 311916
rect 30135 311726 30735 311776
rect 31049 311710 32049 311838
rect 30135 311610 30735 311660
rect 30135 311434 30735 311562
rect 31049 311554 32049 311682
rect 31049 311398 32049 311526
rect 34152 311490 34202 312478
rect 34322 311490 34372 312478
rect 34492 312465 35092 312515
rect 35255 312445 36255 312573
rect 37998 312520 38598 312570
rect 36785 312496 36797 312500
rect 36785 312485 36800 312496
rect 36970 312485 36985 312500
rect 34492 312289 35092 312345
rect 35255 312269 36255 312325
rect 36785 312305 36985 312485
rect 36785 312294 36800 312305
rect 36785 312290 36797 312294
rect 36970 312290 36985 312305
rect 37083 312485 37098 312500
rect 37083 312305 37120 312485
rect 37083 312290 37098 312305
rect 36785 312260 36797 312264
rect 36785 312249 36800 312260
rect 36970 312249 36985 312264
rect 34492 312119 35092 312169
rect 35255 312099 36255 312149
rect 36785 312069 36985 312249
rect 696597 312200 696600 312320
rect 37993 312094 38593 312144
rect 36785 312058 36800 312069
rect 36785 312054 36797 312058
rect 36970 312054 36985 312069
rect 692376 311983 692396 312017
rect 692463 311993 692532 312017
rect 696191 311993 696239 312017
rect 692487 311983 692532 311993
rect 696204 311983 696239 311993
rect 696340 311983 696360 312017
rect 34491 311849 35091 311899
rect 35255 311883 35855 311933
rect 37993 311924 38593 311974
rect 692487 311915 692502 311939
rect 696200 311915 696215 311939
rect 692454 311891 692478 311915
rect 696224 311891 696248 311915
rect 686755 311800 687355 311850
rect 34491 311673 35091 311729
rect 35255 311707 35855 311763
rect 36785 311748 37385 311798
rect 38920 311761 38946 311787
rect 692487 311748 692505 311752
rect 692479 311718 692505 311748
rect 692487 311698 692505 311718
rect 34491 311503 35091 311553
rect 35255 311531 35855 311659
rect 36785 311572 37385 311628
rect 686755 311624 687355 311680
rect 692485 311674 692505 311698
rect 692509 311674 692517 311718
rect 696215 311698 696223 311748
rect 696203 311674 696223 311698
rect 696227 311674 696245 311752
rect 692485 311640 692521 311674
rect 696203 311640 696249 311674
rect 34019 311418 34029 311490
rect 34152 311478 34372 311490
rect 34091 311415 34101 311418
rect 30135 311258 30735 311314
rect 31049 311242 32049 311370
rect 34091 311365 35091 311415
rect 35255 311361 35855 311411
rect 36785 311396 37385 311452
rect 686755 311448 687355 311504
rect 686755 311278 687355 311328
rect 30135 311082 30735 311210
rect 31049 311086 32049 311214
rect 34091 311195 35091 311245
rect 36785 311226 37385 311276
rect 34091 311192 34101 311195
rect 34202 311192 34302 311195
rect 35255 311159 35855 311209
rect 30135 310912 30735 310962
rect 31049 310930 32049 310986
rect 30135 310796 30735 310846
rect 31049 310774 32049 310902
rect 32481 310898 33081 310948
rect 30135 310620 30735 310748
rect 31049 310618 32049 310746
rect 32481 310742 33081 310870
rect 30135 310444 30735 310572
rect 31049 310462 32049 310590
rect 32481 310586 33081 310714
rect 34152 310532 34202 311132
rect 34302 310532 34352 311132
rect 34491 311066 35091 311116
rect 35255 311003 35855 311131
rect 36785 311094 37385 311144
rect 685547 311102 686147 311152
rect 687155 311007 687170 311022
rect 687343 311018 687355 311022
rect 687340 311007 687355 311018
rect 34491 310890 35091 310946
rect 36785 310918 37385 310974
rect 685547 310932 686147 310982
rect 35255 310847 35855 310903
rect 687155 310827 687355 311007
rect 34491 310720 35091 310770
rect 35255 310691 35855 310819
rect 687155 310812 687170 310827
rect 687340 310816 687355 310827
rect 687343 310812 687355 310816
rect 36785 310742 37385 310798
rect 687042 310771 687057 310786
rect 35255 310541 35855 310591
rect 36785 310572 37385 310622
rect 687020 310591 687057 310771
rect 687155 310771 687170 310786
rect 687343 310782 687355 310786
rect 687340 310771 687355 310782
rect 687155 310591 687355 310771
rect 688210 310630 688260 311630
rect 688360 310740 688488 311630
rect 688516 310740 688644 311630
rect 688672 310740 688800 311630
rect 688828 310740 688956 311630
rect 688984 310740 689112 311630
rect 689140 310740 689268 311630
rect 689296 310740 689424 311630
rect 689452 310740 689580 311630
rect 689608 310740 689736 311630
rect 689764 310740 689892 311630
rect 689920 310740 690048 311630
rect 690076 310740 690204 311630
rect 690232 310740 690360 311630
rect 690388 310630 690438 311630
rect 692485 311606 692505 311640
rect 692509 311606 692517 311640
rect 696203 311606 696223 311640
rect 696227 311606 696245 311640
rect 691275 311523 691875 311573
rect 692485 311572 692521 311606
rect 696203 311572 696249 311606
rect 692485 311538 692505 311572
rect 692509 311538 692517 311572
rect 692485 311504 692521 311538
rect 692583 311528 693983 311571
rect 694719 311528 696119 311571
rect 696203 311538 696223 311572
rect 696227 311538 696245 311572
rect 696203 311504 696249 311538
rect 692485 311470 692505 311504
rect 692509 311470 692517 311504
rect 692485 311436 692521 311470
rect 691275 311373 691875 311423
rect 692485 311402 692505 311436
rect 692509 311402 692517 311436
rect 692485 311368 692521 311402
rect 692485 311334 692505 311368
rect 692509 311334 692517 311368
rect 692583 311365 693983 311493
rect 694719 311365 696119 311493
rect 696203 311470 696223 311504
rect 696227 311470 696245 311504
rect 696203 311436 696249 311470
rect 707624 311441 707658 311475
rect 707695 311441 707729 311475
rect 707769 311441 707803 311475
rect 707840 311441 707874 311475
rect 707914 311441 707948 311475
rect 707985 311441 708019 311475
rect 708059 311441 708093 311475
rect 708130 311441 708164 311475
rect 708204 311441 708238 311475
rect 708275 311441 708309 311475
rect 708369 311441 708403 311475
rect 708446 311441 708480 311475
rect 708520 311441 708554 311465
rect 708588 311441 708610 311465
rect 709211 311441 709234 311465
rect 709270 311441 709304 311475
rect 709364 311441 709398 311475
rect 709435 311441 709469 311475
rect 709509 311441 709543 311475
rect 709580 311441 709614 311475
rect 709654 311441 709688 311475
rect 709725 311441 709759 311475
rect 709799 311441 709833 311475
rect 709870 311441 709904 311475
rect 709944 311441 709978 311475
rect 710015 311441 710049 311475
rect 710089 311441 710123 311475
rect 710160 311441 710194 311475
rect 696203 311402 696223 311436
rect 696227 311402 696245 311436
rect 707610 311431 707624 311441
rect 707658 311431 707695 311441
rect 707729 311431 707769 311441
rect 707803 311431 707840 311441
rect 707874 311431 707914 311441
rect 707948 311431 707985 311441
rect 708019 311431 708059 311441
rect 708093 311431 708130 311441
rect 708164 311431 708204 311441
rect 708238 311431 708275 311441
rect 708309 311431 708369 311441
rect 708403 311431 708446 311441
rect 708480 311431 708520 311441
rect 708554 311431 708588 311441
rect 708610 311431 708634 311441
rect 709211 311431 709270 311441
rect 709304 311431 709364 311441
rect 709398 311431 709435 311441
rect 709469 311431 709509 311441
rect 709543 311431 709580 311441
rect 709614 311431 709654 311441
rect 709688 311431 709725 311441
rect 709759 311431 709799 311441
rect 709833 311431 709870 311441
rect 709904 311431 709944 311441
rect 709978 311431 710015 311441
rect 710049 311431 710089 311441
rect 710123 311431 710160 311441
rect 710194 311431 710211 311441
rect 696203 311368 696249 311402
rect 696203 311334 696223 311368
rect 696227 311334 696245 311368
rect 707610 311337 708610 311431
rect 709211 311337 710211 311431
rect 691275 311251 691875 311301
rect 692485 311300 692521 311334
rect 692485 311266 692505 311300
rect 692509 311266 692517 311300
rect 692485 311232 692521 311266
rect 692485 311198 692505 311232
rect 692509 311198 692517 311232
rect 692583 311202 693983 311330
rect 694719 311202 696119 311330
rect 696203 311300 696249 311334
rect 711579 311317 712463 311331
rect 711579 311307 711619 311317
rect 696203 311266 696223 311300
rect 696227 311266 696245 311300
rect 701730 311290 701747 311292
rect 696203 311232 696249 311266
rect 696203 311198 696223 311232
rect 696227 311198 696245 311232
rect 701692 311220 701722 311254
rect 701730 311220 701760 311290
rect 707610 311241 708610 311301
rect 709211 311241 710211 311301
rect 692485 311164 692521 311198
rect 691275 311101 691875 311151
rect 692485 311130 692505 311164
rect 692509 311130 692517 311164
rect 692485 311096 692521 311130
rect 692485 311062 692505 311096
rect 692509 311062 692517 311096
rect 692485 311028 692521 311062
rect 692583 311039 693983 311167
rect 694719 311039 696119 311167
rect 696203 311164 696249 311198
rect 696203 311130 696223 311164
rect 696227 311130 696245 311164
rect 696203 311096 696249 311130
rect 696203 311062 696223 311096
rect 696227 311062 696245 311096
rect 699322 311064 700322 311097
rect 700922 311064 701922 311097
rect 696203 311028 696249 311062
rect 707610 311044 708610 311048
rect 709211 311044 710211 311048
rect 691275 310975 691875 311025
rect 692485 310994 692505 311028
rect 692509 310994 692517 311028
rect 692485 310960 692521 310994
rect 692485 310926 692505 310960
rect 692509 310926 692517 310960
rect 692485 310892 692521 310926
rect 691275 310825 691875 310875
rect 692485 310858 692505 310892
rect 692509 310858 692517 310892
rect 692583 310876 693983 311004
rect 694719 310876 696119 311004
rect 696203 310994 696223 311028
rect 696227 310994 696245 311028
rect 707574 310994 708646 311030
rect 696203 310960 696249 310994
rect 696203 310926 696223 310960
rect 696227 310926 696245 310960
rect 707574 310953 707610 310994
rect 708610 310953 708646 310994
rect 696203 310892 696249 310926
rect 697284 310894 697350 310910
rect 707574 310897 708646 310953
rect 696203 310858 696223 310892
rect 696227 310858 696245 310892
rect 699322 310877 700322 310894
rect 700922 310877 701922 310894
rect 707574 310881 707610 310897
rect 708610 310881 708646 310897
rect 692485 310824 692521 310858
rect 692485 310790 692505 310824
rect 692509 310790 692517 310824
rect 692485 310756 692521 310790
rect 691275 310703 691875 310753
rect 692485 310740 692505 310756
rect 692509 310740 692517 310756
rect 692583 310740 693983 310841
rect 694719 310740 696119 310841
rect 696203 310824 696249 310858
rect 707574 310825 708646 310881
rect 696203 310790 696223 310824
rect 696227 310790 696245 310824
rect 696203 310756 696249 310790
rect 696203 310740 696223 310756
rect 696227 310740 696245 310756
rect 699322 310740 700322 310811
rect 700922 310740 701922 310811
rect 707574 310788 707610 310825
rect 708610 310788 708646 310825
rect 707574 310748 708646 310788
rect 709175 310994 710247 311030
rect 709175 310953 709211 310994
rect 710211 310953 710247 310994
rect 709175 310897 710247 310953
rect 709175 310881 709211 310897
rect 710211 310881 710247 310897
rect 709175 310825 710247 310881
rect 709175 310788 709211 310825
rect 710211 310788 710247 310825
rect 709175 310748 710247 310788
rect 685542 310506 686142 310556
rect 691275 310553 691875 310603
rect 32481 310436 33081 310486
rect 30135 310268 30735 310396
rect 31049 310306 32049 310434
rect 34491 310379 35091 310429
rect 37993 310396 38593 310446
rect 32481 310306 33081 310356
rect 33261 310287 33861 310323
rect 30135 310092 30735 310220
rect 31049 310150 32049 310278
rect 32481 310150 33081 310278
rect 34491 310203 35091 310331
rect 35255 310287 35855 310337
rect 685542 310330 686142 310386
rect 36785 310312 36797 310316
rect 36785 310301 36800 310312
rect 36970 310301 36985 310316
rect 35255 310131 35855 310259
rect 36785 310121 36985 310301
rect 37993 310226 38593 310276
rect 692583 310237 693983 310280
rect 694719 310237 696119 310280
rect 699322 310278 700322 310418
rect 700922 310278 701922 310418
rect 685542 310160 686142 310210
rect 36785 310110 36800 310121
rect 36785 310106 36797 310110
rect 36970 310106 36985 310121
rect 30135 309916 30735 310044
rect 31049 309994 32049 310050
rect 32481 309994 33081 310050
rect 34491 310027 35091 310083
rect 31049 309818 32049 309946
rect 32481 309838 33081 309966
rect 33261 309907 33861 309963
rect 34491 309851 35091 309979
rect 35255 309975 35855 310103
rect 692583 310101 693983 310144
rect 694719 310101 696119 310144
rect 36785 310076 36797 310080
rect 36785 310065 36800 310076
rect 36970 310065 36985 310080
rect 36785 309885 36985 310065
rect 35255 309819 35855 309875
rect 36785 309874 36800 309885
rect 36785 309870 36797 309874
rect 36970 309870 36985 309885
rect 37083 310065 37098 310080
rect 37083 309885 37120 310065
rect 37083 309870 37098 309885
rect 37998 309800 38598 309850
rect 30135 309740 30735 309796
rect 30135 309564 30735 309692
rect 31049 309642 32049 309770
rect 32481 309688 33081 309738
rect 33261 309723 33861 309773
rect 34491 309681 35091 309731
rect 35255 309669 35855 309719
rect 37998 309624 38598 309680
rect 680215 309678 680815 309728
rect 30135 309388 30735 309516
rect 31049 309466 32049 309594
rect 32481 309558 33081 309608
rect 30135 309212 30735 309340
rect 31049 309290 32049 309418
rect 32481 309402 33081 309458
rect 37998 309454 38598 309504
rect 680215 309502 680815 309558
rect 685551 309516 686551 309566
rect 689154 309480 689204 309897
rect 689304 309480 689360 309897
rect 689460 309480 689516 309897
rect 689616 309480 689672 309897
rect 689772 309480 689828 309897
rect 689928 309480 689978 309897
rect 699322 309860 700322 309916
rect 700922 309860 701922 309916
rect 707610 309905 708610 309961
rect 709211 309905 710211 309961
rect 699322 309788 700322 309844
rect 700922 309788 701922 309844
rect 707610 309833 708610 309889
rect 709211 309833 710211 309889
rect 711579 309525 711605 311307
rect 715956 310297 716006 311297
rect 716106 310740 716234 311297
rect 716262 310297 716312 311297
rect 711579 309480 711595 309495
rect 712409 309480 712431 309485
rect 713640 309480 713641 309785
rect 713750 309772 714750 309822
rect 713750 309562 714750 309612
rect 713750 309480 714750 309496
rect 37998 309451 38220 309454
rect 38245 309451 38539 309454
rect 32481 309252 33081 309302
rect 34427 309259 35027 309309
rect 30135 309036 30735 309164
rect 31049 309114 32049 309242
rect 33672 309183 34272 309233
rect 34427 309083 35027 309211
rect 30135 308860 30735 308988
rect 31049 308938 32049 309066
rect 33672 309007 34272 309063
rect 31049 308762 32049 308890
rect 33672 308831 34272 308959
rect 34427 308907 35027 309035
rect 30135 308684 30735 308740
rect 34427 308731 35027 308859
rect 37998 308825 38148 308837
rect 38317 308825 38467 308837
rect 37998 308712 38598 308762
rect 33672 308655 34272 308711
rect 30135 308508 30735 308636
rect 31049 308592 32049 308642
rect 34427 308555 35027 308683
rect 37998 308536 38598 308592
rect 31049 308476 32049 308526
rect 33672 308479 34272 308535
rect 30135 308332 30735 308388
rect 31049 308320 32049 308448
rect 34427 308379 35027 308435
rect 37998 308366 38598 308416
rect 33672 308303 34272 308359
rect 36785 308342 36797 308346
rect 36785 308331 36800 308342
rect 36970 308331 36985 308346
rect 30135 308156 30735 308284
rect 31049 308164 32049 308292
rect 30135 307980 30735 308036
rect 31049 308008 32049 308136
rect 33672 308127 34272 308255
rect 34427 308203 35027 308331
rect 36785 308151 36985 308331
rect 36785 308140 36800 308151
rect 36785 308136 36797 308140
rect 36970 308136 36985 308151
rect 37083 308331 37098 308346
rect 37083 308151 37120 308331
rect 37083 308136 37098 308151
rect 36785 308106 36797 308110
rect 36785 308095 36800 308106
rect 36970 308095 36985 308110
rect 34427 308033 35027 308083
rect 33672 307957 34272 308007
rect 30135 307804 30735 307932
rect 36785 307915 36985 308095
rect 37993 307940 38593 307990
rect 31049 307852 32049 307908
rect 36785 307904 36800 307915
rect 36785 307900 36797 307904
rect 36970 307900 36985 307915
rect 31049 307696 32049 307824
rect 37993 307770 38593 307820
rect 30135 307634 30735 307684
rect 31049 307540 32049 307668
rect 36785 307594 37385 307644
rect 28396 307361 28449 307445
rect 31049 307384 32049 307512
rect 36785 307418 37385 307474
rect 28396 306903 28446 307361
rect 31049 307234 32049 307284
rect 36785 307242 37385 307298
rect 36785 307072 37385 307122
rect 37939 307039 37963 307063
rect 38085 307039 38109 307063
rect 29925 307003 29931 307032
rect 30271 307003 30305 307027
rect 30342 307003 30376 307027
rect 30413 307003 30447 307027
rect 30484 307003 30518 307027
rect 30555 307003 30589 307027
rect 30626 307003 30660 307027
rect 30697 307003 30731 307027
rect 37963 307015 37987 307038
rect 38061 307015 38085 307038
rect 29931 306962 29939 306986
rect 29955 306962 29961 307003
rect 29891 306938 29915 306962
rect 25101 306860 25121 306894
rect 25125 306860 25143 306894
rect 37759 306867 37783 306891
rect 25101 306826 25147 306860
rect 37792 306843 37807 306867
rect 25101 306792 25121 306826
rect 25125 306792 25143 306826
rect 21383 306758 21419 306792
rect 25101 306758 25147 306792
rect 21383 306724 21403 306758
rect 21407 306724 21415 306758
rect 25101 306724 25121 306758
rect 25125 306724 25143 306758
rect 21383 306690 21419 306724
rect 21383 306656 21403 306690
rect 21407 306656 21415 306690
rect 21481 306656 22881 306699
rect 22892 306675 22920 306703
rect 23617 306656 25017 306699
rect 25101 306690 25147 306724
rect 31458 306703 31608 306715
rect 31777 306703 31927 306715
rect 25101 306656 25121 306690
rect 25125 306656 25143 306690
rect 7389 306628 8389 306632
rect 8990 306628 9990 306632
rect 7353 306578 8425 306614
rect 7353 306537 7389 306578
rect 8389 306537 8425 306578
rect 7353 306501 8425 306537
rect 8954 306578 10026 306614
rect 15678 306582 16678 306654
rect 17278 306582 18278 306654
rect 21383 306622 21419 306656
rect 25101 306622 25147 306656
rect 21383 306588 21403 306622
rect 21407 306588 21415 306622
rect 25101 306588 25121 306622
rect 25125 306588 25143 306622
rect 8954 306537 8990 306578
rect 9990 306537 10026 306578
rect 15748 306571 15782 306582
rect 15816 306571 15850 306582
rect 15884 306571 15918 306582
rect 15952 306571 15986 306582
rect 16020 306571 16054 306582
rect 16088 306571 16122 306582
rect 16156 306571 16190 306582
rect 16224 306571 16258 306582
rect 16292 306571 16326 306582
rect 16360 306571 16394 306582
rect 16428 306571 16462 306582
rect 16496 306571 16530 306582
rect 16564 306571 16598 306582
rect 16632 306571 16666 306582
rect 17290 306571 17324 306582
rect 17358 306571 17392 306582
rect 17426 306571 17460 306582
rect 17494 306571 17528 306582
rect 17562 306571 17596 306582
rect 17630 306571 17664 306582
rect 17698 306571 17732 306582
rect 17766 306571 17800 306582
rect 17834 306571 17868 306582
rect 17902 306571 17936 306582
rect 17970 306571 18004 306582
rect 18038 306571 18072 306582
rect 18106 306571 18140 306582
rect 18174 306571 18208 306582
rect 15748 306561 15806 306571
rect 15816 306561 15874 306571
rect 15884 306561 15942 306571
rect 15952 306561 16010 306571
rect 16020 306561 16078 306571
rect 16088 306561 16146 306571
rect 16156 306561 16214 306571
rect 16224 306561 16282 306571
rect 16292 306561 16350 306571
rect 16360 306561 16418 306571
rect 16428 306561 16486 306571
rect 16496 306561 16554 306571
rect 16564 306561 16622 306571
rect 16632 306561 16690 306571
rect 17290 306561 17348 306571
rect 17358 306561 17416 306571
rect 17426 306561 17484 306571
rect 17494 306561 17552 306571
rect 17562 306561 17620 306571
rect 17630 306561 17688 306571
rect 17698 306561 17756 306571
rect 17766 306561 17824 306571
rect 17834 306561 17892 306571
rect 17902 306561 17960 306571
rect 17970 306561 18028 306571
rect 18038 306561 18096 306571
rect 18106 306561 18164 306571
rect 18174 306561 18232 306571
rect 15724 306537 16690 306561
rect 17266 306537 18232 306561
rect 21383 306554 21419 306588
rect 8954 306501 10026 306537
rect 15748 306522 15772 306537
rect 15816 306522 15840 306537
rect 15884 306522 15908 306537
rect 15952 306522 15976 306537
rect 16020 306522 16044 306537
rect 16088 306522 16112 306537
rect 16156 306522 16180 306537
rect 16224 306522 16248 306537
rect 16292 306522 16316 306537
rect 16360 306522 16384 306537
rect 16428 306522 16452 306537
rect 16496 306522 16520 306537
rect 16564 306522 16588 306537
rect 16632 306522 16656 306537
rect 17290 306522 17314 306537
rect 17358 306522 17382 306537
rect 17426 306522 17450 306537
rect 17494 306522 17518 306537
rect 17562 306522 17586 306537
rect 17630 306522 17654 306537
rect 17698 306522 17722 306537
rect 17766 306522 17790 306537
rect 17834 306522 17858 306537
rect 17902 306522 17926 306537
rect 17970 306522 17994 306537
rect 18038 306522 18062 306537
rect 18106 306522 18130 306537
rect 18174 306522 18198 306537
rect 15678 306367 16678 306522
rect 7389 306277 8389 306337
rect 8990 306277 9990 306337
rect 15678 306333 16690 306367
rect 17278 306357 18278 306522
rect 17266 306333 18278 306357
rect 15678 306322 16678 306333
rect 17278 306322 18278 306333
rect 21383 306520 21403 306554
rect 21407 306520 21415 306554
rect 21481 306520 22881 306563
rect 23617 306520 25017 306563
rect 25101 306554 25147 306588
rect 25414 306573 25438 306607
rect 31458 306590 32058 306640
rect 25101 306520 25121 306554
rect 25125 306520 25143 306554
rect 21383 306486 21419 306520
rect 25101 306486 25147 306520
rect 21383 306452 21403 306486
rect 21407 306452 21415 306486
rect 21383 306418 21419 306452
rect 21383 306384 21403 306418
rect 21407 306384 21415 306418
rect 21383 306350 21419 306384
rect 21481 306357 22881 306485
rect 23617 306357 25017 306485
rect 25101 306452 25121 306486
rect 25125 306452 25143 306486
rect 37792 306470 37807 306494
rect 25101 306418 25147 306452
rect 25101 306384 25121 306418
rect 25125 306384 25143 306418
rect 31458 306414 32058 306470
rect 37759 306446 37783 306470
rect 25101 306350 25147 306384
rect 15748 306309 15772 306322
rect 15816 306309 15840 306322
rect 15884 306309 15908 306322
rect 15952 306309 15976 306322
rect 16020 306309 16044 306322
rect 16088 306309 16112 306322
rect 16156 306309 16180 306322
rect 16224 306309 16248 306322
rect 16292 306309 16316 306322
rect 16360 306309 16384 306322
rect 16428 306309 16452 306322
rect 16496 306309 16520 306322
rect 16564 306309 16588 306322
rect 16632 306309 16656 306322
rect 17290 306309 17314 306322
rect 17358 306309 17382 306322
rect 17426 306309 17450 306322
rect 17494 306309 17518 306322
rect 17562 306309 17586 306322
rect 17630 306309 17654 306322
rect 17698 306309 17722 306322
rect 17766 306309 17790 306322
rect 17834 306309 17858 306322
rect 17902 306309 17926 306322
rect 17970 306309 17994 306322
rect 18038 306309 18062 306322
rect 18106 306309 18130 306322
rect 18174 306309 18198 306322
rect 21383 306316 21403 306350
rect 21407 306316 21415 306350
rect 21383 306282 21419 306316
rect 21383 306248 21403 306282
rect 21407 306248 21415 306282
rect 21383 306214 21419 306248
rect 21383 306180 21403 306214
rect 21407 306180 21415 306214
rect 21481 306194 22881 306322
rect 23617 306194 25017 306322
rect 25101 306316 25121 306350
rect 25125 306316 25143 306350
rect 25101 306282 25147 306316
rect 25101 306248 25121 306282
rect 25125 306248 25143 306282
rect 25101 306214 25147 306248
rect 25101 306180 25121 306214
rect 25125 306180 25143 306214
rect 25725 306197 26325 306247
rect 31458 306244 32058 306294
rect 30245 306220 30257 306224
rect 30245 306209 30260 306220
rect 30430 306209 30445 306224
rect 21383 306146 21419 306180
rect 7389 306066 8389 306070
rect 8990 306066 9990 306070
rect 15678 306061 16678 306133
rect 17278 306061 18278 306133
rect 21383 306112 21403 306146
rect 21407 306112 21415 306146
rect 21383 306078 21419 306112
rect 7353 306016 8425 306052
rect 7353 305975 7389 306016
rect 8389 305975 8425 306016
rect 7353 305919 8425 305975
rect 7353 305903 7389 305919
rect 8389 305903 8425 305919
rect 7353 305847 8425 305903
rect 7353 305810 7389 305847
rect 8389 305810 8425 305847
rect 7353 305770 8425 305810
rect 8954 306016 10026 306052
rect 8954 305975 8990 306016
rect 9990 305975 10026 306016
rect 8954 305919 10026 305975
rect 21383 306044 21403 306078
rect 21407 306044 21415 306078
rect 21383 306010 21419 306044
rect 21481 306031 22881 306159
rect 23617 306031 25017 306159
rect 25101 306146 25147 306180
rect 25101 306112 25121 306146
rect 25125 306112 25143 306146
rect 25101 306078 25147 306112
rect 25101 306044 25121 306078
rect 25125 306044 25143 306078
rect 25725 306047 26325 306097
rect 25101 306010 25147 306044
rect 21383 305976 21403 306010
rect 21407 305976 21415 306010
rect 21383 305942 21419 305976
rect 8954 305903 8990 305919
rect 9990 305903 10026 305919
rect 15678 305906 16678 305923
rect 17278 305906 18278 305923
rect 21383 305908 21403 305942
rect 21407 305908 21415 305942
rect 8954 305847 10026 305903
rect 20250 305890 20316 305906
rect 8954 305810 8990 305847
rect 9990 305810 10026 305847
rect 8954 305770 10026 305810
rect 21383 305874 21419 305908
rect 21383 305840 21403 305874
rect 21407 305840 21415 305874
rect 21481 305868 22881 305996
rect 23617 305868 25017 305996
rect 25101 305976 25121 306010
rect 25125 305976 25143 306010
rect 25101 305942 25147 305976
rect 25101 305908 25121 305942
rect 25125 305908 25143 305942
rect 25725 305925 26325 305975
rect 25101 305874 25147 305908
rect 25101 305840 25121 305874
rect 25125 305840 25143 305874
rect 21383 305806 21419 305840
rect 21383 305772 21403 305806
rect 21407 305772 21415 305806
rect 21383 305738 21419 305772
rect 15678 305703 16678 305736
rect 17278 305703 18278 305736
rect 21383 305704 21403 305738
rect 21407 305704 21415 305738
rect 21481 305705 22881 305833
rect 23617 305705 25017 305833
rect 25101 305806 25147 305840
rect 25101 305772 25121 305806
rect 25125 305772 25143 305806
rect 25725 305775 26325 305825
rect 25101 305738 25147 305772
rect 25101 305704 25121 305738
rect 25125 305704 25143 305738
rect 21383 305670 21419 305704
rect 25101 305670 25147 305704
rect 21383 305636 21403 305670
rect 21407 305636 21415 305670
rect 7389 305559 8389 305631
rect 8990 305559 9990 305631
rect 21383 305602 21419 305636
rect 15840 305510 15870 305580
rect 15878 305546 15908 305580
rect 21383 305568 21403 305602
rect 21407 305568 21415 305602
rect 15853 305508 15870 305510
rect 21383 305534 21419 305568
rect 21481 305542 22881 305670
rect 23617 305542 25017 305670
rect 25101 305636 25121 305670
rect 25125 305636 25143 305670
rect 25725 305649 26325 305699
rect 25101 305602 25147 305636
rect 25101 305568 25121 305602
rect 25125 305568 25143 305602
rect 25101 305534 25147 305568
rect 5981 305483 6021 305493
rect 5137 305469 6021 305483
rect 21383 305500 21403 305534
rect 21407 305500 21415 305534
rect 21383 305466 21419 305500
rect 7389 305369 8389 305463
rect 7389 305359 8413 305369
rect 8990 305359 9990 305463
rect 21383 305432 21403 305466
rect 21407 305432 21415 305466
rect 21383 305398 21419 305432
rect 21383 305364 21403 305398
rect 21407 305364 21415 305398
rect 21481 305379 22881 305507
rect 23617 305379 25017 305507
rect 25101 305500 25121 305534
rect 25125 305500 25143 305534
rect 25101 305466 25147 305500
rect 25725 305499 26325 305549
rect 25101 305432 25121 305466
rect 25125 305432 25143 305466
rect 25101 305398 25147 305432
rect 25101 305364 25121 305398
rect 25125 305364 25143 305398
rect 25725 305377 26325 305427
rect 21383 305330 21419 305364
rect 25101 305330 25147 305364
rect 21383 305296 21403 305330
rect 21407 305296 21415 305330
rect 25101 305296 25121 305330
rect 25125 305296 25143 305330
rect 21383 305262 21419 305296
rect 21383 305228 21403 305262
rect 21407 305228 21415 305262
rect 21481 305229 22881 305272
rect 23617 305229 25017 305272
rect 25101 305262 25147 305296
rect 25101 305228 25121 305262
rect 25125 305228 25143 305262
rect 21383 305194 21419 305228
rect 25101 305194 25147 305228
rect 25725 305227 26325 305277
rect 21383 305160 21403 305194
rect 21407 305160 21415 305194
rect 25101 305160 25121 305194
rect 25125 305160 25143 305194
rect 27162 305170 27212 306170
rect 27312 305170 27440 306170
rect 27468 305170 27596 306170
rect 27624 305170 27752 306170
rect 27780 305170 27908 306170
rect 27936 305170 28064 306170
rect 28092 305170 28220 306170
rect 28248 305170 28376 306170
rect 28404 305170 28532 306170
rect 28560 305170 28688 306170
rect 28716 305170 28844 306170
rect 28872 305170 29000 306170
rect 29028 305170 29156 306170
rect 29184 305170 29312 306170
rect 29340 305170 29390 306170
rect 30245 306029 30445 306209
rect 30245 306018 30260 306029
rect 30245 306014 30257 306018
rect 30430 306014 30445 306029
rect 30543 306209 30558 306224
rect 30543 306029 30580 306209
rect 30543 306014 30558 306029
rect 30245 305984 30257 305988
rect 30245 305973 30260 305984
rect 30430 305973 30445 305988
rect 30245 305793 30445 305973
rect 31453 305818 32053 305868
rect 30245 305782 30260 305793
rect 30245 305778 30257 305782
rect 30430 305778 30445 305793
rect 31453 305648 32053 305698
rect 30245 305472 30845 305522
rect 30245 305296 30845 305352
rect 21383 305126 21419 305160
rect 25101 305126 25147 305160
rect 21383 305102 21403 305126
rect 21385 305048 21403 305102
rect 21407 305082 21415 305126
rect 25101 305102 25121 305126
rect 25113 305082 25121 305102
rect 25125 305048 25143 305126
rect 30245 305120 30845 305176
rect 30245 304950 30845 305000
rect 21000 304800 21003 304920
rect 21352 304885 21376 304909
rect 25122 304885 25146 304909
rect 21385 304861 21400 304885
rect 25098 304861 25113 304885
rect 21274 304783 21294 304851
rect 21410 304817 21430 304851
rect 25068 304817 25088 304851
rect 25204 304817 25224 304851
rect 21385 304807 21430 304817
rect 25102 304807 25137 304817
rect 21361 304783 21430 304807
rect 25089 304783 25137 304807
rect 25238 304783 25258 304817
rect 680480 298427 680517 298520
rect 680615 298427 680815 298520
rect 685793 298483 685993 298520
rect 686053 298483 686253 298520
rect 686607 298440 687607 298490
rect 692427 298392 693027 298448
rect 679007 298216 679607 298266
rect 680615 298191 680815 298371
rect 686829 298301 687429 298351
rect 684004 298243 685004 298293
rect 695201 298282 695251 298520
rect 696287 298282 696337 298520
rect 682890 298161 683490 298211
rect 684004 298127 685004 298177
rect 686829 298125 687429 298181
rect 679007 298046 679607 298096
rect 684004 297971 685004 298027
rect 686829 297955 687429 298005
rect 680215 297870 680815 297920
rect 681713 297881 682313 297931
rect 682921 297899 683521 297949
rect 692427 297930 693027 297980
rect 684004 297821 685004 297871
rect 680215 297694 680815 297750
rect 681713 297705 682313 297761
rect 682921 297743 683521 297799
rect 685537 297749 686137 297799
rect 697088 297749 697138 298520
rect 697706 297749 697756 298520
rect 699322 298374 700322 298514
rect 700922 298374 701922 298514
rect 707610 298098 708610 298099
rect 699322 297956 700322 298012
rect 700922 297956 701922 298012
rect 707610 298001 708610 298057
rect 709211 298001 710211 298057
rect 707610 297959 708610 297960
rect 699322 297884 700322 297940
rect 700922 297884 701922 297940
rect 709211 297936 710211 297960
rect 682921 297593 683521 297643
rect 684070 297599 684670 297649
rect 685537 297593 686137 297649
rect 699322 297623 700322 297673
rect 700922 297623 701922 297673
rect 680215 297518 680815 297574
rect 707610 297523 708610 297617
rect 709211 297523 710211 297591
rect 707610 297513 707624 297523
rect 707658 297513 707695 297523
rect 707729 297513 707769 297523
rect 707803 297513 707840 297523
rect 707874 297513 707914 297523
rect 707948 297513 707985 297523
rect 708019 297513 708059 297523
rect 708093 297513 708130 297523
rect 708164 297513 708204 297523
rect 708238 297513 708275 297523
rect 708309 297513 708369 297523
rect 708403 297513 708446 297523
rect 708480 297513 708522 297523
rect 708556 297513 708604 297523
rect 709219 297513 709270 297523
rect 709304 297513 709364 297523
rect 709398 297513 709435 297523
rect 709469 297513 709509 297523
rect 709543 297513 709580 297523
rect 709614 297513 709654 297523
rect 709688 297513 709725 297523
rect 709759 297513 709799 297523
rect 709833 297513 709870 297523
rect 709904 297513 709944 297523
rect 709978 297513 710015 297523
rect 710049 297513 710089 297523
rect 710123 297513 710160 297523
rect 710194 297513 710211 297523
rect 684070 297443 684670 297499
rect 685537 297443 686137 297493
rect 692428 297442 693028 297492
rect 680215 297348 680815 297398
rect 681713 297359 682313 297409
rect 684070 297293 684670 297343
rect 692428 297292 693028 297342
rect 705107 297336 705173 297352
rect 711579 297301 711595 298520
rect 711892 297697 711942 298520
rect 712062 297697 712112 298520
rect 716071 298357 716074 298358
rect 714645 298323 714752 298357
rect 716071 298356 716072 298357
rect 716073 298356 716074 298357
rect 716071 298355 716074 298356
rect 716208 298357 716211 298358
rect 716208 298356 716209 298357
rect 716210 298356 716211 298357
rect 716208 298355 716211 298356
rect 714964 298247 715998 298329
rect 716284 298247 717318 298329
rect 714175 297398 714225 297998
rect 714425 297398 714475 297998
rect 680215 297232 680815 297282
rect 698017 297232 698053 297260
rect 692428 297162 693028 297212
rect 698030 297198 698077 297232
rect 698017 297164 698053 297198
rect 680215 297056 680815 297112
rect 692428 297006 693028 297134
rect 698030 297130 698077 297164
rect 698017 297096 698053 297130
rect 698030 297062 698077 297096
rect 698017 296983 698053 297062
rect 698084 296983 698120 297260
rect 714781 297191 714863 298226
rect 715134 297955 715828 298037
rect 714686 297123 714863 297191
rect 714645 297089 714863 297123
rect 680215 296880 680815 296936
rect 686719 296893 686739 296917
rect 686743 296893 686753 296917
rect 686719 296859 686757 296893
rect 686719 296822 686739 296859
rect 686743 296822 686753 296859
rect 692428 296850 693028 296978
rect 698017 296947 698210 296983
rect 698084 296935 698210 296947
rect 702756 296959 703645 296983
rect 702756 296935 702853 296959
rect 698084 296828 702853 296935
rect 686719 296788 686757 296822
rect 680215 296704 680815 296760
rect 686719 296751 686739 296788
rect 686743 296751 686753 296788
rect 686719 296741 686757 296751
rect 686699 296717 686767 296741
rect 686719 296704 686739 296717
rect 686743 296704 686753 296717
rect 686719 296695 686753 296704
rect 686719 296693 686743 296695
rect 692428 296694 693028 296750
rect 686685 296656 686709 296680
rect 686743 296656 686767 296680
rect 678799 296503 679399 296553
rect 680215 296534 680815 296584
rect 692428 296538 693028 296666
rect 680593 296531 680815 296534
rect 682009 296501 682069 296516
rect 682024 296465 682054 296501
rect 683708 296387 684308 296437
rect 678799 296327 679399 296383
rect 692428 296382 693028 296510
rect 714781 296308 714863 297089
rect 715063 296609 715145 297915
rect 715289 296777 715339 297719
rect 715633 296777 715683 297719
rect 715382 296672 715422 296756
rect 715542 296672 715582 296756
rect 715342 296632 715382 296672
rect 715582 296632 715622 296672
rect 715815 296609 715897 297915
rect 715134 296387 715828 296469
rect 716100 296308 716182 298226
rect 716454 297955 717148 298037
rect 716385 296609 716467 297915
rect 716599 296777 716649 297719
rect 716943 296777 716993 297719
rect 716700 296672 716740 296756
rect 716860 296672 716900 296756
rect 716660 296632 716700 296672
rect 716900 296632 716940 296672
rect 717137 296609 717219 297915
rect 716454 296387 717148 296469
rect 717419 296308 717501 298226
rect 683708 296237 684308 296287
rect 692428 296232 693028 296282
rect 678799 296157 679399 296207
rect 684565 296160 684790 296168
rect 696597 296000 696600 296120
rect 714964 296095 715998 296177
rect 716284 296095 717318 296177
rect 21000 273000 21003 273120
rect 282 272623 1316 272705
rect 1602 272623 2636 272705
rect 32810 272662 33035 272670
rect 38201 272593 38801 272643
rect 24572 272518 25172 272568
rect 33292 272513 33892 272563
rect 99 270574 181 272492
rect 452 272331 1146 272413
rect 381 270885 463 272191
rect 660 272128 700 272168
rect 900 272128 940 272168
rect 700 272044 740 272128
rect 860 272044 900 272128
rect 607 271081 657 272023
rect 951 271081 1001 272023
rect 1133 270885 1215 272191
rect 452 270763 1146 270845
rect 1418 270574 1500 272492
rect 1772 272331 2466 272413
rect 1703 270885 1785 272191
rect 1978 272128 2018 272168
rect 2218 272128 2258 272168
rect 2018 272044 2058 272128
rect 2178 272044 2218 272128
rect 1917 271081 1967 272023
rect 2261 271081 2311 272023
rect 2455 270885 2537 272191
rect 2737 271779 2819 272492
rect 24572 272362 25172 272490
rect 38201 272417 38801 272473
rect 33292 272363 33892 272413
rect 24572 272206 25172 272334
rect 35546 272299 35576 272335
rect 36785 272329 36935 272341
rect 35531 272284 35591 272299
rect 36785 272216 37385 272266
rect 38201 272247 38801 272297
rect 30833 272120 30857 272144
rect 30891 272120 30915 272144
rect 24572 272050 25172 272106
rect 30857 272105 30881 272107
rect 30857 272096 30887 272105
rect 30867 272083 30887 272096
rect 30891 272083 30907 272120
rect 30833 272059 30857 272083
rect 30867 272049 30911 272083
rect 14747 271865 19516 271972
rect 24572 271894 25172 272022
rect 30867 272012 30887 272049
rect 30891 272012 30907 272049
rect 36785 272040 37385 272096
rect 30867 271978 30911 272012
rect 30867 271941 30887 271978
rect 30891 271941 30907 271978
rect 30867 271907 30911 271941
rect 30867 271883 30887 271907
rect 30891 271883 30907 271907
rect 14747 271841 14844 271865
rect 13955 271817 14844 271841
rect 19390 271853 19516 271865
rect 19390 271841 19583 271853
rect 19390 271817 19605 271841
rect 19639 271817 19673 271841
rect 19707 271817 19741 271841
rect 19775 271817 19809 271841
rect 19843 271817 19877 271841
rect 19911 271817 19945 271841
rect 19979 271817 20013 271841
rect 20047 271817 20081 271841
rect 20115 271817 20149 271841
rect 20183 271817 20217 271841
rect 20251 271817 20285 271841
rect 20319 271817 20353 271841
rect 20387 271817 20421 271841
rect 20455 271817 20489 271841
rect 20523 271817 20557 271841
rect 20591 271817 20625 271841
rect 20659 271817 20693 271841
rect 2737 271711 2914 271779
rect 1772 270763 2466 270845
rect 2737 270574 2819 271711
rect 2848 271677 2955 271711
rect 19480 271540 19516 271817
rect 19547 271540 19583 271817
rect 24572 271738 25172 271866
rect 36785 271864 37385 271920
rect 36785 271688 37385 271744
rect 20809 271650 20833 271684
rect 20809 271582 20833 271616
rect 24572 271588 25172 271638
rect 20809 271540 20833 271548
rect 36785 271518 37385 271568
rect 3125 270802 3175 271402
rect 3375 270802 3425 271402
rect 282 270471 1316 270553
rect 1602 270471 2636 270553
rect 1389 270444 1392 270445
rect 1389 270443 1390 270444
rect 1391 270443 1392 270444
rect 1389 270442 1392 270443
rect 1526 270444 1529 270445
rect 1526 270443 1527 270444
rect 1528 270443 1529 270444
rect 2848 270443 2955 270477
rect 1526 270442 1529 270443
rect 5488 270280 5538 271103
rect 5658 270280 5708 271103
rect 6005 270280 6021 271499
rect 12427 271448 12493 271464
rect 24572 271458 25172 271508
rect 32930 271457 33530 271507
rect 35287 271391 35887 271441
rect 36785 271402 37385 271452
rect 24572 271308 25172 271358
rect 31463 271307 32063 271357
rect 32930 271301 33530 271357
rect 7389 271277 7406 271287
rect 7440 271277 7477 271287
rect 7511 271277 7551 271287
rect 7585 271277 7622 271287
rect 7656 271277 7696 271287
rect 7730 271277 7767 271287
rect 7801 271277 7841 271287
rect 7875 271277 7912 271287
rect 7946 271277 7986 271287
rect 8020 271277 8057 271287
rect 8091 271277 8131 271287
rect 8165 271277 8202 271287
rect 8236 271277 8296 271287
rect 8330 271277 8381 271287
rect 8996 271277 9044 271287
rect 9078 271277 9120 271287
rect 9154 271277 9197 271287
rect 9231 271277 9291 271287
rect 9325 271277 9362 271287
rect 9396 271277 9436 271287
rect 9470 271277 9507 271287
rect 9541 271277 9581 271287
rect 9615 271277 9652 271287
rect 9686 271277 9726 271287
rect 9760 271277 9797 271287
rect 9831 271277 9871 271287
rect 9905 271277 9942 271287
rect 9976 271277 9990 271287
rect 7389 271209 8389 271277
rect 8990 271183 9990 271277
rect 36785 271226 37385 271282
rect 15678 271127 16678 271177
rect 17278 271127 18278 271177
rect 31463 271151 32063 271207
rect 32930 271151 33530 271201
rect 34079 271157 34679 271207
rect 7389 270840 8389 270864
rect 15678 270860 16678 270916
rect 17278 270860 18278 270916
rect 8990 270840 9990 270841
rect 7389 270743 8389 270799
rect 8990 270743 9990 270799
rect 15678 270788 16678 270844
rect 17278 270788 18278 270844
rect 8990 270701 9990 270702
rect 15678 270286 16678 270426
rect 17278 270286 18278 270426
rect 19844 270280 19894 271051
rect 20462 270280 20512 271051
rect 31463 271001 32063 271051
rect 34079 271001 34679 271057
rect 35287 271039 35887 271095
rect 36785 271050 37385 271106
rect 32596 270929 33596 270979
rect 24573 270820 25173 270870
rect 34079 270851 34679 270901
rect 35287 270869 35887 270919
rect 36785 270880 37385 270930
rect 30171 270795 30771 270845
rect 32596 270773 33596 270829
rect 37993 270704 38593 270754
rect 30171 270619 30771 270675
rect 32596 270623 33596 270673
rect 34110 270589 34710 270639
rect 21263 270280 21313 270518
rect 22349 270280 22399 270518
rect 32596 270507 33596 270557
rect 30171 270449 30771 270499
rect 36785 270429 36985 270609
rect 37993 270534 38593 270584
rect 24573 270352 25173 270408
rect 29993 270310 30993 270360
rect 31347 270280 31547 270317
rect 31607 270280 31807 270317
rect 36785 270280 36985 270373
rect 37083 270280 37120 270373
rect 696597 264200 696600 264320
rect 692376 263983 692396 264017
rect 692463 263993 692532 264017
rect 696191 263993 696239 264017
rect 692487 263983 692532 263993
rect 696204 263983 696239 263993
rect 696340 263983 696360 264017
rect 692487 263915 692502 263939
rect 696200 263915 696215 263939
rect 692454 263891 692478 263915
rect 696224 263891 696248 263915
rect 686755 263800 687355 263850
rect 692487 263748 692505 263752
rect 692479 263718 692505 263748
rect 692487 263698 692505 263718
rect 686755 263624 687355 263680
rect 692485 263674 692505 263698
rect 692509 263674 692517 263718
rect 696215 263698 696223 263748
rect 696203 263674 696223 263698
rect 696227 263674 696245 263752
rect 692485 263640 692521 263674
rect 696203 263640 696249 263674
rect 686755 263448 687355 263504
rect 686755 263278 687355 263328
rect 685547 263102 686147 263152
rect 687155 263007 687170 263022
rect 687343 263018 687355 263022
rect 687340 263007 687355 263018
rect 685547 262932 686147 262982
rect 687155 262827 687355 263007
rect 687155 262812 687170 262827
rect 687340 262816 687355 262827
rect 687343 262812 687355 262816
rect 687042 262771 687057 262786
rect 687020 262591 687057 262771
rect 687155 262771 687170 262786
rect 687343 262782 687355 262786
rect 687340 262771 687355 262782
rect 687155 262591 687355 262771
rect 688210 262630 688260 263630
rect 688360 262740 688488 263630
rect 688516 262740 688644 263630
rect 688672 262740 688800 263630
rect 688828 262740 688956 263630
rect 688984 262740 689112 263630
rect 689140 262740 689268 263630
rect 689296 262740 689424 263630
rect 689452 262740 689580 263630
rect 689608 262740 689736 263630
rect 689764 262740 689892 263630
rect 689920 262740 690048 263630
rect 690076 262740 690204 263630
rect 690232 262740 690360 263630
rect 690388 262630 690438 263630
rect 692485 263606 692505 263640
rect 692509 263606 692517 263640
rect 696203 263606 696223 263640
rect 696227 263606 696245 263640
rect 691275 263523 691875 263573
rect 692485 263572 692521 263606
rect 696203 263572 696249 263606
rect 692485 263538 692505 263572
rect 692509 263538 692517 263572
rect 692485 263504 692521 263538
rect 692583 263528 693983 263571
rect 694719 263528 696119 263571
rect 696203 263538 696223 263572
rect 696227 263538 696245 263572
rect 696203 263504 696249 263538
rect 692485 263470 692505 263504
rect 692509 263470 692517 263504
rect 692485 263436 692521 263470
rect 691275 263373 691875 263423
rect 692485 263402 692505 263436
rect 692509 263402 692517 263436
rect 692485 263368 692521 263402
rect 692485 263334 692505 263368
rect 692509 263334 692517 263368
rect 692583 263365 693983 263493
rect 694719 263365 696119 263493
rect 696203 263470 696223 263504
rect 696227 263470 696245 263504
rect 696203 263436 696249 263470
rect 707624 263441 707658 263475
rect 707695 263441 707729 263475
rect 707769 263441 707803 263475
rect 707840 263441 707874 263475
rect 707914 263441 707948 263475
rect 707985 263441 708019 263475
rect 708059 263441 708093 263475
rect 708130 263441 708164 263475
rect 708204 263441 708238 263475
rect 708275 263441 708309 263475
rect 708369 263441 708403 263475
rect 708446 263441 708480 263475
rect 708520 263441 708554 263465
rect 708588 263441 708610 263465
rect 709211 263441 709234 263465
rect 709270 263441 709304 263475
rect 709364 263441 709398 263475
rect 709435 263441 709469 263475
rect 709509 263441 709543 263475
rect 709580 263441 709614 263475
rect 709654 263441 709688 263475
rect 709725 263441 709759 263475
rect 709799 263441 709833 263475
rect 709870 263441 709904 263475
rect 709944 263441 709978 263475
rect 710015 263441 710049 263475
rect 710089 263441 710123 263475
rect 710160 263441 710194 263475
rect 696203 263402 696223 263436
rect 696227 263402 696245 263436
rect 707610 263431 707624 263441
rect 707658 263431 707695 263441
rect 707729 263431 707769 263441
rect 707803 263431 707840 263441
rect 707874 263431 707914 263441
rect 707948 263431 707985 263441
rect 708019 263431 708059 263441
rect 708093 263431 708130 263441
rect 708164 263431 708204 263441
rect 708238 263431 708275 263441
rect 708309 263431 708369 263441
rect 708403 263431 708446 263441
rect 708480 263431 708520 263441
rect 708554 263431 708588 263441
rect 708610 263431 708634 263441
rect 709211 263431 709270 263441
rect 709304 263431 709364 263441
rect 709398 263431 709435 263441
rect 709469 263431 709509 263441
rect 709543 263431 709580 263441
rect 709614 263431 709654 263441
rect 709688 263431 709725 263441
rect 709759 263431 709799 263441
rect 709833 263431 709870 263441
rect 709904 263431 709944 263441
rect 709978 263431 710015 263441
rect 710049 263431 710089 263441
rect 710123 263431 710160 263441
rect 710194 263431 710211 263441
rect 696203 263368 696249 263402
rect 696203 263334 696223 263368
rect 696227 263334 696245 263368
rect 707610 263337 708610 263431
rect 709211 263337 710211 263431
rect 691275 263251 691875 263301
rect 692485 263300 692521 263334
rect 692485 263266 692505 263300
rect 692509 263266 692517 263300
rect 692485 263232 692521 263266
rect 692485 263198 692505 263232
rect 692509 263198 692517 263232
rect 692583 263202 693983 263330
rect 694719 263202 696119 263330
rect 696203 263300 696249 263334
rect 711579 263317 712463 263331
rect 711579 263307 711619 263317
rect 696203 263266 696223 263300
rect 696227 263266 696245 263300
rect 701730 263290 701747 263292
rect 696203 263232 696249 263266
rect 696203 263198 696223 263232
rect 696227 263198 696245 263232
rect 701692 263220 701722 263254
rect 701730 263220 701760 263290
rect 707610 263241 708610 263301
rect 709211 263241 710211 263301
rect 692485 263164 692521 263198
rect 691275 263101 691875 263151
rect 692485 263130 692505 263164
rect 692509 263130 692517 263164
rect 692485 263096 692521 263130
rect 692485 263062 692505 263096
rect 692509 263062 692517 263096
rect 692485 263028 692521 263062
rect 692583 263039 693983 263167
rect 694719 263039 696119 263167
rect 696203 263164 696249 263198
rect 696203 263130 696223 263164
rect 696227 263130 696245 263164
rect 696203 263096 696249 263130
rect 696203 263062 696223 263096
rect 696227 263062 696245 263096
rect 699322 263064 700322 263097
rect 700922 263064 701922 263097
rect 696203 263028 696249 263062
rect 707610 263044 708610 263048
rect 709211 263044 710211 263048
rect 691275 262975 691875 263025
rect 692485 262994 692505 263028
rect 692509 262994 692517 263028
rect 692485 262960 692521 262994
rect 692485 262926 692505 262960
rect 692509 262926 692517 262960
rect 692485 262892 692521 262926
rect 691275 262825 691875 262875
rect 692485 262858 692505 262892
rect 692509 262858 692517 262892
rect 692583 262876 693983 263004
rect 694719 262876 696119 263004
rect 696203 262994 696223 263028
rect 696227 262994 696245 263028
rect 707574 262994 708646 263030
rect 696203 262960 696249 262994
rect 696203 262926 696223 262960
rect 696227 262926 696245 262960
rect 707574 262953 707610 262994
rect 708610 262953 708646 262994
rect 696203 262892 696249 262926
rect 697284 262894 697350 262910
rect 707574 262897 708646 262953
rect 696203 262858 696223 262892
rect 696227 262858 696245 262892
rect 699322 262877 700322 262894
rect 700922 262877 701922 262894
rect 707574 262881 707610 262897
rect 708610 262881 708646 262897
rect 692485 262824 692521 262858
rect 692485 262790 692505 262824
rect 692509 262790 692517 262824
rect 692485 262756 692521 262790
rect 691275 262703 691875 262753
rect 692485 262740 692505 262756
rect 692509 262740 692517 262756
rect 692583 262740 693983 262841
rect 694719 262740 696119 262841
rect 696203 262824 696249 262858
rect 707574 262825 708646 262881
rect 696203 262790 696223 262824
rect 696227 262790 696245 262824
rect 696203 262756 696249 262790
rect 696203 262740 696223 262756
rect 696227 262740 696245 262756
rect 699322 262740 700322 262811
rect 700922 262740 701922 262811
rect 707574 262788 707610 262825
rect 708610 262788 708646 262825
rect 707574 262748 708646 262788
rect 709175 262994 710247 263030
rect 709175 262953 709211 262994
rect 710211 262953 710247 262994
rect 709175 262897 710247 262953
rect 709175 262881 709211 262897
rect 710211 262881 710247 262897
rect 709175 262825 710247 262881
rect 709175 262788 709211 262825
rect 710211 262788 710247 262825
rect 709175 262748 710247 262788
rect 685542 262506 686142 262556
rect 691275 262553 691875 262603
rect 685542 262330 686142 262386
rect 692583 262237 693983 262280
rect 694719 262237 696119 262280
rect 699322 262278 700322 262418
rect 700922 262278 701922 262418
rect 685542 262160 686142 262210
rect 692583 262101 693983 262144
rect 694719 262101 696119 262144
rect 680215 261678 680815 261728
rect 680215 261502 680815 261558
rect 685551 261516 686551 261566
rect 689154 261480 689204 261897
rect 689304 261480 689360 261897
rect 689460 261480 689516 261897
rect 689616 261480 689672 261897
rect 689772 261480 689828 261897
rect 689928 261480 689978 261897
rect 699322 261860 700322 261916
rect 700922 261860 701922 261916
rect 707610 261905 708610 261961
rect 709211 261905 710211 261961
rect 699322 261788 700322 261844
rect 700922 261788 701922 261844
rect 707610 261833 708610 261889
rect 709211 261833 710211 261889
rect 711579 261525 711605 263307
rect 715956 262297 716006 263297
rect 716106 262740 716234 263297
rect 716262 262297 716312 263297
rect 711579 261480 711595 261495
rect 712409 261480 712431 261485
rect 713640 261480 713641 261785
rect 713750 261772 714750 261822
rect 713750 261562 714750 261612
rect 713750 261480 714750 261496
rect 2850 259304 3850 259320
rect 2850 259188 3850 259238
rect 2850 258978 3850 259028
rect 3959 259015 3960 259320
rect 5169 259315 5191 259320
rect 6005 259305 6021 259320
rect 1288 257503 1338 258503
rect 1438 257503 1566 258060
rect 1594 257503 1644 258503
rect 5995 257493 6021 259275
rect 7389 258911 8389 258967
rect 8990 258911 9990 258967
rect 15678 258956 16678 259012
rect 17278 258956 18278 259012
rect 7389 258839 8389 258895
rect 8990 258839 9990 258895
rect 15678 258884 16678 258940
rect 17278 258884 18278 258940
rect 27622 258903 27672 259320
rect 27772 258903 27828 259320
rect 27928 258903 27984 259320
rect 28084 258903 28140 259320
rect 28240 258903 28296 259320
rect 28396 258903 28446 259320
rect 31049 259234 32049 259284
rect 36785 259242 37385 259298
rect 36785 259072 37385 259122
rect 21481 258656 22881 258699
rect 23617 258656 25017 258699
rect 31458 258590 32058 258640
rect 15678 258382 16678 258522
rect 17278 258382 18278 258522
rect 21481 258520 22881 258563
rect 23617 258520 25017 258563
rect 31458 258414 32058 258470
rect 25725 258197 26325 258247
rect 31458 258244 32058 258294
rect 7353 258016 8425 258052
rect 7353 257975 7389 258016
rect 8389 257975 8425 258016
rect 7353 257919 8425 257975
rect 7353 257903 7389 257919
rect 8389 257903 8425 257919
rect 7353 257847 8425 257903
rect 7353 257810 7389 257847
rect 8389 257810 8425 257847
rect 7353 257770 8425 257810
rect 8954 258016 10026 258052
rect 8954 257975 8990 258016
rect 9990 257975 10026 258016
rect 8954 257919 10026 257975
rect 21383 258044 21403 258060
rect 21407 258044 21415 258060
rect 21383 258010 21419 258044
rect 21481 258031 22881 258060
rect 23617 258031 25017 258060
rect 25101 258044 25121 258060
rect 25125 258044 25143 258060
rect 25725 258047 26325 258097
rect 25101 258010 25147 258044
rect 21383 257976 21403 258010
rect 21407 257976 21415 258010
rect 21383 257942 21419 257976
rect 8954 257903 8990 257919
rect 9990 257903 10026 257919
rect 15678 257906 16678 257923
rect 17278 257906 18278 257923
rect 21383 257908 21403 257942
rect 21407 257908 21415 257942
rect 8954 257847 10026 257903
rect 20250 257890 20316 257906
rect 8954 257810 8990 257847
rect 9990 257810 10026 257847
rect 8954 257770 10026 257810
rect 21383 257874 21419 257908
rect 21383 257840 21403 257874
rect 21407 257840 21415 257874
rect 21481 257868 22881 257996
rect 23617 257868 25017 257996
rect 25101 257976 25121 258010
rect 25125 257976 25143 258010
rect 25101 257942 25147 257976
rect 25101 257908 25121 257942
rect 25125 257908 25143 257942
rect 25725 257925 26325 257975
rect 25101 257874 25147 257908
rect 25101 257840 25121 257874
rect 25125 257840 25143 257874
rect 21383 257806 21419 257840
rect 21383 257772 21403 257806
rect 21407 257772 21415 257806
rect 21383 257738 21419 257772
rect 15678 257703 16678 257736
rect 17278 257703 18278 257736
rect 21383 257704 21403 257738
rect 21407 257704 21415 257738
rect 21481 257705 22881 257833
rect 23617 257705 25017 257833
rect 25101 257806 25147 257840
rect 25101 257772 25121 257806
rect 25125 257772 25143 257806
rect 25725 257775 26325 257825
rect 25101 257738 25147 257772
rect 25101 257704 25121 257738
rect 25125 257704 25143 257738
rect 21383 257670 21419 257704
rect 25101 257670 25147 257704
rect 21383 257636 21403 257670
rect 21407 257636 21415 257670
rect 7389 257559 8389 257631
rect 8990 257559 9990 257631
rect 21383 257602 21419 257636
rect 15840 257510 15870 257580
rect 15878 257546 15908 257580
rect 21383 257568 21403 257602
rect 21407 257568 21415 257602
rect 15853 257508 15870 257510
rect 21383 257534 21419 257568
rect 21481 257542 22881 257670
rect 23617 257542 25017 257670
rect 25101 257636 25121 257670
rect 25125 257636 25143 257670
rect 25725 257649 26325 257699
rect 25101 257602 25147 257636
rect 25101 257568 25121 257602
rect 25125 257568 25143 257602
rect 25101 257534 25147 257568
rect 5981 257483 6021 257493
rect 5137 257469 6021 257483
rect 21383 257500 21403 257534
rect 21407 257500 21415 257534
rect 21383 257466 21419 257500
rect 7389 257369 8389 257463
rect 7389 257359 8413 257369
rect 8990 257359 9990 257463
rect 21383 257432 21403 257466
rect 21407 257432 21415 257466
rect 21383 257398 21419 257432
rect 21383 257364 21403 257398
rect 21407 257364 21415 257398
rect 21481 257379 22881 257507
rect 23617 257379 25017 257507
rect 25101 257500 25121 257534
rect 25125 257500 25143 257534
rect 25101 257466 25147 257500
rect 25725 257499 26325 257549
rect 25101 257432 25121 257466
rect 25125 257432 25143 257466
rect 25101 257398 25147 257432
rect 25101 257364 25121 257398
rect 25125 257364 25143 257398
rect 25725 257377 26325 257427
rect 21383 257330 21419 257364
rect 25101 257330 25147 257364
rect 21383 257296 21403 257330
rect 21407 257296 21415 257330
rect 25101 257296 25121 257330
rect 25125 257296 25143 257330
rect 21383 257262 21419 257296
rect 21383 257228 21403 257262
rect 21407 257228 21415 257262
rect 21481 257229 22881 257272
rect 23617 257229 25017 257272
rect 25101 257262 25147 257296
rect 25101 257228 25121 257262
rect 25125 257228 25143 257262
rect 21383 257194 21419 257228
rect 25101 257194 25147 257228
rect 25725 257227 26325 257277
rect 21383 257160 21403 257194
rect 21407 257160 21415 257194
rect 25101 257160 25121 257194
rect 25125 257160 25143 257194
rect 27162 257170 27212 258170
rect 27312 257170 27440 258060
rect 27468 257170 27596 258060
rect 27624 257170 27752 258060
rect 27780 257170 27908 258060
rect 27936 257170 28064 258060
rect 28092 257170 28220 258060
rect 28248 257170 28376 258060
rect 28404 257170 28532 258060
rect 28560 257170 28688 258060
rect 28716 257170 28844 258060
rect 28872 257170 29000 258060
rect 29028 257170 29156 258060
rect 29184 257170 29312 258060
rect 29340 257170 29390 258170
rect 30245 258029 30445 258209
rect 30245 258018 30260 258029
rect 30245 258014 30257 258018
rect 30430 258014 30445 258029
rect 30543 258029 30580 258209
rect 30543 258014 30558 258029
rect 30245 257984 30257 257988
rect 30245 257973 30260 257984
rect 30430 257973 30445 257988
rect 30245 257793 30445 257973
rect 31453 257818 32053 257868
rect 30245 257782 30260 257793
rect 30245 257778 30257 257782
rect 30430 257778 30445 257793
rect 31453 257648 32053 257698
rect 30245 257472 30845 257522
rect 30245 257296 30845 257352
rect 21383 257126 21419 257160
rect 25101 257126 25147 257160
rect 21383 257102 21403 257126
rect 21385 257048 21403 257102
rect 21407 257082 21415 257126
rect 25101 257102 25121 257126
rect 25113 257082 25121 257102
rect 25125 257048 25143 257126
rect 30245 257120 30845 257176
rect 30245 256950 30845 257000
rect 21000 256800 21003 256920
rect 21352 256885 21376 256909
rect 25122 256885 25146 256909
rect 21385 256861 21400 256885
rect 25098 256861 25113 256885
rect 21274 256783 21294 256851
rect 21410 256817 21430 256851
rect 25068 256817 25088 256851
rect 25204 256817 25224 256851
rect 21385 256807 21430 256817
rect 25102 256807 25137 256817
rect 21361 256783 21430 256807
rect 25089 256783 25137 256807
rect 25238 256783 25258 256817
rect 680480 250427 680517 250520
rect 680615 250427 680815 250520
rect 685793 250483 685993 250520
rect 686053 250483 686253 250520
rect 686607 250440 687607 250490
rect 692427 250392 693027 250448
rect 679007 250216 679607 250266
rect 680615 250191 680815 250371
rect 686829 250301 687429 250351
rect 684004 250243 685004 250293
rect 695201 250282 695251 250520
rect 696287 250282 696337 250520
rect 682890 250161 683490 250211
rect 684004 250127 685004 250177
rect 686829 250125 687429 250181
rect 679007 250046 679607 250096
rect 684004 249971 685004 250027
rect 686829 249955 687429 250005
rect 680215 249870 680815 249920
rect 681713 249881 682313 249931
rect 682921 249899 683521 249949
rect 692427 249930 693027 249980
rect 684004 249821 685004 249871
rect 680215 249694 680815 249750
rect 681713 249705 682313 249761
rect 682921 249743 683521 249799
rect 685537 249749 686137 249799
rect 697088 249749 697138 250520
rect 697706 249749 697756 250520
rect 699322 250374 700322 250514
rect 700922 250374 701922 250514
rect 707610 250098 708610 250099
rect 699322 249956 700322 250012
rect 700922 249956 701922 250012
rect 707610 250001 708610 250057
rect 709211 250001 710211 250057
rect 707610 249959 708610 249960
rect 699322 249884 700322 249940
rect 700922 249884 701922 249940
rect 709211 249936 710211 249960
rect 682921 249593 683521 249643
rect 684070 249599 684670 249649
rect 685537 249593 686137 249649
rect 699322 249623 700322 249673
rect 700922 249623 701922 249673
rect 680215 249518 680815 249574
rect 707610 249523 708610 249617
rect 709211 249523 710211 249591
rect 707610 249513 707624 249523
rect 707658 249513 707695 249523
rect 707729 249513 707769 249523
rect 707803 249513 707840 249523
rect 707874 249513 707914 249523
rect 707948 249513 707985 249523
rect 708019 249513 708059 249523
rect 708093 249513 708130 249523
rect 708164 249513 708204 249523
rect 708238 249513 708275 249523
rect 708309 249513 708369 249523
rect 708403 249513 708446 249523
rect 708480 249513 708522 249523
rect 708556 249513 708604 249523
rect 709219 249513 709270 249523
rect 709304 249513 709364 249523
rect 709398 249513 709435 249523
rect 709469 249513 709509 249523
rect 709543 249513 709580 249523
rect 709614 249513 709654 249523
rect 709688 249513 709725 249523
rect 709759 249513 709799 249523
rect 709833 249513 709870 249523
rect 709904 249513 709944 249523
rect 709978 249513 710015 249523
rect 710049 249513 710089 249523
rect 710123 249513 710160 249523
rect 710194 249513 710211 249523
rect 684070 249443 684670 249499
rect 685537 249443 686137 249493
rect 692428 249442 693028 249492
rect 680215 249348 680815 249398
rect 681713 249359 682313 249409
rect 684070 249293 684670 249343
rect 692428 249292 693028 249342
rect 705107 249336 705173 249352
rect 711579 249301 711595 250520
rect 711892 249697 711942 250520
rect 712062 249697 712112 250520
rect 716071 250357 716074 250358
rect 714645 250323 714752 250357
rect 716071 250356 716072 250357
rect 716073 250356 716074 250357
rect 716071 250355 716074 250356
rect 716208 250357 716211 250358
rect 716208 250356 716209 250357
rect 716210 250356 716211 250357
rect 716208 250355 716211 250356
rect 714964 250247 715998 250329
rect 716284 250247 717318 250329
rect 714175 249398 714225 249998
rect 714425 249398 714475 249998
rect 680215 249232 680815 249282
rect 698017 249232 698053 249260
rect 692428 249162 693028 249212
rect 698030 249198 698077 249232
rect 698017 249164 698053 249198
rect 680215 249056 680815 249112
rect 692428 249006 693028 249134
rect 698030 249130 698077 249164
rect 698017 249096 698053 249130
rect 698030 249062 698077 249096
rect 698017 248983 698053 249062
rect 698084 248983 698120 249260
rect 714781 249191 714863 250226
rect 715134 249955 715828 250037
rect 714686 249123 714863 249191
rect 714645 249089 714863 249123
rect 680215 248880 680815 248936
rect 686719 248893 686739 248917
rect 686743 248893 686753 248917
rect 686719 248859 686757 248893
rect 686719 248822 686739 248859
rect 686743 248822 686753 248859
rect 692428 248850 693028 248978
rect 698017 248947 698210 248983
rect 698084 248935 698210 248947
rect 702756 248959 703645 248983
rect 702756 248935 702853 248959
rect 698084 248828 702853 248935
rect 686719 248788 686757 248822
rect 680215 248704 680815 248760
rect 686719 248751 686739 248788
rect 686743 248751 686753 248788
rect 686719 248741 686757 248751
rect 686699 248717 686767 248741
rect 686719 248704 686739 248717
rect 686743 248704 686753 248717
rect 686719 248695 686753 248704
rect 686719 248693 686743 248695
rect 692428 248694 693028 248750
rect 686685 248656 686709 248680
rect 686743 248656 686767 248680
rect 678799 248503 679399 248553
rect 680215 248534 680815 248584
rect 692428 248538 693028 248666
rect 680593 248531 680815 248534
rect 682009 248501 682069 248516
rect 682024 248465 682054 248501
rect 683708 248387 684308 248437
rect 678799 248327 679399 248383
rect 692428 248382 693028 248510
rect 714781 248308 714863 249089
rect 715063 248609 715145 249915
rect 715289 248777 715339 249719
rect 715633 248777 715683 249719
rect 715382 248672 715422 248756
rect 715542 248672 715582 248756
rect 715342 248632 715382 248672
rect 715582 248632 715622 248672
rect 715815 248609 715897 249915
rect 715134 248387 715828 248469
rect 716100 248308 716182 250226
rect 716454 249955 717148 250037
rect 716385 248609 716467 249915
rect 716599 248777 716649 249719
rect 716943 248777 716993 249719
rect 716700 248672 716740 248756
rect 716860 248672 716900 248756
rect 716660 248632 716700 248672
rect 716900 248632 716940 248672
rect 717137 248609 717219 249915
rect 716454 248387 717148 248469
rect 717419 248308 717501 250226
rect 683708 248237 684308 248287
rect 692428 248232 693028 248282
rect 678799 248157 679399 248207
rect 684565 248160 684790 248168
rect 696597 248000 696600 248120
rect 714964 248095 715998 248177
rect 716284 248095 717318 248177
rect 21000 221000 21003 221120
rect 282 220623 1316 220705
rect 1602 220623 2636 220705
rect 32810 220662 33035 220670
rect 38201 220593 38801 220643
rect 24572 220518 25172 220568
rect 33292 220513 33892 220563
rect 99 218574 181 220492
rect 452 220331 1146 220413
rect 381 218885 463 220191
rect 660 220128 700 220168
rect 900 220128 940 220168
rect 700 220044 740 220128
rect 860 220044 900 220128
rect 607 219081 657 220023
rect 700 219048 740 219132
rect 860 219048 900 219132
rect 951 219081 1001 220023
rect 660 219008 700 219048
rect 900 219008 940 219048
rect 1133 218885 1215 220191
rect 452 218763 1146 218845
rect 1418 218574 1500 220492
rect 1772 220331 2466 220413
rect 1703 218885 1785 220191
rect 1978 220128 2018 220168
rect 2218 220128 2258 220168
rect 2018 220044 2058 220128
rect 2178 220044 2218 220128
rect 1917 219081 1967 220023
rect 2018 219048 2058 219132
rect 2178 219048 2218 219132
rect 2261 219081 2311 220023
rect 1978 219008 2018 219048
rect 2218 219008 2258 219048
rect 2455 218885 2537 220191
rect 2737 219779 2819 220492
rect 24572 220362 25172 220490
rect 38201 220417 38801 220473
rect 33292 220363 33892 220413
rect 24572 220206 25172 220334
rect 35546 220299 35576 220335
rect 36785 220329 36935 220341
rect 35531 220284 35591 220299
rect 36785 220216 37385 220266
rect 38201 220247 38801 220297
rect 30833 220120 30857 220144
rect 30891 220120 30915 220144
rect 24572 220050 25172 220106
rect 30857 220105 30881 220107
rect 30857 220096 30887 220105
rect 30867 220083 30887 220096
rect 30891 220083 30907 220120
rect 30833 220059 30857 220083
rect 30867 220049 30911 220083
rect 14747 219865 19516 219972
rect 24572 219894 25172 220022
rect 30867 220012 30887 220049
rect 30891 220012 30907 220049
rect 36785 220040 37385 220096
rect 30867 219978 30911 220012
rect 30867 219941 30887 219978
rect 30891 219941 30907 219978
rect 30867 219907 30911 219941
rect 30867 219883 30887 219907
rect 30891 219883 30907 219907
rect 14747 219841 14844 219865
rect 13955 219817 14844 219841
rect 19390 219853 19516 219865
rect 19390 219841 19583 219853
rect 19390 219817 19605 219841
rect 19639 219817 19673 219841
rect 19707 219817 19741 219841
rect 19775 219817 19809 219841
rect 19843 219817 19877 219841
rect 19911 219817 19945 219841
rect 19979 219817 20013 219841
rect 20047 219817 20081 219841
rect 20115 219817 20149 219841
rect 20183 219817 20217 219841
rect 20251 219817 20285 219841
rect 20319 219817 20353 219841
rect 20387 219817 20421 219841
rect 20455 219817 20489 219841
rect 20523 219817 20557 219841
rect 20591 219817 20625 219841
rect 20659 219817 20693 219841
rect 2737 219711 2914 219779
rect 1772 218763 2466 218845
rect 2737 218574 2819 219711
rect 2848 219677 2955 219711
rect 6005 219498 6021 219499
rect 3125 218802 3175 219402
rect 3375 218802 3425 219402
rect 5967 219363 6059 219498
rect 12427 219448 12493 219464
rect 282 218471 1316 218553
rect 1602 218471 2636 218553
rect 2806 218477 2914 218545
rect 1389 218444 1392 218445
rect 1389 218443 1390 218444
rect 1391 218443 1392 218444
rect 1389 218442 1392 218443
rect 1526 218444 1529 218445
rect 1526 218443 1527 218444
rect 1528 218443 1529 218444
rect 2848 218443 2955 218477
rect 1526 218442 1529 218443
rect 5488 218103 5538 219103
rect 5658 218103 5708 219103
rect 183 217602 1183 217652
rect 2850 217632 3850 217682
rect 183 217446 1183 217574
rect 2850 217416 3850 217544
rect 183 217296 1183 217346
rect 183 217180 1183 217230
rect 2850 217200 3850 217328
rect 183 216964 1183 217020
rect 2850 216984 3850 217112
rect 5488 216993 5538 217993
rect 5658 216993 5708 217993
rect 183 216748 1183 216804
rect 2850 216768 3850 216896
rect 183 216592 1183 216720
rect 2850 216552 3850 216608
rect 183 216442 1183 216492
rect 2850 216336 3850 216392
rect 183 216276 1183 216326
rect 2850 216120 3850 216248
rect 183 216060 1183 216116
rect 183 215904 1183 216032
rect 2850 215904 3850 216032
rect 5488 215872 5538 216872
rect 5658 215872 5708 216872
rect 183 215748 1183 215804
rect 183 215592 1183 215720
rect 2850 215688 3850 215816
rect 183 215436 1183 215492
rect 2850 215472 3850 215600
rect 183 215286 1183 215336
rect 2850 215256 3850 215312
rect 583 215170 1183 215220
rect 583 215020 1183 215070
rect 2850 215040 3850 215168
rect 183 214904 1183 214954
rect 2850 214824 3850 214952
rect 183 214748 1183 214804
rect 5488 214751 5538 215751
rect 5658 214751 5708 215751
rect 183 214598 1183 214648
rect 2850 214608 3850 214736
rect 5971 214489 6059 219363
rect 7406 219287 7440 219321
rect 7477 219287 7511 219321
rect 7551 219287 7585 219321
rect 7622 219287 7656 219321
rect 7696 219287 7730 219321
rect 7767 219287 7801 219321
rect 7841 219287 7875 219321
rect 7912 219287 7946 219321
rect 7986 219287 8020 219321
rect 8057 219287 8091 219321
rect 8131 219287 8165 219321
rect 8202 219287 8236 219321
rect 8296 219287 8330 219321
rect 8381 219311 8423 219321
rect 8381 219287 8389 219311
rect 8415 219287 8423 219311
rect 8956 219311 8996 219321
rect 8956 219287 8962 219311
rect 8990 219287 8996 219311
rect 9044 219287 9078 219321
rect 9120 219287 9154 219321
rect 9197 219287 9231 219321
rect 9291 219287 9325 219321
rect 9362 219287 9396 219321
rect 9436 219287 9470 219321
rect 9507 219287 9541 219321
rect 9581 219287 9615 219321
rect 9652 219287 9686 219321
rect 9726 219287 9760 219321
rect 9797 219287 9831 219321
rect 9871 219287 9905 219321
rect 9942 219287 9976 219321
rect 7389 219277 7406 219287
rect 7440 219277 7477 219287
rect 7511 219277 7551 219287
rect 7585 219277 7622 219287
rect 7656 219277 7696 219287
rect 7730 219277 7767 219287
rect 7801 219277 7841 219287
rect 7875 219277 7912 219287
rect 7946 219277 7986 219287
rect 8020 219277 8057 219287
rect 8091 219277 8131 219287
rect 8165 219277 8202 219287
rect 8236 219277 8296 219287
rect 8330 219277 8381 219287
rect 8389 219277 8423 219287
rect 8990 219277 9044 219287
rect 9078 219277 9120 219287
rect 9154 219277 9197 219287
rect 9231 219277 9291 219287
rect 9325 219277 9362 219287
rect 9396 219277 9436 219287
rect 9470 219277 9507 219287
rect 9541 219277 9581 219287
rect 9615 219277 9652 219287
rect 9686 219277 9726 219287
rect 9760 219277 9797 219287
rect 9831 219277 9871 219287
rect 9905 219277 9942 219287
rect 9976 219277 9990 219287
rect 7389 219209 8389 219277
rect 8990 219183 9990 219277
rect 7389 219087 8389 219147
rect 8990 219087 9990 219147
rect 15678 219127 16678 219177
rect 17278 219127 18278 219177
rect 7353 218864 7389 218876
rect 8389 218864 8425 218876
rect 7353 218840 8425 218864
rect 7353 218799 7389 218840
rect 8389 218799 8425 218840
rect 7353 218743 8425 218799
rect 7353 218706 7389 218743
rect 8389 218706 8425 218743
rect 7353 218666 8425 218706
rect 8954 218841 8990 218876
rect 9990 218841 10026 218876
rect 15678 218860 16678 218916
rect 17278 218860 18278 218916
rect 8954 218840 10026 218841
rect 8954 218799 8990 218840
rect 9990 218799 10026 218840
rect 8954 218743 10026 218799
rect 15678 218788 16678 218844
rect 17278 218788 18278 218844
rect 8954 218706 8990 218743
rect 9990 218706 10026 218743
rect 8954 218701 10026 218706
rect 8954 218666 8990 218701
rect 9990 218666 10026 218701
rect 7389 218441 8389 218513
rect 8990 218441 9990 218513
rect 15678 218486 16678 218558
rect 17278 218486 18278 218558
rect 15748 218475 15782 218486
rect 15816 218475 15850 218486
rect 15884 218475 15918 218486
rect 15952 218475 15986 218486
rect 16020 218475 16054 218486
rect 16088 218475 16122 218486
rect 16156 218475 16190 218486
rect 16224 218475 16258 218486
rect 16292 218475 16326 218486
rect 16360 218475 16394 218486
rect 16428 218475 16462 218486
rect 16496 218475 16530 218486
rect 16564 218475 16598 218486
rect 16632 218475 16666 218486
rect 17290 218475 17324 218486
rect 17358 218475 17392 218486
rect 17426 218475 17460 218486
rect 17494 218475 17528 218486
rect 17562 218475 17596 218486
rect 17630 218475 17664 218486
rect 17698 218475 17732 218486
rect 17766 218475 17800 218486
rect 17834 218475 17868 218486
rect 17902 218475 17936 218486
rect 17970 218475 18004 218486
rect 18038 218475 18072 218486
rect 18106 218475 18140 218486
rect 18174 218475 18208 218486
rect 15748 218465 15806 218475
rect 15816 218465 15874 218475
rect 15884 218465 15942 218475
rect 15952 218465 16010 218475
rect 16020 218465 16078 218475
rect 16088 218465 16146 218475
rect 16156 218465 16214 218475
rect 16224 218465 16282 218475
rect 16292 218465 16350 218475
rect 16360 218465 16418 218475
rect 16428 218465 16486 218475
rect 16496 218465 16554 218475
rect 16564 218465 16622 218475
rect 16632 218465 16690 218475
rect 17290 218465 17348 218475
rect 17358 218465 17416 218475
rect 17426 218465 17484 218475
rect 17494 218465 17552 218475
rect 17562 218465 17620 218475
rect 17630 218465 17688 218475
rect 17698 218465 17756 218475
rect 17766 218465 17824 218475
rect 17834 218465 17892 218475
rect 17902 218465 17960 218475
rect 17970 218465 18028 218475
rect 18038 218465 18096 218475
rect 18106 218465 18164 218475
rect 18174 218465 18232 218475
rect 15724 218441 16690 218465
rect 17266 218441 18232 218465
rect 15748 218426 15772 218441
rect 15816 218426 15840 218441
rect 15884 218426 15908 218441
rect 15952 218426 15976 218441
rect 16020 218426 16044 218441
rect 16088 218426 16112 218441
rect 16156 218426 16180 218441
rect 16224 218426 16248 218441
rect 16292 218426 16316 218441
rect 16360 218426 16384 218441
rect 16428 218426 16452 218441
rect 16496 218426 16520 218441
rect 16564 218426 16588 218441
rect 16632 218426 16656 218441
rect 17290 218426 17314 218441
rect 17358 218426 17382 218441
rect 17426 218426 17450 218441
rect 17494 218426 17518 218441
rect 17562 218426 17586 218441
rect 17630 218426 17654 218441
rect 17698 218426 17722 218441
rect 17766 218426 17790 218441
rect 17834 218426 17858 218441
rect 17902 218426 17926 218441
rect 17970 218426 17994 218441
rect 18038 218426 18062 218441
rect 18106 218426 18130 218441
rect 18174 218426 18198 218441
rect 15678 218271 16678 218426
rect 7389 218181 8389 218241
rect 8990 218181 9990 218241
rect 15678 218237 16690 218271
rect 17278 218261 18278 218426
rect 17266 218237 18278 218261
rect 15678 218226 16678 218237
rect 17278 218226 18278 218237
rect 15748 218213 15772 218226
rect 15816 218213 15840 218226
rect 15884 218213 15908 218226
rect 15952 218213 15976 218226
rect 16020 218213 16044 218226
rect 16088 218213 16112 218226
rect 16156 218213 16180 218226
rect 16224 218213 16248 218226
rect 16292 218213 16316 218226
rect 16360 218213 16384 218226
rect 16428 218213 16452 218226
rect 16496 218213 16520 218226
rect 16564 218213 16588 218226
rect 16632 218213 16656 218226
rect 17290 218213 17314 218226
rect 17358 218213 17382 218226
rect 17426 218213 17450 218226
rect 17494 218213 17518 218226
rect 17562 218213 17586 218226
rect 17630 218213 17654 218226
rect 17698 218213 17722 218226
rect 17766 218213 17790 218226
rect 17834 218213 17858 218226
rect 17902 218213 17926 218226
rect 17970 218213 17994 218226
rect 18038 218213 18062 218226
rect 18106 218213 18130 218226
rect 18174 218213 18198 218226
rect 7389 217823 8389 217879
rect 8990 217823 9990 217879
rect 15678 217868 16678 217924
rect 17278 217868 18278 217924
rect 7389 217751 8389 217807
rect 8990 217751 9990 217807
rect 15678 217796 16678 217852
rect 17278 217796 18278 217852
rect 7389 217449 8389 217521
rect 8990 217449 9990 217521
rect 15678 217494 16678 217566
rect 17278 217494 18278 217566
rect 15748 217483 15782 217494
rect 15816 217483 15850 217494
rect 15884 217483 15918 217494
rect 15952 217483 15986 217494
rect 16020 217483 16054 217494
rect 16088 217483 16122 217494
rect 16156 217483 16190 217494
rect 16224 217483 16258 217494
rect 16292 217483 16326 217494
rect 16360 217483 16394 217494
rect 16428 217483 16462 217494
rect 16496 217483 16530 217494
rect 16564 217483 16598 217494
rect 16632 217483 16666 217494
rect 17290 217483 17324 217494
rect 17358 217483 17392 217494
rect 17426 217483 17460 217494
rect 17494 217483 17528 217494
rect 17562 217483 17596 217494
rect 17630 217483 17664 217494
rect 17698 217483 17732 217494
rect 17766 217483 17800 217494
rect 17834 217483 17868 217494
rect 17902 217483 17936 217494
rect 17970 217483 18004 217494
rect 18038 217483 18072 217494
rect 18106 217483 18140 217494
rect 18174 217483 18208 217494
rect 15748 217473 15806 217483
rect 15816 217473 15874 217483
rect 15884 217473 15942 217483
rect 15952 217473 16010 217483
rect 16020 217473 16078 217483
rect 16088 217473 16146 217483
rect 16156 217473 16214 217483
rect 16224 217473 16282 217483
rect 16292 217473 16350 217483
rect 16360 217473 16418 217483
rect 16428 217473 16486 217483
rect 16496 217473 16554 217483
rect 16564 217473 16622 217483
rect 16632 217473 16690 217483
rect 17290 217473 17348 217483
rect 17358 217473 17416 217483
rect 17426 217473 17484 217483
rect 17494 217473 17552 217483
rect 17562 217473 17620 217483
rect 17630 217473 17688 217483
rect 17698 217473 17756 217483
rect 17766 217473 17824 217483
rect 17834 217473 17892 217483
rect 17902 217473 17960 217483
rect 17970 217473 18028 217483
rect 18038 217473 18096 217483
rect 18106 217473 18164 217483
rect 18174 217473 18232 217483
rect 15724 217449 16690 217473
rect 17266 217449 18232 217473
rect 12427 217424 12493 217440
rect 15748 217434 15772 217449
rect 15816 217434 15840 217449
rect 15884 217434 15908 217449
rect 15952 217434 15976 217449
rect 16020 217434 16044 217449
rect 16088 217434 16112 217449
rect 16156 217434 16180 217449
rect 16224 217434 16248 217449
rect 16292 217434 16316 217449
rect 16360 217434 16384 217449
rect 16428 217434 16452 217449
rect 16496 217434 16520 217449
rect 16564 217434 16588 217449
rect 16632 217434 16656 217449
rect 17290 217434 17314 217449
rect 17358 217434 17382 217449
rect 17426 217434 17450 217449
rect 17494 217434 17518 217449
rect 17562 217434 17586 217449
rect 17630 217434 17654 217449
rect 17698 217434 17722 217449
rect 17766 217434 17790 217449
rect 17834 217434 17858 217449
rect 17902 217434 17926 217449
rect 17970 217434 17994 217449
rect 18038 217434 18062 217449
rect 18106 217434 18130 217449
rect 18174 217434 18198 217449
rect 15678 217279 16678 217434
rect 7389 217189 8389 217249
rect 8990 217189 9990 217249
rect 15678 217245 16690 217279
rect 17278 217269 18278 217434
rect 17266 217245 18278 217269
rect 15678 217234 16678 217245
rect 17278 217234 18278 217245
rect 15748 217221 15772 217234
rect 15816 217221 15840 217234
rect 15884 217221 15908 217234
rect 15952 217221 15976 217234
rect 16020 217221 16044 217234
rect 16088 217221 16112 217234
rect 16156 217221 16180 217234
rect 16224 217221 16248 217234
rect 16292 217221 16316 217234
rect 16360 217221 16384 217234
rect 16428 217221 16452 217234
rect 16496 217221 16520 217234
rect 16564 217221 16588 217234
rect 16632 217221 16656 217234
rect 17290 217221 17314 217234
rect 17358 217221 17382 217234
rect 17426 217221 17450 217234
rect 17494 217221 17518 217234
rect 17562 217221 17586 217234
rect 17630 217221 17654 217234
rect 17698 217221 17722 217234
rect 17766 217221 17790 217234
rect 17834 217221 17858 217234
rect 17902 217221 17926 217234
rect 17970 217221 17994 217234
rect 18038 217221 18062 217234
rect 18106 217221 18130 217234
rect 18174 217221 18198 217234
rect 7389 216831 8389 216887
rect 8990 216831 9990 216887
rect 15678 216876 16678 216932
rect 17278 216876 18278 216932
rect 7389 216759 8389 216815
rect 8990 216759 9990 216815
rect 15678 216804 16678 216860
rect 17278 216804 18278 216860
rect 7389 216457 8389 216529
rect 8990 216457 9990 216529
rect 15678 216502 16678 216574
rect 17278 216502 18278 216574
rect 15748 216491 15782 216502
rect 15816 216491 15850 216502
rect 15884 216491 15918 216502
rect 15952 216491 15986 216502
rect 16020 216491 16054 216502
rect 16088 216491 16122 216502
rect 16156 216491 16190 216502
rect 16224 216491 16258 216502
rect 16292 216491 16326 216502
rect 16360 216491 16394 216502
rect 16428 216491 16462 216502
rect 16496 216491 16530 216502
rect 16564 216491 16598 216502
rect 16632 216491 16666 216502
rect 17290 216491 17324 216502
rect 17358 216491 17392 216502
rect 17426 216491 17460 216502
rect 17494 216491 17528 216502
rect 17562 216491 17596 216502
rect 17630 216491 17664 216502
rect 17698 216491 17732 216502
rect 17766 216491 17800 216502
rect 17834 216491 17868 216502
rect 17902 216491 17936 216502
rect 17970 216491 18004 216502
rect 18038 216491 18072 216502
rect 18106 216491 18140 216502
rect 18174 216491 18208 216502
rect 15748 216481 15806 216491
rect 15816 216481 15874 216491
rect 15884 216481 15942 216491
rect 15952 216481 16010 216491
rect 16020 216481 16078 216491
rect 16088 216481 16146 216491
rect 16156 216481 16214 216491
rect 16224 216481 16282 216491
rect 16292 216481 16350 216491
rect 16360 216481 16418 216491
rect 16428 216481 16486 216491
rect 16496 216481 16554 216491
rect 16564 216481 16622 216491
rect 16632 216481 16690 216491
rect 17290 216481 17348 216491
rect 17358 216481 17416 216491
rect 17426 216481 17484 216491
rect 17494 216481 17552 216491
rect 17562 216481 17620 216491
rect 17630 216481 17688 216491
rect 17698 216481 17756 216491
rect 17766 216481 17824 216491
rect 17834 216481 17892 216491
rect 17902 216481 17960 216491
rect 17970 216481 18028 216491
rect 18038 216481 18096 216491
rect 18106 216481 18164 216491
rect 18174 216481 18232 216491
rect 15724 216457 16690 216481
rect 17266 216457 18232 216481
rect 15748 216442 15772 216457
rect 15816 216442 15840 216457
rect 15884 216442 15908 216457
rect 15952 216442 15976 216457
rect 16020 216442 16044 216457
rect 16088 216442 16112 216457
rect 16156 216442 16180 216457
rect 16224 216442 16248 216457
rect 16292 216442 16316 216457
rect 16360 216442 16384 216457
rect 16428 216442 16452 216457
rect 16496 216442 16520 216457
rect 16564 216442 16588 216457
rect 16632 216442 16656 216457
rect 17290 216442 17314 216457
rect 17358 216442 17382 216457
rect 17426 216442 17450 216457
rect 17494 216442 17518 216457
rect 17562 216442 17586 216457
rect 17630 216442 17654 216457
rect 17698 216442 17722 216457
rect 17766 216442 17790 216457
rect 17834 216442 17858 216457
rect 17902 216442 17926 216457
rect 17970 216442 17994 216457
rect 18038 216442 18062 216457
rect 18106 216442 18130 216457
rect 18174 216442 18198 216457
rect 15678 216287 16678 216442
rect 7389 216197 8389 216257
rect 8990 216197 9990 216257
rect 15678 216253 16690 216287
rect 17278 216277 18278 216442
rect 17266 216253 18278 216277
rect 15678 216242 16678 216253
rect 17278 216242 18278 216253
rect 15748 216229 15772 216242
rect 15816 216229 15840 216242
rect 15884 216229 15908 216242
rect 15952 216229 15976 216242
rect 16020 216229 16044 216242
rect 16088 216229 16112 216242
rect 16156 216229 16180 216242
rect 16224 216229 16248 216242
rect 16292 216229 16316 216242
rect 16360 216229 16384 216242
rect 16428 216229 16452 216242
rect 16496 216229 16520 216242
rect 16564 216229 16588 216242
rect 16632 216229 16656 216242
rect 17290 216229 17314 216242
rect 17358 216229 17382 216242
rect 17426 216229 17450 216242
rect 17494 216229 17518 216242
rect 17562 216229 17586 216242
rect 17630 216229 17654 216242
rect 17698 216229 17722 216242
rect 17766 216229 17790 216242
rect 17834 216229 17858 216242
rect 17902 216229 17926 216242
rect 17970 216229 17994 216242
rect 18038 216229 18062 216242
rect 18106 216229 18130 216242
rect 18174 216229 18198 216242
rect 7389 215839 8389 215895
rect 8990 215839 9990 215895
rect 15678 215884 16678 215940
rect 17278 215884 18278 215940
rect 7389 215767 8389 215823
rect 8990 215767 9990 215823
rect 15678 215812 16678 215868
rect 17278 215812 18278 215868
rect 7389 215465 8389 215537
rect 8990 215465 9990 215537
rect 15678 215510 16678 215582
rect 17278 215510 18278 215582
rect 15748 215499 15782 215510
rect 15816 215499 15850 215510
rect 15884 215499 15918 215510
rect 15952 215499 15986 215510
rect 16020 215499 16054 215510
rect 16088 215499 16122 215510
rect 16156 215499 16190 215510
rect 16224 215499 16258 215510
rect 16292 215499 16326 215510
rect 16360 215499 16394 215510
rect 16428 215499 16462 215510
rect 16496 215499 16530 215510
rect 16564 215499 16598 215510
rect 16632 215499 16666 215510
rect 17290 215499 17324 215510
rect 17358 215499 17392 215510
rect 17426 215499 17460 215510
rect 17494 215499 17528 215510
rect 17562 215499 17596 215510
rect 17630 215499 17664 215510
rect 17698 215499 17732 215510
rect 17766 215499 17800 215510
rect 17834 215499 17868 215510
rect 17902 215499 17936 215510
rect 17970 215499 18004 215510
rect 18038 215499 18072 215510
rect 18106 215499 18140 215510
rect 18174 215499 18208 215510
rect 15748 215489 15806 215499
rect 15816 215489 15874 215499
rect 15884 215489 15942 215499
rect 15952 215489 16010 215499
rect 16020 215489 16078 215499
rect 16088 215489 16146 215499
rect 16156 215489 16214 215499
rect 16224 215489 16282 215499
rect 16292 215489 16350 215499
rect 16360 215489 16418 215499
rect 16428 215489 16486 215499
rect 16496 215489 16554 215499
rect 16564 215489 16622 215499
rect 16632 215489 16690 215499
rect 17290 215489 17348 215499
rect 17358 215489 17416 215499
rect 17426 215489 17484 215499
rect 17494 215489 17552 215499
rect 17562 215489 17620 215499
rect 17630 215489 17688 215499
rect 17698 215489 17756 215499
rect 17766 215489 17824 215499
rect 17834 215489 17892 215499
rect 17902 215489 17960 215499
rect 17970 215489 18028 215499
rect 18038 215489 18096 215499
rect 18106 215489 18164 215499
rect 18174 215489 18232 215499
rect 15724 215465 16690 215489
rect 17266 215465 18232 215489
rect 15748 215450 15772 215465
rect 15816 215450 15840 215465
rect 15884 215450 15908 215465
rect 15952 215450 15976 215465
rect 16020 215450 16044 215465
rect 16088 215450 16112 215465
rect 16156 215450 16180 215465
rect 16224 215450 16248 215465
rect 16292 215450 16316 215465
rect 16360 215450 16384 215465
rect 16428 215450 16452 215465
rect 16496 215450 16520 215465
rect 16564 215450 16588 215465
rect 16632 215450 16656 215465
rect 17290 215450 17314 215465
rect 17358 215450 17382 215465
rect 17426 215450 17450 215465
rect 17494 215450 17518 215465
rect 17562 215450 17586 215465
rect 17630 215450 17654 215465
rect 17698 215450 17722 215465
rect 17766 215450 17790 215465
rect 17834 215450 17858 215465
rect 17902 215450 17926 215465
rect 17970 215450 17994 215465
rect 18038 215450 18062 215465
rect 18106 215450 18130 215465
rect 18174 215450 18198 215465
rect 15678 215295 16678 215450
rect 7389 215205 8389 215265
rect 8990 215205 9990 215265
rect 15678 215261 16690 215295
rect 17278 215285 18278 215450
rect 17266 215261 18278 215285
rect 15678 215250 16678 215261
rect 17278 215250 18278 215261
rect 15748 215237 15772 215250
rect 15816 215237 15840 215250
rect 15884 215237 15908 215250
rect 15952 215237 15976 215250
rect 16020 215237 16044 215250
rect 16088 215237 16112 215250
rect 16156 215237 16180 215250
rect 16224 215237 16248 215250
rect 16292 215237 16316 215250
rect 16360 215237 16384 215250
rect 16428 215237 16452 215250
rect 16496 215237 16520 215250
rect 16564 215237 16588 215250
rect 16632 215237 16656 215250
rect 17290 215237 17314 215250
rect 17358 215237 17382 215250
rect 17426 215237 17450 215250
rect 17494 215237 17518 215250
rect 17562 215237 17586 215250
rect 17630 215237 17654 215250
rect 17698 215237 17722 215250
rect 17766 215237 17790 215250
rect 17834 215237 17858 215250
rect 17902 215237 17926 215250
rect 17970 215237 17994 215250
rect 18038 215237 18062 215250
rect 18106 215237 18130 215250
rect 18174 215237 18198 215250
rect 7389 214847 8389 214903
rect 8990 214847 9990 214903
rect 15678 214892 16678 214948
rect 17278 214892 18278 214948
rect 7389 214775 8389 214831
rect 8990 214775 9990 214831
rect 15678 214820 16678 214876
rect 17278 214820 18278 214876
rect 5967 214455 6059 214489
rect 7389 214473 8389 214545
rect 8990 214473 9990 214545
rect 15678 214518 16678 214590
rect 17278 214518 18278 214590
rect 15748 214507 15782 214518
rect 15816 214507 15850 214518
rect 15884 214507 15918 214518
rect 15952 214507 15986 214518
rect 16020 214507 16054 214518
rect 16088 214507 16122 214518
rect 16156 214507 16190 214518
rect 16224 214507 16258 214518
rect 16292 214507 16326 214518
rect 16360 214507 16394 214518
rect 16428 214507 16462 214518
rect 16496 214507 16530 214518
rect 16564 214507 16598 214518
rect 16632 214507 16666 214518
rect 17290 214507 17324 214518
rect 17358 214507 17392 214518
rect 17426 214507 17460 214518
rect 17494 214507 17528 214518
rect 17562 214507 17596 214518
rect 17630 214507 17664 214518
rect 17698 214507 17732 214518
rect 17766 214507 17800 214518
rect 17834 214507 17868 214518
rect 17902 214507 17936 214518
rect 17970 214507 18004 214518
rect 18038 214507 18072 214518
rect 18106 214507 18140 214518
rect 18174 214507 18208 214518
rect 15748 214497 15806 214507
rect 15816 214497 15874 214507
rect 15884 214497 15942 214507
rect 15952 214497 16010 214507
rect 16020 214497 16078 214507
rect 16088 214497 16146 214507
rect 16156 214497 16214 214507
rect 16224 214497 16282 214507
rect 16292 214497 16350 214507
rect 16360 214497 16418 214507
rect 16428 214497 16486 214507
rect 16496 214497 16554 214507
rect 16564 214497 16622 214507
rect 16632 214497 16690 214507
rect 17290 214497 17348 214507
rect 17358 214497 17416 214507
rect 17426 214497 17484 214507
rect 17494 214497 17552 214507
rect 17562 214497 17620 214507
rect 17630 214497 17688 214507
rect 17698 214497 17756 214507
rect 17766 214497 17824 214507
rect 17834 214497 17892 214507
rect 17902 214497 17960 214507
rect 17970 214497 18028 214507
rect 18038 214497 18096 214507
rect 18106 214497 18164 214507
rect 18174 214497 18232 214507
rect 15724 214473 16690 214497
rect 17266 214473 18232 214497
rect 15748 214458 15772 214473
rect 15816 214458 15840 214473
rect 15884 214458 15908 214473
rect 15952 214458 15976 214473
rect 16020 214458 16044 214473
rect 16088 214458 16112 214473
rect 16156 214458 16180 214473
rect 16224 214458 16248 214473
rect 16292 214458 16316 214473
rect 16360 214458 16384 214473
rect 16428 214458 16452 214473
rect 16496 214458 16520 214473
rect 16564 214458 16588 214473
rect 16632 214458 16656 214473
rect 17290 214458 17314 214473
rect 17358 214458 17382 214473
rect 17426 214458 17450 214473
rect 17494 214458 17518 214473
rect 17562 214458 17586 214473
rect 17630 214458 17654 214473
rect 17698 214458 17722 214473
rect 17766 214458 17790 214473
rect 17834 214458 17858 214473
rect 17902 214458 17926 214473
rect 17970 214458 17994 214473
rect 18038 214458 18062 214473
rect 18106 214458 18130 214473
rect 18174 214458 18198 214473
rect 2850 214398 3850 214448
rect 2850 214282 3850 214332
rect 2850 214072 3850 214122
rect 2850 213956 3850 214006
rect 2850 213746 3850 213796
rect 1153 213660 1187 213718
rect 2850 213630 3850 213680
rect 2850 213420 3850 213470
rect 2850 213417 3107 213420
rect 3250 213304 3850 213354
rect 3250 213048 3850 213104
rect 3250 212892 3850 213020
rect 175 212818 1175 212868
rect 175 212662 1175 212790
rect 3250 212736 3850 212792
rect 175 212506 1175 212634
rect 175 212350 1175 212478
rect 175 212194 1175 212322
rect 175 212044 1175 212094
rect 175 211928 1175 211978
rect 175 211772 1175 211828
rect 175 211622 1175 211672
rect 1578 211609 1628 212609
rect 1728 211609 1856 212609
rect 1884 211609 2012 212609
rect 2040 211609 2090 212609
rect 3250 212580 3850 212708
rect 3250 212430 3850 212480
rect 2850 212314 3850 212364
rect 2850 212158 3850 212214
rect 2850 212008 3850 212058
rect 2850 211880 3850 211930
rect 2850 211724 3850 211852
rect 2850 211568 3850 211696
rect 175 211506 1175 211556
rect 175 211350 1175 211478
rect 2850 211412 3850 211468
rect 2850 211256 3850 211384
rect 175 211194 1175 211250
rect 175 211038 1175 211166
rect 175 210888 1175 210938
rect 175 210772 1175 210822
rect 175 210616 1175 210744
rect 1578 210613 1628 211213
rect 1728 210613 1784 211213
rect 1884 210613 1940 211213
rect 2040 210613 2096 211213
rect 2196 210613 2246 211213
rect 2850 211100 3850 211228
rect 2850 210944 3850 211072
rect 2850 210794 3850 210844
rect 2850 210678 3850 210728
rect 2850 210522 3850 210650
rect 175 210460 1175 210516
rect 175 210304 1175 210432
rect 2850 210366 3850 210494
rect 2850 210210 3850 210338
rect 175 210154 1175 210204
rect 803 210151 1175 210154
rect 2850 210054 3850 210110
rect 2850 209898 3850 210026
rect 2850 209742 3850 209870
rect 2850 209586 3850 209642
rect 2850 209436 3850 209486
rect 3926 209455 3960 209491
rect 3967 209339 3989 209455
rect 1638 207869 1688 208869
rect 1848 207869 1976 208869
rect 2064 207869 2114 208869
rect 2850 208275 3050 208287
rect 2850 208162 3850 208212
rect 2850 207946 3850 208074
rect 2850 207730 3850 207786
rect 2850 207514 3850 207642
rect 2850 207304 3850 207354
rect 2850 207188 3850 207238
rect 2850 206978 3850 207028
rect 3926 207015 3960 209339
rect 5169 207315 5191 214429
rect 5488 213194 5538 214194
rect 5658 213194 5708 214194
rect 5488 212073 5538 213073
rect 5658 212073 5708 213073
rect 5488 210952 5538 211952
rect 5658 210952 5708 211952
rect 5488 209842 5538 210842
rect 5658 209842 5708 210842
rect 5488 208721 5538 209721
rect 5658 208721 5708 209721
rect 5488 207600 5538 208600
rect 5658 207600 5708 208600
rect 5971 207386 6059 214455
rect 15678 214303 16678 214458
rect 7389 214213 8389 214273
rect 8990 214213 9990 214273
rect 15678 214269 16690 214303
rect 17278 214293 18278 214458
rect 17266 214269 18278 214293
rect 15678 214258 16678 214269
rect 17278 214258 18278 214269
rect 15748 214245 15772 214258
rect 15816 214245 15840 214258
rect 15884 214245 15908 214258
rect 15952 214245 15976 214258
rect 16020 214245 16044 214258
rect 16088 214245 16112 214258
rect 16156 214245 16180 214258
rect 16224 214245 16248 214258
rect 16292 214245 16316 214258
rect 16360 214245 16384 214258
rect 16428 214245 16452 214258
rect 16496 214245 16520 214258
rect 16564 214245 16588 214258
rect 16632 214245 16656 214258
rect 17290 214245 17314 214258
rect 17358 214245 17382 214258
rect 17426 214245 17450 214258
rect 17494 214245 17518 214258
rect 17562 214245 17586 214258
rect 17630 214245 17654 214258
rect 17698 214245 17722 214258
rect 17766 214245 17790 214258
rect 17834 214245 17858 214258
rect 17902 214245 17926 214258
rect 17970 214245 17994 214258
rect 18038 214245 18062 214258
rect 18106 214245 18130 214258
rect 18174 214245 18198 214258
rect 7389 213855 8389 213911
rect 8990 213855 9990 213911
rect 15678 213900 16678 213956
rect 17278 213900 18278 213956
rect 7389 213783 8389 213839
rect 8990 213783 9990 213839
rect 15678 213828 16678 213884
rect 17278 213828 18278 213884
rect 7389 213481 8389 213553
rect 8990 213481 9990 213553
rect 15678 213526 16678 213598
rect 17278 213526 18278 213598
rect 15748 213515 15782 213526
rect 15816 213515 15850 213526
rect 15884 213515 15918 213526
rect 15952 213515 15986 213526
rect 16020 213515 16054 213526
rect 16088 213515 16122 213526
rect 16156 213515 16190 213526
rect 16224 213515 16258 213526
rect 16292 213515 16326 213526
rect 16360 213515 16394 213526
rect 16428 213515 16462 213526
rect 16496 213515 16530 213526
rect 16564 213515 16598 213526
rect 16632 213515 16666 213526
rect 17290 213515 17324 213526
rect 17358 213515 17392 213526
rect 17426 213515 17460 213526
rect 17494 213515 17528 213526
rect 17562 213515 17596 213526
rect 17630 213515 17664 213526
rect 17698 213515 17732 213526
rect 17766 213515 17800 213526
rect 17834 213515 17868 213526
rect 17902 213515 17936 213526
rect 17970 213515 18004 213526
rect 18038 213515 18072 213526
rect 18106 213515 18140 213526
rect 18174 213515 18208 213526
rect 15748 213505 15806 213515
rect 15816 213505 15874 213515
rect 15884 213505 15942 213515
rect 15952 213505 16010 213515
rect 16020 213505 16078 213515
rect 16088 213505 16146 213515
rect 16156 213505 16214 213515
rect 16224 213505 16282 213515
rect 16292 213505 16350 213515
rect 16360 213505 16418 213515
rect 16428 213505 16486 213515
rect 16496 213505 16554 213515
rect 16564 213505 16622 213515
rect 16632 213505 16690 213515
rect 17290 213505 17348 213515
rect 17358 213505 17416 213515
rect 17426 213505 17484 213515
rect 17494 213505 17552 213515
rect 17562 213505 17620 213515
rect 17630 213505 17688 213515
rect 17698 213505 17756 213515
rect 17766 213505 17824 213515
rect 17834 213505 17892 213515
rect 17902 213505 17960 213515
rect 17970 213505 18028 213515
rect 18038 213505 18096 213515
rect 18106 213505 18164 213515
rect 18174 213505 18232 213515
rect 15724 213481 16690 213505
rect 17266 213481 18232 213505
rect 15748 213466 15772 213481
rect 15816 213466 15840 213481
rect 15884 213466 15908 213481
rect 15952 213466 15976 213481
rect 16020 213466 16044 213481
rect 16088 213466 16112 213481
rect 16156 213466 16180 213481
rect 16224 213466 16248 213481
rect 16292 213466 16316 213481
rect 16360 213466 16384 213481
rect 16428 213466 16452 213481
rect 16496 213466 16520 213481
rect 16564 213466 16588 213481
rect 16632 213466 16656 213481
rect 17290 213466 17314 213481
rect 17358 213466 17382 213481
rect 17426 213466 17450 213481
rect 17494 213466 17518 213481
rect 17562 213466 17586 213481
rect 17630 213466 17654 213481
rect 17698 213466 17722 213481
rect 17766 213466 17790 213481
rect 17834 213466 17858 213481
rect 17902 213466 17926 213481
rect 17970 213466 17994 213481
rect 18038 213466 18062 213481
rect 18106 213466 18130 213481
rect 18174 213466 18198 213481
rect 15678 213311 16678 213466
rect 7389 213221 8389 213281
rect 8990 213221 9990 213281
rect 15678 213277 16690 213311
rect 17278 213301 18278 213466
rect 17266 213277 18278 213301
rect 15678 213266 16678 213277
rect 17278 213266 18278 213277
rect 15748 213253 15772 213266
rect 15816 213253 15840 213266
rect 15884 213253 15908 213266
rect 15952 213253 15976 213266
rect 16020 213253 16044 213266
rect 16088 213253 16112 213266
rect 16156 213253 16180 213266
rect 16224 213253 16248 213266
rect 16292 213253 16316 213266
rect 16360 213253 16384 213266
rect 16428 213253 16452 213266
rect 16496 213253 16520 213266
rect 16564 213253 16588 213266
rect 16632 213253 16656 213266
rect 17290 213253 17314 213266
rect 17358 213253 17382 213266
rect 17426 213253 17450 213266
rect 17494 213253 17518 213266
rect 17562 213253 17586 213266
rect 17630 213253 17654 213266
rect 17698 213253 17722 213266
rect 17766 213253 17790 213266
rect 17834 213253 17858 213266
rect 17902 213253 17926 213266
rect 17970 213253 17994 213266
rect 18038 213253 18062 213266
rect 18106 213253 18130 213266
rect 18174 213253 18198 213266
rect 7389 212863 8389 212919
rect 8990 212863 9990 212919
rect 15678 212908 16678 212964
rect 17278 212908 18278 212964
rect 7389 212791 8389 212847
rect 8990 212791 9990 212847
rect 15678 212836 16678 212892
rect 17278 212836 18278 212892
rect 19480 212867 19516 219817
rect 19547 212867 19583 219817
rect 24572 219738 25172 219866
rect 36785 219864 37385 219920
rect 36785 219688 37385 219744
rect 20809 219650 20833 219684
rect 20809 219582 20833 219616
rect 24572 219588 25172 219638
rect 20809 219514 20833 219548
rect 36785 219518 37385 219568
rect 20809 219446 20833 219480
rect 24572 219458 25172 219508
rect 32930 219457 33530 219507
rect 20809 219378 20833 219412
rect 35287 219391 35887 219441
rect 36785 219402 37385 219452
rect 20809 219310 20833 219344
rect 24572 219308 25172 219358
rect 31463 219307 32063 219357
rect 32930 219301 33530 219357
rect 20809 219242 20833 219276
rect 35287 219215 35887 219343
rect 36785 219226 37385 219282
rect 20809 219174 20833 219208
rect 31463 219151 32063 219207
rect 32930 219151 33530 219201
rect 34079 219157 34679 219207
rect 20809 219106 20833 219140
rect 19844 218051 19894 219051
rect 19994 218051 20122 219051
rect 20150 218051 20278 219051
rect 20306 218051 20434 219051
rect 20462 218051 20512 219051
rect 20809 219038 20833 219072
rect 20809 218970 20833 219004
rect 20973 219000 21007 219024
rect 21041 219000 21075 219024
rect 21109 219000 21143 219024
rect 21177 219000 21211 219024
rect 21245 219000 21279 219024
rect 21313 219000 21347 219024
rect 21381 219000 21415 219024
rect 21449 219000 21483 219024
rect 21517 219000 21551 219024
rect 21585 219000 21619 219024
rect 21653 219000 21687 219024
rect 21721 219000 21755 219024
rect 21789 219000 21823 219024
rect 21857 219000 21891 219024
rect 21925 219000 21959 219024
rect 21993 219000 22027 219024
rect 22061 219000 22095 219024
rect 22129 219000 22163 219024
rect 22197 219000 22210 219024
rect 31463 219001 32063 219051
rect 34079 219001 34679 219057
rect 35287 219039 35887 219095
rect 36785 219050 37385 219106
rect 20809 218902 20833 218936
rect 32596 218929 33596 218979
rect 20809 218834 20833 218868
rect 24573 218820 25173 218870
rect 34079 218851 34679 218901
rect 35287 218869 35887 218919
rect 36785 218880 37385 218930
rect 35287 218866 35559 218869
rect 35716 218866 35887 218869
rect 20809 218766 20833 218800
rect 30171 218795 30771 218845
rect 20809 218698 20833 218732
rect 24573 218664 25173 218792
rect 32596 218773 33596 218829
rect 37993 218704 38593 218754
rect 19844 216521 19894 217921
rect 19994 216521 20122 217921
rect 20150 216521 20278 217921
rect 20306 216521 20434 217921
rect 20462 216521 20512 217921
rect 20809 216219 20833 216253
rect 19844 214759 19894 216159
rect 19994 214759 20122 216159
rect 20150 214759 20278 216159
rect 20306 214759 20434 216159
rect 20462 214759 20512 216159
rect 20809 216151 20833 216185
rect 20809 216083 20833 216117
rect 20809 216015 20833 216049
rect 20809 215947 20833 215981
rect 20809 215879 20833 215913
rect 20809 215811 20833 215845
rect 20809 215743 20833 215777
rect 20809 215675 20833 215709
rect 20809 215607 20833 215641
rect 20809 215539 20833 215573
rect 21263 215518 21313 218518
rect 21413 215518 21541 218518
rect 21569 215518 21697 218518
rect 21725 215518 21853 218518
rect 21881 215518 22009 218518
rect 22037 215518 22165 218518
rect 22193 215518 22321 218518
rect 22349 215518 22399 218518
rect 24573 218508 25173 218636
rect 30171 218619 30771 218675
rect 32596 218623 33596 218673
rect 34110 218589 34710 218639
rect 36785 218620 36797 218624
rect 36785 218609 36800 218620
rect 36970 218609 36985 218624
rect 26348 218530 26372 218564
rect 32596 218507 33596 218557
rect 26348 218461 26372 218495
rect 30171 218449 30771 218499
rect 24573 218352 25173 218408
rect 24573 218196 25173 218324
rect 29993 218310 30993 218360
rect 32596 218351 33596 218479
rect 34110 218433 34710 218561
rect 36785 218429 36985 218609
rect 37993 218534 38593 218584
rect 36785 218418 36800 218429
rect 36785 218414 36797 218418
rect 36970 218414 36985 218429
rect 31347 218317 31362 218332
rect 31535 218328 31547 218332
rect 31532 218317 31547 218328
rect 24573 218040 25173 218168
rect 26490 218122 26690 218172
rect 29993 218160 30993 218210
rect 31347 218137 31547 218317
rect 31347 218122 31362 218137
rect 31532 218126 31547 218137
rect 31535 218122 31547 218126
rect 31607 218317 31622 218332
rect 31795 218328 31807 218332
rect 31792 218317 31807 218328
rect 31607 218137 31807 218317
rect 32596 218195 33596 218323
rect 34110 218277 34710 218405
rect 36785 218384 36797 218388
rect 36785 218373 36800 218384
rect 36970 218373 36985 218388
rect 31607 218122 31622 218137
rect 31792 218126 31807 218137
rect 31795 218122 31807 218126
rect 31347 218081 31362 218096
rect 31535 218092 31547 218096
rect 31532 218081 31547 218092
rect 22906 217855 23212 218025
rect 23406 217855 23712 218025
rect 26490 217966 26690 218022
rect 29993 218001 30993 218051
rect 24573 217890 25173 217940
rect 31347 217901 31547 218081
rect 26490 217816 26690 217866
rect 29993 217851 30993 217901
rect 31347 217886 31362 217901
rect 31532 217890 31547 217901
rect 31535 217886 31547 217890
rect 31607 218081 31622 218096
rect 31795 218092 31807 218096
rect 31792 218081 31807 218092
rect 31607 217901 31807 218081
rect 32596 218039 33596 218167
rect 34110 218121 34710 218249
rect 36785 218193 36985 218373
rect 36785 218182 36800 218193
rect 36785 218178 36797 218182
rect 36970 218178 36985 218193
rect 37083 218373 37098 218388
rect 37083 218193 37120 218373
rect 37083 218178 37098 218193
rect 37998 218108 38598 218158
rect 34110 217971 34710 218021
rect 31607 217886 31622 217901
rect 31792 217890 31807 217901
rect 31795 217886 31807 217890
rect 32596 217883 33596 217939
rect 37998 217932 38598 217988
rect 34110 217855 34710 217905
rect 24573 217760 25173 217810
rect 27691 217682 28291 217732
rect 30253 217721 30268 217736
rect 30441 217732 30453 217736
rect 30438 217721 30453 217732
rect 24573 217610 25173 217660
rect 27691 217532 28291 217582
rect 30253 217541 30453 217721
rect 30253 217526 30268 217541
rect 30438 217530 30453 217541
rect 30441 217526 30453 217530
rect 30513 217721 30528 217736
rect 30701 217732 30713 217736
rect 30698 217721 30713 217732
rect 30513 217541 30713 217721
rect 30513 217526 30528 217541
rect 30698 217530 30713 217541
rect 30701 217526 30713 217530
rect 30773 217721 30788 217736
rect 30961 217732 30973 217736
rect 30958 217721 30973 217732
rect 30773 217541 30973 217721
rect 30773 217526 30788 217541
rect 30958 217530 30973 217541
rect 30961 217526 30973 217530
rect 31087 217721 31102 217736
rect 31275 217732 31287 217736
rect 31272 217721 31287 217732
rect 31087 217541 31287 217721
rect 31087 217526 31102 217541
rect 31272 217530 31287 217541
rect 31275 217526 31287 217530
rect 31347 217721 31362 217736
rect 31535 217732 31547 217736
rect 31532 217721 31547 217732
rect 31347 217541 31547 217721
rect 31347 217526 31362 217541
rect 31532 217530 31547 217541
rect 31535 217526 31547 217530
rect 31607 217721 31622 217736
rect 31795 217732 31807 217736
rect 31792 217721 31807 217732
rect 31607 217541 31807 217721
rect 31607 217526 31622 217541
rect 31792 217530 31807 217541
rect 31795 217526 31807 217530
rect 31867 217721 31882 217736
rect 32055 217732 32067 217736
rect 32052 217721 32067 217732
rect 32596 217727 33596 217855
rect 31867 217541 32067 217721
rect 34110 217699 34710 217827
rect 37998 217762 38598 217812
rect 37998 217759 38220 217762
rect 38245 217759 38539 217762
rect 32596 217571 33596 217699
rect 34110 217543 34710 217671
rect 31867 217526 31882 217541
rect 32052 217530 32067 217541
rect 32055 217526 32067 217530
rect 22619 217446 22647 217474
rect 24573 217438 25173 217488
rect 26490 217416 26690 217466
rect 27691 217402 28291 217452
rect 32596 217415 33596 217543
rect 34110 217387 34710 217515
rect 24573 217288 25173 217338
rect 26490 217260 26690 217316
rect 27691 217246 28291 217374
rect 30253 217361 30268 217376
rect 30441 217372 30453 217376
rect 30438 217361 30453 217372
rect 30253 217331 30453 217361
rect 30253 217316 30268 217331
rect 30438 217320 30453 217331
rect 30441 217316 30453 217320
rect 30513 217361 30528 217376
rect 30701 217372 30713 217376
rect 30698 217361 30713 217372
rect 30513 217331 30713 217361
rect 30513 217316 30528 217331
rect 30698 217320 30713 217331
rect 30701 217316 30713 217320
rect 30773 217361 30788 217376
rect 31347 217361 31362 217376
rect 31535 217372 31547 217376
rect 31532 217361 31547 217372
rect 30773 217331 30793 217361
rect 31347 217331 31547 217361
rect 30773 217316 30788 217331
rect 31347 217316 31362 217331
rect 31532 217320 31547 217331
rect 31535 217316 31547 217320
rect 31607 217361 31622 217376
rect 31795 217372 31807 217376
rect 31792 217361 31807 217372
rect 31607 217331 31807 217361
rect 31607 217316 31622 217331
rect 31792 217320 31807 217331
rect 31795 217316 31807 217320
rect 31867 217361 31882 217376
rect 31867 217331 31921 217361
rect 31867 217316 31882 217331
rect 30253 217275 30268 217290
rect 30441 217286 30453 217290
rect 30438 217275 30453 217286
rect 30253 217245 30453 217275
rect 30253 217230 30268 217245
rect 30438 217234 30453 217245
rect 30441 217230 30453 217234
rect 30513 217275 30528 217290
rect 30701 217286 30713 217290
rect 30698 217275 30713 217286
rect 30513 217245 30713 217275
rect 30513 217230 30528 217245
rect 30698 217234 30713 217245
rect 30701 217230 30713 217234
rect 30773 217275 30788 217290
rect 31347 217275 31362 217290
rect 31535 217286 31547 217290
rect 31532 217275 31547 217286
rect 30773 217245 30793 217275
rect 31347 217245 31547 217275
rect 30773 217230 30788 217245
rect 31347 217230 31362 217245
rect 31532 217234 31547 217245
rect 31535 217230 31547 217234
rect 31607 217275 31622 217290
rect 31795 217286 31807 217290
rect 31792 217275 31807 217286
rect 31607 217245 31807 217275
rect 31607 217230 31622 217245
rect 31792 217234 31807 217245
rect 31795 217230 31807 217234
rect 31867 217275 31882 217290
rect 31867 217245 31921 217275
rect 32596 217265 33596 217315
rect 31867 217230 31882 217245
rect 34110 217231 34710 217287
rect 22906 217055 23212 217225
rect 23406 217055 23712 217225
rect 24573 217158 25173 217208
rect 24573 217002 25173 217130
rect 26490 217107 26690 217160
rect 27691 217090 28291 217218
rect 31823 217084 32061 217118
rect 31481 217080 32061 217084
rect 31481 217068 31797 217080
rect 32596 217063 33596 217113
rect 34110 217075 34710 217203
rect 37998 217133 38148 217145
rect 38317 217133 38467 217145
rect 24573 216846 25173 216974
rect 27691 216934 28291 216990
rect 32596 216907 33596 217035
rect 34110 216919 34710 217047
rect 37998 217020 38598 217070
rect 27691 216778 28291 216906
rect 25286 216758 25310 216762
rect 32596 216751 33596 216879
rect 34110 216763 34710 216891
rect 37998 216844 38598 216900
rect 24573 216690 25173 216746
rect 25286 216687 25310 216721
rect 24573 216534 25173 216662
rect 25286 216615 25310 216649
rect 27691 216622 28291 216750
rect 32596 216595 33596 216723
rect 35287 216695 35487 216707
rect 37998 216674 38598 216724
rect 34110 216607 34710 216663
rect 36785 216650 36797 216654
rect 36785 216639 36800 216650
rect 36970 216639 36985 216654
rect 35134 216582 35734 216632
rect 25286 216543 25310 216577
rect 22906 216255 23212 216425
rect 23406 216255 23712 216425
rect 24573 216378 25173 216506
rect 25286 216471 25310 216505
rect 27691 216472 28291 216522
rect 32596 216439 33596 216567
rect 34110 216451 34710 216507
rect 35134 216432 35734 216482
rect 36785 216459 36985 216639
rect 36785 216448 36800 216459
rect 36785 216444 36797 216448
rect 36970 216444 36985 216459
rect 37083 216639 37098 216654
rect 37083 216459 37120 216639
rect 37083 216444 37098 216459
rect 36785 216414 36797 216418
rect 32596 216283 33596 216411
rect 36785 216403 36800 216414
rect 36970 216403 36985 216418
rect 34110 216295 34710 216351
rect 35134 216316 35734 216366
rect 24573 216228 25173 216278
rect 32596 216127 33596 216255
rect 34110 216145 34710 216195
rect 35134 216160 35734 216288
rect 32596 215971 33596 216099
rect 34110 216029 34710 216079
rect 35134 216004 35734 216132
rect 31481 215862 31797 215880
rect 34110 215873 34710 216001
rect 31823 215828 32061 215860
rect 32596 215821 33596 215871
rect 35134 215848 35734 215976
rect 36071 215805 36098 216295
rect 36785 216223 36985 216403
rect 37993 216248 38593 216298
rect 36785 216212 36800 216223
rect 36785 216208 36797 216212
rect 36970 216208 36985 216223
rect 696597 216200 696600 216320
rect 37993 216078 38593 216128
rect 692376 215983 692396 216017
rect 692463 215993 692532 216017
rect 696191 215993 696239 216017
rect 692487 215983 692532 215993
rect 696204 215983 696239 215993
rect 696340 215983 696360 216017
rect 36785 215902 37385 215952
rect 692487 215915 692502 215939
rect 696200 215915 696215 215939
rect 692454 215891 692478 215915
rect 696224 215891 696248 215915
rect 686755 215800 687355 215850
rect 34110 215717 34710 215773
rect 30253 215701 30268 215716
rect 30441 215712 30453 215716
rect 30438 215701 30453 215712
rect 30253 215671 30453 215701
rect 30253 215656 30268 215671
rect 30438 215660 30453 215671
rect 30441 215656 30453 215660
rect 30513 215701 30528 215716
rect 30701 215712 30713 215716
rect 30698 215701 30713 215712
rect 30513 215671 30713 215701
rect 30513 215656 30528 215671
rect 30698 215660 30713 215671
rect 30701 215656 30713 215660
rect 30773 215701 30788 215716
rect 31347 215701 31362 215716
rect 31535 215712 31547 215716
rect 31532 215701 31547 215712
rect 30773 215671 30793 215701
rect 31347 215671 31547 215701
rect 30773 215656 30788 215671
rect 31347 215656 31362 215671
rect 31532 215660 31547 215671
rect 31535 215656 31547 215660
rect 31607 215701 31622 215716
rect 31795 215712 31807 215716
rect 31792 215701 31807 215712
rect 31607 215671 31807 215701
rect 31607 215656 31622 215671
rect 31792 215660 31807 215671
rect 31795 215656 31807 215660
rect 31867 215701 31882 215716
rect 31867 215671 31921 215701
rect 35134 215698 35734 215770
rect 36785 215726 37385 215782
rect 692487 215748 692505 215752
rect 692479 215718 692505 215748
rect 692487 215698 692505 215718
rect 31867 215656 31882 215671
rect 30253 215615 30268 215630
rect 30441 215626 30453 215630
rect 30438 215615 30453 215626
rect 30253 215585 30453 215615
rect 30253 215570 30268 215585
rect 30438 215574 30453 215585
rect 30441 215570 30453 215574
rect 30513 215615 30528 215630
rect 30701 215626 30713 215630
rect 30698 215615 30713 215626
rect 30513 215585 30713 215615
rect 30513 215570 30528 215585
rect 30698 215574 30713 215585
rect 30701 215570 30713 215574
rect 30773 215615 30788 215630
rect 31347 215615 31362 215630
rect 31535 215626 31547 215630
rect 31532 215615 31547 215626
rect 30773 215585 30793 215615
rect 31347 215585 31547 215615
rect 30773 215570 30788 215585
rect 31347 215570 31362 215585
rect 31532 215574 31547 215585
rect 31535 215570 31547 215574
rect 31607 215615 31622 215630
rect 31795 215626 31807 215630
rect 31792 215615 31807 215626
rect 31607 215585 31807 215615
rect 31607 215570 31622 215585
rect 31792 215574 31807 215585
rect 31795 215570 31807 215574
rect 31867 215615 31882 215630
rect 32546 215619 33546 215669
rect 31867 215585 31921 215615
rect 31867 215570 31882 215585
rect 20809 215471 20833 215505
rect 32546 215463 33546 215591
rect 34110 215561 34710 215689
rect 35134 215645 36134 215695
rect 686755 215624 687355 215680
rect 692485 215674 692505 215698
rect 692509 215674 692517 215718
rect 696215 215698 696223 215748
rect 696203 215674 696223 215698
rect 696227 215674 696245 215752
rect 692485 215640 692521 215674
rect 696203 215640 696249 215674
rect 35134 215489 36134 215617
rect 36785 215550 37385 215606
rect 20809 215403 20833 215437
rect 30253 215405 30268 215420
rect 30441 215416 30453 215420
rect 30438 215405 30453 215416
rect 20809 215335 20833 215369
rect 20809 215267 20833 215301
rect 20809 215199 20833 215233
rect 30253 215225 30453 215405
rect 30253 215210 30268 215225
rect 30438 215214 30453 215225
rect 30441 215210 30453 215214
rect 30513 215405 30528 215420
rect 30701 215416 30713 215420
rect 30698 215405 30713 215416
rect 30513 215225 30713 215405
rect 30513 215210 30528 215225
rect 30698 215214 30713 215225
rect 30701 215210 30713 215214
rect 30773 215405 30788 215420
rect 30961 215416 30973 215420
rect 30958 215405 30973 215416
rect 30773 215225 30973 215405
rect 30773 215210 30788 215225
rect 30958 215214 30973 215225
rect 30961 215210 30973 215214
rect 31087 215405 31102 215420
rect 31275 215416 31287 215420
rect 31272 215405 31287 215416
rect 31087 215225 31287 215405
rect 31087 215210 31102 215225
rect 31272 215214 31287 215225
rect 31275 215210 31287 215214
rect 31347 215405 31362 215420
rect 31535 215416 31547 215420
rect 31532 215405 31547 215416
rect 31347 215225 31547 215405
rect 31347 215210 31362 215225
rect 31532 215214 31547 215225
rect 31535 215210 31547 215214
rect 31607 215405 31622 215420
rect 31795 215416 31807 215420
rect 31792 215405 31807 215416
rect 31607 215225 31807 215405
rect 31607 215210 31622 215225
rect 31792 215214 31807 215225
rect 31795 215210 31807 215214
rect 31867 215405 31882 215420
rect 32055 215416 32067 215420
rect 32052 215405 32067 215416
rect 31867 215225 32067 215405
rect 32546 215307 33546 215435
rect 34110 215411 34710 215461
rect 686755 215448 687355 215504
rect 35134 215339 36134 215389
rect 36785 215380 37385 215430
rect 31867 215210 31882 215225
rect 32052 215214 32067 215225
rect 32055 215210 32067 215214
rect 20809 215131 20833 215165
rect 32546 215151 33546 215279
rect 36785 215248 37385 215298
rect 686755 215278 687355 215328
rect 35285 215162 35319 215172
rect 35353 215162 35387 215172
rect 35421 215162 35455 215172
rect 35489 215162 35523 215172
rect 35564 215162 35598 215172
rect 35632 215162 35666 215172
rect 35700 215162 35734 215172
rect 35768 215162 35802 215172
rect 35836 215162 35870 215172
rect 35904 215162 35938 215172
rect 35972 215162 36006 215172
rect 36040 215162 36074 215172
rect 36108 215162 36142 215172
rect 36176 215162 36210 215172
rect 35255 215126 36255 215138
rect 20809 215063 20833 215097
rect 20940 215085 20983 215103
rect 20940 215069 20949 215085
rect 20974 215069 20983 215085
rect 25113 215069 25349 215093
rect 25383 215069 25417 215093
rect 20974 215051 21008 215069
rect 20809 214995 20833 215029
rect 20974 215028 21003 215051
rect 21361 215045 21409 215069
rect 20949 215027 20983 215028
rect 21385 214991 21409 215045
rect 25113 214991 25137 215069
rect 29993 215045 30993 215095
rect 31347 215045 31362 215060
rect 31535 215056 31547 215060
rect 31532 215045 31547 215056
rect 21361 214967 21409 214991
rect 25089 214967 25137 214991
rect 20809 214927 20833 214961
rect 20809 214859 20833 214893
rect 20809 214791 20833 214825
rect 20809 214723 20833 214757
rect 20809 214655 20833 214689
rect 21413 214638 22813 214681
rect 23685 214638 25085 214681
rect 19844 213229 19894 214629
rect 19994 213229 20122 214629
rect 20150 213229 20278 214629
rect 20306 213229 20434 214629
rect 20462 213229 20512 214629
rect 20809 214587 20833 214621
rect 20809 214519 20833 214553
rect 20809 214451 20833 214485
rect 21413 214475 22813 214603
rect 23685 214475 25085 214603
rect 20809 214383 20833 214417
rect 20809 214315 20833 214349
rect 21413 214312 22813 214440
rect 23685 214312 25085 214440
rect 20809 214247 20833 214281
rect 20809 214179 20833 214213
rect 21413 214149 22813 214277
rect 23685 214149 25085 214277
rect 20809 214111 20833 214145
rect 20809 214043 20833 214077
rect 20809 213975 20833 214009
rect 21413 213986 22813 214114
rect 23685 213986 25085 214114
rect 20809 213907 20833 213941
rect 20809 213839 20833 213873
rect 21413 213823 22813 213951
rect 23685 213823 25085 213951
rect 20809 213771 20833 213805
rect 20809 213703 20833 213737
rect 21413 213673 22813 213716
rect 23685 213673 25085 213716
rect 20809 213635 20833 213669
rect 20809 213567 20833 213601
rect 21361 213552 21419 213586
rect 25089 213552 25147 213586
rect 20809 213499 20833 213533
rect 20809 213431 20833 213465
rect 20809 213363 20833 213397
rect 21361 213373 21419 213397
rect 25089 213373 25147 213397
rect 21385 213363 21419 213373
rect 25113 213363 25147 213373
rect 20809 213295 20833 213329
rect 21385 213291 21419 213325
rect 25113 213291 25147 213325
rect 20809 213227 20833 213261
rect 21385 213219 21419 213253
rect 25113 213219 25147 213253
rect 20809 213159 20833 213193
rect 21385 213171 21419 213181
rect 25113 213171 25147 213181
rect 21361 213147 21419 213171
rect 25089 213147 25147 213171
rect 20809 213091 20833 213125
rect 20809 213023 20833 213057
rect 20809 212955 20833 212989
rect 21361 212969 21409 212993
rect 25089 212969 25137 212993
rect 20809 212887 20833 212921
rect 21385 212915 21409 212969
rect 25113 212915 25137 212969
rect 21361 212891 21409 212915
rect 25089 212891 25137 212915
rect 19480 212831 19583 212867
rect 21413 212754 22813 212804
rect 23685 212754 25085 212804
rect 7389 212489 8389 212561
rect 8990 212489 9990 212561
rect 15678 212534 16678 212606
rect 17278 212534 18278 212606
rect 21413 212591 22813 212719
rect 23685 212591 25085 212719
rect 15748 212523 15782 212534
rect 15816 212523 15850 212534
rect 15884 212523 15918 212534
rect 15952 212523 15986 212534
rect 16020 212523 16054 212534
rect 16088 212523 16122 212534
rect 16156 212523 16190 212534
rect 16224 212523 16258 212534
rect 16292 212523 16326 212534
rect 16360 212523 16394 212534
rect 16428 212523 16462 212534
rect 16496 212523 16530 212534
rect 16564 212523 16598 212534
rect 16632 212523 16666 212534
rect 17290 212523 17324 212534
rect 17358 212523 17392 212534
rect 17426 212523 17460 212534
rect 17494 212523 17528 212534
rect 17562 212523 17596 212534
rect 17630 212523 17664 212534
rect 17698 212523 17732 212534
rect 17766 212523 17800 212534
rect 17834 212523 17868 212534
rect 17902 212523 17936 212534
rect 17970 212523 18004 212534
rect 18038 212523 18072 212534
rect 18106 212523 18140 212534
rect 18174 212523 18208 212534
rect 15748 212513 15806 212523
rect 15816 212513 15874 212523
rect 15884 212513 15942 212523
rect 15952 212513 16010 212523
rect 16020 212513 16078 212523
rect 16088 212513 16146 212523
rect 16156 212513 16214 212523
rect 16224 212513 16282 212523
rect 16292 212513 16350 212523
rect 16360 212513 16418 212523
rect 16428 212513 16486 212523
rect 16496 212513 16554 212523
rect 16564 212513 16622 212523
rect 16632 212513 16690 212523
rect 17290 212513 17348 212523
rect 17358 212513 17416 212523
rect 17426 212513 17484 212523
rect 17494 212513 17552 212523
rect 17562 212513 17620 212523
rect 17630 212513 17688 212523
rect 17698 212513 17756 212523
rect 17766 212513 17824 212523
rect 17834 212513 17892 212523
rect 17902 212513 17960 212523
rect 17970 212513 18028 212523
rect 18038 212513 18096 212523
rect 18106 212513 18164 212523
rect 18174 212513 18232 212523
rect 15724 212489 16690 212513
rect 17266 212489 18232 212513
rect 15748 212474 15772 212489
rect 15816 212474 15840 212489
rect 15884 212474 15908 212489
rect 15952 212474 15976 212489
rect 16020 212474 16044 212489
rect 16088 212474 16112 212489
rect 16156 212474 16180 212489
rect 16224 212474 16248 212489
rect 16292 212474 16316 212489
rect 16360 212474 16384 212489
rect 16428 212474 16452 212489
rect 16496 212474 16520 212489
rect 16564 212474 16588 212489
rect 16632 212474 16656 212489
rect 17290 212474 17314 212489
rect 17358 212474 17382 212489
rect 17426 212474 17450 212489
rect 17494 212474 17518 212489
rect 17562 212474 17586 212489
rect 17630 212474 17654 212489
rect 17698 212474 17722 212489
rect 17766 212474 17790 212489
rect 17834 212474 17858 212489
rect 17902 212474 17926 212489
rect 17970 212474 17994 212489
rect 18038 212474 18062 212489
rect 18106 212474 18130 212489
rect 18174 212474 18198 212489
rect 15678 212319 16678 212474
rect 7389 212229 8389 212289
rect 8990 212229 9990 212289
rect 15678 212285 16690 212319
rect 17278 212309 18278 212474
rect 21413 212428 22813 212556
rect 23685 212428 25085 212556
rect 17266 212285 18278 212309
rect 15678 212274 16678 212285
rect 17278 212274 18278 212285
rect 15748 212261 15772 212274
rect 15816 212261 15840 212274
rect 15884 212261 15908 212274
rect 15952 212261 15976 212274
rect 16020 212261 16044 212274
rect 16088 212261 16112 212274
rect 16156 212261 16180 212274
rect 16224 212261 16248 212274
rect 16292 212261 16316 212274
rect 16360 212261 16384 212274
rect 16428 212261 16452 212274
rect 16496 212261 16520 212274
rect 16564 212261 16588 212274
rect 16632 212261 16656 212274
rect 17290 212261 17314 212274
rect 17358 212261 17382 212274
rect 17426 212261 17450 212274
rect 17494 212261 17518 212274
rect 17562 212261 17586 212274
rect 17630 212261 17654 212274
rect 17698 212261 17722 212274
rect 17766 212261 17790 212274
rect 17834 212261 17858 212274
rect 17902 212261 17926 212274
rect 17970 212261 17994 212274
rect 18038 212261 18062 212274
rect 18106 212261 18130 212274
rect 18174 212261 18198 212274
rect 21413 212265 22813 212393
rect 23685 212265 25085 212393
rect 21413 212102 22813 212230
rect 23685 212102 25085 212230
rect 7389 211871 8389 211927
rect 8990 211871 9990 211927
rect 15678 211916 16678 211972
rect 17278 211916 18278 211972
rect 21413 211952 22813 211995
rect 23685 211952 25085 211995
rect 7389 211799 8389 211855
rect 8990 211799 9990 211855
rect 15678 211844 16678 211900
rect 17278 211844 18278 211900
rect 21406 211865 21430 211889
rect 25068 211865 25092 211889
rect 21382 211841 21385 211865
rect 25113 211841 25116 211865
rect 21382 211763 21396 211787
rect 25102 211763 25116 211787
rect 21348 211739 21372 211763
rect 21406 211739 21430 211763
rect 25068 211739 25092 211763
rect 25126 211739 25150 211763
rect 25524 211703 25548 215001
rect 29993 214895 30993 214945
rect 31347 214865 31547 215045
rect 31347 214850 31362 214865
rect 31532 214854 31547 214865
rect 31535 214850 31547 214854
rect 31607 215045 31622 215060
rect 31795 215056 31807 215060
rect 31792 215045 31807 215056
rect 31607 214865 31807 215045
rect 32546 214995 33546 215123
rect 36785 215072 37385 215128
rect 685547 215102 686147 215152
rect 35255 215019 36255 215069
rect 687155 215007 687170 215022
rect 687343 215018 687355 215022
rect 687340 215007 687355 215018
rect 31607 214850 31622 214865
rect 31792 214854 31807 214865
rect 31795 214850 31807 214854
rect 32546 214839 33546 214967
rect 35255 214843 36255 214971
rect 36785 214896 37385 214952
rect 685547 214932 686147 214982
rect 687155 214827 687355 215007
rect 31347 214809 31362 214824
rect 31535 214820 31547 214824
rect 31532 214809 31547 214820
rect 29993 214736 30993 214786
rect 29993 214586 30993 214636
rect 31347 214629 31547 214809
rect 31347 214614 31362 214629
rect 31532 214618 31547 214629
rect 31535 214614 31547 214618
rect 31607 214809 31622 214824
rect 31795 214820 31807 214824
rect 31792 214809 31807 214820
rect 687155 214812 687170 214827
rect 687340 214816 687355 214827
rect 687343 214812 687355 214816
rect 31607 214629 31807 214809
rect 32546 214683 33546 214811
rect 35255 214667 36255 214795
rect 36785 214726 37385 214776
rect 687042 214771 687057 214786
rect 31607 214614 31622 214629
rect 31792 214618 31807 214629
rect 31795 214614 31807 214618
rect 32546 214527 33546 214655
rect 37993 214550 38593 214600
rect 687020 214591 687057 214771
rect 687155 214771 687170 214786
rect 687343 214782 687355 214786
rect 687340 214771 687355 214782
rect 687155 214591 687355 214771
rect 688210 214630 688260 215630
rect 688360 214740 688488 215630
rect 688516 214740 688644 215630
rect 688672 214740 688800 215630
rect 688828 214740 688956 215630
rect 688984 214740 689112 215630
rect 689140 214740 689268 215630
rect 689296 214740 689424 215630
rect 689452 214740 689580 215630
rect 689608 214740 689736 215630
rect 689764 214740 689892 215630
rect 689920 214740 690048 215630
rect 690076 214740 690204 215630
rect 690232 214740 690360 215630
rect 690388 214630 690438 215630
rect 692485 215606 692505 215640
rect 692509 215606 692517 215640
rect 696203 215606 696223 215640
rect 696227 215606 696245 215640
rect 691275 215523 691875 215573
rect 692485 215572 692521 215606
rect 696203 215572 696249 215606
rect 692485 215538 692505 215572
rect 692509 215538 692517 215572
rect 692485 215504 692521 215538
rect 692583 215528 693983 215571
rect 694719 215528 696119 215571
rect 696203 215538 696223 215572
rect 696227 215538 696245 215572
rect 696203 215504 696249 215538
rect 692485 215470 692505 215504
rect 692509 215470 692517 215504
rect 692485 215436 692521 215470
rect 691275 215373 691875 215423
rect 692485 215402 692505 215436
rect 692509 215402 692517 215436
rect 692485 215368 692521 215402
rect 692485 215334 692505 215368
rect 692509 215334 692517 215368
rect 692583 215365 693983 215493
rect 694719 215365 696119 215493
rect 696203 215470 696223 215504
rect 696227 215470 696245 215504
rect 696203 215436 696249 215470
rect 707624 215441 707658 215475
rect 707695 215441 707729 215475
rect 707769 215441 707803 215475
rect 707840 215441 707874 215475
rect 707914 215441 707948 215475
rect 707985 215441 708019 215475
rect 708059 215441 708093 215475
rect 708130 215441 708164 215475
rect 708204 215441 708238 215475
rect 708275 215441 708309 215475
rect 708369 215441 708403 215475
rect 708446 215441 708480 215475
rect 708520 215441 708554 215465
rect 708588 215441 708610 215465
rect 709211 215441 709234 215465
rect 709270 215441 709304 215475
rect 709364 215441 709398 215475
rect 709435 215441 709469 215475
rect 709509 215441 709543 215475
rect 709580 215441 709614 215475
rect 709654 215441 709688 215475
rect 709725 215441 709759 215475
rect 709799 215441 709833 215475
rect 709870 215441 709904 215475
rect 709944 215441 709978 215475
rect 710015 215441 710049 215475
rect 710089 215441 710123 215475
rect 710160 215441 710194 215475
rect 696203 215402 696223 215436
rect 696227 215402 696245 215436
rect 707610 215431 707624 215441
rect 707658 215431 707695 215441
rect 707729 215431 707769 215441
rect 707803 215431 707840 215441
rect 707874 215431 707914 215441
rect 707948 215431 707985 215441
rect 708019 215431 708059 215441
rect 708093 215431 708130 215441
rect 708164 215431 708204 215441
rect 708238 215431 708275 215441
rect 708309 215431 708369 215441
rect 708403 215431 708446 215441
rect 708480 215431 708520 215441
rect 708554 215431 708588 215441
rect 708610 215431 708634 215441
rect 709211 215431 709270 215441
rect 709304 215431 709364 215441
rect 709398 215431 709435 215441
rect 709469 215431 709509 215441
rect 709543 215431 709580 215441
rect 709614 215431 709654 215441
rect 709688 215431 709725 215441
rect 709759 215431 709799 215441
rect 709833 215431 709870 215441
rect 709904 215431 709944 215441
rect 709978 215431 710015 215441
rect 710049 215431 710089 215441
rect 710123 215431 710160 215441
rect 710194 215431 710211 215441
rect 696203 215368 696249 215402
rect 696203 215334 696223 215368
rect 696227 215334 696245 215368
rect 707610 215337 708610 215431
rect 709211 215337 710211 215431
rect 691275 215251 691875 215301
rect 692485 215300 692521 215334
rect 692485 215266 692505 215300
rect 692509 215266 692517 215300
rect 692485 215232 692521 215266
rect 692485 215198 692505 215232
rect 692509 215198 692517 215232
rect 692583 215202 693983 215330
rect 694719 215202 696119 215330
rect 696203 215300 696249 215334
rect 711579 215317 712463 215331
rect 711579 215307 711619 215317
rect 696203 215266 696223 215300
rect 696227 215266 696245 215300
rect 701730 215290 701747 215292
rect 696203 215232 696249 215266
rect 696203 215198 696223 215232
rect 696227 215198 696245 215232
rect 701692 215220 701722 215254
rect 701730 215220 701760 215290
rect 707610 215241 708610 215301
rect 709211 215241 710211 215301
rect 692485 215164 692521 215198
rect 691275 215101 691875 215151
rect 692485 215130 692505 215164
rect 692509 215130 692517 215164
rect 692485 215096 692521 215130
rect 692485 215062 692505 215096
rect 692509 215062 692517 215096
rect 692485 215028 692521 215062
rect 692583 215039 693983 215167
rect 694719 215039 696119 215167
rect 696203 215164 696249 215198
rect 696203 215130 696223 215164
rect 696227 215130 696245 215164
rect 696203 215096 696249 215130
rect 696203 215062 696223 215096
rect 696227 215062 696245 215096
rect 699322 215064 700322 215097
rect 700922 215064 701922 215097
rect 696203 215028 696249 215062
rect 707610 215044 708610 215048
rect 709211 215044 710211 215048
rect 691275 214975 691875 215025
rect 692485 214994 692505 215028
rect 692509 214994 692517 215028
rect 692485 214960 692521 214994
rect 692485 214926 692505 214960
rect 692509 214926 692517 214960
rect 692485 214892 692521 214926
rect 691275 214825 691875 214875
rect 692485 214858 692505 214892
rect 692509 214858 692517 214892
rect 692583 214876 693983 215004
rect 694719 214876 696119 215004
rect 696203 214994 696223 215028
rect 696227 214994 696245 215028
rect 707574 214994 708646 215030
rect 696203 214960 696249 214994
rect 696203 214926 696223 214960
rect 696227 214926 696245 214960
rect 707574 214953 707610 214994
rect 708610 214953 708646 214994
rect 696203 214892 696249 214926
rect 697284 214894 697350 214910
rect 707574 214897 708646 214953
rect 696203 214858 696223 214892
rect 696227 214858 696245 214892
rect 699322 214877 700322 214894
rect 700922 214877 701922 214894
rect 707574 214881 707610 214897
rect 708610 214881 708646 214897
rect 692485 214824 692521 214858
rect 692485 214790 692505 214824
rect 692509 214790 692517 214824
rect 692485 214756 692521 214790
rect 691275 214703 691875 214753
rect 692485 214740 692505 214756
rect 692509 214740 692517 214756
rect 692583 214740 693983 214841
rect 694719 214740 696119 214841
rect 696203 214824 696249 214858
rect 707574 214825 708646 214881
rect 696203 214790 696223 214824
rect 696227 214790 696245 214824
rect 696203 214756 696249 214790
rect 696203 214740 696223 214756
rect 696227 214740 696245 214756
rect 699322 214740 700322 214811
rect 700922 214740 701922 214811
rect 707574 214788 707610 214825
rect 708610 214788 708646 214825
rect 707574 214748 708646 214788
rect 709175 214994 710247 215030
rect 709175 214953 709211 214994
rect 710211 214953 710247 214994
rect 709175 214897 710247 214953
rect 709175 214881 709211 214897
rect 710211 214881 710247 214897
rect 709175 214825 710247 214881
rect 709175 214788 709211 214825
rect 710211 214788 710247 214825
rect 709175 214748 710247 214788
rect 28647 214450 28671 214477
rect 30171 214447 30771 214497
rect 35255 214491 36255 214547
rect 685542 214506 686142 214556
rect 691275 214553 691875 214603
rect 36785 214466 36797 214470
rect 36785 214455 36800 214466
rect 36970 214455 36985 214470
rect 28683 214397 28717 214431
rect 32546 214377 33546 214427
rect 28683 214328 28717 214362
rect 28683 214259 28717 214293
rect 30171 214271 30771 214327
rect 35255 214321 36255 214371
rect 36785 214275 36985 214455
rect 37993 214380 38593 214430
rect 685542 214330 686142 214386
rect 36785 214264 36800 214275
rect 36785 214260 36797 214264
rect 36970 214260 36985 214275
rect 692583 214237 693983 214280
rect 694719 214237 696119 214280
rect 699322 214278 700322 214418
rect 700922 214278 701922 214418
rect 36785 214230 36797 214234
rect 28683 214190 28717 214224
rect 32596 214175 33596 214225
rect 35359 214156 35375 214222
rect 36143 214156 36159 214222
rect 36785 214219 36800 214230
rect 36970 214219 36985 214234
rect 28683 214121 28717 214155
rect 30171 214101 30771 214151
rect 28683 214052 28717 214086
rect 32596 214019 33596 214147
rect 28683 213983 28717 214017
rect 33959 213994 33975 214060
rect 36143 213994 36159 214060
rect 36785 214039 36985 214219
rect 36785 214028 36800 214039
rect 36785 214024 36797 214028
rect 36970 214024 36985 214039
rect 37083 214219 37098 214234
rect 37083 214039 37120 214219
rect 685542 214160 686142 214210
rect 692583 214101 693983 214144
rect 694719 214101 696119 214144
rect 37083 214024 37098 214039
rect 28683 213914 28717 213948
rect 31463 213895 32063 213945
rect 28683 213845 28717 213879
rect 32596 213863 33596 213991
rect 37998 213954 38598 214004
rect 28683 213776 28717 213810
rect 28683 213707 28717 213741
rect 31463 213739 32063 213795
rect 32596 213707 33596 213835
rect 33959 213832 33975 213898
rect 36143 213832 36159 213898
rect 37998 213778 38598 213834
rect 28683 213638 28717 213672
rect 28683 213569 28717 213603
rect 31463 213589 32063 213639
rect 32596 213551 33596 213679
rect 35359 213670 35375 213736
rect 36143 213670 36159 213736
rect 680215 213678 680815 213728
rect 37998 213608 38598 213658
rect 37998 213605 38220 213608
rect 38245 213605 38539 213608
rect 28683 213500 28717 213534
rect 28683 213431 28717 213465
rect 28683 213362 28717 213396
rect 32596 213395 33596 213523
rect 35255 213521 36255 213571
rect 680215 213502 680815 213558
rect 685551 213516 686551 213566
rect 689154 213480 689204 213897
rect 689304 213480 689360 213897
rect 689460 213480 689516 213897
rect 689616 213480 689672 213897
rect 689772 213480 689828 213897
rect 689928 213480 689978 213897
rect 699322 213860 700322 213916
rect 700922 213860 701922 213916
rect 707610 213905 708610 213961
rect 709211 213905 710211 213961
rect 699322 213788 700322 213844
rect 700922 213788 701922 213844
rect 707610 213833 708610 213889
rect 709211 213833 710211 213889
rect 711579 213525 711605 215307
rect 715956 214297 716006 215297
rect 716106 214740 716234 215297
rect 716262 214297 716312 215297
rect 711579 213480 711595 213495
rect 712409 213480 712431 213485
rect 713640 213480 713641 213785
rect 713750 213772 714750 213822
rect 713750 213562 714750 213612
rect 713750 213480 714750 213496
rect 28683 213293 28717 213327
rect 28683 213224 28717 213258
rect 30015 213256 30718 213272
rect 30015 213246 30721 213256
rect 28683 213155 28717 213189
rect 28683 213086 28717 213120
rect 28683 213017 28717 213051
rect 28683 212948 28717 212982
rect 28683 212879 28717 212913
rect 28683 212810 28717 212844
rect 28683 212741 28717 212775
rect 28683 212672 28717 212706
rect 28683 212603 28717 212637
rect 28683 212534 28717 212568
rect 28683 212465 28717 212499
rect 28683 212396 28717 212430
rect 28682 212361 28683 212366
rect 28682 212332 28717 212361
rect 28647 212303 28671 212332
rect 28647 212234 28671 212268
rect 28647 212165 28671 212199
rect 28647 212096 28671 212130
rect 28647 212027 28671 212061
rect 28647 211958 28671 211992
rect 28647 211889 28671 211923
rect 28647 211820 28671 211854
rect 28647 211751 28671 211785
rect 28647 211682 28671 211716
rect 29778 211695 29802 211719
rect 29802 211671 29826 211683
rect 29880 211681 29914 211715
rect 25524 211635 25548 211669
rect 7389 211497 8389 211569
rect 8990 211497 9990 211569
rect 15678 211542 16678 211614
rect 17278 211542 18278 211614
rect 28647 211613 28671 211647
rect 29778 211635 29802 211659
rect 21361 211586 21409 211610
rect 25089 211586 25137 211610
rect 15748 211531 15782 211542
rect 15816 211531 15850 211542
rect 15884 211531 15918 211542
rect 15952 211531 15986 211542
rect 16020 211531 16054 211542
rect 16088 211531 16122 211542
rect 16156 211531 16190 211542
rect 16224 211531 16258 211542
rect 16292 211531 16326 211542
rect 16360 211531 16394 211542
rect 16428 211531 16462 211542
rect 16496 211531 16530 211542
rect 16564 211531 16598 211542
rect 16632 211531 16666 211542
rect 17290 211531 17324 211542
rect 17358 211531 17392 211542
rect 17426 211531 17460 211542
rect 17494 211531 17528 211542
rect 17562 211531 17596 211542
rect 17630 211531 17664 211542
rect 17698 211531 17732 211542
rect 17766 211531 17800 211542
rect 17834 211531 17868 211542
rect 17902 211531 17936 211542
rect 17970 211531 18004 211542
rect 18038 211531 18072 211542
rect 18106 211531 18140 211542
rect 18174 211531 18208 211542
rect 21385 211532 21409 211586
rect 25113 211532 25137 211586
rect 28647 211544 28671 211578
rect 15748 211521 15806 211531
rect 15816 211521 15874 211531
rect 15884 211521 15942 211531
rect 15952 211521 16010 211531
rect 16020 211521 16078 211531
rect 16088 211521 16146 211531
rect 16156 211521 16214 211531
rect 16224 211521 16282 211531
rect 16292 211521 16350 211531
rect 16360 211521 16418 211531
rect 16428 211521 16486 211531
rect 16496 211521 16554 211531
rect 16564 211521 16622 211531
rect 16632 211521 16690 211531
rect 17290 211521 17348 211531
rect 17358 211521 17416 211531
rect 17426 211521 17484 211531
rect 17494 211521 17552 211531
rect 17562 211521 17620 211531
rect 17630 211521 17688 211531
rect 17698 211521 17756 211531
rect 17766 211521 17824 211531
rect 17834 211521 17892 211531
rect 17902 211521 17960 211531
rect 17970 211521 18028 211531
rect 18038 211521 18096 211531
rect 18106 211521 18164 211531
rect 18174 211521 18232 211531
rect 15724 211497 16690 211521
rect 17266 211497 18232 211521
rect 21361 211508 21409 211532
rect 25089 211508 25137 211532
rect 15748 211482 15772 211497
rect 15816 211482 15840 211497
rect 15884 211482 15908 211497
rect 15952 211482 15976 211497
rect 16020 211482 16044 211497
rect 16088 211482 16112 211497
rect 16156 211482 16180 211497
rect 16224 211482 16248 211497
rect 16292 211482 16316 211497
rect 16360 211482 16384 211497
rect 16428 211482 16452 211497
rect 16496 211482 16520 211497
rect 16564 211482 16588 211497
rect 16632 211482 16656 211497
rect 17290 211482 17314 211497
rect 17358 211482 17382 211497
rect 17426 211482 17450 211497
rect 17494 211482 17518 211497
rect 17562 211482 17586 211497
rect 17630 211482 17654 211497
rect 17698 211482 17722 211497
rect 17766 211482 17790 211497
rect 17834 211482 17858 211497
rect 17902 211482 17926 211497
rect 17970 211482 17994 211497
rect 18038 211482 18062 211497
rect 18106 211482 18130 211497
rect 18174 211482 18198 211497
rect 7389 211237 8389 211297
rect 8990 211237 9990 211297
rect 12559 211273 12865 211375
rect 15678 211327 16678 211482
rect 15678 211293 16690 211327
rect 17278 211317 18278 211482
rect 28647 211475 28671 211509
rect 28647 211406 28671 211440
rect 28647 211337 28671 211371
rect 17266 211293 18278 211317
rect 15678 211282 16678 211293
rect 17278 211282 18278 211293
rect 12543 211257 12881 211273
rect 15748 211269 15772 211282
rect 15816 211269 15840 211282
rect 15884 211269 15908 211282
rect 15952 211269 15976 211282
rect 16020 211269 16044 211282
rect 16088 211269 16112 211282
rect 16156 211269 16180 211282
rect 16224 211269 16248 211282
rect 16292 211269 16316 211282
rect 16360 211269 16384 211282
rect 16428 211269 16452 211282
rect 16496 211269 16520 211282
rect 16564 211269 16588 211282
rect 16632 211269 16656 211282
rect 17290 211269 17314 211282
rect 17358 211269 17382 211282
rect 17426 211269 17450 211282
rect 17494 211269 17518 211282
rect 17562 211269 17586 211282
rect 17630 211269 17654 211282
rect 17698 211269 17722 211282
rect 17766 211269 17790 211282
rect 17834 211269 17858 211282
rect 17902 211269 17926 211282
rect 17970 211269 17994 211282
rect 18038 211269 18062 211282
rect 18106 211269 18130 211282
rect 18174 211269 18198 211282
rect 19980 211048 20286 211218
rect 7389 210879 8389 210935
rect 8990 210879 9990 210935
rect 15678 210924 16678 210980
rect 17278 210924 18278 210980
rect 7389 210807 8389 210863
rect 8990 210807 9990 210863
rect 15678 210852 16678 210908
rect 17278 210852 18278 210908
rect 20945 210796 25553 211332
rect 28647 211268 28671 211302
rect 28647 211199 28671 211233
rect 28647 211154 28671 211164
rect 21413 210706 22813 210796
rect 23685 210706 25085 210796
rect 7389 210505 8389 210577
rect 8990 210505 9990 210577
rect 15678 210550 16678 210622
rect 17278 210550 18278 210622
rect 15748 210539 15782 210550
rect 15816 210539 15850 210550
rect 15884 210539 15918 210550
rect 15952 210539 15986 210550
rect 16020 210539 16054 210550
rect 16088 210539 16122 210550
rect 16156 210539 16190 210550
rect 16224 210539 16258 210550
rect 16292 210539 16326 210550
rect 16360 210539 16394 210550
rect 16428 210539 16462 210550
rect 16496 210539 16530 210550
rect 16564 210539 16598 210550
rect 16632 210539 16666 210550
rect 17290 210539 17324 210550
rect 17358 210539 17392 210550
rect 17426 210539 17460 210550
rect 17494 210539 17528 210550
rect 17562 210539 17596 210550
rect 17630 210539 17664 210550
rect 17698 210539 17732 210550
rect 17766 210539 17800 210550
rect 17834 210539 17868 210550
rect 17902 210539 17936 210550
rect 17970 210539 18004 210550
rect 18038 210539 18072 210550
rect 18106 210539 18140 210550
rect 18174 210539 18208 210550
rect 21413 210543 22813 210671
rect 23685 210543 25085 210671
rect 15748 210529 15806 210539
rect 15816 210529 15874 210539
rect 15884 210529 15942 210539
rect 15952 210529 16010 210539
rect 16020 210529 16078 210539
rect 16088 210529 16146 210539
rect 16156 210529 16214 210539
rect 16224 210529 16282 210539
rect 16292 210529 16350 210539
rect 16360 210529 16418 210539
rect 16428 210529 16486 210539
rect 16496 210529 16554 210539
rect 16564 210529 16622 210539
rect 16632 210529 16690 210539
rect 17290 210529 17348 210539
rect 17358 210529 17416 210539
rect 17426 210529 17484 210539
rect 17494 210529 17552 210539
rect 17562 210529 17620 210539
rect 17630 210529 17688 210539
rect 17698 210529 17756 210539
rect 17766 210529 17824 210539
rect 17834 210529 17892 210539
rect 17902 210529 17960 210539
rect 17970 210529 18028 210539
rect 18038 210529 18096 210539
rect 18106 210529 18164 210539
rect 18174 210529 18232 210539
rect 15724 210505 16690 210529
rect 17266 210505 18232 210529
rect 15748 210490 15772 210505
rect 15816 210490 15840 210505
rect 15884 210490 15908 210505
rect 15952 210490 15976 210505
rect 16020 210490 16044 210505
rect 16088 210490 16112 210505
rect 16156 210490 16180 210505
rect 16224 210490 16248 210505
rect 16292 210490 16316 210505
rect 16360 210490 16384 210505
rect 16428 210490 16452 210505
rect 16496 210490 16520 210505
rect 16564 210490 16588 210505
rect 16632 210490 16656 210505
rect 17290 210490 17314 210505
rect 17358 210490 17382 210505
rect 17426 210490 17450 210505
rect 17494 210490 17518 210505
rect 17562 210490 17586 210505
rect 17630 210490 17654 210505
rect 17698 210490 17722 210505
rect 17766 210490 17790 210505
rect 17834 210490 17858 210505
rect 17902 210490 17926 210505
rect 17970 210490 17994 210505
rect 18038 210490 18062 210505
rect 18106 210490 18130 210505
rect 18174 210490 18198 210505
rect 15678 210335 16678 210490
rect 7389 210245 8389 210305
rect 8990 210245 9990 210305
rect 15678 210301 16690 210335
rect 17278 210325 18278 210490
rect 21413 210380 22813 210508
rect 23685 210380 25085 210508
rect 17266 210301 18278 210325
rect 15678 210290 16678 210301
rect 17278 210290 18278 210301
rect 15748 210277 15772 210290
rect 15816 210277 15840 210290
rect 15884 210277 15908 210290
rect 15952 210277 15976 210290
rect 16020 210277 16044 210290
rect 16088 210277 16112 210290
rect 16156 210277 16180 210290
rect 16224 210277 16248 210290
rect 16292 210277 16316 210290
rect 16360 210277 16384 210290
rect 16428 210277 16452 210290
rect 16496 210277 16520 210290
rect 16564 210277 16588 210290
rect 16632 210277 16656 210290
rect 17290 210277 17314 210290
rect 17358 210277 17382 210290
rect 17426 210277 17450 210290
rect 17494 210277 17518 210290
rect 17562 210277 17586 210290
rect 17630 210277 17654 210290
rect 17698 210277 17722 210290
rect 17766 210277 17790 210290
rect 17834 210277 17858 210290
rect 17902 210277 17926 210290
rect 17970 210277 17994 210290
rect 18038 210277 18062 210290
rect 18106 210277 18130 210290
rect 18174 210277 18198 210290
rect 21413 210217 22813 210345
rect 23685 210217 25085 210345
rect 21413 210054 22813 210182
rect 23685 210054 25085 210182
rect 25936 210132 26936 210182
rect 27274 210033 27358 210036
rect 13899 209998 14059 210002
rect 7389 209887 8389 209943
rect 8990 209887 9990 209943
rect 15678 209932 16678 209988
rect 17278 209932 18278 209988
rect 7389 209815 8389 209871
rect 8990 209815 9990 209871
rect 15678 209860 16678 209916
rect 17278 209860 18278 209916
rect 21413 209891 22813 210019
rect 23685 209891 25085 210019
rect 25936 209976 26936 210032
rect 27158 209983 27358 210033
rect 13899 209852 14059 209856
rect 25936 209820 26936 209876
rect 27158 209807 27358 209935
rect 21413 209741 22813 209784
rect 23685 209741 25085 209784
rect 25936 209664 26936 209720
rect 7389 209513 8389 209585
rect 8990 209513 9990 209585
rect 15678 209558 16678 209630
rect 17278 209558 18278 209630
rect 21413 209605 22813 209648
rect 23685 209605 25085 209648
rect 27158 209631 27358 209687
rect 15748 209547 15782 209558
rect 15816 209547 15850 209558
rect 15884 209547 15918 209558
rect 15952 209547 15986 209558
rect 16020 209547 16054 209558
rect 16088 209547 16122 209558
rect 16156 209547 16190 209558
rect 16224 209547 16258 209558
rect 16292 209547 16326 209558
rect 16360 209547 16394 209558
rect 16428 209547 16462 209558
rect 16496 209547 16530 209558
rect 16564 209547 16598 209558
rect 16632 209547 16666 209558
rect 17290 209547 17324 209558
rect 17358 209547 17392 209558
rect 17426 209547 17460 209558
rect 17494 209547 17528 209558
rect 17562 209547 17596 209558
rect 17630 209547 17664 209558
rect 17698 209547 17732 209558
rect 17766 209547 17800 209558
rect 17834 209547 17868 209558
rect 17902 209547 17936 209558
rect 17970 209547 18004 209558
rect 18038 209547 18072 209558
rect 18106 209547 18140 209558
rect 18174 209547 18208 209558
rect 15748 209537 15806 209547
rect 15816 209537 15874 209547
rect 15884 209537 15942 209547
rect 15952 209537 16010 209547
rect 16020 209537 16078 209547
rect 16088 209537 16146 209547
rect 16156 209537 16214 209547
rect 16224 209537 16282 209547
rect 16292 209537 16350 209547
rect 16360 209537 16418 209547
rect 16428 209537 16486 209547
rect 16496 209537 16554 209547
rect 16564 209537 16622 209547
rect 16632 209537 16690 209547
rect 17290 209537 17348 209547
rect 17358 209537 17416 209547
rect 17426 209537 17484 209547
rect 17494 209537 17552 209547
rect 17562 209537 17620 209547
rect 17630 209537 17688 209547
rect 17698 209537 17756 209547
rect 17766 209537 17824 209547
rect 17834 209537 17892 209547
rect 17902 209537 17960 209547
rect 17970 209537 18028 209547
rect 18038 209537 18096 209547
rect 18106 209537 18164 209547
rect 18174 209537 18232 209547
rect 15724 209513 16690 209537
rect 17266 209513 18232 209537
rect 15748 209498 15772 209513
rect 15816 209498 15840 209513
rect 15884 209498 15908 209513
rect 15952 209498 15976 209513
rect 16020 209498 16044 209513
rect 16088 209498 16112 209513
rect 16156 209498 16180 209513
rect 16224 209498 16248 209513
rect 16292 209498 16316 209513
rect 16360 209498 16384 209513
rect 16428 209498 16452 209513
rect 16496 209498 16520 209513
rect 16564 209498 16588 209513
rect 16632 209498 16656 209513
rect 17290 209498 17314 209513
rect 17358 209498 17382 209513
rect 17426 209498 17450 209513
rect 17494 209498 17518 209513
rect 17562 209498 17586 209513
rect 17630 209498 17654 209513
rect 17698 209498 17722 209513
rect 17766 209498 17790 209513
rect 17834 209498 17858 209513
rect 17902 209498 17926 209513
rect 17970 209498 17994 209513
rect 18038 209498 18062 209513
rect 18106 209498 18130 209513
rect 18174 209498 18198 209513
rect 15678 209343 16678 209498
rect 7389 209253 8389 209313
rect 8990 209253 9990 209313
rect 15678 209309 16690 209343
rect 17278 209333 18278 209498
rect 21413 209442 22813 209570
rect 23685 209442 25085 209570
rect 25936 209514 26936 209564
rect 26393 209511 26477 209514
rect 26726 209511 26810 209514
rect 27158 209455 27358 209583
rect 17266 209309 18278 209333
rect 15678 209298 16678 209309
rect 17278 209298 18278 209309
rect 15748 209285 15772 209298
rect 15816 209285 15840 209298
rect 15884 209285 15908 209298
rect 15952 209285 15976 209298
rect 16020 209285 16044 209298
rect 16088 209285 16112 209298
rect 16156 209285 16180 209298
rect 16224 209285 16248 209298
rect 16292 209285 16316 209298
rect 16360 209285 16384 209298
rect 16428 209285 16452 209298
rect 16496 209285 16520 209298
rect 16564 209285 16588 209298
rect 16632 209285 16656 209298
rect 17290 209285 17314 209298
rect 17358 209285 17382 209298
rect 17426 209285 17450 209298
rect 17494 209285 17518 209298
rect 17562 209285 17586 209298
rect 17630 209285 17654 209298
rect 17698 209285 17722 209298
rect 17766 209285 17790 209298
rect 17834 209285 17858 209298
rect 17902 209285 17926 209298
rect 17970 209285 17994 209298
rect 18038 209285 18062 209298
rect 18106 209285 18130 209298
rect 18174 209285 18198 209298
rect 21413 209279 22813 209407
rect 23685 209279 25085 209407
rect 27158 209279 27358 209335
rect 21413 209116 22813 209244
rect 23685 209116 25085 209244
rect 27158 209103 27358 209231
rect 26393 209100 26477 209103
rect 26726 209100 26810 209103
rect 12543 209069 12881 209085
rect 12559 208967 12865 209069
rect 7389 208895 8389 208951
rect 8990 208895 9990 208951
rect 15678 208940 16678 208996
rect 17278 208940 18278 208996
rect 21413 208953 22813 209081
rect 23685 208953 25085 209081
rect 25936 209050 26936 209100
rect 27622 209095 27672 210095
rect 27772 209095 27828 210095
rect 27928 209095 27984 210095
rect 28084 209095 28140 210095
rect 28240 209095 28296 210095
rect 28396 209637 28446 210095
rect 28396 209553 28449 209637
rect 28396 209305 28446 209553
rect 29778 209320 29802 209344
rect 28396 209221 28449 209305
rect 29802 209296 29826 209309
rect 29880 209299 29914 209333
rect 29778 209261 29802 209285
rect 29890 209275 29914 209299
rect 28396 209095 28446 209221
rect 7389 208823 8389 208879
rect 8990 208823 9990 208879
rect 15678 208868 16678 208924
rect 17278 208868 18278 208924
rect 21413 208790 22813 208918
rect 23685 208790 25085 208918
rect 25936 208894 26936 208950
rect 27158 208927 27358 208983
rect 13899 208656 14059 208660
rect 7389 208521 8389 208593
rect 8990 208521 9990 208593
rect 15678 208566 16678 208638
rect 17278 208566 18278 208638
rect 21413 208627 22813 208755
rect 23685 208627 25085 208755
rect 25936 208738 26936 208794
rect 27158 208751 27358 208879
rect 27912 208757 27962 208873
rect 27909 208673 27962 208757
rect 28082 208673 28210 208873
rect 28258 208673 28314 208873
rect 28434 208673 28562 208873
rect 28610 208673 28660 208873
rect 27917 208669 27951 208673
rect 29880 208672 29914 208706
rect 25936 208582 26936 208638
rect 27158 208581 27358 208631
rect 27274 208578 27358 208581
rect 15748 208555 15782 208566
rect 15816 208555 15850 208566
rect 15884 208555 15918 208566
rect 15952 208555 15986 208566
rect 16020 208555 16054 208566
rect 16088 208555 16122 208566
rect 16156 208555 16190 208566
rect 16224 208555 16258 208566
rect 16292 208555 16326 208566
rect 16360 208555 16394 208566
rect 16428 208555 16462 208566
rect 16496 208555 16530 208566
rect 16564 208555 16598 208566
rect 16632 208555 16666 208566
rect 17290 208555 17324 208566
rect 17358 208555 17392 208566
rect 17426 208555 17460 208566
rect 17494 208555 17528 208566
rect 17562 208555 17596 208566
rect 17630 208555 17664 208566
rect 17698 208555 17732 208566
rect 17766 208555 17800 208566
rect 17834 208555 17868 208566
rect 17902 208555 17936 208566
rect 17970 208555 18004 208566
rect 18038 208555 18072 208566
rect 18106 208555 18140 208566
rect 18174 208555 18208 208566
rect 15748 208545 15806 208555
rect 15816 208545 15874 208555
rect 15884 208545 15942 208555
rect 15952 208545 16010 208555
rect 16020 208545 16078 208555
rect 16088 208545 16146 208555
rect 16156 208545 16214 208555
rect 16224 208545 16282 208555
rect 16292 208545 16350 208555
rect 16360 208545 16418 208555
rect 16428 208545 16486 208555
rect 16496 208545 16554 208555
rect 16564 208545 16622 208555
rect 16632 208545 16690 208555
rect 17290 208545 17348 208555
rect 17358 208545 17416 208555
rect 17426 208545 17484 208555
rect 17494 208545 17552 208555
rect 17562 208545 17620 208555
rect 17630 208545 17688 208555
rect 17698 208545 17756 208555
rect 17766 208545 17824 208555
rect 17834 208545 17892 208555
rect 17902 208545 17960 208555
rect 17970 208545 18028 208555
rect 18038 208545 18096 208555
rect 18106 208545 18164 208555
rect 18174 208545 18232 208555
rect 15724 208521 16690 208545
rect 17266 208521 18232 208545
rect 13901 208510 14061 208514
rect 15748 208506 15772 208521
rect 15816 208506 15840 208521
rect 15884 208506 15908 208521
rect 15952 208506 15976 208521
rect 16020 208506 16044 208521
rect 16088 208506 16112 208521
rect 16156 208506 16180 208521
rect 16224 208506 16248 208521
rect 16292 208506 16316 208521
rect 16360 208506 16384 208521
rect 16428 208506 16452 208521
rect 16496 208506 16520 208521
rect 16564 208506 16588 208521
rect 16632 208506 16656 208521
rect 17290 208506 17314 208521
rect 17358 208506 17382 208521
rect 17426 208506 17450 208521
rect 17494 208506 17518 208521
rect 17562 208506 17586 208521
rect 17630 208506 17654 208521
rect 17698 208506 17722 208521
rect 17766 208506 17790 208521
rect 17834 208506 17858 208521
rect 17902 208506 17926 208521
rect 17970 208506 17994 208521
rect 18038 208506 18062 208521
rect 18106 208506 18130 208521
rect 18174 208506 18198 208521
rect 15678 208351 16678 208506
rect 7389 208261 8389 208321
rect 8990 208261 9990 208321
rect 15678 208317 16690 208351
rect 17278 208341 18278 208506
rect 21413 208470 22813 208520
rect 23685 208470 25085 208520
rect 25936 208432 26936 208482
rect 21349 208390 21373 208414
rect 21407 208390 21431 208414
rect 25067 208390 25091 208414
rect 25125 208390 25149 208414
rect 21383 208356 21397 208390
rect 25101 208356 25115 208390
rect 17266 208317 18278 208341
rect 21349 208332 21373 208356
rect 21407 208332 21431 208356
rect 25067 208332 25091 208356
rect 25125 208332 25149 208356
rect 27917 208325 27951 208329
rect 15678 208306 16678 208317
rect 17278 208306 18278 208317
rect 15748 208293 15772 208306
rect 15816 208293 15840 208306
rect 15884 208293 15908 208306
rect 15952 208293 15976 208306
rect 16020 208293 16044 208306
rect 16088 208293 16112 208306
rect 16156 208293 16180 208306
rect 16224 208293 16248 208306
rect 16292 208293 16316 208306
rect 16360 208293 16384 208306
rect 16428 208293 16452 208306
rect 16496 208293 16520 208306
rect 16564 208293 16588 208306
rect 16632 208293 16656 208306
rect 17290 208293 17314 208306
rect 17358 208293 17382 208306
rect 17426 208293 17450 208306
rect 17494 208293 17518 208306
rect 17562 208293 17586 208306
rect 17630 208293 17654 208306
rect 17698 208293 17722 208306
rect 17766 208293 17790 208306
rect 17834 208293 17858 208306
rect 17902 208293 17926 208306
rect 17970 208293 17994 208306
rect 18038 208293 18062 208306
rect 18106 208293 18130 208306
rect 18174 208293 18198 208306
rect 27909 208241 27962 208325
rect 21634 208101 24864 208203
rect 27912 208125 27962 208241
rect 28082 208125 28210 208325
rect 28258 208125 28314 208325
rect 28434 208125 28562 208325
rect 28610 208125 28660 208325
rect 21186 208047 21210 208071
rect 25288 208047 25312 208071
rect 21162 208023 21186 208037
rect 25312 208023 25336 208037
rect 7389 207903 8389 207959
rect 8990 207903 9990 207959
rect 15678 207948 16678 208004
rect 17278 207948 18278 208004
rect 21072 207989 21084 208013
rect 21186 207989 21210 208013
rect 25288 207989 25312 208013
rect 25414 207989 25426 208013
rect 21385 207944 21403 207948
rect 7389 207831 8389 207887
rect 8990 207831 9990 207887
rect 15678 207876 16678 207932
rect 17278 207876 18278 207932
rect 20250 207914 20316 207930
rect 21377 207914 21403 207944
rect 21385 207904 21403 207914
rect 21383 207880 21403 207904
rect 21407 207880 21415 207914
rect 25113 207904 25121 207944
rect 25101 207880 25121 207904
rect 25125 207880 25143 207948
rect 21383 207846 21419 207880
rect 25101 207846 25147 207880
rect 21383 207812 21403 207846
rect 21407 207812 21415 207846
rect 21383 207778 21419 207812
rect 21481 207784 22881 207834
rect 23617 207784 25017 207834
rect 25101 207812 25121 207846
rect 25125 207812 25143 207846
rect 25101 207778 25147 207812
rect 21383 207744 21403 207778
rect 21407 207744 21415 207778
rect 21383 207710 21419 207744
rect 21383 207676 21403 207710
rect 21407 207676 21415 207710
rect 7389 207529 8389 207601
rect 8990 207529 9990 207601
rect 15678 207574 16678 207646
rect 17278 207574 18278 207646
rect 21383 207642 21419 207676
rect 21383 207608 21403 207642
rect 21407 207608 21415 207642
rect 21481 207621 22881 207749
rect 23617 207621 25017 207749
rect 25101 207744 25121 207778
rect 25125 207744 25143 207778
rect 25101 207710 25147 207744
rect 25101 207676 25121 207710
rect 25125 207676 25143 207710
rect 25101 207642 25147 207676
rect 25101 207608 25121 207642
rect 25125 207608 25143 207642
rect 21383 207574 21419 207608
rect 15748 207563 15782 207574
rect 15816 207563 15850 207574
rect 15884 207563 15918 207574
rect 15952 207563 15986 207574
rect 16020 207563 16054 207574
rect 16088 207563 16122 207574
rect 16156 207563 16190 207574
rect 16224 207563 16258 207574
rect 16292 207563 16326 207574
rect 16360 207563 16394 207574
rect 16428 207563 16462 207574
rect 16496 207563 16530 207574
rect 16564 207563 16598 207574
rect 16632 207563 16666 207574
rect 17290 207563 17324 207574
rect 17358 207563 17392 207574
rect 17426 207563 17460 207574
rect 17494 207563 17528 207574
rect 17562 207563 17596 207574
rect 17630 207563 17664 207574
rect 17698 207563 17732 207574
rect 17766 207563 17800 207574
rect 17834 207563 17868 207574
rect 17902 207563 17936 207574
rect 17970 207563 18004 207574
rect 18038 207563 18072 207574
rect 18106 207563 18140 207574
rect 18174 207563 18208 207574
rect 15748 207553 15806 207563
rect 15816 207553 15874 207563
rect 15884 207553 15942 207563
rect 15952 207553 16010 207563
rect 16020 207553 16078 207563
rect 16088 207553 16146 207563
rect 16156 207553 16214 207563
rect 16224 207553 16282 207563
rect 16292 207553 16350 207563
rect 16360 207553 16418 207563
rect 16428 207553 16486 207563
rect 16496 207553 16554 207563
rect 16564 207553 16622 207563
rect 16632 207553 16690 207563
rect 17290 207553 17348 207563
rect 17358 207553 17416 207563
rect 17426 207553 17484 207563
rect 17494 207553 17552 207563
rect 17562 207553 17620 207563
rect 17630 207553 17688 207563
rect 17698 207553 17756 207563
rect 17766 207553 17824 207563
rect 17834 207553 17892 207563
rect 17902 207553 17960 207563
rect 17970 207553 18028 207563
rect 18038 207553 18096 207563
rect 18106 207553 18164 207563
rect 18174 207553 18232 207563
rect 15724 207529 16690 207553
rect 17266 207529 18232 207553
rect 21383 207540 21403 207574
rect 21407 207540 21415 207574
rect 15748 207514 15772 207529
rect 15816 207514 15840 207529
rect 15884 207514 15908 207529
rect 15952 207514 15976 207529
rect 16020 207514 16044 207529
rect 16088 207514 16112 207529
rect 16156 207514 16180 207529
rect 16224 207514 16248 207529
rect 16292 207514 16316 207529
rect 16360 207514 16384 207529
rect 16428 207514 16452 207529
rect 16496 207514 16520 207529
rect 16564 207514 16588 207529
rect 16632 207514 16656 207529
rect 17290 207514 17314 207529
rect 17358 207514 17382 207529
rect 17426 207514 17450 207529
rect 17494 207514 17518 207529
rect 17562 207514 17586 207529
rect 17630 207514 17654 207529
rect 17698 207514 17722 207529
rect 17766 207514 17790 207529
rect 17834 207514 17858 207529
rect 17902 207514 17926 207529
rect 17970 207514 17994 207529
rect 18038 207514 18062 207529
rect 18106 207514 18130 207529
rect 18174 207514 18198 207529
rect 5937 207318 6089 207386
rect 15678 207359 16678 207514
rect 6005 207315 6089 207318
rect 5967 207305 6059 207315
rect 6005 207275 6021 207305
rect 1288 205503 1338 206503
rect 1438 205503 1566 206503
rect 1594 205503 1644 206503
rect 5995 205493 6021 207275
rect 7389 207269 8389 207329
rect 8990 207269 9990 207329
rect 15678 207325 16690 207359
rect 17278 207349 18278 207514
rect 17266 207325 18278 207349
rect 15678 207314 16678 207325
rect 17278 207314 18278 207325
rect 21383 207506 21419 207540
rect 21383 207472 21403 207506
rect 21407 207472 21415 207506
rect 21383 207438 21419 207472
rect 21481 207458 22881 207586
rect 23617 207458 25017 207586
rect 25101 207574 25147 207608
rect 25101 207540 25121 207574
rect 25125 207540 25143 207574
rect 25101 207506 25147 207540
rect 25101 207472 25121 207506
rect 25125 207472 25143 207506
rect 25101 207438 25147 207472
rect 21383 207404 21403 207438
rect 21407 207404 21415 207438
rect 21383 207370 21419 207404
rect 21383 207336 21403 207370
rect 21407 207336 21415 207370
rect 15748 207301 15772 207314
rect 15816 207301 15840 207314
rect 15884 207301 15908 207314
rect 15952 207301 15976 207314
rect 16020 207301 16044 207314
rect 16088 207301 16112 207314
rect 16156 207301 16180 207314
rect 16224 207301 16248 207314
rect 16292 207301 16316 207314
rect 16360 207301 16384 207314
rect 16428 207301 16452 207314
rect 16496 207301 16520 207314
rect 16564 207301 16588 207314
rect 16632 207301 16656 207314
rect 17290 207301 17314 207314
rect 17358 207301 17382 207314
rect 17426 207301 17450 207314
rect 17494 207301 17518 207314
rect 17562 207301 17586 207314
rect 17630 207301 17654 207314
rect 17698 207301 17722 207314
rect 17766 207301 17790 207314
rect 17834 207301 17858 207314
rect 17902 207301 17926 207314
rect 17970 207301 17994 207314
rect 18038 207301 18062 207314
rect 18106 207301 18130 207314
rect 18174 207301 18198 207314
rect 21383 207302 21419 207336
rect 21383 207268 21403 207302
rect 21407 207268 21415 207302
rect 21481 207295 22881 207423
rect 23617 207295 25017 207423
rect 25101 207404 25121 207438
rect 25125 207404 25143 207438
rect 25101 207370 25147 207404
rect 25101 207336 25121 207370
rect 25125 207336 25143 207370
rect 25101 207302 25147 207336
rect 25101 207268 25121 207302
rect 25125 207268 25143 207302
rect 21383 207234 21419 207268
rect 21383 207200 21403 207234
rect 21407 207200 21415 207234
rect 21383 207166 21419 207200
rect 21383 207132 21403 207166
rect 21407 207132 21415 207166
rect 21481 207132 22881 207260
rect 23617 207132 25017 207260
rect 25101 207234 25147 207268
rect 25101 207200 25121 207234
rect 25125 207200 25143 207234
rect 25101 207166 25147 207200
rect 25101 207132 25121 207166
rect 25125 207132 25143 207166
rect 21383 207098 21419 207132
rect 25101 207098 25147 207132
rect 21383 207064 21403 207098
rect 21407 207064 21415 207098
rect 21383 207030 21419 207064
rect 7389 206911 8389 206967
rect 8990 206911 9990 206967
rect 15678 206956 16678 207012
rect 17278 206956 18278 207012
rect 21383 206996 21403 207030
rect 21407 206996 21415 207030
rect 21383 206962 21419 206996
rect 21481 206969 22881 207097
rect 23617 206969 25017 207097
rect 25101 207064 25121 207098
rect 25125 207064 25143 207098
rect 25101 207030 25147 207064
rect 25101 206996 25121 207030
rect 25125 206996 25143 207030
rect 25101 206962 25147 206996
rect 26478 206985 26648 207291
rect 7389 206839 8389 206895
rect 8990 206839 9990 206895
rect 15678 206884 16678 206940
rect 17278 206884 18278 206940
rect 21383 206928 21403 206962
rect 21407 206928 21415 206962
rect 21383 206894 21419 206928
rect 21383 206860 21403 206894
rect 21407 206860 21415 206894
rect 21383 206826 21419 206860
rect 21383 206792 21403 206826
rect 21407 206792 21415 206826
rect 21481 206806 22881 206934
rect 23617 206806 25017 206934
rect 25101 206928 25121 206962
rect 25125 206928 25143 206962
rect 25101 206894 25147 206928
rect 27622 206903 27672 207903
rect 27772 206903 27828 207903
rect 27928 206903 27984 207903
rect 28084 206903 28140 207903
rect 28240 206903 28296 207903
rect 28396 207777 28446 207903
rect 28396 207693 28449 207777
rect 28396 207445 28446 207693
rect 30015 207523 30027 213246
rect 32596 213239 33596 213367
rect 35255 213345 36255 213401
rect 30135 213062 30735 213112
rect 31049 213042 32049 213092
rect 32596 213083 33596 213211
rect 35255 213169 36255 213297
rect 35255 212993 36255 213121
rect 30135 212886 30735 212942
rect 31049 212886 32049 212942
rect 32596 212927 33596 212983
rect 37998 212979 38148 212991
rect 38317 212979 38467 212991
rect 30135 212716 30735 212766
rect 31049 212736 32049 212786
rect 32596 212777 33596 212827
rect 35255 212823 36255 212873
rect 37998 212866 38598 212916
rect 35255 212754 36255 212766
rect 37998 212690 38598 212746
rect 30135 212600 30735 212650
rect 31049 212600 32049 212650
rect 32596 212575 33196 212625
rect 35255 212621 36255 212671
rect 30135 212424 30735 212480
rect 31049 212444 32049 212500
rect 30135 212248 30735 212376
rect 31049 212288 32049 212344
rect 30135 212072 30735 212200
rect 31049 212132 32049 212188
rect 32596 212141 33196 212191
rect 30135 211896 30735 212024
rect 31049 211982 32049 212032
rect 31049 211866 32049 211916
rect 30135 211726 30735 211776
rect 31049 211710 32049 211838
rect 30135 211610 30735 211660
rect 30135 211434 30735 211562
rect 31049 211554 32049 211682
rect 31049 211398 32049 211526
rect 34152 211490 34202 212478
rect 34322 211490 34372 212478
rect 34492 212465 35092 212515
rect 35255 212445 36255 212573
rect 37998 212520 38598 212570
rect 36785 212496 36797 212500
rect 36785 212485 36800 212496
rect 36970 212485 36985 212500
rect 34492 212289 35092 212345
rect 35255 212269 36255 212325
rect 36785 212305 36985 212485
rect 36785 212294 36800 212305
rect 36785 212290 36797 212294
rect 36970 212290 36985 212305
rect 37083 212485 37098 212500
rect 37083 212305 37120 212485
rect 37083 212290 37098 212305
rect 36785 212260 36797 212264
rect 36785 212249 36800 212260
rect 36970 212249 36985 212264
rect 34492 212119 35092 212169
rect 35255 212099 36255 212149
rect 36785 212069 36985 212249
rect 37993 212094 38593 212144
rect 36785 212058 36800 212069
rect 36785 212054 36797 212058
rect 36970 212054 36985 212069
rect 34491 211849 35091 211899
rect 35255 211883 35855 211933
rect 37993 211924 38593 211974
rect 34491 211673 35091 211729
rect 35255 211707 35855 211763
rect 36785 211748 37385 211798
rect 38920 211761 38946 211787
rect 34491 211503 35091 211553
rect 35255 211531 35855 211659
rect 36785 211572 37385 211628
rect 34019 211418 34029 211490
rect 34152 211478 34372 211490
rect 34091 211415 34101 211418
rect 30135 211258 30735 211314
rect 31049 211242 32049 211370
rect 34091 211365 35091 211415
rect 35255 211361 35855 211411
rect 36785 211396 37385 211452
rect 30135 211082 30735 211210
rect 31049 211086 32049 211214
rect 34091 211195 35091 211245
rect 36785 211226 37385 211276
rect 34091 211192 34101 211195
rect 34202 211192 34302 211195
rect 35255 211159 35855 211209
rect 30135 210912 30735 210962
rect 31049 210930 32049 210986
rect 30135 210796 30735 210846
rect 31049 210774 32049 210902
rect 32481 210898 33081 210948
rect 30135 210620 30735 210748
rect 31049 210618 32049 210746
rect 32481 210742 33081 210870
rect 30135 210444 30735 210572
rect 31049 210462 32049 210590
rect 32481 210586 33081 210714
rect 34152 210532 34202 211132
rect 34302 210532 34352 211132
rect 34491 211066 35091 211116
rect 35255 211003 35855 211131
rect 36785 211094 37385 211144
rect 34491 210890 35091 210946
rect 36785 210918 37385 210974
rect 35255 210847 35855 210903
rect 34491 210720 35091 210770
rect 35255 210691 35855 210819
rect 36785 210742 37385 210798
rect 35255 210541 35855 210591
rect 36785 210572 37385 210622
rect 32481 210436 33081 210486
rect 30135 210268 30735 210396
rect 31049 210306 32049 210434
rect 34491 210379 35091 210429
rect 37993 210396 38593 210446
rect 32481 210306 33081 210356
rect 33261 210287 33861 210323
rect 30135 210092 30735 210220
rect 31049 210150 32049 210278
rect 32481 210150 33081 210278
rect 34491 210203 35091 210331
rect 35255 210287 35855 210337
rect 36785 210312 36797 210316
rect 36785 210301 36800 210312
rect 36970 210301 36985 210316
rect 35255 210131 35855 210259
rect 36785 210121 36985 210301
rect 37993 210226 38593 210276
rect 36785 210110 36800 210121
rect 36785 210106 36797 210110
rect 36970 210106 36985 210121
rect 30135 209916 30735 210044
rect 31049 209994 32049 210050
rect 32481 209994 33081 210050
rect 34491 210027 35091 210083
rect 31049 209818 32049 209946
rect 32481 209838 33081 209966
rect 33261 209907 33861 209963
rect 34491 209851 35091 209979
rect 35255 209975 35855 210103
rect 36785 210076 36797 210080
rect 36785 210065 36800 210076
rect 36970 210065 36985 210080
rect 36785 209885 36985 210065
rect 35255 209819 35855 209875
rect 36785 209874 36800 209885
rect 36785 209870 36797 209874
rect 36970 209870 36985 209885
rect 37083 210065 37098 210080
rect 37083 209885 37120 210065
rect 37083 209870 37098 209885
rect 37998 209800 38598 209850
rect 30135 209740 30735 209796
rect 30135 209564 30735 209692
rect 31049 209642 32049 209770
rect 32481 209688 33081 209738
rect 33261 209723 33861 209773
rect 34491 209681 35091 209731
rect 35255 209669 35855 209719
rect 37998 209624 38598 209680
rect 30135 209388 30735 209516
rect 31049 209466 32049 209594
rect 32481 209558 33081 209608
rect 30135 209212 30735 209340
rect 31049 209290 32049 209418
rect 32481 209402 33081 209458
rect 37998 209454 38598 209504
rect 37998 209451 38220 209454
rect 38245 209451 38539 209454
rect 32481 209252 33081 209302
rect 34427 209259 35027 209309
rect 30135 209036 30735 209164
rect 31049 209114 32049 209242
rect 33672 209183 34272 209233
rect 34427 209083 35027 209211
rect 30135 208860 30735 208988
rect 31049 208938 32049 209066
rect 33672 209007 34272 209063
rect 31049 208762 32049 208890
rect 33672 208831 34272 208959
rect 34427 208907 35027 209035
rect 30135 208684 30735 208740
rect 34427 208731 35027 208859
rect 37998 208825 38148 208837
rect 38317 208825 38467 208837
rect 37998 208712 38598 208762
rect 33672 208655 34272 208711
rect 30135 208508 30735 208636
rect 31049 208592 32049 208642
rect 34427 208555 35027 208683
rect 37998 208536 38598 208592
rect 31049 208476 32049 208526
rect 33672 208479 34272 208535
rect 30135 208332 30735 208388
rect 31049 208320 32049 208448
rect 34427 208379 35027 208435
rect 37998 208366 38598 208416
rect 33672 208303 34272 208359
rect 36785 208342 36797 208346
rect 36785 208331 36800 208342
rect 36970 208331 36985 208346
rect 30135 208156 30735 208284
rect 31049 208164 32049 208292
rect 30135 207980 30735 208036
rect 31049 208008 32049 208136
rect 33672 208127 34272 208255
rect 34427 208203 35027 208331
rect 36785 208151 36985 208331
rect 36785 208140 36800 208151
rect 36785 208136 36797 208140
rect 36970 208136 36985 208151
rect 37083 208331 37098 208346
rect 37083 208151 37120 208331
rect 37083 208136 37098 208151
rect 36785 208106 36797 208110
rect 36785 208095 36800 208106
rect 36970 208095 36985 208110
rect 34427 208033 35027 208083
rect 33672 207957 34272 208007
rect 30135 207804 30735 207932
rect 36785 207915 36985 208095
rect 37993 207940 38593 207990
rect 31049 207852 32049 207908
rect 36785 207904 36800 207915
rect 36785 207900 36797 207904
rect 36970 207900 36985 207915
rect 31049 207696 32049 207824
rect 37993 207770 38593 207820
rect 30135 207634 30735 207684
rect 31049 207540 32049 207668
rect 36785 207594 37385 207644
rect 28396 207361 28449 207445
rect 31049 207384 32049 207512
rect 36785 207418 37385 207474
rect 28396 206903 28446 207361
rect 31049 207234 32049 207284
rect 36785 207242 37385 207298
rect 36785 207072 37385 207122
rect 37939 207039 37963 207063
rect 38085 207039 38109 207063
rect 29925 207003 29931 207032
rect 30271 207003 30305 207027
rect 30342 207003 30376 207027
rect 30413 207003 30447 207027
rect 30484 207003 30518 207027
rect 30555 207003 30589 207027
rect 30626 207003 30660 207027
rect 30697 207003 30731 207027
rect 37963 207015 37987 207038
rect 38061 207015 38085 207038
rect 29931 206962 29939 206986
rect 29955 206962 29961 207003
rect 29891 206938 29915 206962
rect 25101 206860 25121 206894
rect 25125 206860 25143 206894
rect 37759 206867 37783 206891
rect 25101 206826 25147 206860
rect 37792 206843 37807 206867
rect 25101 206792 25121 206826
rect 25125 206792 25143 206826
rect 21383 206758 21419 206792
rect 25101 206758 25147 206792
rect 21383 206724 21403 206758
rect 21407 206724 21415 206758
rect 25101 206724 25121 206758
rect 25125 206724 25143 206758
rect 21383 206690 21419 206724
rect 21383 206656 21403 206690
rect 21407 206656 21415 206690
rect 21481 206656 22881 206699
rect 22892 206675 22920 206703
rect 23617 206656 25017 206699
rect 25101 206690 25147 206724
rect 31458 206703 31608 206715
rect 31777 206703 31927 206715
rect 25101 206656 25121 206690
rect 25125 206656 25143 206690
rect 7389 206628 8389 206632
rect 8990 206628 9990 206632
rect 7353 206578 8425 206614
rect 7353 206537 7389 206578
rect 8389 206537 8425 206578
rect 7353 206501 8425 206537
rect 8954 206578 10026 206614
rect 15678 206582 16678 206654
rect 17278 206582 18278 206654
rect 21383 206622 21419 206656
rect 25101 206622 25147 206656
rect 21383 206588 21403 206622
rect 21407 206588 21415 206622
rect 25101 206588 25121 206622
rect 25125 206588 25143 206622
rect 8954 206537 8990 206578
rect 9990 206537 10026 206578
rect 15748 206571 15782 206582
rect 15816 206571 15850 206582
rect 15884 206571 15918 206582
rect 15952 206571 15986 206582
rect 16020 206571 16054 206582
rect 16088 206571 16122 206582
rect 16156 206571 16190 206582
rect 16224 206571 16258 206582
rect 16292 206571 16326 206582
rect 16360 206571 16394 206582
rect 16428 206571 16462 206582
rect 16496 206571 16530 206582
rect 16564 206571 16598 206582
rect 16632 206571 16666 206582
rect 17290 206571 17324 206582
rect 17358 206571 17392 206582
rect 17426 206571 17460 206582
rect 17494 206571 17528 206582
rect 17562 206571 17596 206582
rect 17630 206571 17664 206582
rect 17698 206571 17732 206582
rect 17766 206571 17800 206582
rect 17834 206571 17868 206582
rect 17902 206571 17936 206582
rect 17970 206571 18004 206582
rect 18038 206571 18072 206582
rect 18106 206571 18140 206582
rect 18174 206571 18208 206582
rect 15748 206561 15806 206571
rect 15816 206561 15874 206571
rect 15884 206561 15942 206571
rect 15952 206561 16010 206571
rect 16020 206561 16078 206571
rect 16088 206561 16146 206571
rect 16156 206561 16214 206571
rect 16224 206561 16282 206571
rect 16292 206561 16350 206571
rect 16360 206561 16418 206571
rect 16428 206561 16486 206571
rect 16496 206561 16554 206571
rect 16564 206561 16622 206571
rect 16632 206561 16690 206571
rect 17290 206561 17348 206571
rect 17358 206561 17416 206571
rect 17426 206561 17484 206571
rect 17494 206561 17552 206571
rect 17562 206561 17620 206571
rect 17630 206561 17688 206571
rect 17698 206561 17756 206571
rect 17766 206561 17824 206571
rect 17834 206561 17892 206571
rect 17902 206561 17960 206571
rect 17970 206561 18028 206571
rect 18038 206561 18096 206571
rect 18106 206561 18164 206571
rect 18174 206561 18232 206571
rect 15724 206537 16690 206561
rect 17266 206537 18232 206561
rect 21383 206554 21419 206588
rect 8954 206501 10026 206537
rect 15748 206522 15772 206537
rect 15816 206522 15840 206537
rect 15884 206522 15908 206537
rect 15952 206522 15976 206537
rect 16020 206522 16044 206537
rect 16088 206522 16112 206537
rect 16156 206522 16180 206537
rect 16224 206522 16248 206537
rect 16292 206522 16316 206537
rect 16360 206522 16384 206537
rect 16428 206522 16452 206537
rect 16496 206522 16520 206537
rect 16564 206522 16588 206537
rect 16632 206522 16656 206537
rect 17290 206522 17314 206537
rect 17358 206522 17382 206537
rect 17426 206522 17450 206537
rect 17494 206522 17518 206537
rect 17562 206522 17586 206537
rect 17630 206522 17654 206537
rect 17698 206522 17722 206537
rect 17766 206522 17790 206537
rect 17834 206522 17858 206537
rect 17902 206522 17926 206537
rect 17970 206522 17994 206537
rect 18038 206522 18062 206537
rect 18106 206522 18130 206537
rect 18174 206522 18198 206537
rect 15678 206367 16678 206522
rect 7389 206277 8389 206337
rect 8990 206277 9990 206337
rect 15678 206333 16690 206367
rect 17278 206357 18278 206522
rect 17266 206333 18278 206357
rect 15678 206322 16678 206333
rect 17278 206322 18278 206333
rect 21383 206520 21403 206554
rect 21407 206520 21415 206554
rect 21481 206520 22881 206563
rect 23617 206520 25017 206563
rect 25101 206554 25147 206588
rect 25414 206573 25438 206607
rect 31458 206590 32058 206640
rect 25101 206520 25121 206554
rect 25125 206520 25143 206554
rect 21383 206486 21419 206520
rect 25101 206486 25147 206520
rect 21383 206452 21403 206486
rect 21407 206452 21415 206486
rect 21383 206418 21419 206452
rect 21383 206384 21403 206418
rect 21407 206384 21415 206418
rect 21383 206350 21419 206384
rect 21481 206357 22881 206485
rect 23617 206357 25017 206485
rect 25101 206452 25121 206486
rect 25125 206452 25143 206486
rect 37792 206470 37807 206494
rect 25101 206418 25147 206452
rect 25101 206384 25121 206418
rect 25125 206384 25143 206418
rect 31458 206414 32058 206470
rect 37759 206446 37783 206470
rect 25101 206350 25147 206384
rect 15748 206309 15772 206322
rect 15816 206309 15840 206322
rect 15884 206309 15908 206322
rect 15952 206309 15976 206322
rect 16020 206309 16044 206322
rect 16088 206309 16112 206322
rect 16156 206309 16180 206322
rect 16224 206309 16248 206322
rect 16292 206309 16316 206322
rect 16360 206309 16384 206322
rect 16428 206309 16452 206322
rect 16496 206309 16520 206322
rect 16564 206309 16588 206322
rect 16632 206309 16656 206322
rect 17290 206309 17314 206322
rect 17358 206309 17382 206322
rect 17426 206309 17450 206322
rect 17494 206309 17518 206322
rect 17562 206309 17586 206322
rect 17630 206309 17654 206322
rect 17698 206309 17722 206322
rect 17766 206309 17790 206322
rect 17834 206309 17858 206322
rect 17902 206309 17926 206322
rect 17970 206309 17994 206322
rect 18038 206309 18062 206322
rect 18106 206309 18130 206322
rect 18174 206309 18198 206322
rect 21383 206316 21403 206350
rect 21407 206316 21415 206350
rect 21383 206282 21419 206316
rect 21383 206248 21403 206282
rect 21407 206248 21415 206282
rect 21383 206214 21419 206248
rect 21383 206180 21403 206214
rect 21407 206180 21415 206214
rect 21481 206194 22881 206322
rect 23617 206194 25017 206322
rect 25101 206316 25121 206350
rect 25125 206316 25143 206350
rect 25101 206282 25147 206316
rect 25101 206248 25121 206282
rect 25125 206248 25143 206282
rect 25101 206214 25147 206248
rect 25101 206180 25121 206214
rect 25125 206180 25143 206214
rect 25725 206197 26325 206247
rect 31458 206244 32058 206294
rect 30245 206220 30257 206224
rect 30245 206209 30260 206220
rect 30430 206209 30445 206224
rect 21383 206146 21419 206180
rect 7389 206066 8389 206070
rect 8990 206066 9990 206070
rect 15678 206061 16678 206133
rect 17278 206061 18278 206133
rect 21383 206112 21403 206146
rect 21407 206112 21415 206146
rect 21383 206078 21419 206112
rect 7353 206016 8425 206052
rect 7353 205975 7389 206016
rect 8389 205975 8425 206016
rect 7353 205919 8425 205975
rect 7353 205903 7389 205919
rect 8389 205903 8425 205919
rect 7353 205847 8425 205903
rect 7353 205810 7389 205847
rect 8389 205810 8425 205847
rect 7353 205770 8425 205810
rect 8954 206016 10026 206052
rect 8954 205975 8990 206016
rect 9990 205975 10026 206016
rect 8954 205919 10026 205975
rect 21383 206044 21403 206078
rect 21407 206044 21415 206078
rect 21383 206010 21419 206044
rect 21481 206031 22881 206159
rect 23617 206031 25017 206159
rect 25101 206146 25147 206180
rect 25101 206112 25121 206146
rect 25125 206112 25143 206146
rect 25101 206078 25147 206112
rect 25101 206044 25121 206078
rect 25125 206044 25143 206078
rect 25725 206047 26325 206097
rect 25101 206010 25147 206044
rect 21383 205976 21403 206010
rect 21407 205976 21415 206010
rect 21383 205942 21419 205976
rect 8954 205903 8990 205919
rect 9990 205903 10026 205919
rect 15678 205906 16678 205923
rect 17278 205906 18278 205923
rect 21383 205908 21403 205942
rect 21407 205908 21415 205942
rect 8954 205847 10026 205903
rect 20250 205890 20316 205906
rect 8954 205810 8990 205847
rect 9990 205810 10026 205847
rect 8954 205770 10026 205810
rect 21383 205874 21419 205908
rect 21383 205840 21403 205874
rect 21407 205840 21415 205874
rect 21481 205868 22881 205996
rect 23617 205868 25017 205996
rect 25101 205976 25121 206010
rect 25125 205976 25143 206010
rect 25101 205942 25147 205976
rect 25101 205908 25121 205942
rect 25125 205908 25143 205942
rect 25725 205925 26325 205975
rect 25101 205874 25147 205908
rect 25101 205840 25121 205874
rect 25125 205840 25143 205874
rect 21383 205806 21419 205840
rect 21383 205772 21403 205806
rect 21407 205772 21415 205806
rect 21383 205738 21419 205772
rect 15678 205703 16678 205736
rect 17278 205703 18278 205736
rect 21383 205704 21403 205738
rect 21407 205704 21415 205738
rect 21481 205705 22881 205833
rect 23617 205705 25017 205833
rect 25101 205806 25147 205840
rect 25101 205772 25121 205806
rect 25125 205772 25143 205806
rect 25725 205775 26325 205825
rect 25101 205738 25147 205772
rect 25101 205704 25121 205738
rect 25125 205704 25143 205738
rect 21383 205670 21419 205704
rect 25101 205670 25147 205704
rect 21383 205636 21403 205670
rect 21407 205636 21415 205670
rect 7389 205559 8389 205631
rect 8990 205559 9990 205631
rect 21383 205602 21419 205636
rect 15840 205510 15870 205580
rect 15878 205546 15908 205580
rect 21383 205568 21403 205602
rect 21407 205568 21415 205602
rect 15853 205508 15870 205510
rect 21383 205534 21419 205568
rect 21481 205542 22881 205670
rect 23617 205542 25017 205670
rect 25101 205636 25121 205670
rect 25125 205636 25143 205670
rect 25725 205649 26325 205699
rect 25101 205602 25147 205636
rect 25101 205568 25121 205602
rect 25125 205568 25143 205602
rect 25101 205534 25147 205568
rect 5981 205483 6021 205493
rect 5137 205469 6021 205483
rect 21383 205500 21403 205534
rect 21407 205500 21415 205534
rect 21383 205466 21419 205500
rect 7389 205369 8389 205463
rect 7389 205359 8413 205369
rect 8990 205359 9990 205463
rect 21383 205432 21403 205466
rect 21407 205432 21415 205466
rect 21383 205398 21419 205432
rect 21383 205364 21403 205398
rect 21407 205364 21415 205398
rect 21481 205379 22881 205507
rect 23617 205379 25017 205507
rect 25101 205500 25121 205534
rect 25125 205500 25143 205534
rect 25101 205466 25147 205500
rect 25725 205499 26325 205549
rect 25101 205432 25121 205466
rect 25125 205432 25143 205466
rect 25101 205398 25147 205432
rect 25101 205364 25121 205398
rect 25125 205364 25143 205398
rect 25725 205377 26325 205427
rect 21383 205330 21419 205364
rect 25101 205330 25147 205364
rect 21383 205296 21403 205330
rect 21407 205296 21415 205330
rect 25101 205296 25121 205330
rect 25125 205296 25143 205330
rect 21383 205262 21419 205296
rect 21383 205228 21403 205262
rect 21407 205228 21415 205262
rect 21481 205229 22881 205272
rect 23617 205229 25017 205272
rect 25101 205262 25147 205296
rect 25101 205228 25121 205262
rect 25125 205228 25143 205262
rect 21383 205194 21419 205228
rect 25101 205194 25147 205228
rect 25725 205227 26325 205277
rect 21383 205160 21403 205194
rect 21407 205160 21415 205194
rect 25101 205160 25121 205194
rect 25125 205160 25143 205194
rect 27162 205170 27212 206170
rect 27312 205170 27440 206170
rect 27468 205170 27596 206170
rect 27624 205170 27752 206170
rect 27780 205170 27908 206170
rect 27936 205170 28064 206170
rect 28092 205170 28220 206170
rect 28248 205170 28376 206170
rect 28404 205170 28532 206170
rect 28560 205170 28688 206170
rect 28716 205170 28844 206170
rect 28872 205170 29000 206170
rect 29028 205170 29156 206170
rect 29184 205170 29312 206170
rect 29340 205170 29390 206170
rect 30245 206029 30445 206209
rect 30245 206018 30260 206029
rect 30245 206014 30257 206018
rect 30430 206014 30445 206029
rect 30543 206209 30558 206224
rect 30543 206029 30580 206209
rect 30543 206014 30558 206029
rect 30245 205984 30257 205988
rect 30245 205973 30260 205984
rect 30430 205973 30445 205988
rect 30245 205793 30445 205973
rect 31453 205818 32053 205868
rect 30245 205782 30260 205793
rect 30245 205778 30257 205782
rect 30430 205778 30445 205793
rect 31453 205648 32053 205698
rect 30245 205472 30845 205522
rect 30245 205296 30845 205352
rect 21383 205126 21419 205160
rect 25101 205126 25147 205160
rect 21383 205102 21403 205126
rect 21385 205048 21403 205102
rect 21407 205082 21415 205126
rect 25101 205102 25121 205126
rect 25113 205082 25121 205102
rect 25125 205048 25143 205126
rect 30245 205120 30845 205176
rect 30245 204950 30845 205000
rect 21000 204800 21003 204920
rect 21352 204885 21376 204909
rect 25122 204885 25146 204909
rect 21385 204861 21400 204885
rect 25098 204861 25113 204885
rect 21274 204783 21294 204851
rect 21410 204817 21430 204851
rect 25068 204817 25088 204851
rect 25204 204817 25224 204851
rect 21385 204807 21430 204817
rect 25102 204807 25137 204817
rect 21361 204783 21430 204807
rect 25089 204783 25137 204807
rect 25238 204783 25258 204817
rect 684180 202243 685004 202293
rect 684180 202127 685004 202177
rect 684180 201971 685004 202027
rect 684180 201821 685004 201871
rect 684180 201600 684670 201649
rect 682921 201593 683521 201600
rect 684070 201599 684670 201600
rect 685537 201593 686137 201600
rect 680215 201518 680815 201574
rect 707610 201523 708610 201600
rect 709211 201523 710211 201591
rect 707610 201513 707624 201523
rect 707658 201513 707695 201523
rect 707729 201513 707769 201523
rect 707803 201513 707840 201523
rect 707874 201513 707914 201523
rect 707948 201513 707985 201523
rect 708019 201513 708059 201523
rect 708093 201513 708130 201523
rect 708164 201513 708204 201523
rect 708238 201513 708275 201523
rect 708309 201513 708369 201523
rect 708403 201513 708446 201523
rect 708480 201513 708522 201523
rect 708556 201513 708604 201523
rect 709219 201513 709270 201523
rect 709304 201513 709364 201523
rect 709398 201513 709435 201523
rect 709469 201513 709509 201523
rect 709543 201513 709580 201523
rect 709614 201513 709654 201523
rect 709688 201513 709725 201523
rect 709759 201513 709799 201523
rect 709833 201513 709870 201523
rect 709904 201513 709944 201523
rect 709978 201513 710015 201523
rect 710049 201513 710089 201523
rect 710123 201513 710160 201523
rect 710194 201513 710211 201523
rect 684070 201443 684670 201499
rect 685537 201443 686137 201493
rect 692428 201442 693028 201492
rect 680215 201348 680815 201398
rect 681713 201359 682313 201409
rect 684070 201293 684670 201343
rect 692428 201292 693028 201342
rect 705107 201336 705173 201352
rect 711579 201301 711595 201600
rect 714175 201398 714225 201600
rect 714425 201398 714475 201600
rect 680215 201232 680815 201282
rect 698017 201232 698053 201260
rect 692428 201162 693028 201212
rect 698030 201198 698077 201232
rect 698017 201164 698053 201198
rect 680215 201056 680815 201112
rect 692428 201006 693028 201134
rect 698030 201130 698077 201164
rect 698017 201096 698053 201130
rect 698030 201062 698077 201096
rect 698017 200983 698053 201062
rect 698084 200983 698120 201260
rect 714781 201191 714863 201600
rect 714686 201123 714863 201191
rect 714645 201089 714863 201123
rect 680215 200880 680815 200936
rect 686719 200893 686739 200917
rect 686743 200893 686753 200917
rect 686719 200859 686757 200893
rect 686719 200822 686739 200859
rect 686743 200822 686753 200859
rect 692428 200850 693028 200978
rect 698017 200947 698210 200983
rect 698084 200935 698210 200947
rect 702756 200959 703645 200983
rect 702756 200935 702853 200959
rect 698084 200828 702853 200935
rect 686719 200788 686757 200822
rect 680215 200704 680815 200760
rect 686719 200751 686739 200788
rect 686743 200751 686753 200788
rect 686719 200741 686757 200751
rect 686699 200717 686767 200741
rect 686719 200704 686739 200717
rect 686743 200704 686753 200717
rect 686719 200695 686753 200704
rect 686719 200693 686743 200695
rect 692428 200694 693028 200750
rect 686685 200656 686709 200680
rect 686743 200656 686767 200680
rect 678799 200503 679399 200553
rect 680215 200534 680815 200584
rect 692428 200538 693028 200666
rect 680593 200531 680815 200534
rect 682009 200501 682069 200516
rect 682024 200465 682054 200501
rect 683708 200387 684308 200437
rect 678799 200327 679399 200383
rect 692428 200382 693028 200510
rect 714781 200308 714863 201089
rect 715063 200609 715145 201600
rect 715289 200777 715339 201600
rect 715633 200777 715683 201600
rect 715382 200672 715422 200756
rect 715542 200672 715582 200756
rect 715342 200632 715382 200672
rect 715582 200632 715622 200672
rect 715815 200609 715897 201600
rect 715134 200387 715828 200469
rect 716100 200308 716182 201600
rect 716385 200609 716467 201600
rect 716599 200777 716649 201600
rect 716943 200777 716993 201600
rect 716700 200672 716740 200756
rect 716860 200672 716900 200756
rect 716660 200632 716700 200672
rect 716900 200632 716940 200672
rect 717137 200609 717219 201600
rect 716454 200387 717148 200469
rect 717419 200308 717501 201600
rect 683708 200237 684308 200287
rect 692428 200232 693028 200282
rect 678799 200157 679399 200207
rect 684565 200160 684790 200168
rect 696597 200000 696600 200120
rect 714964 200095 715998 200177
rect 716284 200095 717318 200177
rect 21000 173000 21003 173120
rect 282 172623 1316 172705
rect 1602 172623 2636 172705
rect 32810 172662 33035 172670
rect 38201 172593 38801 172643
rect 24572 172518 25172 172568
rect 33292 172513 33892 172563
rect 99 170574 181 172492
rect 452 172331 1146 172413
rect 381 170885 463 172191
rect 660 172128 700 172168
rect 900 172128 940 172168
rect 700 172044 740 172128
rect 860 172044 900 172128
rect 607 171081 657 172023
rect 951 171081 1001 172023
rect 1133 170885 1215 172191
rect 452 170763 1146 170845
rect 1418 170574 1500 172492
rect 1772 172331 2466 172413
rect 1703 170885 1785 172191
rect 1978 172128 2018 172168
rect 2218 172128 2258 172168
rect 2018 172044 2058 172128
rect 2178 172044 2218 172128
rect 1917 171081 1967 172023
rect 2261 171081 2311 172023
rect 2455 170885 2537 172191
rect 2737 171779 2819 172492
rect 24572 172362 25172 172490
rect 38201 172417 38801 172473
rect 33292 172363 33892 172413
rect 24572 172206 25172 172334
rect 35546 172299 35576 172335
rect 36785 172329 36935 172341
rect 35531 172284 35591 172299
rect 36785 172216 37385 172266
rect 38201 172247 38801 172297
rect 30833 172120 30857 172144
rect 30891 172120 30915 172144
rect 24572 172050 25172 172106
rect 30857 172105 30881 172107
rect 30857 172096 30887 172105
rect 30867 172083 30887 172096
rect 30891 172083 30907 172120
rect 30833 172059 30857 172083
rect 30867 172049 30911 172083
rect 14747 171865 19516 171972
rect 24572 171894 25172 172022
rect 30867 172012 30887 172049
rect 30891 172012 30907 172049
rect 36785 172040 37385 172096
rect 30867 171978 30911 172012
rect 30867 171941 30887 171978
rect 30891 171941 30907 171978
rect 30867 171907 30911 171941
rect 30867 171883 30887 171907
rect 30891 171883 30907 171907
rect 14747 171841 14844 171865
rect 13955 171817 14844 171841
rect 19390 171853 19516 171865
rect 19390 171841 19583 171853
rect 19390 171817 19605 171841
rect 19639 171817 19673 171841
rect 19707 171817 19741 171841
rect 19775 171817 19809 171841
rect 19843 171817 19877 171841
rect 19911 171817 19945 171841
rect 19979 171817 20013 171841
rect 20047 171817 20081 171841
rect 20115 171817 20149 171841
rect 20183 171817 20217 171841
rect 20251 171817 20285 171841
rect 20319 171817 20353 171841
rect 20387 171817 20421 171841
rect 20455 171817 20489 171841
rect 20523 171817 20557 171841
rect 20591 171817 20625 171841
rect 20659 171817 20693 171841
rect 2737 171711 2914 171779
rect 1772 170763 2466 170845
rect 2737 170574 2819 171711
rect 2848 171677 2955 171711
rect 19480 171540 19516 171817
rect 19547 171540 19583 171817
rect 24572 171738 25172 171866
rect 36785 171864 37385 171920
rect 36785 171688 37385 171744
rect 20809 171650 20833 171684
rect 20809 171582 20833 171616
rect 24572 171588 25172 171638
rect 20809 171540 20833 171548
rect 36785 171518 37385 171568
rect 3125 170802 3175 171402
rect 3375 170802 3425 171402
rect 282 170471 1316 170553
rect 1602 170471 2636 170553
rect 1389 170444 1392 170445
rect 1389 170443 1390 170444
rect 1391 170443 1392 170444
rect 1389 170442 1392 170443
rect 1526 170444 1529 170445
rect 1526 170443 1527 170444
rect 1528 170443 1529 170444
rect 2848 170443 2955 170477
rect 1526 170442 1529 170443
rect 5488 170280 5538 171103
rect 5658 170280 5708 171103
rect 6005 170280 6021 171499
rect 12427 171448 12493 171464
rect 24572 171458 25172 171508
rect 32930 171457 33530 171507
rect 35287 171391 35887 171441
rect 36785 171402 37385 171452
rect 24572 171308 25172 171358
rect 31463 171307 32063 171357
rect 32930 171301 33530 171357
rect 7389 171277 7406 171287
rect 7440 171277 7477 171287
rect 7511 171277 7551 171287
rect 7585 171277 7622 171287
rect 7656 171277 7696 171287
rect 7730 171277 7767 171287
rect 7801 171277 7841 171287
rect 7875 171277 7912 171287
rect 7946 171277 7986 171287
rect 8020 171277 8057 171287
rect 8091 171277 8131 171287
rect 8165 171277 8202 171287
rect 8236 171277 8296 171287
rect 8330 171277 8381 171287
rect 8996 171277 9044 171287
rect 9078 171277 9120 171287
rect 9154 171277 9197 171287
rect 9231 171277 9291 171287
rect 9325 171277 9362 171287
rect 9396 171277 9436 171287
rect 9470 171277 9507 171287
rect 9541 171277 9581 171287
rect 9615 171277 9652 171287
rect 9686 171277 9726 171287
rect 9760 171277 9797 171287
rect 9831 171277 9871 171287
rect 9905 171277 9942 171287
rect 9976 171277 9990 171287
rect 7389 171209 8389 171277
rect 8990 171183 9990 171277
rect 36785 171226 37385 171282
rect 15678 171127 16678 171177
rect 17278 171127 18278 171177
rect 31463 171151 32063 171207
rect 32930 171151 33530 171201
rect 34079 171157 34679 171207
rect 7389 170840 8389 170864
rect 15678 170860 16678 170916
rect 17278 170860 18278 170916
rect 8990 170840 9990 170841
rect 7389 170743 8389 170799
rect 8990 170743 9990 170799
rect 15678 170788 16678 170844
rect 17278 170788 18278 170844
rect 8990 170701 9990 170702
rect 15678 170286 16678 170426
rect 17278 170286 18278 170426
rect 19844 170280 19894 171051
rect 20462 170280 20512 171051
rect 31463 171001 32063 171051
rect 34079 171001 34679 171057
rect 35287 171039 35887 171095
rect 36785 171050 37385 171106
rect 32596 170929 33596 170979
rect 24573 170820 25173 170870
rect 34079 170851 34679 170901
rect 35287 170869 35887 170919
rect 36785 170880 37385 170930
rect 30171 170795 30771 170845
rect 32596 170773 33596 170829
rect 37993 170704 38593 170754
rect 30171 170619 30771 170675
rect 32596 170623 33596 170673
rect 34110 170589 34710 170639
rect 21263 170280 21313 170518
rect 22349 170280 22399 170518
rect 32596 170507 33596 170557
rect 30171 170449 30771 170499
rect 36785 170429 36985 170609
rect 37993 170534 38593 170584
rect 24573 170352 25173 170408
rect 29993 170310 30993 170360
rect 31347 170280 31547 170317
rect 31607 170280 31807 170317
rect 36785 170280 36985 170373
rect 37083 170280 37120 170373
rect 696597 168200 696600 168320
rect 692376 167983 692396 168017
rect 692463 167993 692532 168017
rect 696191 167993 696239 168017
rect 692487 167983 692532 167993
rect 696204 167983 696239 167993
rect 696340 167983 696360 168017
rect 692487 167915 692502 167939
rect 696200 167915 696215 167939
rect 692454 167891 692478 167915
rect 696224 167891 696248 167915
rect 686755 167800 687355 167850
rect 692487 167748 692505 167752
rect 692479 167718 692505 167748
rect 692487 167698 692505 167718
rect 686755 167624 687355 167680
rect 692485 167674 692505 167698
rect 692509 167674 692517 167718
rect 696215 167698 696223 167748
rect 696203 167674 696223 167698
rect 696227 167674 696245 167752
rect 692485 167640 692521 167674
rect 696203 167640 696249 167674
rect 686755 167448 687355 167504
rect 686755 167278 687355 167328
rect 685547 167102 686147 167152
rect 687155 167007 687170 167022
rect 687343 167018 687355 167022
rect 687340 167007 687355 167018
rect 685547 166932 686147 166982
rect 687155 166827 687355 167007
rect 687155 166812 687170 166827
rect 687340 166816 687355 166827
rect 687343 166812 687355 166816
rect 687042 166771 687057 166786
rect 687020 166591 687057 166771
rect 687155 166771 687170 166786
rect 687343 166782 687355 166786
rect 687340 166771 687355 166782
rect 687155 166591 687355 166771
rect 688210 166630 688260 167630
rect 688360 166740 688488 167630
rect 688516 166740 688644 167630
rect 688672 166740 688800 167630
rect 688828 166740 688956 167630
rect 688984 166740 689112 167630
rect 689140 166740 689268 167630
rect 689296 166740 689424 167630
rect 689452 166740 689580 167630
rect 689608 166740 689736 167630
rect 689764 166740 689892 167630
rect 689920 166740 690048 167630
rect 690076 166740 690204 167630
rect 690232 166740 690360 167630
rect 690388 166630 690438 167630
rect 692485 167606 692505 167640
rect 692509 167606 692517 167640
rect 696203 167606 696223 167640
rect 696227 167606 696245 167640
rect 691275 167523 691875 167573
rect 692485 167572 692521 167606
rect 696203 167572 696249 167606
rect 692485 167538 692505 167572
rect 692509 167538 692517 167572
rect 692485 167504 692521 167538
rect 692583 167528 693983 167571
rect 694719 167528 696119 167571
rect 696203 167538 696223 167572
rect 696227 167538 696245 167572
rect 696203 167504 696249 167538
rect 692485 167470 692505 167504
rect 692509 167470 692517 167504
rect 692485 167436 692521 167470
rect 691275 167373 691875 167423
rect 692485 167402 692505 167436
rect 692509 167402 692517 167436
rect 692485 167368 692521 167402
rect 692485 167334 692505 167368
rect 692509 167334 692517 167368
rect 692583 167365 693983 167493
rect 694719 167365 696119 167493
rect 696203 167470 696223 167504
rect 696227 167470 696245 167504
rect 696203 167436 696249 167470
rect 707624 167441 707658 167475
rect 707695 167441 707729 167475
rect 707769 167441 707803 167475
rect 707840 167441 707874 167475
rect 707914 167441 707948 167475
rect 707985 167441 708019 167475
rect 708059 167441 708093 167475
rect 708130 167441 708164 167475
rect 708204 167441 708238 167475
rect 708275 167441 708309 167475
rect 708369 167441 708403 167475
rect 708446 167441 708480 167475
rect 708520 167441 708554 167465
rect 708588 167441 708610 167465
rect 709211 167441 709234 167465
rect 709270 167441 709304 167475
rect 709364 167441 709398 167475
rect 709435 167441 709469 167475
rect 709509 167441 709543 167475
rect 709580 167441 709614 167475
rect 709654 167441 709688 167475
rect 709725 167441 709759 167475
rect 709799 167441 709833 167475
rect 709870 167441 709904 167475
rect 709944 167441 709978 167475
rect 710015 167441 710049 167475
rect 710089 167441 710123 167475
rect 710160 167441 710194 167475
rect 696203 167402 696223 167436
rect 696227 167402 696245 167436
rect 707610 167431 707624 167441
rect 707658 167431 707695 167441
rect 707729 167431 707769 167441
rect 707803 167431 707840 167441
rect 707874 167431 707914 167441
rect 707948 167431 707985 167441
rect 708019 167431 708059 167441
rect 708093 167431 708130 167441
rect 708164 167431 708204 167441
rect 708238 167431 708275 167441
rect 708309 167431 708369 167441
rect 708403 167431 708446 167441
rect 708480 167431 708520 167441
rect 708554 167431 708588 167441
rect 708610 167431 708634 167441
rect 709211 167431 709270 167441
rect 709304 167431 709364 167441
rect 709398 167431 709435 167441
rect 709469 167431 709509 167441
rect 709543 167431 709580 167441
rect 709614 167431 709654 167441
rect 709688 167431 709725 167441
rect 709759 167431 709799 167441
rect 709833 167431 709870 167441
rect 709904 167431 709944 167441
rect 709978 167431 710015 167441
rect 710049 167431 710089 167441
rect 710123 167431 710160 167441
rect 710194 167431 710211 167441
rect 696203 167368 696249 167402
rect 696203 167334 696223 167368
rect 696227 167334 696245 167368
rect 707610 167337 708610 167431
rect 709211 167337 710211 167431
rect 691275 167251 691875 167301
rect 692485 167300 692521 167334
rect 692485 167266 692505 167300
rect 692509 167266 692517 167300
rect 692485 167232 692521 167266
rect 692485 167198 692505 167232
rect 692509 167198 692517 167232
rect 692583 167202 693983 167330
rect 694719 167202 696119 167330
rect 696203 167300 696249 167334
rect 711579 167317 712463 167331
rect 711579 167307 711619 167317
rect 696203 167266 696223 167300
rect 696227 167266 696245 167300
rect 701730 167290 701747 167292
rect 696203 167232 696249 167266
rect 696203 167198 696223 167232
rect 696227 167198 696245 167232
rect 701692 167220 701722 167254
rect 701730 167220 701760 167290
rect 707610 167241 708610 167301
rect 709211 167241 710211 167301
rect 692485 167164 692521 167198
rect 691275 167101 691875 167151
rect 692485 167130 692505 167164
rect 692509 167130 692517 167164
rect 692485 167096 692521 167130
rect 692485 167062 692505 167096
rect 692509 167062 692517 167096
rect 692485 167028 692521 167062
rect 692583 167039 693983 167167
rect 694719 167039 696119 167167
rect 696203 167164 696249 167198
rect 696203 167130 696223 167164
rect 696227 167130 696245 167164
rect 696203 167096 696249 167130
rect 696203 167062 696223 167096
rect 696227 167062 696245 167096
rect 699322 167064 700322 167097
rect 700922 167064 701922 167097
rect 696203 167028 696249 167062
rect 707610 167044 708610 167048
rect 709211 167044 710211 167048
rect 691275 166975 691875 167025
rect 692485 166994 692505 167028
rect 692509 166994 692517 167028
rect 692485 166960 692521 166994
rect 692485 166926 692505 166960
rect 692509 166926 692517 166960
rect 692485 166892 692521 166926
rect 691275 166825 691875 166875
rect 692485 166858 692505 166892
rect 692509 166858 692517 166892
rect 692583 166876 693983 167004
rect 694719 166876 696119 167004
rect 696203 166994 696223 167028
rect 696227 166994 696245 167028
rect 707574 166994 708646 167030
rect 696203 166960 696249 166994
rect 696203 166926 696223 166960
rect 696227 166926 696245 166960
rect 707574 166953 707610 166994
rect 708610 166953 708646 166994
rect 696203 166892 696249 166926
rect 697284 166894 697350 166910
rect 707574 166897 708646 166953
rect 696203 166858 696223 166892
rect 696227 166858 696245 166892
rect 699322 166877 700322 166894
rect 700922 166877 701922 166894
rect 707574 166881 707610 166897
rect 708610 166881 708646 166897
rect 692485 166824 692521 166858
rect 692485 166790 692505 166824
rect 692509 166790 692517 166824
rect 692485 166756 692521 166790
rect 691275 166703 691875 166753
rect 692485 166740 692505 166756
rect 692509 166740 692517 166756
rect 692583 166740 693983 166841
rect 694719 166740 696119 166841
rect 696203 166824 696249 166858
rect 707574 166825 708646 166881
rect 696203 166790 696223 166824
rect 696227 166790 696245 166824
rect 696203 166756 696249 166790
rect 696203 166740 696223 166756
rect 696227 166740 696245 166756
rect 699322 166740 700322 166811
rect 700922 166740 701922 166811
rect 707574 166788 707610 166825
rect 708610 166788 708646 166825
rect 707574 166748 708646 166788
rect 709175 166994 710247 167030
rect 709175 166953 709211 166994
rect 710211 166953 710247 166994
rect 709175 166897 710247 166953
rect 709175 166881 709211 166897
rect 710211 166881 710247 166897
rect 709175 166825 710247 166881
rect 709175 166788 709211 166825
rect 710211 166788 710247 166825
rect 709175 166748 710247 166788
rect 685542 166506 686142 166556
rect 691275 166553 691875 166603
rect 685542 166330 686142 166386
rect 692583 166237 693983 166280
rect 694719 166237 696119 166280
rect 699322 166278 700322 166418
rect 700922 166278 701922 166418
rect 685542 166160 686142 166210
rect 692583 166101 693983 166144
rect 694719 166101 696119 166144
rect 680215 165678 680815 165728
rect 680215 165502 680815 165558
rect 685551 165516 686551 165566
rect 689154 165480 689204 165897
rect 689304 165480 689360 165897
rect 689460 165480 689516 165897
rect 689616 165480 689672 165897
rect 689772 165480 689828 165897
rect 689928 165480 689978 165897
rect 699322 165860 700322 165916
rect 700922 165860 701922 165916
rect 707610 165905 708610 165961
rect 709211 165905 710211 165961
rect 699322 165788 700322 165844
rect 700922 165788 701922 165844
rect 707610 165833 708610 165889
rect 709211 165833 710211 165889
rect 711579 165525 711605 167307
rect 715956 166297 716006 167297
rect 716106 166740 716234 167297
rect 716262 166297 716312 167297
rect 711579 165480 711595 165495
rect 712409 165480 712431 165485
rect 713640 165480 713641 165785
rect 713750 165772 714750 165822
rect 713750 165562 714750 165612
rect 713750 165480 714750 165496
rect 2850 159304 3850 159320
rect 2850 159188 3850 159238
rect 2850 158978 3850 159028
rect 3959 159015 3960 159320
rect 5169 159315 5191 159320
rect 6005 159305 6021 159320
rect 1288 157503 1338 158503
rect 1438 157503 1566 158060
rect 1594 157503 1644 158503
rect 5995 157493 6021 159275
rect 7389 158911 8389 158967
rect 8990 158911 9990 158967
rect 15678 158956 16678 159012
rect 17278 158956 18278 159012
rect 7389 158839 8389 158895
rect 8990 158839 9990 158895
rect 15678 158884 16678 158940
rect 17278 158884 18278 158940
rect 27622 158903 27672 159320
rect 27772 158903 27828 159320
rect 27928 158903 27984 159320
rect 28084 158903 28140 159320
rect 28240 158903 28296 159320
rect 28396 158903 28446 159320
rect 31049 159234 32049 159284
rect 36785 159242 37385 159298
rect 36785 159072 37385 159122
rect 21481 158656 22881 158699
rect 23617 158656 25017 158699
rect 31458 158590 32058 158640
rect 15678 158382 16678 158522
rect 17278 158382 18278 158522
rect 21481 158520 22881 158563
rect 23617 158520 25017 158563
rect 31458 158414 32058 158470
rect 25725 158197 26325 158247
rect 31458 158244 32058 158294
rect 7353 158016 8425 158052
rect 7353 157975 7389 158016
rect 8389 157975 8425 158016
rect 7353 157919 8425 157975
rect 7353 157903 7389 157919
rect 8389 157903 8425 157919
rect 7353 157847 8425 157903
rect 7353 157810 7389 157847
rect 8389 157810 8425 157847
rect 7353 157770 8425 157810
rect 8954 158016 10026 158052
rect 8954 157975 8990 158016
rect 9990 157975 10026 158016
rect 8954 157919 10026 157975
rect 21383 158044 21403 158060
rect 21407 158044 21415 158060
rect 21383 158010 21419 158044
rect 21481 158031 22881 158060
rect 23617 158031 25017 158060
rect 25101 158044 25121 158060
rect 25125 158044 25143 158060
rect 25725 158047 26325 158097
rect 25101 158010 25147 158044
rect 21383 157976 21403 158010
rect 21407 157976 21415 158010
rect 21383 157942 21419 157976
rect 8954 157903 8990 157919
rect 9990 157903 10026 157919
rect 15678 157906 16678 157923
rect 17278 157906 18278 157923
rect 21383 157908 21403 157942
rect 21407 157908 21415 157942
rect 8954 157847 10026 157903
rect 20250 157890 20316 157906
rect 8954 157810 8990 157847
rect 9990 157810 10026 157847
rect 8954 157770 10026 157810
rect 21383 157874 21419 157908
rect 21383 157840 21403 157874
rect 21407 157840 21415 157874
rect 21481 157868 22881 157996
rect 23617 157868 25017 157996
rect 25101 157976 25121 158010
rect 25125 157976 25143 158010
rect 25101 157942 25147 157976
rect 25101 157908 25121 157942
rect 25125 157908 25143 157942
rect 25725 157925 26325 157975
rect 25101 157874 25147 157908
rect 25101 157840 25121 157874
rect 25125 157840 25143 157874
rect 21383 157806 21419 157840
rect 21383 157772 21403 157806
rect 21407 157772 21415 157806
rect 21383 157738 21419 157772
rect 15678 157703 16678 157736
rect 17278 157703 18278 157736
rect 21383 157704 21403 157738
rect 21407 157704 21415 157738
rect 21481 157705 22881 157833
rect 23617 157705 25017 157833
rect 25101 157806 25147 157840
rect 25101 157772 25121 157806
rect 25125 157772 25143 157806
rect 25725 157775 26325 157825
rect 25101 157738 25147 157772
rect 25101 157704 25121 157738
rect 25125 157704 25143 157738
rect 21383 157670 21419 157704
rect 25101 157670 25147 157704
rect 21383 157636 21403 157670
rect 21407 157636 21415 157670
rect 7389 157559 8389 157631
rect 8990 157559 9990 157631
rect 21383 157602 21419 157636
rect 15840 157510 15870 157580
rect 15878 157546 15908 157580
rect 21383 157568 21403 157602
rect 21407 157568 21415 157602
rect 15853 157508 15870 157510
rect 21383 157534 21419 157568
rect 21481 157542 22881 157670
rect 23617 157542 25017 157670
rect 25101 157636 25121 157670
rect 25125 157636 25143 157670
rect 25725 157649 26325 157699
rect 25101 157602 25147 157636
rect 25101 157568 25121 157602
rect 25125 157568 25143 157602
rect 25101 157534 25147 157568
rect 5981 157483 6021 157493
rect 5137 157469 6021 157483
rect 21383 157500 21403 157534
rect 21407 157500 21415 157534
rect 21383 157466 21419 157500
rect 7389 157369 8389 157463
rect 7389 157359 8413 157369
rect 8990 157359 9990 157463
rect 21383 157432 21403 157466
rect 21407 157432 21415 157466
rect 21383 157398 21419 157432
rect 21383 157364 21403 157398
rect 21407 157364 21415 157398
rect 21481 157379 22881 157507
rect 23617 157379 25017 157507
rect 25101 157500 25121 157534
rect 25125 157500 25143 157534
rect 25101 157466 25147 157500
rect 25725 157499 26325 157549
rect 25101 157432 25121 157466
rect 25125 157432 25143 157466
rect 25101 157398 25147 157432
rect 25101 157364 25121 157398
rect 25125 157364 25143 157398
rect 25725 157377 26325 157427
rect 21383 157330 21419 157364
rect 25101 157330 25147 157364
rect 21383 157296 21403 157330
rect 21407 157296 21415 157330
rect 25101 157296 25121 157330
rect 25125 157296 25143 157330
rect 21383 157262 21419 157296
rect 21383 157228 21403 157262
rect 21407 157228 21415 157262
rect 21481 157229 22881 157272
rect 23617 157229 25017 157272
rect 25101 157262 25147 157296
rect 25101 157228 25121 157262
rect 25125 157228 25143 157262
rect 21383 157194 21419 157228
rect 25101 157194 25147 157228
rect 25725 157227 26325 157277
rect 21383 157160 21403 157194
rect 21407 157160 21415 157194
rect 25101 157160 25121 157194
rect 25125 157160 25143 157194
rect 27162 157170 27212 158170
rect 27312 157170 27440 158060
rect 27468 157170 27596 158060
rect 27624 157170 27752 158060
rect 27780 157170 27908 158060
rect 27936 157170 28064 158060
rect 28092 157170 28220 158060
rect 28248 157170 28376 158060
rect 28404 157170 28532 158060
rect 28560 157170 28688 158060
rect 28716 157170 28844 158060
rect 28872 157170 29000 158060
rect 29028 157170 29156 158060
rect 29184 157170 29312 158060
rect 29340 157170 29390 158170
rect 30245 158029 30445 158209
rect 30245 158018 30260 158029
rect 30245 158014 30257 158018
rect 30430 158014 30445 158029
rect 30543 158029 30580 158209
rect 30543 158014 30558 158029
rect 30245 157984 30257 157988
rect 30245 157973 30260 157984
rect 30430 157973 30445 157988
rect 30245 157793 30445 157973
rect 31453 157818 32053 157868
rect 30245 157782 30260 157793
rect 30245 157778 30257 157782
rect 30430 157778 30445 157793
rect 31453 157648 32053 157698
rect 30245 157472 30845 157522
rect 30245 157296 30845 157352
rect 21383 157126 21419 157160
rect 25101 157126 25147 157160
rect 21383 157102 21403 157126
rect 21385 157048 21403 157102
rect 21407 157082 21415 157126
rect 25101 157102 25121 157126
rect 25113 157082 25121 157102
rect 25125 157048 25143 157126
rect 30245 157120 30845 157176
rect 30245 156950 30845 157000
rect 21000 156800 21003 156920
rect 21352 156885 21376 156909
rect 25122 156885 25146 156909
rect 21385 156861 21400 156885
rect 25098 156861 25113 156885
rect 21274 156783 21294 156851
rect 21410 156817 21430 156851
rect 25068 156817 25088 156851
rect 25204 156817 25224 156851
rect 21385 156807 21430 156817
rect 25102 156807 25137 156817
rect 21361 156783 21430 156807
rect 25089 156783 25137 156807
rect 25238 156783 25258 156817
rect 680480 154427 680517 154520
rect 680615 154427 680815 154520
rect 685793 154483 685993 154520
rect 686053 154483 686253 154520
rect 686607 154440 687607 154490
rect 692427 154392 693027 154448
rect 679007 154216 679607 154266
rect 680615 154191 680815 154371
rect 686829 154301 687429 154351
rect 684004 154243 685004 154293
rect 695201 154282 695251 154520
rect 696287 154282 696337 154520
rect 682890 154161 683490 154211
rect 684004 154127 685004 154177
rect 686829 154125 687429 154181
rect 679007 154046 679607 154096
rect 684004 153971 685004 154027
rect 686829 153955 687429 154005
rect 680215 153870 680815 153920
rect 681713 153881 682313 153931
rect 682921 153899 683521 153949
rect 692427 153930 693027 153980
rect 684004 153821 685004 153871
rect 680215 153694 680815 153750
rect 681713 153705 682313 153761
rect 682921 153743 683521 153799
rect 685537 153749 686137 153799
rect 697088 153749 697138 154520
rect 697706 153749 697756 154520
rect 699322 154374 700322 154514
rect 700922 154374 701922 154514
rect 707610 154098 708610 154099
rect 699322 153956 700322 154012
rect 700922 153956 701922 154012
rect 707610 154001 708610 154057
rect 709211 154001 710211 154057
rect 707610 153959 708610 153960
rect 699322 153884 700322 153940
rect 700922 153884 701922 153940
rect 709211 153936 710211 153960
rect 682921 153593 683521 153643
rect 684070 153599 684670 153649
rect 685537 153593 686137 153649
rect 699322 153623 700322 153673
rect 700922 153623 701922 153673
rect 680215 153518 680815 153574
rect 707610 153523 708610 153617
rect 709211 153523 710211 153591
rect 707610 153513 707624 153523
rect 707658 153513 707695 153523
rect 707729 153513 707769 153523
rect 707803 153513 707840 153523
rect 707874 153513 707914 153523
rect 707948 153513 707985 153523
rect 708019 153513 708059 153523
rect 708093 153513 708130 153523
rect 708164 153513 708204 153523
rect 708238 153513 708275 153523
rect 708309 153513 708369 153523
rect 708403 153513 708446 153523
rect 708480 153513 708522 153523
rect 708556 153513 708604 153523
rect 709219 153513 709270 153523
rect 709304 153513 709364 153523
rect 709398 153513 709435 153523
rect 709469 153513 709509 153523
rect 709543 153513 709580 153523
rect 709614 153513 709654 153523
rect 709688 153513 709725 153523
rect 709759 153513 709799 153523
rect 709833 153513 709870 153523
rect 709904 153513 709944 153523
rect 709978 153513 710015 153523
rect 710049 153513 710089 153523
rect 710123 153513 710160 153523
rect 710194 153513 710211 153523
rect 684070 153443 684670 153499
rect 685537 153443 686137 153493
rect 692428 153442 693028 153492
rect 680215 153348 680815 153398
rect 681713 153359 682313 153409
rect 684070 153293 684670 153343
rect 692428 153292 693028 153342
rect 705107 153336 705173 153352
rect 711579 153301 711595 154520
rect 711892 153697 711942 154520
rect 712062 153697 712112 154520
rect 716071 154357 716074 154358
rect 714645 154323 714752 154357
rect 716071 154356 716072 154357
rect 716073 154356 716074 154357
rect 716071 154355 716074 154356
rect 716208 154357 716211 154358
rect 716208 154356 716209 154357
rect 716210 154356 716211 154357
rect 716208 154355 716211 154356
rect 714964 154247 715998 154329
rect 716284 154247 717318 154329
rect 714175 153398 714225 153998
rect 714425 153398 714475 153998
rect 680215 153232 680815 153282
rect 698017 153232 698053 153260
rect 692428 153162 693028 153212
rect 698030 153198 698077 153232
rect 698017 153164 698053 153198
rect 680215 153056 680815 153112
rect 692428 153006 693028 153134
rect 698030 153130 698077 153164
rect 698017 153096 698053 153130
rect 698030 153062 698077 153096
rect 698017 152983 698053 153062
rect 698084 152983 698120 153260
rect 714781 153191 714863 154226
rect 715134 153955 715828 154037
rect 714686 153123 714863 153191
rect 714645 153089 714863 153123
rect 680215 152880 680815 152936
rect 686719 152893 686739 152917
rect 686743 152893 686753 152917
rect 686719 152859 686757 152893
rect 686719 152822 686739 152859
rect 686743 152822 686753 152859
rect 692428 152850 693028 152978
rect 698017 152947 698210 152983
rect 698084 152935 698210 152947
rect 702756 152959 703645 152983
rect 702756 152935 702853 152959
rect 698084 152828 702853 152935
rect 686719 152788 686757 152822
rect 680215 152704 680815 152760
rect 686719 152751 686739 152788
rect 686743 152751 686753 152788
rect 686719 152741 686757 152751
rect 686699 152717 686767 152741
rect 686719 152704 686739 152717
rect 686743 152704 686753 152717
rect 686719 152695 686753 152704
rect 686719 152693 686743 152695
rect 692428 152694 693028 152750
rect 686685 152656 686709 152680
rect 686743 152656 686767 152680
rect 678799 152503 679399 152553
rect 680215 152534 680815 152584
rect 692428 152538 693028 152666
rect 680593 152531 680815 152534
rect 682009 152501 682069 152516
rect 682024 152465 682054 152501
rect 683708 152387 684308 152437
rect 678799 152327 679399 152383
rect 692428 152382 693028 152510
rect 714781 152308 714863 153089
rect 715063 152609 715145 153915
rect 715289 152777 715339 153719
rect 715633 152777 715683 153719
rect 715382 152672 715422 152756
rect 715542 152672 715582 152756
rect 715342 152632 715382 152672
rect 715582 152632 715622 152672
rect 715815 152609 715897 153915
rect 715134 152387 715828 152469
rect 716100 152308 716182 154226
rect 716454 153955 717148 154037
rect 716385 152609 716467 153915
rect 716599 152777 716649 153719
rect 716943 152777 716993 153719
rect 716700 152672 716740 152756
rect 716860 152672 716900 152756
rect 716660 152632 716700 152672
rect 716900 152632 716940 152672
rect 717137 152609 717219 153915
rect 716454 152387 717148 152469
rect 717419 152308 717501 154226
rect 683708 152237 684308 152287
rect 692428 152232 693028 152282
rect 678799 152157 679399 152207
rect 684565 152160 684790 152168
rect 696597 152000 696600 152120
rect 714964 152095 715998 152177
rect 716284 152095 717318 152177
rect 21000 125000 21003 125120
rect 282 124623 1316 124705
rect 1602 124623 2636 124705
rect 32810 124662 33035 124670
rect 38201 124593 38801 124643
rect 24572 124518 25172 124568
rect 33292 124513 33892 124563
rect 99 122574 181 124492
rect 452 124331 1146 124413
rect 381 122885 463 124191
rect 660 124128 700 124168
rect 900 124128 940 124168
rect 700 124044 740 124128
rect 860 124044 900 124128
rect 607 123081 657 124023
rect 951 123081 1001 124023
rect 1133 122885 1215 124191
rect 452 122763 1146 122845
rect 1418 122574 1500 124492
rect 1772 124331 2466 124413
rect 1703 122885 1785 124191
rect 1978 124128 2018 124168
rect 2218 124128 2258 124168
rect 2018 124044 2058 124128
rect 2178 124044 2218 124128
rect 1917 123081 1967 124023
rect 2261 123081 2311 124023
rect 2455 122885 2537 124191
rect 2737 123779 2819 124492
rect 24572 124362 25172 124490
rect 38201 124417 38801 124473
rect 33292 124363 33892 124413
rect 24572 124206 25172 124334
rect 35546 124299 35576 124335
rect 36785 124329 36935 124341
rect 35531 124284 35591 124299
rect 36785 124216 37385 124266
rect 38201 124247 38801 124297
rect 30833 124120 30857 124144
rect 30891 124120 30915 124144
rect 24572 124050 25172 124106
rect 30857 124105 30881 124107
rect 30857 124096 30887 124105
rect 30867 124083 30887 124096
rect 30891 124083 30907 124120
rect 30833 124059 30857 124083
rect 30867 124049 30911 124083
rect 14747 123865 19516 123972
rect 24572 123894 25172 124022
rect 30867 124012 30887 124049
rect 30891 124012 30907 124049
rect 36785 124040 37385 124096
rect 30867 123978 30911 124012
rect 30867 123941 30887 123978
rect 30891 123941 30907 123978
rect 30867 123907 30911 123941
rect 30867 123883 30887 123907
rect 30891 123883 30907 123907
rect 14747 123841 14844 123865
rect 13955 123817 14844 123841
rect 19390 123853 19516 123865
rect 19390 123841 19583 123853
rect 19390 123817 19605 123841
rect 19639 123817 19673 123841
rect 19707 123817 19741 123841
rect 19775 123817 19809 123841
rect 19843 123817 19877 123841
rect 19911 123817 19945 123841
rect 19979 123817 20013 123841
rect 20047 123817 20081 123841
rect 20115 123817 20149 123841
rect 20183 123817 20217 123841
rect 20251 123817 20285 123841
rect 20319 123817 20353 123841
rect 20387 123817 20421 123841
rect 20455 123817 20489 123841
rect 20523 123817 20557 123841
rect 20591 123817 20625 123841
rect 20659 123817 20693 123841
rect 2737 123711 2914 123779
rect 1772 122763 2466 122845
rect 2737 122574 2819 123711
rect 2848 123677 2955 123711
rect 19480 123540 19516 123817
rect 19547 123540 19583 123817
rect 24572 123738 25172 123866
rect 36785 123864 37385 123920
rect 36785 123688 37385 123744
rect 20809 123650 20833 123684
rect 20809 123582 20833 123616
rect 24572 123588 25172 123638
rect 20809 123540 20833 123548
rect 36785 123518 37385 123568
rect 3125 122802 3175 123402
rect 3375 122802 3425 123402
rect 282 122471 1316 122553
rect 1602 122471 2636 122553
rect 1389 122444 1392 122445
rect 1389 122443 1390 122444
rect 1391 122443 1392 122444
rect 1389 122442 1392 122443
rect 1526 122444 1529 122445
rect 1526 122443 1527 122444
rect 1528 122443 1529 122444
rect 2848 122443 2955 122477
rect 1526 122442 1529 122443
rect 5488 122280 5538 123103
rect 5658 122280 5708 123103
rect 6005 122280 6021 123499
rect 12427 123448 12493 123464
rect 24572 123458 25172 123508
rect 32930 123457 33530 123507
rect 35287 123391 35887 123441
rect 36785 123402 37385 123452
rect 24572 123308 25172 123358
rect 31463 123307 32063 123357
rect 32930 123301 33530 123357
rect 7389 123277 7406 123287
rect 7440 123277 7477 123287
rect 7511 123277 7551 123287
rect 7585 123277 7622 123287
rect 7656 123277 7696 123287
rect 7730 123277 7767 123287
rect 7801 123277 7841 123287
rect 7875 123277 7912 123287
rect 7946 123277 7986 123287
rect 8020 123277 8057 123287
rect 8091 123277 8131 123287
rect 8165 123277 8202 123287
rect 8236 123277 8296 123287
rect 8330 123277 8381 123287
rect 8996 123277 9044 123287
rect 9078 123277 9120 123287
rect 9154 123277 9197 123287
rect 9231 123277 9291 123287
rect 9325 123277 9362 123287
rect 9396 123277 9436 123287
rect 9470 123277 9507 123287
rect 9541 123277 9581 123287
rect 9615 123277 9652 123287
rect 9686 123277 9726 123287
rect 9760 123277 9797 123287
rect 9831 123277 9871 123287
rect 9905 123277 9942 123287
rect 9976 123277 9990 123287
rect 7389 123209 8389 123277
rect 8990 123183 9990 123277
rect 36785 123226 37385 123282
rect 15678 123127 16678 123177
rect 17278 123127 18278 123177
rect 31463 123151 32063 123207
rect 32930 123151 33530 123201
rect 34079 123157 34679 123207
rect 7389 122840 8389 122864
rect 15678 122860 16678 122916
rect 17278 122860 18278 122916
rect 8990 122840 9990 122841
rect 7389 122743 8389 122799
rect 8990 122743 9990 122799
rect 15678 122788 16678 122844
rect 17278 122788 18278 122844
rect 8990 122701 9990 122702
rect 15678 122286 16678 122426
rect 17278 122286 18278 122426
rect 19844 122280 19894 123051
rect 20462 122280 20512 123051
rect 31463 123001 32063 123051
rect 34079 123001 34679 123057
rect 35287 123039 35887 123095
rect 36785 123050 37385 123106
rect 32596 122929 33596 122979
rect 24573 122820 25173 122870
rect 34079 122851 34679 122901
rect 35287 122869 35887 122919
rect 36785 122880 37385 122930
rect 30171 122795 30771 122845
rect 32596 122773 33596 122829
rect 37993 122704 38593 122754
rect 30171 122619 30771 122675
rect 32596 122623 33596 122673
rect 34110 122589 34710 122639
rect 21263 122280 21313 122518
rect 22349 122280 22399 122518
rect 32596 122507 33596 122557
rect 30171 122449 30771 122499
rect 36785 122429 36985 122609
rect 37993 122534 38593 122584
rect 24573 122352 25173 122408
rect 29993 122310 30993 122360
rect 31347 122280 31547 122317
rect 31607 122280 31807 122317
rect 36785 122280 36985 122373
rect 37083 122280 37120 122373
rect 696597 120200 696600 120320
rect 692376 119983 692396 120017
rect 692463 119993 692532 120017
rect 696191 119993 696239 120017
rect 692487 119983 692532 119993
rect 696204 119983 696239 119993
rect 696340 119983 696360 120017
rect 692487 119915 692502 119939
rect 696200 119915 696215 119939
rect 692454 119891 692478 119915
rect 696224 119891 696248 119915
rect 686755 119800 687355 119850
rect 692487 119748 692505 119752
rect 692479 119718 692505 119748
rect 692487 119698 692505 119718
rect 686755 119624 687355 119680
rect 692485 119674 692505 119698
rect 692509 119674 692517 119718
rect 696215 119698 696223 119748
rect 696203 119674 696223 119698
rect 696227 119674 696245 119752
rect 692485 119640 692521 119674
rect 696203 119640 696249 119674
rect 686755 119448 687355 119504
rect 686755 119278 687355 119328
rect 685547 119102 686147 119152
rect 687155 119007 687170 119022
rect 687343 119018 687355 119022
rect 687340 119007 687355 119018
rect 685547 118932 686147 118982
rect 687155 118827 687355 119007
rect 687155 118812 687170 118827
rect 687340 118816 687355 118827
rect 687343 118812 687355 118816
rect 687042 118771 687057 118786
rect 687020 118591 687057 118771
rect 687042 118576 687057 118591
rect 687155 118771 687170 118786
rect 687343 118782 687355 118786
rect 687340 118771 687355 118782
rect 687155 118591 687355 118771
rect 688210 118630 688260 119630
rect 688360 118630 688488 119630
rect 688516 118630 688644 119630
rect 688672 118630 688800 119630
rect 688828 118630 688956 119630
rect 688984 118630 689112 119630
rect 689140 118630 689268 119630
rect 689296 118630 689424 119630
rect 689452 118630 689580 119630
rect 689608 118630 689736 119630
rect 689764 118630 689892 119630
rect 689920 118630 690048 119630
rect 690076 118630 690204 119630
rect 690232 118630 690360 119630
rect 690388 118630 690438 119630
rect 692485 119606 692505 119640
rect 692509 119606 692517 119640
rect 696203 119606 696223 119640
rect 696227 119606 696245 119640
rect 691275 119523 691875 119573
rect 692485 119572 692521 119606
rect 696203 119572 696249 119606
rect 692485 119538 692505 119572
rect 692509 119538 692517 119572
rect 692485 119504 692521 119538
rect 692583 119528 693983 119571
rect 694719 119528 696119 119571
rect 696203 119538 696223 119572
rect 696227 119538 696245 119572
rect 696203 119504 696249 119538
rect 692485 119470 692505 119504
rect 692509 119470 692517 119504
rect 692485 119436 692521 119470
rect 691275 119373 691875 119423
rect 692485 119402 692505 119436
rect 692509 119402 692517 119436
rect 692485 119368 692521 119402
rect 692485 119334 692505 119368
rect 692509 119334 692517 119368
rect 692583 119365 693983 119493
rect 694719 119365 696119 119493
rect 696203 119470 696223 119504
rect 696227 119470 696245 119504
rect 696203 119436 696249 119470
rect 707624 119441 707658 119475
rect 707695 119441 707729 119475
rect 707769 119441 707803 119475
rect 707840 119441 707874 119475
rect 707914 119441 707948 119475
rect 707985 119441 708019 119475
rect 708059 119441 708093 119475
rect 708130 119441 708164 119475
rect 708204 119441 708238 119475
rect 708275 119441 708309 119475
rect 708369 119441 708403 119475
rect 708446 119441 708480 119475
rect 708520 119441 708554 119465
rect 708588 119441 708610 119465
rect 709211 119441 709234 119465
rect 709270 119441 709304 119475
rect 709364 119441 709398 119475
rect 709435 119441 709469 119475
rect 709509 119441 709543 119475
rect 709580 119441 709614 119475
rect 709654 119441 709688 119475
rect 709725 119441 709759 119475
rect 709799 119441 709833 119475
rect 709870 119441 709904 119475
rect 709944 119441 709978 119475
rect 710015 119441 710049 119475
rect 710089 119441 710123 119475
rect 710160 119441 710194 119475
rect 696203 119402 696223 119436
rect 696227 119402 696245 119436
rect 707610 119431 707624 119441
rect 707658 119431 707695 119441
rect 707729 119431 707769 119441
rect 707803 119431 707840 119441
rect 707874 119431 707914 119441
rect 707948 119431 707985 119441
rect 708019 119431 708059 119441
rect 708093 119431 708130 119441
rect 708164 119431 708204 119441
rect 708238 119431 708275 119441
rect 708309 119431 708369 119441
rect 708403 119431 708446 119441
rect 708480 119431 708520 119441
rect 708554 119431 708588 119441
rect 708610 119431 708634 119441
rect 709211 119431 709270 119441
rect 709304 119431 709364 119441
rect 709398 119431 709435 119441
rect 709469 119431 709509 119441
rect 709543 119431 709580 119441
rect 709614 119431 709654 119441
rect 709688 119431 709725 119441
rect 709759 119431 709799 119441
rect 709833 119431 709870 119441
rect 709904 119431 709944 119441
rect 709978 119431 710015 119441
rect 710049 119431 710089 119441
rect 710123 119431 710160 119441
rect 710194 119431 710211 119441
rect 696203 119368 696249 119402
rect 696203 119334 696223 119368
rect 696227 119334 696245 119368
rect 707610 119337 708610 119431
rect 709211 119337 710211 119431
rect 691275 119251 691875 119301
rect 692485 119300 692521 119334
rect 692485 119266 692505 119300
rect 692509 119266 692517 119300
rect 692485 119232 692521 119266
rect 692485 119198 692505 119232
rect 692509 119198 692517 119232
rect 692583 119202 693983 119330
rect 694719 119202 696119 119330
rect 696203 119300 696249 119334
rect 711579 119317 712463 119331
rect 711579 119307 711619 119317
rect 696203 119266 696223 119300
rect 696227 119266 696245 119300
rect 701730 119290 701747 119292
rect 696203 119232 696249 119266
rect 696203 119198 696223 119232
rect 696227 119198 696245 119232
rect 701692 119220 701722 119254
rect 701730 119220 701760 119290
rect 707610 119241 708610 119301
rect 709211 119241 710211 119301
rect 692485 119164 692521 119198
rect 691275 119101 691875 119151
rect 692485 119130 692505 119164
rect 692509 119130 692517 119164
rect 692485 119096 692521 119130
rect 692485 119062 692505 119096
rect 692509 119062 692517 119096
rect 692485 119028 692521 119062
rect 692583 119039 693983 119167
rect 694719 119039 696119 119167
rect 696203 119164 696249 119198
rect 696203 119130 696223 119164
rect 696227 119130 696245 119164
rect 696203 119096 696249 119130
rect 696203 119062 696223 119096
rect 696227 119062 696245 119096
rect 699322 119064 700322 119097
rect 700922 119064 701922 119097
rect 696203 119028 696249 119062
rect 707610 119044 708610 119048
rect 709211 119044 710211 119048
rect 691275 118975 691875 119025
rect 692485 118994 692505 119028
rect 692509 118994 692517 119028
rect 692485 118960 692521 118994
rect 692485 118926 692505 118960
rect 692509 118926 692517 118960
rect 692485 118892 692521 118926
rect 691275 118825 691875 118875
rect 692485 118858 692505 118892
rect 692509 118858 692517 118892
rect 692583 118876 693983 119004
rect 694719 118876 696119 119004
rect 696203 118994 696223 119028
rect 696227 118994 696245 119028
rect 707574 118994 708646 119030
rect 696203 118960 696249 118994
rect 696203 118926 696223 118960
rect 696227 118926 696245 118960
rect 707574 118953 707610 118994
rect 708610 118953 708646 118994
rect 696203 118892 696249 118926
rect 697284 118894 697350 118910
rect 707574 118897 708646 118953
rect 696203 118858 696223 118892
rect 696227 118858 696245 118892
rect 699322 118877 700322 118894
rect 700922 118877 701922 118894
rect 707574 118881 707610 118897
rect 708610 118881 708646 118897
rect 692485 118824 692521 118858
rect 692485 118790 692505 118824
rect 692509 118790 692517 118824
rect 692485 118756 692521 118790
rect 691275 118703 691875 118753
rect 692485 118722 692505 118756
rect 692509 118722 692517 118756
rect 692485 118688 692521 118722
rect 692583 118713 693983 118841
rect 694719 118713 696119 118841
rect 696203 118824 696249 118858
rect 707574 118825 708646 118881
rect 696203 118790 696223 118824
rect 696227 118790 696245 118824
rect 696203 118756 696249 118790
rect 696203 118722 696223 118756
rect 696227 118722 696245 118756
rect 699322 118739 700322 118811
rect 700922 118739 701922 118811
rect 707574 118788 707610 118825
rect 708610 118788 708646 118825
rect 707574 118748 708646 118788
rect 709175 118994 710247 119030
rect 709175 118953 709211 118994
rect 710211 118953 710247 118994
rect 709175 118897 710247 118953
rect 709175 118881 709211 118897
rect 710211 118881 710247 118897
rect 709175 118825 710247 118881
rect 709175 118788 709211 118825
rect 710211 118788 710247 118825
rect 709175 118748 710247 118788
rect 696203 118688 696249 118722
rect 692485 118654 692505 118688
rect 692509 118654 692517 118688
rect 692485 118620 692521 118654
rect 687155 118576 687170 118591
rect 687340 118580 687355 118591
rect 687343 118576 687355 118580
rect 685542 118506 686142 118556
rect 691275 118553 691875 118603
rect 692485 118586 692505 118620
rect 692509 118586 692517 118620
rect 692485 118552 692521 118586
rect 692485 118518 692505 118552
rect 692509 118518 692517 118552
rect 692583 118550 693983 118678
rect 694719 118550 696119 118678
rect 696203 118654 696223 118688
rect 696227 118654 696245 118688
rect 696203 118620 696249 118654
rect 696203 118586 696223 118620
rect 696227 118586 696245 118620
rect 696203 118552 696249 118586
rect 696203 118518 696223 118552
rect 696227 118518 696245 118552
rect 692485 118484 692521 118518
rect 692485 118450 692505 118484
rect 692509 118450 692517 118484
rect 692485 118416 692521 118450
rect 679817 118330 679841 118354
rect 685542 118330 686142 118386
rect 692485 118382 692505 118416
rect 692509 118382 692517 118416
rect 692583 118387 693983 118515
rect 694719 118387 696119 118515
rect 696203 118484 696249 118518
rect 696203 118450 696223 118484
rect 696227 118450 696245 118484
rect 699322 118478 700322 118550
rect 700922 118478 701922 118550
rect 707610 118523 708610 118595
rect 709211 118523 710211 118595
rect 699392 118467 699426 118478
rect 699460 118467 699494 118478
rect 699528 118467 699562 118478
rect 699596 118467 699630 118478
rect 699664 118467 699698 118478
rect 699732 118467 699766 118478
rect 699800 118467 699834 118478
rect 699868 118467 699902 118478
rect 699936 118467 699970 118478
rect 700004 118467 700038 118478
rect 700072 118467 700106 118478
rect 700140 118467 700174 118478
rect 700208 118467 700242 118478
rect 700276 118467 700310 118478
rect 700934 118467 700968 118478
rect 701002 118467 701036 118478
rect 701070 118467 701104 118478
rect 701138 118467 701172 118478
rect 701206 118467 701240 118478
rect 701274 118467 701308 118478
rect 701342 118467 701376 118478
rect 701410 118467 701444 118478
rect 701478 118467 701512 118478
rect 701546 118467 701580 118478
rect 701614 118467 701648 118478
rect 701682 118467 701716 118478
rect 701750 118467 701784 118478
rect 701818 118467 701852 118478
rect 699392 118457 699450 118467
rect 699460 118457 699518 118467
rect 699528 118457 699586 118467
rect 699596 118457 699654 118467
rect 699664 118457 699722 118467
rect 699732 118457 699790 118467
rect 699800 118457 699858 118467
rect 699868 118457 699926 118467
rect 699936 118457 699994 118467
rect 700004 118457 700062 118467
rect 700072 118457 700130 118467
rect 700140 118457 700198 118467
rect 700208 118457 700266 118467
rect 700276 118457 700334 118467
rect 700934 118457 700992 118467
rect 701002 118457 701060 118467
rect 701070 118457 701128 118467
rect 701138 118457 701196 118467
rect 701206 118457 701264 118467
rect 701274 118457 701332 118467
rect 701342 118457 701400 118467
rect 701410 118457 701468 118467
rect 701478 118457 701536 118467
rect 701546 118457 701604 118467
rect 701614 118457 701672 118467
rect 701682 118457 701740 118467
rect 701750 118457 701808 118467
rect 701818 118457 701876 118467
rect 696203 118416 696249 118450
rect 699368 118433 700334 118457
rect 700910 118433 701876 118457
rect 699392 118418 699416 118433
rect 699460 118418 699484 118433
rect 699528 118418 699552 118433
rect 699596 118418 699620 118433
rect 699664 118418 699688 118433
rect 699732 118418 699756 118433
rect 699800 118418 699824 118433
rect 699868 118418 699892 118433
rect 699936 118418 699960 118433
rect 700004 118418 700028 118433
rect 700072 118418 700096 118433
rect 700140 118418 700164 118433
rect 700208 118418 700232 118433
rect 700276 118418 700300 118433
rect 700934 118418 700958 118433
rect 701002 118418 701026 118433
rect 701070 118418 701094 118433
rect 701138 118418 701162 118433
rect 701206 118418 701230 118433
rect 701274 118418 701298 118433
rect 701342 118418 701366 118433
rect 701410 118418 701434 118433
rect 701478 118418 701502 118433
rect 701546 118418 701570 118433
rect 701614 118418 701638 118433
rect 701682 118418 701706 118433
rect 701750 118418 701774 118433
rect 701818 118418 701842 118433
rect 696203 118382 696223 118416
rect 696227 118382 696245 118416
rect 692485 118348 692521 118382
rect 696203 118348 696249 118382
rect 679549 118307 679573 118330
rect 679793 118306 679808 118330
rect 692485 118314 692505 118348
rect 692509 118314 692517 118348
rect 696203 118314 696223 118348
rect 696227 118314 696245 118348
rect 692485 118280 692521 118314
rect 696203 118280 696249 118314
rect 679549 118237 679573 118271
rect 692485 118246 692505 118280
rect 692509 118246 692517 118280
rect 692485 118212 692521 118246
rect 692583 118237 693983 118280
rect 694719 118237 696119 118280
rect 696203 118246 696223 118280
rect 696227 118246 696245 118280
rect 699322 118263 700322 118418
rect 696203 118212 696249 118246
rect 699322 118229 700334 118263
rect 700922 118253 701922 118418
rect 700910 118229 701922 118253
rect 699322 118218 700322 118229
rect 700922 118218 701922 118229
rect 707574 118263 708646 118299
rect 707574 118226 707610 118263
rect 708610 118226 708646 118263
rect 679549 118167 679573 118201
rect 685542 118160 686142 118210
rect 685601 118157 685895 118160
rect 685920 118157 686142 118160
rect 692485 118178 692505 118212
rect 692509 118178 692517 118212
rect 696203 118178 696223 118212
rect 696227 118178 696245 118212
rect 699392 118205 699416 118218
rect 699460 118205 699484 118218
rect 699528 118205 699552 118218
rect 699596 118205 699620 118218
rect 699664 118205 699688 118218
rect 699732 118205 699756 118218
rect 699800 118205 699824 118218
rect 699868 118205 699892 118218
rect 699936 118205 699960 118218
rect 700004 118205 700028 118218
rect 700072 118205 700096 118218
rect 700140 118205 700164 118218
rect 700208 118205 700232 118218
rect 700276 118205 700300 118218
rect 700934 118205 700958 118218
rect 701002 118205 701026 118218
rect 701070 118205 701094 118218
rect 701138 118205 701162 118218
rect 701206 118205 701230 118218
rect 701274 118205 701298 118218
rect 701342 118205 701366 118218
rect 701410 118205 701434 118218
rect 701478 118205 701502 118218
rect 701546 118205 701570 118218
rect 701614 118205 701638 118218
rect 701682 118205 701706 118218
rect 701750 118205 701774 118218
rect 701818 118205 701842 118218
rect 707574 118186 708646 118226
rect 709175 118263 710247 118299
rect 709175 118226 709211 118263
rect 710211 118226 710247 118263
rect 709175 118186 710247 118226
rect 692485 118144 692521 118178
rect 696203 118144 696249 118178
rect 679549 118097 679573 118131
rect 692485 118110 692505 118144
rect 692509 118110 692517 118144
rect 692485 118076 692521 118110
rect 692583 118101 693983 118144
rect 694719 118101 696119 118144
rect 696203 118110 696223 118144
rect 696227 118110 696245 118144
rect 696203 118076 696249 118110
rect 679549 118027 679573 118061
rect 692485 118042 692505 118076
rect 692509 118042 692517 118076
rect 692485 118008 692521 118042
rect 679549 117957 679573 117991
rect 692485 117974 692505 118008
rect 692509 117974 692517 118008
rect 679793 117933 679808 117957
rect 692485 117940 692521 117974
rect 679817 117909 679841 117933
rect 692485 117906 692505 117940
rect 692509 117906 692517 117940
rect 692583 117938 693983 118066
rect 694719 117938 696119 118066
rect 696203 118042 696223 118076
rect 696227 118042 696245 118076
rect 696203 118008 696249 118042
rect 696203 117974 696223 118008
rect 696227 117974 696245 118008
rect 696203 117940 696249 117974
rect 696203 117906 696223 117940
rect 696227 117906 696245 117940
rect 687685 117838 687709 117862
rect 687661 117814 687675 117838
rect 687669 117797 687675 117814
rect 679515 117762 679539 117785
rect 679613 117762 679637 117785
rect 679491 117737 679515 117761
rect 679637 117737 679661 117761
rect 680215 117678 680815 117728
rect 680215 117502 680815 117558
rect 685551 117516 686551 117566
rect 680215 117326 680815 117382
rect 685551 117360 686551 117488
rect 689154 117439 689204 117897
rect 689151 117355 689204 117439
rect 680215 117156 680815 117206
rect 685551 117204 686551 117332
rect 685551 117048 686551 117176
rect 686865 117116 687465 117166
rect 679007 116980 679607 117030
rect 680615 116885 680630 116900
rect 680803 116896 680815 116900
rect 680800 116885 680815 116896
rect 685551 116892 686551 116948
rect 686865 116940 687465 117068
rect 679007 116810 679607 116860
rect 680615 116705 680815 116885
rect 683328 116793 683928 116843
rect 682573 116717 683173 116767
rect 680615 116690 680630 116705
rect 680800 116694 680815 116705
rect 680803 116690 680815 116694
rect 680502 116649 680517 116664
rect 680480 116469 680517 116649
rect 680502 116454 680517 116469
rect 680615 116649 680630 116664
rect 680803 116660 680815 116664
rect 680800 116649 680815 116660
rect 680615 116469 680815 116649
rect 682573 116541 683173 116669
rect 683328 116617 683928 116745
rect 685551 116736 686551 116864
rect 686865 116764 687465 116820
rect 685551 116580 686551 116708
rect 686865 116588 687465 116716
rect 680615 116454 680630 116469
rect 680800 116458 680815 116469
rect 680803 116454 680815 116458
rect 683328 116441 683928 116497
rect 679002 116384 679602 116434
rect 685551 116424 686551 116552
rect 682573 116365 683173 116421
rect 686865 116412 687465 116468
rect 679002 116208 679602 116264
rect 682573 116189 683173 116317
rect 683328 116265 683928 116321
rect 685551 116274 686551 116324
rect 686865 116236 687465 116364
rect 685551 116158 686551 116208
rect 678680 116123 678704 116157
rect 678680 116055 678704 116089
rect 679002 116038 679602 116088
rect 679061 116035 679355 116038
rect 679380 116035 679602 116038
rect 678680 115987 678704 116021
rect 682573 116013 683173 116141
rect 683328 116089 683928 116145
rect 678680 115919 678704 115953
rect 678680 115851 678704 115885
rect 682573 115837 683173 115965
rect 683328 115913 683928 116041
rect 685551 115982 686551 116110
rect 686865 116060 687465 116116
rect 678680 115783 678704 115817
rect 685551 115806 686551 115934
rect 686865 115884 687465 116012
rect 678680 115715 678704 115749
rect 678680 115647 678704 115681
rect 682573 115661 683173 115789
rect 683328 115737 683928 115793
rect 685551 115630 686551 115758
rect 686865 115708 687465 115836
rect 678680 115579 678704 115613
rect 683328 115567 683928 115617
rect 678680 115511 678704 115545
rect 682573 115491 683173 115541
rect 684519 115498 685119 115548
rect 678680 115443 678704 115477
rect 685551 115454 686551 115582
rect 686865 115532 687465 115660
rect 679133 115409 679283 115421
rect 679452 115409 679602 115421
rect 678680 115375 678704 115409
rect 678680 115307 678704 115341
rect 679002 115296 679602 115346
rect 684519 115342 685119 115398
rect 685551 115278 686551 115406
rect 686865 115356 687465 115484
rect 678680 115239 678704 115273
rect 678680 115171 678704 115205
rect 684519 115192 685119 115242
rect 678680 115103 678704 115137
rect 679002 115120 679602 115176
rect 681745 115081 682345 115131
rect 682509 115069 683109 115119
rect 678680 115035 678704 115069
rect 683739 115027 684339 115077
rect 684519 115062 685119 115112
rect 685551 115102 686551 115230
rect 686865 115180 687465 115308
rect 678680 114967 678704 115001
rect 679002 114950 679602 115000
rect 678680 114899 678704 114933
rect 680502 114915 680517 114930
rect 678680 114831 678704 114865
rect 678680 114763 678704 114797
rect 680480 114735 680517 114915
rect 678680 114695 678704 114729
rect 680502 114720 680517 114735
rect 680615 114915 680630 114930
rect 680803 114926 680815 114930
rect 680800 114915 680815 114926
rect 681745 114925 682345 114981
rect 680615 114735 680815 114915
rect 681745 114769 682345 114897
rect 682509 114893 683109 115021
rect 684519 114906 685119 115034
rect 685551 114926 686551 115054
rect 686865 115004 687465 115060
rect 683739 114837 684339 114893
rect 686865 114828 687465 114956
rect 680615 114720 680630 114735
rect 680800 114724 680815 114735
rect 680803 114720 680815 114724
rect 680615 114679 680630 114694
rect 680803 114690 680815 114694
rect 680800 114679 680815 114690
rect 678680 114627 678704 114661
rect 678680 114559 678704 114593
rect 678680 114491 678704 114525
rect 679007 114524 679607 114574
rect 680615 114499 680815 114679
rect 681745 114613 682345 114741
rect 682509 114717 683109 114773
rect 684519 114750 685119 114806
rect 685551 114750 686551 114806
rect 682509 114541 683109 114669
rect 684519 114594 685119 114722
rect 685551 114594 686551 114722
rect 686865 114652 687465 114780
rect 680615 114484 680630 114499
rect 680800 114488 680815 114499
rect 680803 114484 680815 114488
rect 681745 114463 682345 114513
rect 683739 114477 684339 114513
rect 678680 114423 678704 114457
rect 684519 114444 685119 114494
rect 685551 114438 686551 114566
rect 686865 114476 687465 114604
rect 678680 114355 678704 114389
rect 679007 114354 679607 114404
rect 682509 114371 683109 114421
rect 678680 114287 678704 114321
rect 684519 114314 685119 114364
rect 678680 114219 678704 114253
rect 678680 114151 678704 114185
rect 680215 114178 680815 114228
rect 681745 114209 682345 114259
rect 678680 114083 678704 114117
rect 678680 114015 678704 114049
rect 680215 114002 680815 114058
rect 681745 114053 682345 114181
rect 682509 114030 683109 114080
rect 678680 113947 678704 113981
rect 678680 113879 678704 113913
rect 681745 113897 682345 113953
rect 678680 113811 678704 113845
rect 680215 113826 680815 113882
rect 678680 113743 678704 113777
rect 681745 113741 682345 113869
rect 682509 113854 683109 113910
rect 678680 113675 678704 113709
rect 680215 113656 680815 113706
rect 682509 113684 683109 113734
rect 683248 113680 683298 114268
rect 683398 113680 683448 114268
rect 684519 114158 685119 114286
rect 685551 114282 686551 114410
rect 686865 114300 687465 114428
rect 684519 114002 685119 114130
rect 685551 114126 686551 114254
rect 686865 114124 687465 114252
rect 685551 113970 686551 114098
rect 686865 113954 687465 114004
rect 684519 113852 685119 113902
rect 685551 113814 686551 113870
rect 686865 113838 687465 113888
rect 683248 113668 683448 113680
rect 685551 113658 686551 113786
rect 686865 113662 687465 113790
rect 678680 113607 678704 113641
rect 681745 113591 682345 113641
rect 683571 113605 683581 113646
rect 678680 113539 678704 113573
rect 680215 113524 680815 113574
rect 682509 113555 683509 113605
rect 678680 113471 678704 113505
rect 685551 113502 686551 113630
rect 686865 113486 687465 113542
rect 678680 113403 678704 113437
rect 678680 113335 678704 113369
rect 680215 113348 680815 113404
rect 681745 113389 682345 113439
rect 682509 113385 683509 113435
rect 683278 113382 683398 113385
rect 683571 113382 683581 113385
rect 685551 113346 686551 113474
rect 678680 113267 678704 113301
rect 678680 113199 678704 113233
rect 680215 113172 680815 113228
rect 681745 113213 682345 113341
rect 682509 113247 683109 113297
rect 678680 113131 678704 113165
rect 678680 113063 678704 113097
rect 678654 113013 678680 113039
rect 680215 113002 680815 113052
rect 681745 113037 682345 113093
rect 682509 113071 683109 113127
rect 678680 112929 678704 112963
rect 678680 112861 678704 112895
rect 678680 112793 678704 112827
rect 679007 112826 679607 112876
rect 681745 112867 682345 112917
rect 682509 112901 683109 112951
rect 678680 112725 678704 112759
rect 680615 112731 680630 112746
rect 680803 112742 680815 112746
rect 680800 112731 680815 112742
rect 678680 112657 678704 112691
rect 679007 112656 679607 112706
rect 678680 112589 678704 112623
rect 678680 112521 678704 112555
rect 680615 112551 680815 112731
rect 681345 112651 682345 112701
rect 682508 112631 683108 112681
rect 680615 112536 680630 112551
rect 680800 112540 680815 112551
rect 680803 112536 680815 112540
rect 680502 112495 680517 112510
rect 678680 112453 678704 112487
rect 678680 112385 678704 112419
rect 678680 112317 678704 112351
rect 680480 112315 680517 112495
rect 680502 112300 680517 112315
rect 680615 112495 680630 112510
rect 680803 112506 680815 112510
rect 680800 112495 680815 112506
rect 680615 112315 680815 112495
rect 681345 112475 682345 112531
rect 682508 112455 683108 112511
rect 680615 112300 680630 112315
rect 680800 112304 680815 112315
rect 680803 112300 680815 112304
rect 681345 112299 682345 112427
rect 682508 112285 683108 112335
rect 683228 112322 683278 113322
rect 683398 112322 683448 113322
rect 685551 113190 686551 113318
rect 686865 113310 687465 113438
rect 685551 113034 686551 113162
rect 686865 113140 687465 113190
rect 686865 113024 687465 113074
rect 685551 112884 686551 112934
rect 686865 112848 687465 112976
rect 685551 112768 686551 112818
rect 686865 112672 687465 112800
rect 684404 112609 685004 112659
rect 685551 112612 686551 112668
rect 685551 112456 686551 112512
rect 686865 112496 687465 112624
rect 685551 112300 686551 112356
rect 686865 112320 687465 112376
rect 678680 112249 678704 112283
rect 679002 112230 679602 112280
rect 678680 112181 678704 112215
rect 678680 112113 678704 112147
rect 681345 112129 682345 112179
rect 684404 112175 685004 112225
rect 685551 112150 686551 112200
rect 686865 112150 687465 112200
rect 678680 112045 678704 112079
rect 679002 112054 679602 112110
rect 681390 112070 681424 112080
rect 681458 112070 681492 112080
rect 681526 112070 681560 112080
rect 681594 112070 681628 112080
rect 681662 112070 681696 112080
rect 681730 112070 681764 112080
rect 681798 112070 681832 112080
rect 681866 112070 681900 112080
rect 681934 112070 681968 112080
rect 682002 112070 682036 112080
rect 682077 112070 682111 112080
rect 682145 112070 682179 112080
rect 682213 112070 682247 112080
rect 682281 112070 682315 112080
rect 681345 112034 682345 112046
rect 678680 111977 678704 112011
rect 678680 111909 678704 111943
rect 679002 111884 679602 111934
rect 681345 111927 682345 111977
rect 684004 111973 685004 112023
rect 685551 112014 686551 112064
rect 686865 112034 687465 112084
rect 679061 111881 679355 111884
rect 679380 111881 679602 111884
rect 678680 111841 678704 111875
rect 678680 111773 678704 111807
rect 681345 111751 682345 111879
rect 684004 111817 685004 111873
rect 685551 111858 686551 111914
rect 686865 111858 687465 111914
rect 686686 111812 686714 111840
rect 678680 111705 678704 111739
rect 678680 111637 678704 111671
rect 678680 111569 678704 111603
rect 681345 111575 682345 111703
rect 684004 111661 685004 111789
rect 685551 111708 686551 111758
rect 686865 111688 687465 111738
rect 678680 111501 678704 111535
rect 684004 111505 685004 111633
rect 687573 111554 687585 117277
rect 689154 117107 689204 117355
rect 689151 117023 689204 117107
rect 689154 116897 689204 117023
rect 689304 116897 689360 117897
rect 689460 116897 689516 117897
rect 689616 116897 689672 117897
rect 689772 116897 689828 117897
rect 689928 116897 689978 117897
rect 692485 117872 692521 117906
rect 692485 117838 692505 117872
rect 692509 117838 692517 117872
rect 690952 117509 691122 117815
rect 692485 117804 692521 117838
rect 692485 117770 692505 117804
rect 692509 117770 692517 117804
rect 692583 117775 693983 117903
rect 694719 117775 696119 117903
rect 696203 117872 696249 117906
rect 696203 117838 696223 117872
rect 696227 117838 696245 117872
rect 699322 117860 700322 117916
rect 700922 117860 701922 117916
rect 707610 117905 708610 117961
rect 709211 117905 710211 117961
rect 696203 117804 696249 117838
rect 696203 117770 696223 117804
rect 696227 117770 696245 117804
rect 699322 117788 700322 117844
rect 700922 117788 701922 117844
rect 707610 117833 708610 117889
rect 709211 117833 710211 117889
rect 692485 117736 692521 117770
rect 692485 117702 692505 117736
rect 692509 117702 692517 117736
rect 692485 117668 692521 117702
rect 692485 117634 692505 117668
rect 692509 117634 692517 117668
rect 692485 117600 692521 117634
rect 692583 117612 693983 117740
rect 694719 117612 696119 117740
rect 696203 117736 696249 117770
rect 696203 117702 696223 117736
rect 696227 117702 696245 117736
rect 696203 117668 696249 117702
rect 696203 117634 696223 117668
rect 696227 117634 696245 117668
rect 696203 117600 696249 117634
rect 692485 117566 692505 117600
rect 692509 117566 692517 117600
rect 692485 117532 692521 117566
rect 692485 117498 692505 117532
rect 692509 117498 692517 117532
rect 692485 117464 692521 117498
rect 692485 117430 692505 117464
rect 692509 117430 692517 117464
rect 692583 117449 693983 117577
rect 694719 117449 696119 117577
rect 696203 117566 696223 117600
rect 696227 117566 696245 117600
rect 696203 117532 696249 117566
rect 696203 117498 696223 117532
rect 696227 117498 696245 117532
rect 696203 117464 696249 117498
rect 699322 117486 700322 117558
rect 700922 117486 701922 117558
rect 707610 117531 708610 117603
rect 709211 117531 710211 117603
rect 711579 117553 711605 119307
rect 715956 118297 716006 119297
rect 716106 118297 716234 119297
rect 716262 118297 716312 119297
rect 699392 117475 699426 117486
rect 699460 117475 699494 117486
rect 699528 117475 699562 117486
rect 699596 117475 699630 117486
rect 699664 117475 699698 117486
rect 699732 117475 699766 117486
rect 699800 117475 699834 117486
rect 699868 117475 699902 117486
rect 699936 117475 699970 117486
rect 700004 117475 700038 117486
rect 700072 117475 700106 117486
rect 700140 117475 700174 117486
rect 700208 117475 700242 117486
rect 700276 117475 700310 117486
rect 700934 117475 700968 117486
rect 701002 117475 701036 117486
rect 701070 117475 701104 117486
rect 701138 117475 701172 117486
rect 701206 117475 701240 117486
rect 701274 117475 701308 117486
rect 701342 117475 701376 117486
rect 701410 117475 701444 117486
rect 701478 117475 701512 117486
rect 701546 117475 701580 117486
rect 701614 117475 701648 117486
rect 701682 117475 701716 117486
rect 701750 117475 701784 117486
rect 701818 117475 701852 117486
rect 711511 117485 711663 117553
rect 712447 117501 712557 117511
rect 711579 117482 711663 117485
rect 699392 117465 699450 117475
rect 699460 117465 699518 117475
rect 699528 117465 699586 117475
rect 699596 117465 699654 117475
rect 699664 117465 699722 117475
rect 699732 117465 699790 117475
rect 699800 117465 699858 117475
rect 699868 117465 699926 117475
rect 699936 117465 699994 117475
rect 700004 117465 700062 117475
rect 700072 117465 700130 117475
rect 700140 117465 700198 117475
rect 700208 117465 700266 117475
rect 700276 117465 700334 117475
rect 700934 117465 700992 117475
rect 701002 117465 701060 117475
rect 701070 117465 701128 117475
rect 701138 117465 701196 117475
rect 701206 117465 701264 117475
rect 701274 117465 701332 117475
rect 701342 117465 701400 117475
rect 701410 117465 701468 117475
rect 701478 117465 701536 117475
rect 701546 117465 701604 117475
rect 701614 117465 701672 117475
rect 701682 117465 701740 117475
rect 701750 117465 701808 117475
rect 701818 117465 701876 117475
rect 696203 117430 696223 117464
rect 696227 117430 696245 117464
rect 699368 117441 700334 117465
rect 700910 117441 701876 117465
rect 711541 117461 711633 117482
rect 692485 117396 692521 117430
rect 692485 117362 692505 117396
rect 692509 117362 692517 117396
rect 692485 117328 692521 117362
rect 692485 117294 692505 117328
rect 692509 117294 692517 117328
rect 692485 117260 692521 117294
rect 692583 117286 693983 117414
rect 694719 117286 696119 117414
rect 696203 117396 696249 117430
rect 699392 117426 699416 117441
rect 699460 117426 699484 117441
rect 699528 117426 699552 117441
rect 699596 117426 699620 117441
rect 699664 117426 699688 117441
rect 699732 117426 699756 117441
rect 699800 117426 699824 117441
rect 699868 117426 699892 117441
rect 699936 117426 699960 117441
rect 700004 117426 700028 117441
rect 700072 117426 700096 117441
rect 700140 117426 700164 117441
rect 700208 117426 700232 117441
rect 700276 117426 700300 117441
rect 700934 117426 700958 117441
rect 701002 117426 701026 117441
rect 701070 117426 701094 117441
rect 701138 117426 701162 117441
rect 701206 117426 701230 117441
rect 701274 117426 701298 117441
rect 701342 117426 701366 117441
rect 701410 117426 701434 117441
rect 701478 117426 701502 117441
rect 701546 117426 701570 117441
rect 701614 117426 701638 117441
rect 701682 117426 701706 117441
rect 701750 117426 701774 117441
rect 701818 117426 701842 117441
rect 696203 117362 696223 117396
rect 696227 117362 696245 117396
rect 696203 117328 696249 117362
rect 696203 117294 696223 117328
rect 696227 117294 696245 117328
rect 696203 117260 696249 117294
rect 699322 117271 700322 117426
rect 692485 117226 692505 117260
rect 692509 117226 692517 117260
rect 692485 117192 692521 117226
rect 692485 117158 692505 117192
rect 692509 117158 692517 117192
rect 692485 117124 692521 117158
rect 692485 117090 692505 117124
rect 692509 117090 692517 117124
rect 692583 117123 693983 117251
rect 694719 117123 696119 117251
rect 696203 117226 696223 117260
rect 696227 117226 696245 117260
rect 699322 117237 700334 117271
rect 700922 117261 701922 117426
rect 707610 117271 708610 117331
rect 709211 117271 710211 117331
rect 700910 117237 701922 117261
rect 699322 117226 700322 117237
rect 700922 117226 701922 117237
rect 696203 117192 696249 117226
rect 699392 117213 699416 117226
rect 699460 117213 699484 117226
rect 699528 117213 699552 117226
rect 699596 117213 699620 117226
rect 699664 117213 699688 117226
rect 699732 117213 699756 117226
rect 699800 117213 699824 117226
rect 699868 117213 699892 117226
rect 699936 117213 699960 117226
rect 700004 117213 700028 117226
rect 700072 117213 700096 117226
rect 700140 117213 700164 117226
rect 700208 117213 700232 117226
rect 700276 117213 700300 117226
rect 700934 117213 700958 117226
rect 701002 117213 701026 117226
rect 701070 117213 701094 117226
rect 701138 117213 701162 117226
rect 701206 117213 701230 117226
rect 701274 117213 701298 117226
rect 701342 117213 701366 117226
rect 701410 117213 701434 117226
rect 701478 117213 701502 117226
rect 701546 117213 701570 117226
rect 701614 117213 701638 117226
rect 701682 117213 701706 117226
rect 701750 117213 701774 117226
rect 701818 117213 701842 117226
rect 696203 117158 696223 117192
rect 696227 117158 696245 117192
rect 696203 117124 696249 117158
rect 696203 117090 696223 117124
rect 696227 117090 696245 117124
rect 692485 117056 692521 117090
rect 696203 117056 696249 117090
rect 692485 117022 692505 117056
rect 692509 117022 692517 117056
rect 696203 117022 696223 117056
rect 696227 117022 696245 117056
rect 692485 116988 692521 117022
rect 692485 116954 692505 116988
rect 692509 116954 692517 116988
rect 692583 116966 693983 117016
rect 694719 116966 696119 117016
rect 696203 116988 696249 117022
rect 696203 116954 696223 116988
rect 696227 116954 696245 116988
rect 692485 116920 692521 116954
rect 696203 116920 696249 116954
rect 692485 116896 692505 116920
rect 692487 116852 692505 116896
rect 692509 116886 692517 116920
rect 696203 116896 696223 116920
rect 696215 116886 696223 116896
rect 696227 116852 696245 116920
rect 697284 116870 697350 116886
rect 699322 116868 700322 116924
rect 700922 116868 701922 116924
rect 707610 116913 708610 116969
rect 709211 116913 710211 116969
rect 692174 116787 692186 116811
rect 692288 116787 692312 116811
rect 696390 116787 696414 116811
rect 696516 116787 696528 116811
rect 699322 116796 700322 116852
rect 700922 116796 701922 116852
rect 707610 116841 708610 116897
rect 709211 116841 710211 116897
rect 692264 116763 692288 116777
rect 696414 116763 696438 116777
rect 692288 116729 692312 116753
rect 696390 116729 696414 116753
rect 688940 116475 688990 116675
rect 689110 116475 689238 116675
rect 689286 116475 689342 116675
rect 689462 116475 689590 116675
rect 689638 116559 689688 116675
rect 692736 116597 695966 116699
rect 689638 116475 689691 116559
rect 699322 116494 700322 116566
rect 700922 116494 701922 116566
rect 707610 116539 708610 116611
rect 709211 116539 710211 116611
rect 699392 116483 699426 116494
rect 699460 116483 699494 116494
rect 699528 116483 699562 116494
rect 699596 116483 699630 116494
rect 699664 116483 699698 116494
rect 699732 116483 699766 116494
rect 699800 116483 699834 116494
rect 699868 116483 699902 116494
rect 699936 116483 699970 116494
rect 700004 116483 700038 116494
rect 700072 116483 700106 116494
rect 700140 116483 700174 116494
rect 700208 116483 700242 116494
rect 700276 116483 700310 116494
rect 700934 116483 700968 116494
rect 701002 116483 701036 116494
rect 701070 116483 701104 116494
rect 701138 116483 701172 116494
rect 701206 116483 701240 116494
rect 701274 116483 701308 116494
rect 701342 116483 701376 116494
rect 701410 116483 701444 116494
rect 701478 116483 701512 116494
rect 701546 116483 701580 116494
rect 701614 116483 701648 116494
rect 701682 116483 701716 116494
rect 701750 116483 701784 116494
rect 701818 116483 701852 116494
rect 689649 116471 689683 116475
rect 699392 116473 699450 116483
rect 699460 116473 699518 116483
rect 699528 116473 699586 116483
rect 699596 116473 699654 116483
rect 699664 116473 699722 116483
rect 699732 116473 699790 116483
rect 699800 116473 699858 116483
rect 699868 116473 699926 116483
rect 699936 116473 699994 116483
rect 700004 116473 700062 116483
rect 700072 116473 700130 116483
rect 700140 116473 700198 116483
rect 700208 116473 700266 116483
rect 700276 116473 700334 116483
rect 700934 116473 700992 116483
rect 701002 116473 701060 116483
rect 701070 116473 701128 116483
rect 701138 116473 701196 116483
rect 701206 116473 701264 116483
rect 701274 116473 701332 116483
rect 701342 116473 701400 116483
rect 701410 116473 701468 116483
rect 701478 116473 701536 116483
rect 701546 116473 701604 116483
rect 701614 116473 701672 116483
rect 701682 116473 701740 116483
rect 701750 116473 701808 116483
rect 701818 116473 701876 116483
rect 692451 116444 692475 116468
rect 692509 116444 692533 116468
rect 696169 116444 696193 116468
rect 696227 116444 696251 116468
rect 699368 116449 700334 116473
rect 700910 116449 701876 116473
rect 692485 116410 692499 116444
rect 696203 116410 696217 116444
rect 699392 116434 699416 116449
rect 699460 116434 699484 116449
rect 699528 116434 699552 116449
rect 699596 116434 699620 116449
rect 699664 116434 699688 116449
rect 699732 116434 699756 116449
rect 699800 116434 699824 116449
rect 699868 116434 699892 116449
rect 699936 116434 699960 116449
rect 700004 116434 700028 116449
rect 700072 116434 700096 116449
rect 700140 116434 700164 116449
rect 700208 116434 700232 116449
rect 700276 116434 700300 116449
rect 700934 116434 700958 116449
rect 701002 116434 701026 116449
rect 701070 116434 701094 116449
rect 701138 116434 701162 116449
rect 701206 116434 701230 116449
rect 701274 116434 701298 116449
rect 701342 116434 701366 116449
rect 701410 116434 701434 116449
rect 701478 116434 701502 116449
rect 701546 116434 701570 116449
rect 701614 116434 701638 116449
rect 701682 116434 701706 116449
rect 701750 116434 701774 116449
rect 701818 116434 701842 116449
rect 692451 116386 692475 116410
rect 692509 116386 692533 116410
rect 696169 116386 696193 116410
rect 696227 116386 696251 116410
rect 690664 116318 691664 116368
rect 692515 116280 693915 116330
rect 694787 116280 696187 116330
rect 699322 116279 700322 116434
rect 699322 116245 700334 116279
rect 700922 116269 701922 116434
rect 703539 116286 703699 116290
rect 707610 116279 708610 116339
rect 709211 116279 710211 116339
rect 700910 116245 701922 116269
rect 690242 116219 690326 116222
rect 690242 116214 690442 116219
rect 690238 116180 690442 116214
rect 690242 116169 690442 116180
rect 690664 116162 691664 116218
rect 687686 116128 687720 116162
rect 687686 116104 687710 116128
rect 689649 116127 689683 116131
rect 688940 115927 688990 116127
rect 689110 115927 689238 116127
rect 689286 115927 689342 116127
rect 689462 115927 689590 116127
rect 689638 116043 689691 116127
rect 689638 115927 689688 116043
rect 690242 115993 690442 116121
rect 692515 116117 693915 116245
rect 694787 116117 696187 116245
rect 699322 116234 700322 116245
rect 700922 116234 701922 116245
rect 699392 116221 699416 116234
rect 699460 116221 699484 116234
rect 699528 116221 699552 116234
rect 699596 116221 699620 116234
rect 699664 116221 699688 116234
rect 699732 116221 699756 116234
rect 699800 116221 699824 116234
rect 699868 116221 699892 116234
rect 699936 116221 699960 116234
rect 700004 116221 700028 116234
rect 700072 116221 700096 116234
rect 700140 116221 700164 116234
rect 700208 116221 700232 116234
rect 700276 116221 700300 116234
rect 700934 116221 700958 116234
rect 701002 116221 701026 116234
rect 701070 116221 701094 116234
rect 701138 116221 701162 116234
rect 701206 116221 701230 116234
rect 701274 116221 701298 116234
rect 701342 116221 701366 116234
rect 701410 116221 701434 116234
rect 701478 116221 701502 116234
rect 701546 116221 701570 116234
rect 701614 116221 701638 116234
rect 701682 116221 701706 116234
rect 701750 116221 701774 116234
rect 701818 116221 701842 116234
rect 703541 116140 703701 116144
rect 690664 116006 691664 116062
rect 692515 115954 693915 116082
rect 694787 115954 696187 116082
rect 690242 115817 690442 115873
rect 690664 115850 691664 115906
rect 692515 115791 693915 115919
rect 694787 115791 696187 115919
rect 699322 115876 700322 115932
rect 700922 115876 701922 115932
rect 707610 115921 708610 115977
rect 709211 115921 710211 115977
rect 699322 115804 700322 115860
rect 700922 115804 701922 115860
rect 707610 115849 708610 115905
rect 709211 115849 710211 115905
rect 689154 115579 689204 115705
rect 687686 115501 687720 115535
rect 687798 115515 687822 115539
rect 687774 115491 687798 115504
rect 689151 115495 689204 115579
rect 687798 115456 687822 115480
rect 689154 115247 689204 115495
rect 689151 115163 689204 115247
rect 689154 114705 689204 115163
rect 689304 114705 689360 115705
rect 689460 114705 689516 115705
rect 689616 114705 689672 115705
rect 689772 114705 689828 115705
rect 689928 114705 689978 115705
rect 690242 115641 690442 115769
rect 690664 115700 691664 115750
rect 690790 115697 690874 115700
rect 691123 115697 691207 115700
rect 692515 115628 693915 115756
rect 694787 115628 696187 115756
rect 704735 115731 705041 115833
rect 704719 115715 705057 115731
rect 690242 115465 690442 115521
rect 692515 115465 693915 115593
rect 694787 115465 696187 115593
rect 699322 115502 700322 115574
rect 700922 115502 701922 115574
rect 707610 115547 708610 115619
rect 709211 115547 710211 115619
rect 699392 115491 699426 115502
rect 699460 115491 699494 115502
rect 699528 115491 699562 115502
rect 699596 115491 699630 115502
rect 699664 115491 699698 115502
rect 699732 115491 699766 115502
rect 699800 115491 699834 115502
rect 699868 115491 699902 115502
rect 699936 115491 699970 115502
rect 700004 115491 700038 115502
rect 700072 115491 700106 115502
rect 700140 115491 700174 115502
rect 700208 115491 700242 115502
rect 700276 115491 700310 115502
rect 700934 115491 700968 115502
rect 701002 115491 701036 115502
rect 701070 115491 701104 115502
rect 701138 115491 701172 115502
rect 701206 115491 701240 115502
rect 701274 115491 701308 115502
rect 701342 115491 701376 115502
rect 701410 115491 701444 115502
rect 701478 115491 701512 115502
rect 701546 115491 701580 115502
rect 701614 115491 701648 115502
rect 701682 115491 701716 115502
rect 701750 115491 701784 115502
rect 701818 115491 701852 115502
rect 699392 115481 699450 115491
rect 699460 115481 699518 115491
rect 699528 115481 699586 115491
rect 699596 115481 699654 115491
rect 699664 115481 699722 115491
rect 699732 115481 699790 115491
rect 699800 115481 699858 115491
rect 699868 115481 699926 115491
rect 699936 115481 699994 115491
rect 700004 115481 700062 115491
rect 700072 115481 700130 115491
rect 700140 115481 700198 115491
rect 700208 115481 700266 115491
rect 700276 115481 700334 115491
rect 700934 115481 700992 115491
rect 701002 115481 701060 115491
rect 701070 115481 701128 115491
rect 701138 115481 701196 115491
rect 701206 115481 701264 115491
rect 701274 115481 701332 115491
rect 701342 115481 701400 115491
rect 701410 115481 701468 115491
rect 701478 115481 701536 115491
rect 701546 115481 701604 115491
rect 701614 115481 701672 115491
rect 701682 115481 701740 115491
rect 701750 115481 701808 115491
rect 701818 115481 701876 115491
rect 699368 115457 700334 115481
rect 700910 115457 701876 115481
rect 699392 115442 699416 115457
rect 699460 115442 699484 115457
rect 699528 115442 699552 115457
rect 699596 115442 699620 115457
rect 699664 115442 699688 115457
rect 699732 115442 699756 115457
rect 699800 115442 699824 115457
rect 699868 115442 699892 115457
rect 699936 115442 699960 115457
rect 700004 115442 700028 115457
rect 700072 115442 700096 115457
rect 700140 115442 700164 115457
rect 700208 115442 700232 115457
rect 700276 115442 700300 115457
rect 700934 115442 700958 115457
rect 701002 115442 701026 115457
rect 701070 115442 701094 115457
rect 701138 115442 701162 115457
rect 701206 115442 701230 115457
rect 701274 115442 701298 115457
rect 701342 115442 701366 115457
rect 701410 115442 701434 115457
rect 701478 115442 701502 115457
rect 701546 115442 701570 115457
rect 701614 115442 701638 115457
rect 701682 115442 701706 115457
rect 701750 115442 701774 115457
rect 701818 115442 701842 115457
rect 690242 115289 690442 115417
rect 692515 115302 693915 115430
rect 694787 115302 696187 115430
rect 690790 115286 690874 115289
rect 691123 115286 691207 115289
rect 699322 115287 700322 115442
rect 690664 115236 691664 115286
rect 699322 115253 700334 115287
rect 700922 115277 701922 115442
rect 707610 115287 708610 115347
rect 709211 115287 710211 115347
rect 700910 115253 701922 115277
rect 699322 115242 700322 115253
rect 700922 115242 701922 115253
rect 699392 115229 699416 115242
rect 699460 115229 699484 115242
rect 699528 115229 699552 115242
rect 699596 115229 699620 115242
rect 699664 115229 699688 115242
rect 699732 115229 699756 115242
rect 699800 115229 699824 115242
rect 699868 115229 699892 115242
rect 699936 115229 699960 115242
rect 700004 115229 700028 115242
rect 700072 115229 700096 115242
rect 700140 115229 700164 115242
rect 700208 115229 700232 115242
rect 700276 115229 700300 115242
rect 700934 115229 700958 115242
rect 701002 115229 701026 115242
rect 701070 115229 701094 115242
rect 701138 115229 701162 115242
rect 701206 115229 701230 115242
rect 701274 115229 701298 115242
rect 701342 115229 701366 115242
rect 701410 115229 701434 115242
rect 701478 115229 701502 115242
rect 701546 115229 701570 115242
rect 701614 115229 701638 115242
rect 701682 115229 701706 115242
rect 701750 115229 701774 115242
rect 701818 115229 701842 115242
rect 690242 115113 690442 115169
rect 692515 115152 693915 115195
rect 694787 115152 696187 115195
rect 690664 115080 691664 115136
rect 690242 114937 690442 115065
rect 692515 115016 693915 115059
rect 694787 115016 696187 115059
rect 690664 114924 691664 114980
rect 692515 114853 693915 114981
rect 694787 114853 696187 114981
rect 703541 114944 703701 114948
rect 699322 114884 700322 114940
rect 700922 114884 701922 114940
rect 707610 114929 708610 114985
rect 709211 114929 710211 114985
rect 690242 114806 690442 114817
rect 690238 114772 690442 114806
rect 690242 114767 690442 114772
rect 690664 114768 691664 114824
rect 690242 114764 690326 114767
rect 692515 114690 693915 114818
rect 694787 114690 696187 114818
rect 699322 114812 700322 114868
rect 700922 114812 701922 114868
rect 707610 114857 708610 114913
rect 709211 114857 710211 114913
rect 703541 114798 703701 114802
rect 690664 114618 691664 114668
rect 692515 114527 693915 114655
rect 694787 114527 696187 114655
rect 699322 114510 700322 114582
rect 700922 114510 701922 114582
rect 707610 114555 708610 114627
rect 709211 114555 710211 114627
rect 699392 114499 699426 114510
rect 699460 114499 699494 114510
rect 699528 114499 699562 114510
rect 699596 114499 699630 114510
rect 699664 114499 699698 114510
rect 699732 114499 699766 114510
rect 699800 114499 699834 114510
rect 699868 114499 699902 114510
rect 699936 114499 699970 114510
rect 700004 114499 700038 114510
rect 700072 114499 700106 114510
rect 700140 114499 700174 114510
rect 700208 114499 700242 114510
rect 700276 114499 700310 114510
rect 700934 114499 700968 114510
rect 701002 114499 701036 114510
rect 701070 114499 701104 114510
rect 701138 114499 701172 114510
rect 701206 114499 701240 114510
rect 701274 114499 701308 114510
rect 701342 114499 701376 114510
rect 701410 114499 701444 114510
rect 701478 114499 701512 114510
rect 701546 114499 701580 114510
rect 701614 114499 701648 114510
rect 701682 114499 701716 114510
rect 701750 114499 701784 114510
rect 701818 114499 701852 114510
rect 692515 114364 693915 114492
rect 694787 114364 696187 114492
rect 699392 114489 699450 114499
rect 699460 114489 699518 114499
rect 699528 114489 699586 114499
rect 699596 114489 699654 114499
rect 699664 114489 699722 114499
rect 699732 114489 699790 114499
rect 699800 114489 699858 114499
rect 699868 114489 699926 114499
rect 699936 114489 699994 114499
rect 700004 114489 700062 114499
rect 700072 114489 700130 114499
rect 700140 114489 700198 114499
rect 700208 114489 700266 114499
rect 700276 114489 700334 114499
rect 700934 114489 700992 114499
rect 701002 114489 701060 114499
rect 701070 114489 701128 114499
rect 701138 114489 701196 114499
rect 701206 114489 701264 114499
rect 701274 114489 701332 114499
rect 701342 114489 701400 114499
rect 701410 114489 701468 114499
rect 701478 114489 701536 114499
rect 701546 114489 701604 114499
rect 701614 114489 701672 114499
rect 701682 114489 701740 114499
rect 701750 114489 701808 114499
rect 701818 114489 701876 114499
rect 699368 114465 700334 114489
rect 700910 114465 701876 114489
rect 699392 114450 699416 114465
rect 699460 114450 699484 114465
rect 699528 114450 699552 114465
rect 699596 114450 699620 114465
rect 699664 114450 699688 114465
rect 699732 114450 699756 114465
rect 699800 114450 699824 114465
rect 699868 114450 699892 114465
rect 699936 114450 699960 114465
rect 700004 114450 700028 114465
rect 700072 114450 700096 114465
rect 700140 114450 700164 114465
rect 700208 114450 700232 114465
rect 700276 114450 700300 114465
rect 700934 114450 700958 114465
rect 701002 114450 701026 114465
rect 701070 114450 701094 114465
rect 701138 114450 701162 114465
rect 701206 114450 701230 114465
rect 701274 114450 701298 114465
rect 701342 114450 701366 114465
rect 701410 114450 701434 114465
rect 701478 114450 701502 114465
rect 701546 114450 701570 114465
rect 701614 114450 701638 114465
rect 701682 114450 701706 114465
rect 701750 114450 701774 114465
rect 701818 114450 701842 114465
rect 692515 114201 693915 114329
rect 694787 114201 696187 114329
rect 699322 114295 700322 114450
rect 699322 114261 700334 114295
rect 700922 114285 701922 114450
rect 707610 114295 708610 114355
rect 709211 114295 710211 114355
rect 700910 114261 701922 114285
rect 699322 114250 700322 114261
rect 700922 114250 701922 114261
rect 699392 114237 699416 114250
rect 699460 114237 699484 114250
rect 699528 114237 699552 114250
rect 699596 114237 699620 114250
rect 699664 114237 699688 114250
rect 699732 114237 699756 114250
rect 699800 114237 699824 114250
rect 699868 114237 699892 114250
rect 699936 114237 699960 114250
rect 700004 114237 700028 114250
rect 700072 114237 700096 114250
rect 700140 114237 700164 114250
rect 700208 114237 700232 114250
rect 700276 114237 700300 114250
rect 700934 114237 700958 114250
rect 701002 114237 701026 114250
rect 701070 114237 701094 114250
rect 701138 114237 701162 114250
rect 701206 114237 701230 114250
rect 701274 114237 701298 114250
rect 701342 114237 701366 114250
rect 701410 114237 701434 114250
rect 701478 114237 701502 114250
rect 701546 114237 701570 114250
rect 701614 114237 701638 114250
rect 701682 114237 701706 114250
rect 701750 114237 701774 114250
rect 701818 114237 701842 114250
rect 692515 114038 693915 114166
rect 694787 114038 696187 114166
rect 692047 113468 696655 114004
rect 699322 113892 700322 113948
rect 700922 113892 701922 113948
rect 707610 113937 708610 113993
rect 709211 113937 710211 113993
rect 699322 113820 700322 113876
rect 700922 113820 701922 113876
rect 707610 113865 708610 113921
rect 709211 113865 710211 113921
rect 697314 113582 697620 113752
rect 699322 113518 700322 113590
rect 700922 113518 701922 113590
rect 707610 113563 708610 113635
rect 709211 113563 710211 113635
rect 704719 113527 705057 113543
rect 699392 113507 699426 113518
rect 699460 113507 699494 113518
rect 699528 113507 699562 113518
rect 699596 113507 699630 113518
rect 699664 113507 699698 113518
rect 699732 113507 699766 113518
rect 699800 113507 699834 113518
rect 699868 113507 699902 113518
rect 699936 113507 699970 113518
rect 700004 113507 700038 113518
rect 700072 113507 700106 113518
rect 700140 113507 700174 113518
rect 700208 113507 700242 113518
rect 700276 113507 700310 113518
rect 700934 113507 700968 113518
rect 701002 113507 701036 113518
rect 701070 113507 701104 113518
rect 701138 113507 701172 113518
rect 701206 113507 701240 113518
rect 701274 113507 701308 113518
rect 701342 113507 701376 113518
rect 701410 113507 701444 113518
rect 701478 113507 701512 113518
rect 701546 113507 701580 113518
rect 701614 113507 701648 113518
rect 701682 113507 701716 113518
rect 701750 113507 701784 113518
rect 701818 113507 701852 113518
rect 699392 113497 699450 113507
rect 699460 113497 699518 113507
rect 699528 113497 699586 113507
rect 699596 113497 699654 113507
rect 699664 113497 699722 113507
rect 699732 113497 699790 113507
rect 699800 113497 699858 113507
rect 699868 113497 699926 113507
rect 699936 113497 699994 113507
rect 700004 113497 700062 113507
rect 700072 113497 700130 113507
rect 700140 113497 700198 113507
rect 700208 113497 700266 113507
rect 700276 113497 700334 113507
rect 700934 113497 700992 113507
rect 701002 113497 701060 113507
rect 701070 113497 701128 113507
rect 701138 113497 701196 113507
rect 701206 113497 701264 113507
rect 701274 113497 701332 113507
rect 701342 113497 701400 113507
rect 701410 113497 701468 113507
rect 701478 113497 701536 113507
rect 701546 113497 701604 113507
rect 701614 113497 701672 113507
rect 701682 113497 701740 113507
rect 701750 113497 701808 113507
rect 701818 113497 701876 113507
rect 699368 113473 700334 113497
rect 700910 113473 701876 113497
rect 699392 113458 699416 113473
rect 699460 113458 699484 113473
rect 699528 113458 699552 113473
rect 699596 113458 699620 113473
rect 699664 113458 699688 113473
rect 699732 113458 699756 113473
rect 699800 113458 699824 113473
rect 699868 113458 699892 113473
rect 699936 113458 699960 113473
rect 700004 113458 700028 113473
rect 700072 113458 700096 113473
rect 700140 113458 700164 113473
rect 700208 113458 700232 113473
rect 700276 113458 700300 113473
rect 700934 113458 700958 113473
rect 701002 113458 701026 113473
rect 701070 113458 701094 113473
rect 701138 113458 701162 113473
rect 701206 113458 701230 113473
rect 701274 113458 701298 113473
rect 701342 113458 701366 113473
rect 701410 113458 701434 113473
rect 701478 113458 701502 113473
rect 701546 113458 701570 113473
rect 701614 113458 701638 113473
rect 701682 113458 701706 113473
rect 701750 113458 701774 113473
rect 701818 113458 701842 113473
rect 699322 113303 700322 113458
rect 692463 113268 692511 113292
rect 696191 113268 696239 113292
rect 692487 113214 692511 113268
rect 696215 113214 696239 113268
rect 699322 113269 700334 113303
rect 700922 113293 701922 113458
rect 704735 113425 705041 113527
rect 707610 113303 708610 113363
rect 709211 113303 710211 113363
rect 700910 113269 701922 113293
rect 699322 113258 700322 113269
rect 700922 113258 701922 113269
rect 699392 113245 699416 113258
rect 699460 113245 699484 113258
rect 699528 113245 699552 113258
rect 699596 113245 699620 113258
rect 699664 113245 699688 113258
rect 699732 113245 699756 113258
rect 699800 113245 699824 113258
rect 699868 113245 699892 113258
rect 699936 113245 699960 113258
rect 700004 113245 700028 113258
rect 700072 113245 700096 113258
rect 700140 113245 700164 113258
rect 700208 113245 700232 113258
rect 700276 113245 700300 113258
rect 700934 113245 700958 113258
rect 701002 113245 701026 113258
rect 701070 113245 701094 113258
rect 701138 113245 701162 113258
rect 701206 113245 701230 113258
rect 701274 113245 701298 113258
rect 701342 113245 701366 113258
rect 701410 113245 701434 113258
rect 701478 113245 701502 113258
rect 701546 113245 701570 113258
rect 701614 113245 701638 113258
rect 701682 113245 701706 113258
rect 701750 113245 701774 113258
rect 701818 113245 701842 113258
rect 692463 113190 692511 113214
rect 696191 113190 696239 113214
rect 687686 113119 687720 113153
rect 687798 113141 687822 113165
rect 687686 113095 687710 113119
rect 687774 113117 687798 113129
rect 687798 113081 687822 113105
rect 692450 113037 692474 113061
rect 692508 113037 692532 113061
rect 696170 113037 696194 113061
rect 696228 113037 696252 113061
rect 692484 113013 692498 113037
rect 696204 113013 696218 113037
rect 692484 112935 692487 112959
rect 696215 112935 696218 112959
rect 692508 112911 692532 112935
rect 696170 112911 696194 112935
rect 699322 112900 700322 112956
rect 700922 112900 701922 112956
rect 707610 112945 708610 113001
rect 709211 112945 710211 113001
rect 692515 112805 693915 112848
rect 694787 112805 696187 112848
rect 699322 112828 700322 112884
rect 700922 112828 701922 112884
rect 707610 112873 708610 112929
rect 709211 112873 710211 112929
rect 692515 112642 693915 112770
rect 694787 112642 696187 112770
rect 688883 112473 688918 112502
rect 692515 112479 693915 112607
rect 694787 112479 696187 112607
rect 699322 112526 700322 112598
rect 700922 112526 701922 112598
rect 707610 112571 708610 112643
rect 709211 112571 710211 112643
rect 699392 112515 699426 112526
rect 699460 112515 699494 112526
rect 699528 112515 699562 112526
rect 699596 112515 699630 112526
rect 699664 112515 699698 112526
rect 699732 112515 699766 112526
rect 699800 112515 699834 112526
rect 699868 112515 699902 112526
rect 699936 112515 699970 112526
rect 700004 112515 700038 112526
rect 700072 112515 700106 112526
rect 700140 112515 700174 112526
rect 700208 112515 700242 112526
rect 700276 112515 700310 112526
rect 700934 112515 700968 112526
rect 701002 112515 701036 112526
rect 701070 112515 701104 112526
rect 701138 112515 701172 112526
rect 701206 112515 701240 112526
rect 701274 112515 701308 112526
rect 701342 112515 701376 112526
rect 701410 112515 701444 112526
rect 701478 112515 701512 112526
rect 701546 112515 701580 112526
rect 701614 112515 701648 112526
rect 701682 112515 701716 112526
rect 701750 112515 701784 112526
rect 701818 112515 701852 112526
rect 699392 112505 699450 112515
rect 699460 112505 699518 112515
rect 699528 112505 699586 112515
rect 699596 112505 699654 112515
rect 699664 112505 699722 112515
rect 699732 112505 699790 112515
rect 699800 112505 699858 112515
rect 699868 112505 699926 112515
rect 699936 112505 699994 112515
rect 700004 112505 700062 112515
rect 700072 112505 700130 112515
rect 700140 112505 700198 112515
rect 700208 112505 700266 112515
rect 700276 112505 700334 112515
rect 700934 112505 700992 112515
rect 701002 112505 701060 112515
rect 701070 112505 701128 112515
rect 701138 112505 701196 112515
rect 701206 112505 701264 112515
rect 701274 112505 701332 112515
rect 701342 112505 701400 112515
rect 701410 112505 701468 112515
rect 701478 112505 701536 112515
rect 701546 112505 701604 112515
rect 701614 112505 701672 112515
rect 701682 112505 701740 112515
rect 701750 112505 701808 112515
rect 701818 112505 701876 112515
rect 699368 112481 700334 112505
rect 700910 112481 701876 112505
rect 688883 112468 688884 112473
rect 688917 112468 688918 112473
rect 688917 112439 688951 112468
rect 699392 112466 699416 112481
rect 699460 112466 699484 112481
rect 699528 112466 699552 112481
rect 699596 112466 699620 112481
rect 699664 112466 699688 112481
rect 699732 112466 699756 112481
rect 699800 112466 699824 112481
rect 699868 112466 699892 112481
rect 699936 112466 699960 112481
rect 700004 112466 700028 112481
rect 700072 112466 700096 112481
rect 700140 112466 700164 112481
rect 700208 112466 700232 112481
rect 700276 112466 700300 112481
rect 700934 112466 700958 112481
rect 701002 112466 701026 112481
rect 701070 112466 701094 112481
rect 701138 112466 701162 112481
rect 701206 112466 701230 112481
rect 701274 112466 701298 112481
rect 701342 112466 701366 112481
rect 701410 112466 701434 112481
rect 701478 112466 701502 112481
rect 701546 112466 701570 112481
rect 701614 112466 701638 112481
rect 701682 112466 701706 112481
rect 701750 112466 701774 112481
rect 701818 112466 701842 112481
rect 688917 112370 688951 112404
rect 688917 112301 688951 112335
rect 692515 112316 693915 112444
rect 694787 112316 696187 112444
rect 699322 112311 700322 112466
rect 688917 112232 688951 112266
rect 688917 112163 688951 112197
rect 692515 112153 693915 112281
rect 694787 112153 696187 112281
rect 699322 112277 700334 112311
rect 700922 112301 701922 112466
rect 707610 112311 708610 112371
rect 709211 112311 710211 112371
rect 700910 112277 701922 112301
rect 699322 112266 700322 112277
rect 700922 112266 701922 112277
rect 699392 112253 699416 112266
rect 699460 112253 699484 112266
rect 699528 112253 699552 112266
rect 699596 112253 699620 112266
rect 699664 112253 699688 112266
rect 699732 112253 699756 112266
rect 699800 112253 699824 112266
rect 699868 112253 699892 112266
rect 699936 112253 699960 112266
rect 700004 112253 700028 112266
rect 700072 112253 700096 112266
rect 700140 112253 700164 112266
rect 700208 112253 700232 112266
rect 700276 112253 700300 112266
rect 700934 112253 700958 112266
rect 701002 112253 701026 112266
rect 701070 112253 701094 112266
rect 701138 112253 701162 112266
rect 701206 112253 701230 112266
rect 701274 112253 701298 112266
rect 701342 112253 701366 112266
rect 701410 112253 701434 112266
rect 701478 112253 701502 112266
rect 701546 112253 701570 112266
rect 701614 112253 701638 112266
rect 701682 112253 701706 112266
rect 701750 112253 701774 112266
rect 701818 112253 701842 112266
rect 688917 112094 688951 112128
rect 688917 112025 688951 112059
rect 692515 111996 693915 112046
rect 694787 111996 696187 112046
rect 688917 111956 688951 111990
rect 698017 111933 698120 111969
rect 688917 111887 688951 111921
rect 692463 111885 692511 111909
rect 696191 111885 696239 111909
rect 688917 111818 688951 111852
rect 692487 111831 692511 111885
rect 696215 111831 696239 111885
rect 698017 111858 698053 111933
rect 692463 111807 692511 111831
rect 696191 111807 696239 111831
rect 698030 111824 698077 111858
rect 698017 111790 698053 111824
rect 688917 111749 688951 111783
rect 698030 111756 698077 111790
rect 698017 111722 698053 111756
rect 688917 111680 688951 111714
rect 698030 111688 698077 111722
rect 698017 111654 698053 111688
rect 688917 111611 688951 111645
rect 692463 111629 692521 111653
rect 696191 111629 696249 111653
rect 692487 111619 692521 111629
rect 696215 111619 696249 111629
rect 698030 111620 698077 111654
rect 698017 111586 698053 111620
rect 686879 111544 687585 111554
rect 686882 111528 687585 111544
rect 688917 111542 688951 111576
rect 692487 111547 692521 111581
rect 696215 111547 696249 111581
rect 678680 111433 678704 111467
rect 681345 111399 682345 111455
rect 678680 111365 678704 111399
rect 684004 111349 685004 111477
rect 688917 111473 688951 111507
rect 692487 111475 692521 111509
rect 696215 111475 696249 111509
rect 688917 111404 688951 111438
rect 692487 111427 692521 111437
rect 696215 111427 696249 111437
rect 692463 111403 692521 111427
rect 696191 111403 696249 111427
rect 688917 111335 688951 111369
rect 2850 111304 3850 111320
rect 2850 111188 3850 111238
rect 2850 110978 3850 111028
rect 3959 111015 3960 111320
rect 5169 111315 5191 111320
rect 6005 111305 6021 111320
rect 1288 109503 1338 110503
rect 1438 109503 1566 110060
rect 1594 109503 1644 110503
rect 5995 109493 6021 111275
rect 7389 110911 8389 110967
rect 8990 110911 9990 110967
rect 15678 110956 16678 111012
rect 17278 110956 18278 111012
rect 7389 110839 8389 110895
rect 8990 110839 9990 110895
rect 15678 110884 16678 110940
rect 17278 110884 18278 110940
rect 27622 110903 27672 111320
rect 27772 110903 27828 111320
rect 27928 110903 27984 111320
rect 28084 110903 28140 111320
rect 28240 110903 28296 111320
rect 28396 110903 28446 111320
rect 31049 111234 32049 111284
rect 36785 111242 37385 111298
rect 678680 111297 678704 111331
rect 678680 111229 678704 111263
rect 679133 111255 679283 111267
rect 679452 111255 679602 111267
rect 681345 111229 682345 111279
rect 678680 111161 678704 111195
rect 684004 111193 685004 111321
rect 688917 111266 688951 111300
rect 679002 111142 679602 111192
rect 36785 111072 37385 111122
rect 678680 111093 678704 111127
rect 681441 111064 681457 111130
rect 682225 111064 682241 111130
rect 678680 111025 678704 111059
rect 684004 111037 685004 111165
rect 685537 111161 686137 111211
rect 688917 111197 688951 111231
rect 692463 111214 692521 111248
rect 696191 111214 696249 111248
rect 688917 111128 688951 111162
rect 678680 110957 678704 110991
rect 679002 110966 679602 111022
rect 678680 110889 678704 110923
rect 681441 110902 681457 110968
rect 683625 110902 683641 110968
rect 684004 110881 685004 111009
rect 685537 111005 686137 111061
rect 688917 111059 688951 111093
rect 692515 111084 693915 111127
rect 694787 111084 696187 111127
rect 688917 110990 688951 111024
rect 688917 110921 688951 110955
rect 692515 110921 693915 111049
rect 694787 110921 696187 111049
rect 685537 110855 686137 110905
rect 678680 110821 678704 110855
rect 679002 110796 679602 110846
rect 678680 110753 678704 110787
rect 680502 110761 680517 110776
rect 21481 110656 22881 110699
rect 23617 110656 25017 110699
rect 678680 110685 678704 110719
rect 31458 110590 32058 110640
rect 678680 110617 678704 110651
rect 15678 110382 16678 110522
rect 17278 110382 18278 110522
rect 21481 110520 22881 110563
rect 23617 110520 25017 110563
rect 678680 110549 678704 110583
rect 680480 110581 680517 110761
rect 680502 110566 680517 110581
rect 680615 110761 680630 110776
rect 680803 110772 680815 110776
rect 680800 110761 680815 110772
rect 680615 110581 680815 110761
rect 681441 110740 681457 110806
rect 683625 110740 683641 110806
rect 684004 110725 685004 110853
rect 688917 110852 688951 110886
rect 688917 110783 688951 110817
rect 692515 110758 693915 110886
rect 694787 110758 696187 110886
rect 688917 110714 688951 110748
rect 686829 110649 687429 110699
rect 688917 110645 688951 110679
rect 680615 110566 680630 110581
rect 680800 110570 680815 110581
rect 681441 110578 681457 110644
rect 682225 110578 682241 110644
rect 684004 110575 685004 110625
rect 688917 110576 688951 110610
rect 692515 110595 693915 110723
rect 694787 110595 696187 110723
rect 680803 110566 680815 110570
rect 680615 110525 680630 110540
rect 680803 110536 680815 110540
rect 680800 110525 680815 110536
rect 678680 110481 678704 110515
rect 31458 110414 32058 110470
rect 678680 110413 678704 110447
rect 678680 110345 678704 110379
rect 679007 110370 679607 110420
rect 680615 110345 680815 110525
rect 681345 110429 682345 110479
rect 686829 110473 687429 110529
rect 688917 110507 688951 110541
rect 688917 110438 688951 110472
rect 692515 110432 693915 110560
rect 694787 110432 696187 110560
rect 684054 110373 685054 110423
rect 688917 110393 688951 110403
rect 688893 110369 688951 110393
rect 680615 110330 680630 110345
rect 680800 110334 680815 110345
rect 680803 110330 680815 110334
rect 25725 110197 26325 110247
rect 31458 110244 32058 110294
rect 678680 110277 678704 110311
rect 681345 110253 682345 110309
rect 678680 110209 678704 110243
rect 7353 110016 8425 110052
rect 7353 109975 7389 110016
rect 8389 109975 8425 110016
rect 7353 109919 8425 109975
rect 7353 109903 7389 109919
rect 8389 109903 8425 109919
rect 7353 109847 8425 109903
rect 7353 109810 7389 109847
rect 8389 109810 8425 109847
rect 7353 109770 8425 109810
rect 8954 110016 10026 110052
rect 8954 109975 8990 110016
rect 9990 109975 10026 110016
rect 8954 109919 10026 109975
rect 21383 110044 21403 110060
rect 21407 110044 21415 110060
rect 21383 110010 21419 110044
rect 21481 110031 22881 110060
rect 23617 110031 25017 110060
rect 25101 110044 25121 110060
rect 25125 110044 25143 110060
rect 25725 110047 26325 110097
rect 25101 110010 25147 110044
rect 21383 109976 21403 110010
rect 21407 109976 21415 110010
rect 21383 109942 21419 109976
rect 8954 109903 8990 109919
rect 9990 109903 10026 109919
rect 15678 109906 16678 109923
rect 17278 109906 18278 109923
rect 21383 109908 21403 109942
rect 21407 109908 21415 109942
rect 8954 109847 10026 109903
rect 20250 109890 20316 109906
rect 8954 109810 8990 109847
rect 9990 109810 10026 109847
rect 8954 109770 10026 109810
rect 21383 109874 21419 109908
rect 21383 109840 21403 109874
rect 21407 109840 21415 109874
rect 21481 109868 22881 109996
rect 23617 109868 25017 109996
rect 25101 109976 25121 110010
rect 25125 109976 25143 110010
rect 25101 109942 25147 109976
rect 25101 109908 25121 109942
rect 25125 109908 25143 109942
rect 25725 109925 26325 109975
rect 25101 109874 25147 109908
rect 25101 109840 25121 109874
rect 25125 109840 25143 109874
rect 21383 109806 21419 109840
rect 21383 109772 21403 109806
rect 21407 109772 21415 109806
rect 21383 109738 21419 109772
rect 15678 109703 16678 109736
rect 17278 109703 18278 109736
rect 21383 109704 21403 109738
rect 21407 109704 21415 109738
rect 21481 109705 22881 109833
rect 23617 109705 25017 109833
rect 25101 109806 25147 109840
rect 25101 109772 25121 109806
rect 25125 109772 25143 109806
rect 25725 109775 26325 109825
rect 25101 109738 25147 109772
rect 25101 109704 25121 109738
rect 25125 109704 25143 109738
rect 21383 109670 21419 109704
rect 25101 109670 25147 109704
rect 21383 109636 21403 109670
rect 21407 109636 21415 109670
rect 7389 109559 8389 109631
rect 8990 109559 9990 109631
rect 21383 109602 21419 109636
rect 15840 109510 15870 109580
rect 15878 109546 15908 109580
rect 21383 109568 21403 109602
rect 21407 109568 21415 109602
rect 15853 109508 15870 109510
rect 21383 109534 21419 109568
rect 21481 109542 22881 109670
rect 23617 109542 25017 109670
rect 25101 109636 25121 109670
rect 25125 109636 25143 109670
rect 25725 109649 26325 109699
rect 25101 109602 25147 109636
rect 25101 109568 25121 109602
rect 25125 109568 25143 109602
rect 25101 109534 25147 109568
rect 5981 109483 6021 109493
rect 5137 109469 6021 109483
rect 21383 109500 21403 109534
rect 21407 109500 21415 109534
rect 21383 109466 21419 109500
rect 7389 109369 8389 109463
rect 7389 109359 8413 109369
rect 8990 109359 9990 109463
rect 21383 109432 21403 109466
rect 21407 109432 21415 109466
rect 21383 109398 21419 109432
rect 21383 109364 21403 109398
rect 21407 109364 21415 109398
rect 21481 109379 22881 109507
rect 23617 109379 25017 109507
rect 25101 109500 25121 109534
rect 25125 109500 25143 109534
rect 25101 109466 25147 109500
rect 25725 109499 26325 109549
rect 25101 109432 25121 109466
rect 25125 109432 25143 109466
rect 25101 109398 25147 109432
rect 25101 109364 25121 109398
rect 25125 109364 25143 109398
rect 25725 109377 26325 109427
rect 21383 109330 21419 109364
rect 25101 109330 25147 109364
rect 21383 109296 21403 109330
rect 21407 109296 21415 109330
rect 25101 109296 25121 109330
rect 25125 109296 25143 109330
rect 21383 109262 21419 109296
rect 21383 109228 21403 109262
rect 21407 109228 21415 109262
rect 21481 109229 22881 109272
rect 23617 109229 25017 109272
rect 25101 109262 25147 109296
rect 25101 109228 25121 109262
rect 25125 109228 25143 109262
rect 21383 109194 21419 109228
rect 25101 109194 25147 109228
rect 25725 109227 26325 109277
rect 21383 109160 21403 109194
rect 21407 109160 21415 109194
rect 25101 109160 25121 109194
rect 25125 109160 25143 109194
rect 27162 109170 27212 110170
rect 27312 109170 27440 110060
rect 27468 109170 27596 110060
rect 27624 109170 27752 110060
rect 27780 109170 27908 110060
rect 27936 109170 28064 110060
rect 28092 109170 28220 110060
rect 28248 109170 28376 110060
rect 28404 109170 28532 110060
rect 28560 109170 28688 110060
rect 28716 109170 28844 110060
rect 28872 109170 29000 110060
rect 29028 109170 29156 110060
rect 29184 109170 29312 110060
rect 29340 109170 29390 110170
rect 30245 110029 30445 110209
rect 30245 110018 30260 110029
rect 30245 110014 30257 110018
rect 30430 110014 30445 110029
rect 30543 110029 30580 110209
rect 679007 110200 679607 110250
rect 684054 110217 685054 110345
rect 686829 110303 687429 110353
rect 692515 110269 693915 110397
rect 694787 110269 696187 110397
rect 678680 110141 678704 110175
rect 678680 110073 678704 110107
rect 681345 110077 682345 110205
rect 30543 110014 30558 110029
rect 678680 110005 678704 110039
rect 680215 110024 680815 110074
rect 684054 110061 685054 110189
rect 685793 110182 685805 110186
rect 685793 110171 685808 110182
rect 685978 110171 685993 110186
rect 30245 109984 30257 109988
rect 30245 109973 30260 109984
rect 30430 109973 30445 109988
rect 30245 109793 30445 109973
rect 678680 109937 678704 109971
rect 678680 109869 678704 109903
rect 31453 109818 32053 109868
rect 680215 109848 680815 109904
rect 681345 109901 682345 110029
rect 684054 109905 685054 110033
rect 685793 109991 685993 110171
rect 685793 109980 685808 109991
rect 685793 109976 685805 109980
rect 685978 109976 685993 109991
rect 686053 110182 686065 110186
rect 686053 110171 686068 110182
rect 686238 110171 686253 110186
rect 686053 109991 686253 110171
rect 686607 110164 687607 110214
rect 697088 110171 697138 111571
rect 697238 110171 697366 111571
rect 697394 110171 697522 111571
rect 697550 110171 697678 111571
rect 697706 110171 697756 111571
rect 698030 111552 698077 111586
rect 698017 111518 698053 111552
rect 698030 111484 698077 111518
rect 698017 111450 698053 111484
rect 698030 111416 698077 111450
rect 698017 111382 698053 111416
rect 698030 111348 698077 111382
rect 698017 111314 698053 111348
rect 698030 111280 698077 111314
rect 698017 111246 698053 111280
rect 698030 111212 698077 111246
rect 698017 111178 698053 111212
rect 698030 111144 698077 111178
rect 698017 111110 698053 111144
rect 698030 111076 698077 111110
rect 698017 111042 698053 111076
rect 698030 111008 698077 111042
rect 698017 110974 698053 111008
rect 698030 110940 698077 110974
rect 698017 110906 698053 110940
rect 698030 110872 698077 110906
rect 698017 110838 698053 110872
rect 698030 110804 698077 110838
rect 698017 110770 698053 110804
rect 698030 110736 698077 110770
rect 698017 110702 698053 110736
rect 698030 110668 698077 110702
rect 698017 110634 698053 110668
rect 698030 110600 698077 110634
rect 698017 110566 698053 110600
rect 698030 110532 698077 110566
rect 698017 110498 698053 110532
rect 698030 110464 698077 110498
rect 698017 110430 698053 110464
rect 698030 110396 698077 110430
rect 698017 110362 698053 110396
rect 698030 110328 698077 110362
rect 698017 110294 698053 110328
rect 698030 110260 698077 110294
rect 698017 110226 698053 110260
rect 698030 110192 698077 110226
rect 692515 110119 693915 110162
rect 694787 110119 696187 110162
rect 698017 110158 698053 110192
rect 698030 110124 698077 110158
rect 698017 110090 698053 110124
rect 686607 110014 687607 110064
rect 698030 110056 698077 110090
rect 686053 109980 686068 109991
rect 686053 109976 686065 109980
rect 686238 109976 686253 109991
rect 685793 109946 685805 109950
rect 685793 109935 685808 109946
rect 685978 109935 685993 109950
rect 678680 109801 678704 109835
rect 30245 109782 30260 109793
rect 30245 109778 30257 109782
rect 30430 109778 30445 109793
rect 678680 109733 678704 109767
rect 681345 109731 682345 109781
rect 684054 109749 685054 109877
rect 685793 109755 685993 109935
rect 685793 109744 685808 109755
rect 685793 109740 685805 109744
rect 685978 109740 685993 109755
rect 686053 109946 686065 109950
rect 686053 109935 686068 109946
rect 686238 109935 686253 109950
rect 686053 109755 686253 109935
rect 686607 109855 687607 109905
rect 692463 109809 692511 109833
rect 696191 109809 696239 109833
rect 686053 109744 686068 109755
rect 686053 109740 686065 109744
rect 686238 109740 686253 109755
rect 31453 109648 32053 109698
rect 678680 109665 678704 109699
rect 680215 109672 680815 109728
rect 681345 109662 682345 109674
rect 678680 109597 678704 109631
rect 684054 109593 685054 109721
rect 686607 109705 687607 109755
rect 692487 109731 692511 109809
rect 696215 109755 696239 109809
rect 696191 109731 696239 109755
rect 696617 109772 696651 109773
rect 696617 109749 696626 109772
rect 696617 109731 696675 109749
rect 696651 109715 696675 109731
rect 696651 109647 696675 109681
rect 685533 109586 685545 109590
rect 685533 109575 685548 109586
rect 685718 109575 685733 109590
rect 678680 109529 678704 109563
rect 30245 109472 30845 109522
rect 680215 109502 680815 109552
rect 678680 109461 678704 109495
rect 678680 109393 678704 109427
rect 680215 109370 680815 109420
rect 681466 109411 682466 109461
rect 684054 109437 685054 109565
rect 30245 109296 30845 109352
rect 678680 109325 678704 109359
rect 678680 109257 678704 109291
rect 681466 109255 682466 109383
rect 682890 109339 683490 109389
rect 678680 109189 678704 109223
rect 680215 109194 680815 109250
rect 682890 109183 683490 109311
rect 684054 109281 685054 109409
rect 685533 109395 685733 109575
rect 685533 109384 685548 109395
rect 685533 109380 685545 109384
rect 685718 109380 685733 109395
rect 685793 109586 685805 109590
rect 685793 109575 685808 109586
rect 685978 109575 685993 109590
rect 685793 109395 685993 109575
rect 685793 109384 685808 109395
rect 685793 109380 685805 109384
rect 685978 109380 685993 109395
rect 686053 109586 686065 109590
rect 686053 109575 686068 109586
rect 686238 109575 686253 109590
rect 686053 109395 686253 109575
rect 686053 109384 686068 109395
rect 686053 109380 686065 109384
rect 686238 109380 686253 109395
rect 686313 109586 686325 109590
rect 686313 109575 686328 109586
rect 686498 109575 686513 109590
rect 686313 109395 686513 109575
rect 686313 109384 686328 109395
rect 686313 109380 686325 109384
rect 686498 109380 686513 109395
rect 686627 109586 686639 109590
rect 686627 109575 686642 109586
rect 686812 109575 686827 109590
rect 686627 109395 686827 109575
rect 686627 109384 686642 109395
rect 686627 109380 686639 109384
rect 686812 109380 686827 109395
rect 686887 109586 686899 109590
rect 686887 109575 686902 109586
rect 687072 109575 687087 109590
rect 686887 109395 687087 109575
rect 686887 109384 686902 109395
rect 686887 109380 686899 109384
rect 687072 109380 687087 109395
rect 687147 109586 687159 109590
rect 687147 109575 687162 109586
rect 687332 109575 687347 109590
rect 696651 109579 696675 109613
rect 687147 109395 687347 109575
rect 696651 109511 696675 109545
rect 696651 109443 696675 109477
rect 687147 109384 687162 109395
rect 687147 109380 687159 109384
rect 687332 109380 687347 109395
rect 696651 109375 696675 109409
rect 696651 109307 696675 109341
rect 685718 109215 685733 109230
rect 685679 109185 685733 109215
rect 21383 109126 21419 109160
rect 25101 109126 25147 109160
rect 21383 109102 21403 109126
rect 21385 109048 21403 109102
rect 21407 109082 21415 109126
rect 25101 109102 25121 109126
rect 25113 109082 25121 109102
rect 25125 109048 25143 109126
rect 30245 109120 30845 109176
rect 678680 109121 678704 109155
rect 681466 109105 682466 109155
rect 684054 109131 685054 109181
rect 685718 109170 685733 109185
rect 685793 109226 685805 109230
rect 685793 109215 685808 109226
rect 685978 109215 685993 109230
rect 685793 109185 685993 109215
rect 685793 109174 685808 109185
rect 685793 109170 685805 109174
rect 685978 109170 685993 109185
rect 686053 109226 686065 109230
rect 686053 109215 686068 109226
rect 686238 109215 686253 109230
rect 686812 109215 686827 109230
rect 686053 109185 686253 109215
rect 686807 109185 686827 109215
rect 686053 109174 686068 109185
rect 686053 109170 686065 109174
rect 686238 109170 686253 109185
rect 686812 109170 686827 109185
rect 686887 109226 686899 109230
rect 686887 109215 686902 109226
rect 687072 109215 687087 109230
rect 686887 109185 687087 109215
rect 686887 109174 686902 109185
rect 686887 109170 686899 109174
rect 687072 109170 687087 109185
rect 687147 109226 687159 109230
rect 687147 109215 687162 109226
rect 687332 109215 687347 109230
rect 687147 109185 687347 109215
rect 687147 109174 687162 109185
rect 687147 109170 687159 109174
rect 687332 109170 687347 109185
rect 685718 109129 685733 109144
rect 681794 109102 682466 109105
rect 685679 109099 685733 109129
rect 678680 109053 678704 109087
rect 685718 109084 685733 109099
rect 685793 109140 685805 109144
rect 685793 109129 685808 109140
rect 685978 109129 685993 109144
rect 685793 109099 685993 109129
rect 685793 109088 685808 109099
rect 685793 109084 685805 109088
rect 685978 109084 685993 109099
rect 686053 109140 686065 109144
rect 686053 109129 686068 109140
rect 686238 109129 686253 109144
rect 686812 109129 686827 109144
rect 686053 109099 686253 109129
rect 686807 109099 686827 109129
rect 686053 109088 686068 109099
rect 686053 109084 686065 109088
rect 686238 109084 686253 109099
rect 686812 109084 686827 109099
rect 686887 109140 686899 109144
rect 686887 109129 686902 109140
rect 687072 109129 687087 109144
rect 686887 109099 687087 109129
rect 686887 109088 686902 109099
rect 686887 109084 686899 109088
rect 687072 109084 687087 109099
rect 687147 109140 687159 109144
rect 687147 109129 687162 109140
rect 687332 109129 687347 109144
rect 687147 109099 687347 109129
rect 687147 109088 687162 109099
rect 687147 109084 687159 109088
rect 687332 109084 687347 109099
rect 30245 108950 30845 109000
rect 678680 108985 678704 109019
rect 680215 109018 680815 109074
rect 682890 109027 683490 109083
rect 21000 108800 21003 108920
rect 678680 108917 678704 108951
rect 21352 108885 21376 108909
rect 25122 108885 25146 108909
rect 21385 108861 21400 108885
rect 25098 108861 25113 108885
rect 21274 108783 21294 108851
rect 21410 108817 21430 108851
rect 25068 108817 25088 108851
rect 25204 108817 25224 108851
rect 678680 108849 678704 108883
rect 680215 108848 680815 108898
rect 21385 108807 21430 108817
rect 25102 108807 25137 108817
rect 21361 108783 21430 108807
rect 25089 108783 25137 108807
rect 25238 108783 25258 108817
rect 678680 108781 678704 108815
rect 678680 108713 678704 108747
rect 678680 108645 678704 108679
rect 679007 108672 679607 108722
rect 678680 108577 678704 108611
rect 680615 108577 680630 108592
rect 680803 108588 680815 108592
rect 680800 108577 680815 108588
rect 678680 108509 678704 108543
rect 679007 108502 679607 108552
rect 678680 108441 678704 108475
rect 678680 108373 678704 108407
rect 680615 108397 680815 108577
rect 681502 108505 681529 108995
rect 681866 108896 682466 109024
rect 682890 108871 683490 108999
rect 684004 108929 685004 108979
rect 685539 108940 685777 108972
rect 685803 108920 686119 108938
rect 681866 108740 682466 108868
rect 684004 108773 685004 108901
rect 682890 108721 683490 108771
rect 681866 108584 682466 108712
rect 682890 108605 683490 108655
rect 684004 108617 685004 108745
rect 681866 108434 682466 108484
rect 682890 108449 683490 108505
rect 684004 108461 685004 108589
rect 692427 108522 693027 108572
rect 680615 108382 680630 108397
rect 680800 108386 680815 108397
rect 680803 108382 680815 108386
rect 680502 108341 680517 108356
rect 678680 108305 678704 108339
rect 678680 108237 678704 108271
rect 678680 108169 678704 108203
rect 680480 108161 680517 108341
rect 680502 108146 680517 108161
rect 680615 108341 680630 108356
rect 680803 108352 680815 108356
rect 680800 108341 680815 108352
rect 680615 108161 680815 108341
rect 681866 108318 682466 108368
rect 682890 108293 683490 108349
rect 684004 108305 685004 108433
rect 692427 108366 693027 108494
rect 693888 108375 694194 108545
rect 694388 108375 694694 108545
rect 689309 108278 689909 108328
rect 681866 108168 682466 108218
rect 682041 108165 682385 108168
rect 680615 108146 680630 108161
rect 680800 108150 680815 108161
rect 680803 108146 680815 108150
rect 682890 108137 683490 108193
rect 684004 108149 685004 108277
rect 678680 108101 678704 108135
rect 679002 108076 679602 108126
rect 689309 108122 689909 108250
rect 692427 108210 693027 108338
rect 678680 108033 678704 108067
rect 678680 107965 678704 107999
rect 682890 107981 683490 108109
rect 684004 107993 685004 108121
rect 689309 107966 689909 108094
rect 692427 108054 693027 108110
rect 678680 107897 678704 107931
rect 679002 107900 679602 107956
rect 678680 107829 678704 107863
rect 682890 107825 683490 107953
rect 684004 107837 685004 107965
rect 692427 107898 693027 108026
rect 689309 107810 689909 107866
rect 678680 107761 678704 107795
rect 679002 107730 679602 107780
rect 679061 107727 679355 107730
rect 679380 107727 679602 107730
rect 678680 107693 678704 107727
rect 682890 107669 683490 107797
rect 684004 107687 685004 107737
rect 685803 107720 686119 107732
rect 685539 107716 686119 107720
rect 685513 107682 685537 107716
rect 685539 107682 685777 107716
rect 678680 107625 678704 107659
rect 689309 107654 689909 107782
rect 690910 107754 691110 107765
rect 692427 107742 693027 107870
rect 690910 107640 691110 107690
rect 678680 107557 678704 107591
rect 678680 107489 678704 107523
rect 682890 107513 683490 107569
rect 685718 107555 685733 107570
rect 684004 107485 685004 107535
rect 685679 107525 685733 107555
rect 685718 107510 685733 107525
rect 685793 107566 685805 107570
rect 685793 107555 685808 107566
rect 685978 107555 685993 107570
rect 685793 107525 685993 107555
rect 685793 107514 685808 107525
rect 685793 107510 685805 107514
rect 685978 107510 685993 107525
rect 686053 107566 686065 107570
rect 686053 107555 686068 107566
rect 686238 107555 686253 107570
rect 686812 107555 686827 107570
rect 686053 107525 686253 107555
rect 686807 107525 686827 107555
rect 686053 107514 686068 107525
rect 686053 107510 686065 107514
rect 686238 107510 686253 107525
rect 686812 107510 686827 107525
rect 686887 107566 686899 107570
rect 686887 107555 686902 107566
rect 687072 107555 687087 107570
rect 686887 107525 687087 107555
rect 686887 107514 686902 107525
rect 686887 107510 686899 107514
rect 687072 107510 687087 107525
rect 687147 107566 687159 107570
rect 687147 107555 687162 107566
rect 687332 107555 687347 107570
rect 687147 107525 687347 107555
rect 687147 107514 687162 107525
rect 687147 107510 687159 107514
rect 687332 107510 687347 107525
rect 689309 107498 689909 107626
rect 692427 107592 693027 107642
rect 693888 107575 694194 107745
rect 694388 107575 694694 107745
rect 678680 107421 678704 107455
rect 678680 107353 678704 107387
rect 682890 107357 683490 107485
rect 690910 107484 691110 107540
rect 685718 107469 685733 107484
rect 684004 107329 685004 107457
rect 685679 107439 685733 107469
rect 685718 107424 685733 107439
rect 685793 107480 685805 107484
rect 685793 107469 685808 107480
rect 685978 107469 685993 107484
rect 685793 107439 685993 107469
rect 685793 107428 685808 107439
rect 685793 107424 685805 107428
rect 685978 107424 685993 107439
rect 686053 107480 686065 107484
rect 686053 107469 686068 107480
rect 686238 107469 686253 107484
rect 686812 107469 686827 107484
rect 686053 107439 686253 107469
rect 686807 107439 686827 107469
rect 686053 107428 686068 107439
rect 686053 107424 686065 107428
rect 686238 107424 686253 107439
rect 686812 107424 686827 107439
rect 686887 107480 686899 107484
rect 686887 107469 686902 107480
rect 687072 107469 687087 107484
rect 686887 107439 687087 107469
rect 686887 107428 686902 107439
rect 686887 107424 686899 107428
rect 687072 107424 687087 107439
rect 687147 107480 687159 107484
rect 687147 107469 687162 107480
rect 687332 107469 687347 107484
rect 687147 107439 687347 107469
rect 692427 107462 693027 107512
rect 687147 107428 687162 107439
rect 687147 107424 687159 107428
rect 687332 107424 687347 107439
rect 689309 107348 689909 107398
rect 690910 107334 691110 107384
rect 678680 107285 678704 107319
rect 678680 107217 678704 107251
rect 682890 107201 683490 107329
rect 692427 107312 693027 107362
rect 678680 107149 678704 107183
rect 684004 107173 685004 107301
rect 685533 107270 685545 107274
rect 685533 107259 685548 107270
rect 685718 107259 685733 107274
rect 678680 107081 678704 107115
rect 679133 107101 679283 107113
rect 679452 107101 679602 107113
rect 678680 107013 678704 107047
rect 682890 107045 683490 107173
rect 679002 106988 679602 107038
rect 684004 107017 685004 107145
rect 685533 107079 685733 107259
rect 685533 107068 685548 107079
rect 685533 107064 685545 107068
rect 685718 107064 685733 107079
rect 685793 107270 685805 107274
rect 685793 107259 685808 107270
rect 685978 107259 685993 107274
rect 685793 107079 685993 107259
rect 685793 107068 685808 107079
rect 685793 107064 685805 107068
rect 685978 107064 685993 107079
rect 686053 107270 686065 107274
rect 686053 107259 686068 107270
rect 686238 107259 686253 107274
rect 686053 107079 686253 107259
rect 686053 107068 686068 107079
rect 686053 107064 686065 107068
rect 686238 107064 686253 107079
rect 686313 107270 686325 107274
rect 686313 107259 686328 107270
rect 686498 107259 686513 107274
rect 686313 107079 686513 107259
rect 686313 107068 686328 107079
rect 686313 107064 686325 107068
rect 686498 107064 686513 107079
rect 686627 107270 686639 107274
rect 686627 107259 686642 107270
rect 686812 107259 686827 107274
rect 686627 107079 686827 107259
rect 686627 107068 686642 107079
rect 686627 107064 686639 107068
rect 686812 107064 686827 107079
rect 686887 107270 686899 107274
rect 686887 107259 686902 107270
rect 687072 107259 687087 107274
rect 686887 107079 687087 107259
rect 686887 107068 686902 107079
rect 686887 107064 686899 107068
rect 687072 107064 687087 107079
rect 687147 107270 687159 107274
rect 687147 107259 687162 107270
rect 687332 107259 687347 107274
rect 687147 107079 687347 107259
rect 689309 107218 689909 107268
rect 692427 107140 693027 107190
rect 687147 107068 687162 107079
rect 687147 107064 687159 107068
rect 687332 107064 687347 107079
rect 689309 107068 689909 107118
rect 692427 106990 693027 107040
rect 678680 106945 678704 106979
rect 678680 106877 678704 106911
rect 682890 106895 683490 106945
rect 678680 106809 678704 106843
rect 679002 106812 679602 106868
rect 684004 106861 685004 106917
rect 685793 106910 685805 106914
rect 685793 106899 685808 106910
rect 685978 106899 685993 106914
rect 682890 106779 683490 106829
rect 678680 106741 678704 106775
rect 678680 106673 678704 106707
rect 679002 106642 679602 106692
rect 678680 106605 678704 106639
rect 682890 106623 683490 106751
rect 684004 106705 685004 106833
rect 685793 106719 685993 106899
rect 685793 106708 685808 106719
rect 685793 106704 685805 106708
rect 685978 106704 685993 106719
rect 686053 106910 686065 106914
rect 686053 106899 686068 106910
rect 686238 106899 686253 106914
rect 686607 106899 687607 106949
rect 690910 106934 691110 106984
rect 686053 106719 686253 106899
rect 692427 106860 693027 106910
rect 686607 106749 687607 106799
rect 690910 106778 691110 106834
rect 686053 106708 686068 106719
rect 686053 106704 686065 106708
rect 686238 106704 686253 106719
rect 692427 106704 693027 106832
rect 693888 106775 694194 106945
rect 694388 106775 694694 106945
rect 680502 106607 680517 106622
rect 678680 106537 678704 106571
rect 678680 106469 678704 106503
rect 678680 106401 678704 106435
rect 680480 106427 680517 106607
rect 680502 106412 680517 106427
rect 680615 106607 680630 106622
rect 680803 106618 680815 106622
rect 680800 106607 680815 106618
rect 680615 106427 680815 106607
rect 682890 106467 683490 106595
rect 684004 106549 685004 106677
rect 685793 106674 685805 106678
rect 685793 106663 685808 106674
rect 685978 106663 685993 106678
rect 680615 106412 680630 106427
rect 680800 106416 680815 106427
rect 680803 106412 680815 106416
rect 680615 106371 680630 106386
rect 680803 106382 680815 106386
rect 680800 106371 680815 106382
rect 678680 106333 678704 106367
rect 678680 106265 678704 106299
rect 678680 106197 678704 106231
rect 679007 106216 679607 106266
rect 680615 106191 680815 106371
rect 682890 106311 683490 106439
rect 684004 106393 685004 106521
rect 685793 106483 685993 106663
rect 685793 106472 685808 106483
rect 685793 106468 685805 106472
rect 685978 106468 685993 106483
rect 686053 106674 686065 106678
rect 686053 106663 686068 106674
rect 686238 106663 686253 106678
rect 686053 106483 686253 106663
rect 686607 106590 687607 106640
rect 690910 106628 691110 106678
rect 692427 106548 693027 106676
rect 686053 106472 686068 106483
rect 686053 106468 686065 106472
rect 686238 106468 686253 106483
rect 686607 106440 687607 106490
rect 692427 106392 693027 106448
rect 686829 106301 687429 106351
rect 684004 106243 685004 106293
rect 692427 106236 693027 106364
rect 695201 106282 695251 109282
rect 695351 106282 695479 109282
rect 695507 106282 695635 109282
rect 695663 106282 695791 109282
rect 695819 106282 695947 109282
rect 695975 106282 696103 109282
rect 696131 106282 696259 109282
rect 696287 106282 696337 109282
rect 696651 109239 696675 109273
rect 696651 109171 696675 109205
rect 696651 109103 696675 109137
rect 696651 109035 696675 109069
rect 696651 108967 696675 109001
rect 696651 108899 696675 108933
rect 696651 108831 696675 108865
rect 696651 108763 696675 108797
rect 696651 108695 696675 108729
rect 696651 108627 696675 108661
rect 697088 108641 697138 110041
rect 697238 108641 697366 110041
rect 697394 108641 697522 110041
rect 697550 108641 697678 110041
rect 697706 108641 697756 110041
rect 698017 110022 698053 110056
rect 698030 109988 698077 110022
rect 698017 109954 698053 109988
rect 698030 109920 698077 109954
rect 698017 109886 698053 109920
rect 698030 109852 698077 109886
rect 698017 109818 698053 109852
rect 698030 109784 698077 109818
rect 698017 109750 698053 109784
rect 698030 109716 698077 109750
rect 698017 109682 698053 109716
rect 698030 109648 698077 109682
rect 698017 109614 698053 109648
rect 698030 109580 698077 109614
rect 698017 109546 698053 109580
rect 698030 109512 698077 109546
rect 698017 109478 698053 109512
rect 698030 109444 698077 109478
rect 698017 109410 698053 109444
rect 698030 109376 698077 109410
rect 698017 109342 698053 109376
rect 698030 109308 698077 109342
rect 698017 109274 698053 109308
rect 698030 109240 698077 109274
rect 698017 109206 698053 109240
rect 698030 109172 698077 109206
rect 698017 109138 698053 109172
rect 698030 109104 698077 109138
rect 698017 109070 698053 109104
rect 698030 109036 698077 109070
rect 698017 109002 698053 109036
rect 698030 108968 698077 109002
rect 698017 108934 698053 108968
rect 698030 108900 698077 108934
rect 698017 108866 698053 108900
rect 698030 108832 698077 108866
rect 698017 108798 698053 108832
rect 698030 108764 698077 108798
rect 698017 108730 698053 108764
rect 698030 108696 698077 108730
rect 698017 108662 698053 108696
rect 698030 108628 698077 108662
rect 698017 108594 698053 108628
rect 696651 108559 696675 108593
rect 698030 108560 698077 108594
rect 698017 108526 698053 108560
rect 696651 108491 696675 108525
rect 698030 108492 698077 108526
rect 696651 108423 696675 108457
rect 698017 108428 698053 108492
rect 698030 108394 698077 108428
rect 696651 108355 696675 108389
rect 698017 108360 698053 108394
rect 698030 108326 698077 108360
rect 696651 108287 696675 108321
rect 698017 108292 698053 108326
rect 696651 108219 696675 108253
rect 696651 108151 696675 108185
rect 696651 108083 696675 108117
rect 696651 108015 696675 108049
rect 696651 107947 696675 107981
rect 696651 107879 696675 107913
rect 696651 107811 696675 107845
rect 696651 107743 696675 107777
rect 696651 107675 696675 107709
rect 696651 107607 696675 107641
rect 696651 107539 696675 107573
rect 696651 107471 696675 107505
rect 696651 107403 696675 107437
rect 696651 107335 696675 107369
rect 696651 107267 696675 107301
rect 696651 107199 696675 107233
rect 696651 107131 696675 107165
rect 696651 107063 696675 107097
rect 696651 106995 696675 107029
rect 696651 106927 696675 106961
rect 696651 106859 696675 106893
rect 697088 106879 697138 108279
rect 697238 106879 697366 108279
rect 697394 106879 697522 108279
rect 697550 106879 697678 108279
rect 697706 106879 697756 108279
rect 698030 108258 698077 108292
rect 698017 108224 698053 108258
rect 698030 108190 698077 108224
rect 698017 108156 698053 108190
rect 698030 108122 698077 108156
rect 698017 108088 698053 108122
rect 698030 108054 698077 108088
rect 698017 108020 698053 108054
rect 698030 107986 698077 108020
rect 698017 107952 698053 107986
rect 698030 107918 698077 107952
rect 698017 107884 698053 107918
rect 698030 107850 698077 107884
rect 698017 107816 698053 107850
rect 698030 107782 698077 107816
rect 698017 107748 698053 107782
rect 698030 107714 698077 107748
rect 698017 107680 698053 107714
rect 698030 107646 698077 107680
rect 698017 107612 698053 107646
rect 698030 107578 698077 107612
rect 698017 107544 698053 107578
rect 698030 107510 698077 107544
rect 698017 107476 698053 107510
rect 698030 107442 698077 107476
rect 698017 107408 698053 107442
rect 698030 107374 698077 107408
rect 698017 107340 698053 107374
rect 698030 107306 698077 107340
rect 698017 107272 698053 107306
rect 698030 107238 698077 107272
rect 698017 107204 698053 107238
rect 698030 107170 698077 107204
rect 698017 107136 698053 107170
rect 698030 107102 698077 107136
rect 698017 107068 698053 107102
rect 698030 107034 698077 107068
rect 698017 107000 698053 107034
rect 698030 106966 698077 107000
rect 698017 106932 698053 106966
rect 698030 106898 698077 106932
rect 698017 106864 698053 106898
rect 698030 106830 698077 106864
rect 696651 106791 696675 106825
rect 698017 106796 698053 106830
rect 698030 106762 698077 106796
rect 696651 106723 696675 106757
rect 696651 106655 696675 106689
rect 696651 106587 696675 106621
rect 696651 106519 696675 106553
rect 696651 106451 696675 106485
rect 696651 106383 696675 106417
rect 696651 106315 696675 106349
rect 696651 106247 696675 106281
rect 680615 106176 680630 106191
rect 680800 106180 680815 106191
rect 680803 106176 680815 106180
rect 678680 106129 678704 106163
rect 682890 106161 683490 106211
rect 684004 106127 685004 106177
rect 686829 106125 687429 106181
rect 678680 106061 678704 106095
rect 679007 106046 679607 106096
rect 692427 106080 693027 106208
rect 696651 106179 696675 106213
rect 696651 106111 696675 106145
rect 696651 106043 696675 106077
rect 678680 105993 678704 106027
rect 681664 106002 681812 106006
rect 681641 105994 681812 106002
rect 682113 105994 682313 106006
rect 684004 105971 685004 106027
rect 678680 105925 678704 105959
rect 686829 105955 687429 106005
rect 678680 105857 678704 105891
rect 680215 105870 680815 105920
rect 681713 105881 682313 105931
rect 682921 105899 683521 105949
rect 692427 105930 693027 105980
rect 696651 105975 696675 106009
rect 696651 105907 696675 105941
rect 678680 105789 678704 105823
rect 684004 105821 685004 105871
rect 678680 105721 678704 105755
rect 680215 105694 680815 105750
rect 681713 105705 682313 105761
rect 682921 105743 683521 105799
rect 685537 105749 686137 105799
rect 697088 105749 697138 106749
rect 697238 105749 697366 106749
rect 697394 105749 697522 106749
rect 697550 105749 697678 106749
rect 697706 105749 697756 106749
rect 698017 106728 698053 106762
rect 698030 106694 698077 106728
rect 698017 106660 698053 106694
rect 698030 106626 698077 106660
rect 698017 106592 698053 106626
rect 698030 106558 698077 106592
rect 698017 106524 698053 106558
rect 698030 106490 698077 106524
rect 698017 106456 698053 106490
rect 698030 106422 698077 106456
rect 698017 106388 698053 106422
rect 698030 106354 698077 106388
rect 698017 106320 698053 106354
rect 698030 106286 698077 106320
rect 698017 106252 698053 106286
rect 698030 106218 698077 106252
rect 698017 106184 698053 106218
rect 698030 106150 698077 106184
rect 698017 106116 698053 106150
rect 698030 106082 698077 106116
rect 698017 106048 698053 106082
rect 698030 106014 698077 106048
rect 698017 105980 698053 106014
rect 698030 105946 698077 105980
rect 698017 105912 698053 105946
rect 698030 105878 698077 105912
rect 698017 105844 698053 105878
rect 698030 105810 698077 105844
rect 698017 105776 698053 105810
rect 698030 105742 698077 105776
rect 698017 105708 698053 105742
rect 678680 105653 678704 105687
rect 698030 105674 698077 105708
rect 678680 105585 678704 105619
rect 680215 105518 680815 105574
rect 681713 105529 682313 105657
rect 682921 105593 683521 105643
rect 684070 105599 684670 105649
rect 685537 105593 686137 105649
rect 698017 105640 698053 105674
rect 698030 105606 698077 105640
rect 698017 105572 698053 105606
rect 698030 105538 698077 105572
rect 698017 105504 698053 105538
rect 684070 105443 684670 105499
rect 685537 105443 686137 105493
rect 692428 105442 693028 105492
rect 698030 105470 698077 105504
rect 698017 105436 698053 105470
rect 680215 105348 680815 105398
rect 681713 105359 682313 105409
rect 698030 105402 698077 105436
rect 698017 105368 698053 105402
rect 684070 105293 684670 105343
rect 692428 105292 693028 105342
rect 698030 105334 698077 105368
rect 698017 105300 698053 105334
rect 680215 105232 680815 105282
rect 698030 105266 698077 105300
rect 698017 105232 698053 105266
rect 692428 105162 693028 105212
rect 698030 105198 698077 105232
rect 698017 105164 698053 105198
rect 680215 105056 680815 105112
rect 692428 105006 693028 105134
rect 698030 105130 698077 105164
rect 698017 105096 698053 105130
rect 698030 105062 698077 105096
rect 698017 104983 698053 105062
rect 698084 104983 698120 111933
rect 699322 111908 700322 111964
rect 700922 111908 701922 111964
rect 707610 111953 708610 112009
rect 709211 111953 710211 112009
rect 699322 111836 700322 111892
rect 700922 111836 701922 111892
rect 707610 111881 708610 111937
rect 709211 111881 710211 111937
rect 699322 111534 700322 111606
rect 700922 111534 701922 111606
rect 707610 111579 708610 111651
rect 709211 111579 710211 111651
rect 699392 111523 699426 111534
rect 699460 111523 699494 111534
rect 699528 111523 699562 111534
rect 699596 111523 699630 111534
rect 699664 111523 699698 111534
rect 699732 111523 699766 111534
rect 699800 111523 699834 111534
rect 699868 111523 699902 111534
rect 699936 111523 699970 111534
rect 700004 111523 700038 111534
rect 700072 111523 700106 111534
rect 700140 111523 700174 111534
rect 700208 111523 700242 111534
rect 700276 111523 700310 111534
rect 700934 111523 700968 111534
rect 701002 111523 701036 111534
rect 701070 111523 701104 111534
rect 701138 111523 701172 111534
rect 701206 111523 701240 111534
rect 701274 111523 701308 111534
rect 701342 111523 701376 111534
rect 701410 111523 701444 111534
rect 701478 111523 701512 111534
rect 701546 111523 701580 111534
rect 701614 111523 701648 111534
rect 701682 111523 701716 111534
rect 701750 111523 701784 111534
rect 701818 111523 701852 111534
rect 699392 111513 699450 111523
rect 699460 111513 699518 111523
rect 699528 111513 699586 111523
rect 699596 111513 699654 111523
rect 699664 111513 699722 111523
rect 699732 111513 699790 111523
rect 699800 111513 699858 111523
rect 699868 111513 699926 111523
rect 699936 111513 699994 111523
rect 700004 111513 700062 111523
rect 700072 111513 700130 111523
rect 700140 111513 700198 111523
rect 700208 111513 700266 111523
rect 700276 111513 700334 111523
rect 700934 111513 700992 111523
rect 701002 111513 701060 111523
rect 701070 111513 701128 111523
rect 701138 111513 701196 111523
rect 701206 111513 701264 111523
rect 701274 111513 701332 111523
rect 701342 111513 701400 111523
rect 701410 111513 701468 111523
rect 701478 111513 701536 111523
rect 701546 111513 701604 111523
rect 701614 111513 701672 111523
rect 701682 111513 701740 111523
rect 701750 111513 701808 111523
rect 701818 111513 701876 111523
rect 699368 111489 700334 111513
rect 700910 111489 701876 111513
rect 699392 111474 699416 111489
rect 699460 111474 699484 111489
rect 699528 111474 699552 111489
rect 699596 111474 699620 111489
rect 699664 111474 699688 111489
rect 699732 111474 699756 111489
rect 699800 111474 699824 111489
rect 699868 111474 699892 111489
rect 699936 111474 699960 111489
rect 700004 111474 700028 111489
rect 700072 111474 700096 111489
rect 700140 111474 700164 111489
rect 700208 111474 700232 111489
rect 700276 111474 700300 111489
rect 700934 111474 700958 111489
rect 701002 111474 701026 111489
rect 701070 111474 701094 111489
rect 701138 111474 701162 111489
rect 701206 111474 701230 111489
rect 701274 111474 701298 111489
rect 701342 111474 701366 111489
rect 701410 111474 701434 111489
rect 701478 111474 701502 111489
rect 701546 111474 701570 111489
rect 701614 111474 701638 111489
rect 701682 111474 701706 111489
rect 701750 111474 701774 111489
rect 701818 111474 701842 111489
rect 699322 111319 700322 111474
rect 699322 111285 700334 111319
rect 700922 111309 701922 111474
rect 707610 111319 708610 111379
rect 709211 111319 710211 111379
rect 700910 111285 701922 111309
rect 699322 111274 700322 111285
rect 700922 111274 701922 111285
rect 699392 111261 699416 111274
rect 699460 111261 699484 111274
rect 699528 111261 699552 111274
rect 699596 111261 699620 111274
rect 699664 111261 699688 111274
rect 699732 111261 699756 111274
rect 699800 111261 699824 111274
rect 699868 111261 699892 111274
rect 699936 111261 699960 111274
rect 700004 111261 700028 111274
rect 700072 111261 700096 111274
rect 700140 111261 700164 111274
rect 700208 111261 700232 111274
rect 700276 111261 700300 111274
rect 700934 111261 700958 111274
rect 701002 111261 701026 111274
rect 701070 111261 701094 111274
rect 701138 111261 701162 111274
rect 701206 111261 701230 111274
rect 701274 111261 701298 111274
rect 701342 111261 701366 111274
rect 701410 111261 701434 111274
rect 701478 111261 701502 111274
rect 701546 111261 701570 111274
rect 701614 111261 701638 111274
rect 701682 111261 701706 111274
rect 701750 111261 701774 111274
rect 701818 111261 701842 111274
rect 699322 110916 700322 110972
rect 700922 110916 701922 110972
rect 707610 110961 708610 111017
rect 709211 110961 710211 111017
rect 699322 110844 700322 110900
rect 700922 110844 701922 110900
rect 707610 110889 708610 110945
rect 709211 110889 710211 110945
rect 699322 110542 700322 110614
rect 700922 110542 701922 110614
rect 707610 110587 708610 110659
rect 709211 110587 710211 110659
rect 699392 110531 699426 110542
rect 699460 110531 699494 110542
rect 699528 110531 699562 110542
rect 699596 110531 699630 110542
rect 699664 110531 699698 110542
rect 699732 110531 699766 110542
rect 699800 110531 699834 110542
rect 699868 110531 699902 110542
rect 699936 110531 699970 110542
rect 700004 110531 700038 110542
rect 700072 110531 700106 110542
rect 700140 110531 700174 110542
rect 700208 110531 700242 110542
rect 700276 110531 700310 110542
rect 700934 110531 700968 110542
rect 701002 110531 701036 110542
rect 701070 110531 701104 110542
rect 701138 110531 701172 110542
rect 701206 110531 701240 110542
rect 701274 110531 701308 110542
rect 701342 110531 701376 110542
rect 701410 110531 701444 110542
rect 701478 110531 701512 110542
rect 701546 110531 701580 110542
rect 701614 110531 701648 110542
rect 701682 110531 701716 110542
rect 701750 110531 701784 110542
rect 701818 110531 701852 110542
rect 699392 110521 699450 110531
rect 699460 110521 699518 110531
rect 699528 110521 699586 110531
rect 699596 110521 699654 110531
rect 699664 110521 699722 110531
rect 699732 110521 699790 110531
rect 699800 110521 699858 110531
rect 699868 110521 699926 110531
rect 699936 110521 699994 110531
rect 700004 110521 700062 110531
rect 700072 110521 700130 110531
rect 700140 110521 700198 110531
rect 700208 110521 700266 110531
rect 700276 110521 700334 110531
rect 700934 110521 700992 110531
rect 701002 110521 701060 110531
rect 701070 110521 701128 110531
rect 701138 110521 701196 110531
rect 701206 110521 701264 110531
rect 701274 110521 701332 110531
rect 701342 110521 701400 110531
rect 701410 110521 701468 110531
rect 701478 110521 701536 110531
rect 701546 110521 701604 110531
rect 701614 110521 701672 110531
rect 701682 110521 701740 110531
rect 701750 110521 701808 110531
rect 701818 110521 701876 110531
rect 699368 110497 700334 110521
rect 700910 110497 701876 110521
rect 699392 110482 699416 110497
rect 699460 110482 699484 110497
rect 699528 110482 699552 110497
rect 699596 110482 699620 110497
rect 699664 110482 699688 110497
rect 699732 110482 699756 110497
rect 699800 110482 699824 110497
rect 699868 110482 699892 110497
rect 699936 110482 699960 110497
rect 700004 110482 700028 110497
rect 700072 110482 700096 110497
rect 700140 110482 700164 110497
rect 700208 110482 700232 110497
rect 700276 110482 700300 110497
rect 700934 110482 700958 110497
rect 701002 110482 701026 110497
rect 701070 110482 701094 110497
rect 701138 110482 701162 110497
rect 701206 110482 701230 110497
rect 701274 110482 701298 110497
rect 701342 110482 701366 110497
rect 701410 110482 701434 110497
rect 701478 110482 701502 110497
rect 701546 110482 701570 110497
rect 701614 110482 701638 110497
rect 701682 110482 701706 110497
rect 701750 110482 701774 110497
rect 701818 110482 701842 110497
rect 699322 110327 700322 110482
rect 699322 110293 700334 110327
rect 700922 110317 701922 110482
rect 707610 110327 708610 110387
rect 709211 110327 710211 110387
rect 711541 110345 711629 117461
rect 711892 116200 711942 117200
rect 712062 116200 712112 117200
rect 711892 115079 711942 116079
rect 712062 115079 712112 116079
rect 711892 113958 711942 114958
rect 712062 113958 712112 114958
rect 711892 112848 711942 113848
rect 712062 112848 712112 113848
rect 711892 111727 711942 112727
rect 712062 111727 712112 112727
rect 711892 110606 711942 111606
rect 712062 110606 712112 111606
rect 712409 110371 712431 117485
rect 712469 117459 712487 117501
rect 712499 117459 712505 117467
rect 712499 117455 712511 117459
rect 712539 117455 712557 117501
rect 713640 115461 713674 117785
rect 713750 117772 714750 117822
rect 717367 117820 717413 117853
rect 717367 117819 717379 117820
rect 717401 117819 717413 117820
rect 717401 117809 717600 117819
rect 717401 117786 717413 117809
rect 713750 117562 714750 117612
rect 713750 117446 714750 117496
rect 713750 117230 714750 117358
rect 713750 117014 714750 117070
rect 713750 116798 714750 116926
rect 713750 116588 714750 116638
rect 714478 116585 714750 116588
rect 715486 115931 715536 116931
rect 715696 115931 715824 116931
rect 715912 115931 715962 116931
rect 713641 115345 713663 115461
rect 713640 115309 713674 115345
rect 713750 115314 714750 115364
rect 713750 115158 714750 115214
rect 713750 115002 714750 115130
rect 713750 114846 714750 114974
rect 713750 114690 714750 114746
rect 716425 114709 716725 114721
rect 713750 114534 714750 114662
rect 716425 114596 717425 114646
rect 713750 114378 714750 114506
rect 716425 114440 717425 114568
rect 713750 114222 714750 114350
rect 716425 114284 717425 114340
rect 713750 114072 714750 114122
rect 713750 113956 714750 114006
rect 713750 113800 714750 113928
rect 713750 113644 714750 113772
rect 713750 113488 714750 113616
rect 715354 113587 715404 114187
rect 715504 113587 715560 114187
rect 715660 113587 715716 114187
rect 715816 113587 715872 114187
rect 715972 113587 716022 114187
rect 716425 114128 717425 114256
rect 716425 113978 717425 114028
rect 716425 113862 717425 113912
rect 716425 113706 717425 113834
rect 716425 113550 717425 113606
rect 716425 113394 717425 113522
rect 713750 113332 714750 113388
rect 713750 113176 714750 113304
rect 716425 113244 717425 113294
rect 713750 113020 714750 113148
rect 713750 112870 714750 112920
rect 713750 112742 714750 112792
rect 713750 112586 714750 112642
rect 713750 112436 714750 112486
rect 713750 112320 714350 112370
rect 713750 112164 714350 112292
rect 715510 112191 715560 113191
rect 715660 112191 715788 113191
rect 715816 112191 715944 113191
rect 715972 112191 716022 113191
rect 716425 113128 717425 113178
rect 716425 112972 717425 113028
rect 716425 112822 717425 112872
rect 716425 112706 717425 112756
rect 716425 112550 717425 112678
rect 716425 112394 717425 112522
rect 716425 112238 717425 112366
rect 716425 112082 717425 112210
rect 713750 112008 714350 112064
rect 713750 111852 714350 111980
rect 716425 111932 717425 111982
rect 713750 111696 714350 111752
rect 713750 111446 714350 111496
rect 714565 111443 714765 111455
rect 713750 111330 714750 111380
rect 713750 111120 714750 111170
rect 716413 111092 716447 111150
rect 713750 111004 714750 111054
rect 713750 110794 714750 110844
rect 713750 110678 714750 110728
rect 713750 110468 714750 110518
rect 713750 110352 714750 110402
rect 700910 110293 701922 110317
rect 699322 110282 700322 110293
rect 700922 110282 701922 110293
rect 711541 110311 711633 110345
rect 699392 110269 699416 110282
rect 699460 110269 699484 110282
rect 699528 110269 699552 110282
rect 699596 110269 699620 110282
rect 699664 110269 699688 110282
rect 699732 110269 699756 110282
rect 699800 110269 699824 110282
rect 699868 110269 699892 110282
rect 699936 110269 699960 110282
rect 700004 110269 700028 110282
rect 700072 110269 700096 110282
rect 700140 110269 700164 110282
rect 700208 110269 700232 110282
rect 700276 110269 700300 110282
rect 700934 110269 700958 110282
rect 701002 110269 701026 110282
rect 701070 110269 701094 110282
rect 701138 110269 701162 110282
rect 701206 110269 701230 110282
rect 701274 110269 701298 110282
rect 701342 110269 701366 110282
rect 701410 110269 701434 110282
rect 701478 110269 701502 110282
rect 701546 110269 701570 110282
rect 701614 110269 701638 110282
rect 701682 110269 701706 110282
rect 701750 110269 701774 110282
rect 701818 110269 701842 110282
rect 699322 109924 700322 109980
rect 700922 109924 701922 109980
rect 707610 109969 708610 110025
rect 709211 109969 710211 110025
rect 699322 109852 700322 109908
rect 700922 109852 701922 109908
rect 707610 109897 708610 109953
rect 709211 109897 710211 109953
rect 699322 109550 700322 109622
rect 700922 109550 701922 109622
rect 707610 109595 708610 109667
rect 709211 109595 710211 109667
rect 699392 109539 699426 109550
rect 699460 109539 699494 109550
rect 699528 109539 699562 109550
rect 699596 109539 699630 109550
rect 699664 109539 699698 109550
rect 699732 109539 699766 109550
rect 699800 109539 699834 109550
rect 699868 109539 699902 109550
rect 699936 109539 699970 109550
rect 700004 109539 700038 109550
rect 700072 109539 700106 109550
rect 700140 109539 700174 109550
rect 700208 109539 700242 109550
rect 700276 109539 700310 109550
rect 700934 109539 700968 109550
rect 701002 109539 701036 109550
rect 701070 109539 701104 109550
rect 701138 109539 701172 109550
rect 701206 109539 701240 109550
rect 701274 109539 701308 109550
rect 701342 109539 701376 109550
rect 701410 109539 701444 109550
rect 701478 109539 701512 109550
rect 701546 109539 701580 109550
rect 701614 109539 701648 109550
rect 701682 109539 701716 109550
rect 701750 109539 701784 109550
rect 701818 109539 701852 109550
rect 699392 109529 699450 109539
rect 699460 109529 699518 109539
rect 699528 109529 699586 109539
rect 699596 109529 699654 109539
rect 699664 109529 699722 109539
rect 699732 109529 699790 109539
rect 699800 109529 699858 109539
rect 699868 109529 699926 109539
rect 699936 109529 699994 109539
rect 700004 109529 700062 109539
rect 700072 109529 700130 109539
rect 700140 109529 700198 109539
rect 700208 109529 700266 109539
rect 700276 109529 700334 109539
rect 700934 109529 700992 109539
rect 701002 109529 701060 109539
rect 701070 109529 701128 109539
rect 701138 109529 701196 109539
rect 701206 109529 701264 109539
rect 701274 109529 701332 109539
rect 701342 109529 701400 109539
rect 701410 109529 701468 109539
rect 701478 109529 701536 109539
rect 701546 109529 701604 109539
rect 701614 109529 701672 109539
rect 701682 109529 701740 109539
rect 701750 109529 701808 109539
rect 701818 109529 701876 109539
rect 699368 109505 700334 109529
rect 700910 109505 701876 109529
rect 699392 109490 699416 109505
rect 699460 109490 699484 109505
rect 699528 109490 699552 109505
rect 699596 109490 699620 109505
rect 699664 109490 699688 109505
rect 699732 109490 699756 109505
rect 699800 109490 699824 109505
rect 699868 109490 699892 109505
rect 699936 109490 699960 109505
rect 700004 109490 700028 109505
rect 700072 109490 700096 109505
rect 700140 109490 700164 109505
rect 700208 109490 700232 109505
rect 700276 109490 700300 109505
rect 700934 109490 700958 109505
rect 701002 109490 701026 109505
rect 701070 109490 701094 109505
rect 701138 109490 701162 109505
rect 701206 109490 701230 109505
rect 701274 109490 701298 109505
rect 701342 109490 701366 109505
rect 701410 109490 701434 109505
rect 701478 109490 701502 109505
rect 701546 109490 701570 109505
rect 701614 109490 701638 109505
rect 701682 109490 701706 109505
rect 701750 109490 701774 109505
rect 701818 109490 701842 109505
rect 699322 109335 700322 109490
rect 699322 109301 700334 109335
rect 700922 109325 701922 109490
rect 707610 109335 708610 109395
rect 709211 109335 710211 109395
rect 700910 109301 701922 109325
rect 699322 109290 700322 109301
rect 700922 109290 701922 109301
rect 699392 109277 699416 109290
rect 699460 109277 699484 109290
rect 699528 109277 699552 109290
rect 699596 109277 699620 109290
rect 699664 109277 699688 109290
rect 699732 109277 699756 109290
rect 699800 109277 699824 109290
rect 699868 109277 699892 109290
rect 699936 109277 699960 109290
rect 700004 109277 700028 109290
rect 700072 109277 700096 109290
rect 700140 109277 700164 109290
rect 700208 109277 700232 109290
rect 700276 109277 700300 109290
rect 700934 109277 700958 109290
rect 701002 109277 701026 109290
rect 701070 109277 701094 109290
rect 701138 109277 701162 109290
rect 701206 109277 701230 109290
rect 701274 109277 701298 109290
rect 701342 109277 701366 109290
rect 701410 109277 701434 109290
rect 701478 109277 701502 109290
rect 701546 109277 701570 109290
rect 701614 109277 701638 109290
rect 701682 109277 701706 109290
rect 701750 109277 701774 109290
rect 701818 109277 701842 109290
rect 699322 108932 700322 108988
rect 700922 108932 701922 108988
rect 707610 108977 708610 109033
rect 709211 108977 710211 109033
rect 699322 108860 700322 108916
rect 700922 108860 701922 108916
rect 707610 108905 708610 108961
rect 709211 108905 710211 108961
rect 699322 108558 700322 108630
rect 700922 108558 701922 108630
rect 707610 108603 708610 108675
rect 709211 108603 710211 108675
rect 699392 108547 699426 108558
rect 699460 108547 699494 108558
rect 699528 108547 699562 108558
rect 699596 108547 699630 108558
rect 699664 108547 699698 108558
rect 699732 108547 699766 108558
rect 699800 108547 699834 108558
rect 699868 108547 699902 108558
rect 699936 108547 699970 108558
rect 700004 108547 700038 108558
rect 700072 108547 700106 108558
rect 700140 108547 700174 108558
rect 700208 108547 700242 108558
rect 700276 108547 700310 108558
rect 700934 108547 700968 108558
rect 701002 108547 701036 108558
rect 701070 108547 701104 108558
rect 701138 108547 701172 108558
rect 701206 108547 701240 108558
rect 701274 108547 701308 108558
rect 701342 108547 701376 108558
rect 701410 108547 701444 108558
rect 701478 108547 701512 108558
rect 701546 108547 701580 108558
rect 701614 108547 701648 108558
rect 701682 108547 701716 108558
rect 701750 108547 701784 108558
rect 701818 108547 701852 108558
rect 699392 108537 699450 108547
rect 699460 108537 699518 108547
rect 699528 108537 699586 108547
rect 699596 108537 699654 108547
rect 699664 108537 699722 108547
rect 699732 108537 699790 108547
rect 699800 108537 699858 108547
rect 699868 108537 699926 108547
rect 699936 108537 699994 108547
rect 700004 108537 700062 108547
rect 700072 108537 700130 108547
rect 700140 108537 700198 108547
rect 700208 108537 700266 108547
rect 700276 108537 700334 108547
rect 700934 108537 700992 108547
rect 701002 108537 701060 108547
rect 701070 108537 701128 108547
rect 701138 108537 701196 108547
rect 701206 108537 701264 108547
rect 701274 108537 701332 108547
rect 701342 108537 701400 108547
rect 701410 108537 701468 108547
rect 701478 108537 701536 108547
rect 701546 108537 701604 108547
rect 701614 108537 701672 108547
rect 701682 108537 701740 108547
rect 701750 108537 701808 108547
rect 701818 108537 701876 108547
rect 699368 108513 700334 108537
rect 700910 108513 701876 108537
rect 699392 108498 699416 108513
rect 699460 108498 699484 108513
rect 699528 108498 699552 108513
rect 699596 108498 699620 108513
rect 699664 108498 699688 108513
rect 699732 108498 699756 108513
rect 699800 108498 699824 108513
rect 699868 108498 699892 108513
rect 699936 108498 699960 108513
rect 700004 108498 700028 108513
rect 700072 108498 700096 108513
rect 700140 108498 700164 108513
rect 700208 108498 700232 108513
rect 700276 108498 700300 108513
rect 700934 108498 700958 108513
rect 701002 108498 701026 108513
rect 701070 108498 701094 108513
rect 701138 108498 701162 108513
rect 701206 108498 701230 108513
rect 701274 108498 701298 108513
rect 701342 108498 701366 108513
rect 701410 108498 701434 108513
rect 701478 108498 701502 108513
rect 701546 108498 701570 108513
rect 701614 108498 701638 108513
rect 701682 108498 701706 108513
rect 701750 108498 701774 108513
rect 701818 108498 701842 108513
rect 699322 108343 700322 108498
rect 699322 108309 700334 108343
rect 700922 108333 701922 108498
rect 707610 108343 708610 108403
rect 709211 108343 710211 108403
rect 700910 108309 701922 108333
rect 699322 108298 700322 108309
rect 700922 108298 701922 108309
rect 699392 108285 699416 108298
rect 699460 108285 699484 108298
rect 699528 108285 699552 108298
rect 699596 108285 699620 108298
rect 699664 108285 699688 108298
rect 699732 108285 699756 108298
rect 699800 108285 699824 108298
rect 699868 108285 699892 108298
rect 699936 108285 699960 108298
rect 700004 108285 700028 108298
rect 700072 108285 700096 108298
rect 700140 108285 700164 108298
rect 700208 108285 700232 108298
rect 700276 108285 700300 108298
rect 700934 108285 700958 108298
rect 701002 108285 701026 108298
rect 701070 108285 701094 108298
rect 701138 108285 701162 108298
rect 701206 108285 701230 108298
rect 701274 108285 701298 108298
rect 701342 108285 701366 108298
rect 701410 108285 701434 108298
rect 701478 108285 701502 108298
rect 701546 108285 701570 108298
rect 701614 108285 701638 108298
rect 701682 108285 701706 108298
rect 701750 108285 701774 108298
rect 701818 108285 701842 108298
rect 699322 107940 700322 107996
rect 700922 107940 701922 107996
rect 707610 107985 708610 108041
rect 709211 107985 710211 108041
rect 699322 107868 700322 107924
rect 700922 107868 701922 107924
rect 707610 107913 708610 107969
rect 709211 107913 710211 107969
rect 699322 107566 700322 107638
rect 700922 107566 701922 107638
rect 707610 107611 708610 107683
rect 709211 107611 710211 107683
rect 699392 107555 699426 107566
rect 699460 107555 699494 107566
rect 699528 107555 699562 107566
rect 699596 107555 699630 107566
rect 699664 107555 699698 107566
rect 699732 107555 699766 107566
rect 699800 107555 699834 107566
rect 699868 107555 699902 107566
rect 699936 107555 699970 107566
rect 700004 107555 700038 107566
rect 700072 107555 700106 107566
rect 700140 107555 700174 107566
rect 700208 107555 700242 107566
rect 700276 107555 700310 107566
rect 700934 107555 700968 107566
rect 701002 107555 701036 107566
rect 701070 107555 701104 107566
rect 701138 107555 701172 107566
rect 701206 107555 701240 107566
rect 701274 107555 701308 107566
rect 701342 107555 701376 107566
rect 701410 107555 701444 107566
rect 701478 107555 701512 107566
rect 701546 107555 701580 107566
rect 701614 107555 701648 107566
rect 701682 107555 701716 107566
rect 701750 107555 701784 107566
rect 701818 107555 701852 107566
rect 699392 107545 699450 107555
rect 699460 107545 699518 107555
rect 699528 107545 699586 107555
rect 699596 107545 699654 107555
rect 699664 107545 699722 107555
rect 699732 107545 699790 107555
rect 699800 107545 699858 107555
rect 699868 107545 699926 107555
rect 699936 107545 699994 107555
rect 700004 107545 700062 107555
rect 700072 107545 700130 107555
rect 700140 107545 700198 107555
rect 700208 107545 700266 107555
rect 700276 107545 700334 107555
rect 700934 107545 700992 107555
rect 701002 107545 701060 107555
rect 701070 107545 701128 107555
rect 701138 107545 701196 107555
rect 701206 107545 701264 107555
rect 701274 107545 701332 107555
rect 701342 107545 701400 107555
rect 701410 107545 701468 107555
rect 701478 107545 701536 107555
rect 701546 107545 701604 107555
rect 701614 107545 701672 107555
rect 701682 107545 701740 107555
rect 701750 107545 701808 107555
rect 701818 107545 701876 107555
rect 699368 107521 700334 107545
rect 700910 107521 701876 107545
rect 699392 107506 699416 107521
rect 699460 107506 699484 107521
rect 699528 107506 699552 107521
rect 699596 107506 699620 107521
rect 699664 107506 699688 107521
rect 699732 107506 699756 107521
rect 699800 107506 699824 107521
rect 699868 107506 699892 107521
rect 699936 107506 699960 107521
rect 700004 107506 700028 107521
rect 700072 107506 700096 107521
rect 700140 107506 700164 107521
rect 700208 107506 700232 107521
rect 700276 107506 700300 107521
rect 700934 107506 700958 107521
rect 701002 107506 701026 107521
rect 701070 107506 701094 107521
rect 701138 107506 701162 107521
rect 701206 107506 701230 107521
rect 701274 107506 701298 107521
rect 701342 107506 701366 107521
rect 701410 107506 701434 107521
rect 701478 107506 701502 107521
rect 701546 107506 701570 107521
rect 701614 107506 701638 107521
rect 701682 107506 701706 107521
rect 701750 107506 701774 107521
rect 701818 107506 701842 107521
rect 699322 107351 700322 107506
rect 699322 107317 700334 107351
rect 700922 107341 701922 107506
rect 705107 107360 705173 107376
rect 707610 107351 708610 107411
rect 709211 107351 710211 107411
rect 700910 107317 701922 107341
rect 699322 107306 700322 107317
rect 700922 107306 701922 107317
rect 699392 107293 699416 107306
rect 699460 107293 699484 107306
rect 699528 107293 699552 107306
rect 699596 107293 699620 107306
rect 699664 107293 699688 107306
rect 699732 107293 699756 107306
rect 699800 107293 699824 107306
rect 699868 107293 699892 107306
rect 699936 107293 699960 107306
rect 700004 107293 700028 107306
rect 700072 107293 700096 107306
rect 700140 107293 700164 107306
rect 700208 107293 700232 107306
rect 700276 107293 700300 107306
rect 700934 107293 700958 107306
rect 701002 107293 701026 107306
rect 701070 107293 701094 107306
rect 701138 107293 701162 107306
rect 701206 107293 701230 107306
rect 701274 107293 701298 107306
rect 701342 107293 701366 107306
rect 701410 107293 701434 107306
rect 701478 107293 701502 107306
rect 701546 107293 701570 107306
rect 701614 107293 701638 107306
rect 701682 107293 701706 107306
rect 701750 107293 701774 107306
rect 701818 107293 701842 107306
rect 699322 106948 700322 107004
rect 700922 106948 701922 107004
rect 707610 106993 708610 107049
rect 709211 106993 710211 107049
rect 699322 106876 700322 106932
rect 700922 106876 701922 106932
rect 707610 106921 708610 106977
rect 709211 106921 710211 106977
rect 699322 106574 700322 106646
rect 700922 106574 701922 106646
rect 707610 106619 708610 106691
rect 709211 106619 710211 106691
rect 699392 106563 699426 106574
rect 699460 106563 699494 106574
rect 699528 106563 699562 106574
rect 699596 106563 699630 106574
rect 699664 106563 699698 106574
rect 699732 106563 699766 106574
rect 699800 106563 699834 106574
rect 699868 106563 699902 106574
rect 699936 106563 699970 106574
rect 700004 106563 700038 106574
rect 700072 106563 700106 106574
rect 700140 106563 700174 106574
rect 700208 106563 700242 106574
rect 700276 106563 700310 106574
rect 700934 106563 700968 106574
rect 701002 106563 701036 106574
rect 701070 106563 701104 106574
rect 701138 106563 701172 106574
rect 701206 106563 701240 106574
rect 701274 106563 701308 106574
rect 701342 106563 701376 106574
rect 701410 106563 701444 106574
rect 701478 106563 701512 106574
rect 701546 106563 701580 106574
rect 701614 106563 701648 106574
rect 701682 106563 701716 106574
rect 701750 106563 701784 106574
rect 701818 106563 701852 106574
rect 699392 106553 699450 106563
rect 699460 106553 699518 106563
rect 699528 106553 699586 106563
rect 699596 106553 699654 106563
rect 699664 106553 699722 106563
rect 699732 106553 699790 106563
rect 699800 106553 699858 106563
rect 699868 106553 699926 106563
rect 699936 106553 699994 106563
rect 700004 106553 700062 106563
rect 700072 106553 700130 106563
rect 700140 106553 700198 106563
rect 700208 106553 700266 106563
rect 700276 106553 700334 106563
rect 700934 106553 700992 106563
rect 701002 106553 701060 106563
rect 701070 106553 701128 106563
rect 701138 106553 701196 106563
rect 701206 106553 701264 106563
rect 701274 106553 701332 106563
rect 701342 106553 701400 106563
rect 701410 106553 701468 106563
rect 701478 106553 701536 106563
rect 701546 106553 701604 106563
rect 701614 106553 701672 106563
rect 701682 106553 701740 106563
rect 701750 106553 701808 106563
rect 701818 106553 701876 106563
rect 699368 106529 700334 106553
rect 700910 106529 701876 106553
rect 699392 106514 699416 106529
rect 699460 106514 699484 106529
rect 699528 106514 699552 106529
rect 699596 106514 699620 106529
rect 699664 106514 699688 106529
rect 699732 106514 699756 106529
rect 699800 106514 699824 106529
rect 699868 106514 699892 106529
rect 699936 106514 699960 106529
rect 700004 106514 700028 106529
rect 700072 106514 700096 106529
rect 700140 106514 700164 106529
rect 700208 106514 700232 106529
rect 700276 106514 700300 106529
rect 700934 106514 700958 106529
rect 701002 106514 701026 106529
rect 701070 106514 701094 106529
rect 701138 106514 701162 106529
rect 701206 106514 701230 106529
rect 701274 106514 701298 106529
rect 701342 106514 701366 106529
rect 701410 106514 701434 106529
rect 701478 106514 701502 106529
rect 701546 106514 701570 106529
rect 701614 106514 701638 106529
rect 701682 106514 701706 106529
rect 701750 106514 701774 106529
rect 701818 106514 701842 106529
rect 699322 106359 700322 106514
rect 699322 106325 700334 106359
rect 700922 106349 701922 106514
rect 707610 106359 708610 106419
rect 709211 106359 710211 106419
rect 700910 106325 701922 106349
rect 699322 106314 700322 106325
rect 700922 106314 701922 106325
rect 699392 106301 699416 106314
rect 699460 106301 699484 106314
rect 699528 106301 699552 106314
rect 699596 106301 699620 106314
rect 699664 106301 699688 106314
rect 699732 106301 699756 106314
rect 699800 106301 699824 106314
rect 699868 106301 699892 106314
rect 699936 106301 699960 106314
rect 700004 106301 700028 106314
rect 700072 106301 700096 106314
rect 700140 106301 700164 106314
rect 700208 106301 700232 106314
rect 700276 106301 700300 106314
rect 700934 106301 700958 106314
rect 701002 106301 701026 106314
rect 701070 106301 701094 106314
rect 701138 106301 701162 106314
rect 701206 106301 701230 106314
rect 701274 106301 701298 106314
rect 701342 106301 701366 106314
rect 701410 106301 701434 106314
rect 701478 106301 701502 106314
rect 701546 106301 701570 106314
rect 701614 106301 701638 106314
rect 701682 106301 701706 106314
rect 701750 106301 701774 106314
rect 701818 106301 701842 106314
rect 709211 106148 710211 106152
rect 707574 106099 707610 106134
rect 708610 106099 708646 106134
rect 707574 106098 708646 106099
rect 707574 106057 707610 106098
rect 708610 106057 708646 106098
rect 699322 105956 700322 106012
rect 700922 105956 701922 106012
rect 707574 106001 708646 106057
rect 707574 105964 707610 106001
rect 708610 105964 708646 106001
rect 707574 105959 708646 105964
rect 699322 105884 700322 105940
rect 700922 105884 701922 105940
rect 707574 105924 707610 105959
rect 708610 105924 708646 105959
rect 709175 106098 710247 106134
rect 709175 106057 709211 106098
rect 710211 106057 710247 106098
rect 709175 106001 710247 106057
rect 709175 105964 709211 106001
rect 710211 105964 710247 106001
rect 709175 105936 710247 105964
rect 709175 105924 709211 105936
rect 710211 105924 710247 105936
rect 707610 105713 708610 105785
rect 709211 105713 710211 105785
rect 699322 105623 700322 105673
rect 700922 105623 701922 105673
rect 707610 105523 708610 105617
rect 707610 105513 708644 105523
rect 709211 105513 710211 105591
rect 711541 105437 711629 110311
rect 713750 110136 714750 110264
rect 716417 110152 717417 110202
rect 711892 109049 711942 110049
rect 712062 109049 712112 110049
rect 713750 109920 714750 110048
rect 716417 109996 717417 110052
rect 716417 109846 717417 109896
rect 713750 109704 714750 109832
rect 716417 109730 717017 109780
rect 716417 109580 717017 109630
rect 713750 109488 714750 109544
rect 716417 109464 717417 109514
rect 713750 109272 714750 109400
rect 716417 109308 717417 109364
rect 713750 109056 714750 109184
rect 716417 109152 717417 109280
rect 716417 108996 717417 109052
rect 711892 107928 711942 108928
rect 712062 107928 712112 108928
rect 713750 108840 714750 108968
rect 716417 108840 717417 108968
rect 713750 108624 714750 108752
rect 716417 108684 717417 108740
rect 716417 108474 717417 108524
rect 713750 108408 714750 108464
rect 716417 108308 717417 108358
rect 713750 108192 714750 108248
rect 716417 108152 717417 108280
rect 713750 107976 714750 108104
rect 716417 107996 717417 108052
rect 711892 106807 711942 107807
rect 712062 106807 712112 107807
rect 713750 107760 714750 107888
rect 716417 107780 717417 107836
rect 713750 107544 714750 107672
rect 716417 107570 717417 107620
rect 713750 107328 714750 107456
rect 716417 107454 717417 107504
rect 716417 107298 717417 107426
rect 713750 107118 714750 107168
rect 716417 107148 717417 107198
rect 711892 105697 711942 106697
rect 712062 105697 712112 106697
rect 714686 106357 714794 106424
rect 714645 106323 714794 106357
rect 716071 106357 716074 106358
rect 716071 106356 716072 106357
rect 716073 106356 716074 106357
rect 716071 106355 716074 106356
rect 716208 106357 716211 106358
rect 716208 106356 716209 106357
rect 716210 106356 716211 106357
rect 716208 106355 716211 106356
rect 714964 106247 715998 106329
rect 716284 106247 717318 106329
rect 705107 105336 705173 105352
rect 711541 105302 711633 105437
rect 714175 105398 714225 105998
rect 714425 105398 714475 105998
rect 711579 105301 711595 105302
rect 714781 105191 714863 106226
rect 715134 105955 715828 106037
rect 714686 105123 714863 105191
rect 714645 105089 714863 105123
rect 680215 104880 680815 104936
rect 686719 104893 686739 104917
rect 686743 104893 686753 104917
rect 686719 104859 686757 104893
rect 686719 104822 686739 104859
rect 686743 104822 686753 104859
rect 692428 104850 693028 104978
rect 698017 104947 698210 104983
rect 698084 104935 698210 104947
rect 702756 104959 703645 104983
rect 702756 104935 702853 104959
rect 698084 104828 702853 104935
rect 686719 104788 686757 104822
rect 680215 104704 680815 104760
rect 686719 104751 686739 104788
rect 686743 104751 686753 104788
rect 686719 104741 686757 104751
rect 686699 104717 686767 104741
rect 686719 104704 686739 104717
rect 686743 104704 686753 104717
rect 686719 104695 686753 104704
rect 686719 104693 686743 104695
rect 692428 104694 693028 104750
rect 686685 104656 686709 104680
rect 686743 104656 686767 104680
rect 678799 104503 679399 104553
rect 680215 104534 680815 104584
rect 692428 104538 693028 104666
rect 680593 104531 680815 104534
rect 682009 104501 682069 104516
rect 682024 104465 682054 104501
rect 683708 104387 684308 104437
rect 678799 104327 679399 104383
rect 692428 104382 693028 104510
rect 714781 104308 714863 105089
rect 715063 104609 715145 105915
rect 715342 105752 715382 105792
rect 715582 105752 715622 105792
rect 715289 104777 715339 105719
rect 715382 105668 715422 105752
rect 715542 105668 715582 105752
rect 715633 104777 715683 105719
rect 715382 104672 715422 104756
rect 715542 104672 715582 104756
rect 715342 104632 715382 104672
rect 715582 104632 715622 104672
rect 715815 104609 715897 105915
rect 715134 104387 715828 104469
rect 716100 104308 716182 106226
rect 716454 105955 717148 106037
rect 716385 104609 716467 105915
rect 716660 105752 716700 105792
rect 716900 105752 716940 105792
rect 716599 104777 716649 105719
rect 716700 105668 716740 105752
rect 716860 105668 716900 105752
rect 716943 104777 716993 105719
rect 716700 104672 716740 104756
rect 716860 104672 716900 104756
rect 716660 104632 716700 104672
rect 716900 104632 716940 104672
rect 717137 104609 717219 105915
rect 716454 104387 717148 104469
rect 717419 104308 717501 106226
rect 683708 104237 684308 104287
rect 692428 104232 693028 104282
rect 678799 104157 679399 104207
rect 684565 104160 684790 104168
rect 696597 104000 696600 104120
rect 714964 104095 715998 104177
rect 716284 104095 717318 104177
rect 21000 77000 21003 77120
rect 282 76623 1316 76705
rect 1602 76623 2636 76705
rect 32810 76662 33035 76670
rect 38201 76593 38801 76643
rect 24572 76518 25172 76568
rect 33292 76513 33892 76563
rect 99 74574 181 76492
rect 452 76331 1146 76413
rect 381 74885 463 76191
rect 660 76128 700 76168
rect 900 76128 940 76168
rect 700 76044 740 76128
rect 860 76044 900 76128
rect 607 75081 657 76023
rect 700 75048 740 75132
rect 860 75048 900 75132
rect 951 75081 1001 76023
rect 660 75008 700 75048
rect 900 75008 940 75048
rect 1133 74885 1215 76191
rect 452 74763 1146 74845
rect 1418 74574 1500 76492
rect 1772 76331 2466 76413
rect 1703 74885 1785 76191
rect 1978 76128 2018 76168
rect 2218 76128 2258 76168
rect 2018 76044 2058 76128
rect 2178 76044 2218 76128
rect 1917 75081 1967 76023
rect 2018 75048 2058 75132
rect 2178 75048 2218 75132
rect 2261 75081 2311 76023
rect 1978 75008 2018 75048
rect 2218 75008 2258 75048
rect 2455 74885 2537 76191
rect 2737 75779 2819 76492
rect 24572 76362 25172 76490
rect 38201 76417 38801 76473
rect 33292 76363 33892 76413
rect 24572 76206 25172 76334
rect 35546 76299 35576 76335
rect 36785 76329 36935 76341
rect 35531 76284 35591 76299
rect 36785 76216 37385 76266
rect 38201 76247 38801 76297
rect 30833 76120 30857 76144
rect 30891 76120 30915 76144
rect 24572 76050 25172 76106
rect 30857 76105 30881 76107
rect 30857 76096 30887 76105
rect 30867 76083 30887 76096
rect 30891 76083 30907 76120
rect 30833 76059 30857 76083
rect 30867 76049 30911 76083
rect 14747 75865 19516 75972
rect 24572 75894 25172 76022
rect 30867 76012 30887 76049
rect 30891 76012 30907 76049
rect 36785 76040 37385 76096
rect 30867 75978 30911 76012
rect 30867 75941 30887 75978
rect 30891 75941 30907 75978
rect 30867 75907 30911 75941
rect 30867 75883 30887 75907
rect 30891 75883 30907 75907
rect 14747 75841 14844 75865
rect 13955 75817 14844 75841
rect 19390 75853 19516 75865
rect 19390 75841 19583 75853
rect 19390 75817 19605 75841
rect 19639 75817 19673 75841
rect 19707 75817 19741 75841
rect 19775 75817 19809 75841
rect 19843 75817 19877 75841
rect 19911 75817 19945 75841
rect 19979 75817 20013 75841
rect 20047 75817 20081 75841
rect 20115 75817 20149 75841
rect 20183 75817 20217 75841
rect 20251 75817 20285 75841
rect 20319 75817 20353 75841
rect 20387 75817 20421 75841
rect 20455 75817 20489 75841
rect 20523 75817 20557 75841
rect 20591 75817 20625 75841
rect 20659 75817 20693 75841
rect 2737 75711 2914 75779
rect 1772 74763 2466 74845
rect 2737 74574 2819 75711
rect 2848 75677 2955 75711
rect 6005 75498 6021 75499
rect 3125 74802 3175 75402
rect 3375 74802 3425 75402
rect 5967 75363 6059 75498
rect 12427 75448 12493 75464
rect 282 74471 1316 74553
rect 1602 74471 2636 74553
rect 2806 74477 2914 74545
rect 1389 74444 1392 74445
rect 1389 74443 1390 74444
rect 1391 74443 1392 74444
rect 1389 74442 1392 74443
rect 1526 74444 1529 74445
rect 1526 74443 1527 74444
rect 1528 74443 1529 74444
rect 2848 74443 2955 74477
rect 1526 74442 1529 74443
rect 5488 74103 5538 75103
rect 5658 74103 5708 75103
rect 183 73602 1183 73652
rect 2850 73632 3850 73682
rect 183 73446 1183 73574
rect 2850 73416 3850 73544
rect 183 73296 1183 73346
rect 183 73180 1183 73230
rect 2850 73200 3850 73328
rect 183 72964 1183 73020
rect 2850 72984 3850 73112
rect 5488 72993 5538 73993
rect 5658 72993 5708 73993
rect 183 72748 1183 72804
rect 2850 72768 3850 72896
rect 183 72592 1183 72720
rect 2850 72552 3850 72608
rect 183 72442 1183 72492
rect 2850 72336 3850 72392
rect 183 72276 1183 72326
rect 2850 72120 3850 72248
rect 183 72060 1183 72116
rect 183 71904 1183 72032
rect 2850 71904 3850 72032
rect 5488 71872 5538 72872
rect 5658 71872 5708 72872
rect 183 71748 1183 71804
rect 183 71592 1183 71720
rect 2850 71688 3850 71816
rect 183 71436 1183 71492
rect 2850 71472 3850 71600
rect 183 71286 1183 71336
rect 2850 71256 3850 71312
rect 583 71170 1183 71220
rect 583 71020 1183 71070
rect 2850 71040 3850 71168
rect 183 70904 1183 70954
rect 2850 70824 3850 70952
rect 183 70748 1183 70804
rect 5488 70751 5538 71751
rect 5658 70751 5708 71751
rect 183 70598 1183 70648
rect 2850 70608 3850 70736
rect 5971 70489 6059 75363
rect 7406 75287 7440 75321
rect 7477 75287 7511 75321
rect 7551 75287 7585 75321
rect 7622 75287 7656 75321
rect 7696 75287 7730 75321
rect 7767 75287 7801 75321
rect 7841 75287 7875 75321
rect 7912 75287 7946 75321
rect 7986 75287 8020 75321
rect 8057 75287 8091 75321
rect 8131 75287 8165 75321
rect 8202 75287 8236 75321
rect 8296 75287 8330 75321
rect 8381 75311 8423 75321
rect 8381 75287 8389 75311
rect 8415 75287 8423 75311
rect 8956 75311 8996 75321
rect 8956 75287 8962 75311
rect 8990 75287 8996 75311
rect 9044 75287 9078 75321
rect 9120 75287 9154 75321
rect 9197 75287 9231 75321
rect 9291 75287 9325 75321
rect 9362 75287 9396 75321
rect 9436 75287 9470 75321
rect 9507 75287 9541 75321
rect 9581 75287 9615 75321
rect 9652 75287 9686 75321
rect 9726 75287 9760 75321
rect 9797 75287 9831 75321
rect 9871 75287 9905 75321
rect 9942 75287 9976 75321
rect 7389 75277 7406 75287
rect 7440 75277 7477 75287
rect 7511 75277 7551 75287
rect 7585 75277 7622 75287
rect 7656 75277 7696 75287
rect 7730 75277 7767 75287
rect 7801 75277 7841 75287
rect 7875 75277 7912 75287
rect 7946 75277 7986 75287
rect 8020 75277 8057 75287
rect 8091 75277 8131 75287
rect 8165 75277 8202 75287
rect 8236 75277 8296 75287
rect 8330 75277 8381 75287
rect 8389 75277 8423 75287
rect 8990 75277 9044 75287
rect 9078 75277 9120 75287
rect 9154 75277 9197 75287
rect 9231 75277 9291 75287
rect 9325 75277 9362 75287
rect 9396 75277 9436 75287
rect 9470 75277 9507 75287
rect 9541 75277 9581 75287
rect 9615 75277 9652 75287
rect 9686 75277 9726 75287
rect 9760 75277 9797 75287
rect 9831 75277 9871 75287
rect 9905 75277 9942 75287
rect 9976 75277 9990 75287
rect 7389 75209 8389 75277
rect 8990 75183 9990 75277
rect 7389 75087 8389 75147
rect 8990 75087 9990 75147
rect 15678 75127 16678 75177
rect 17278 75127 18278 75177
rect 7353 74864 7389 74876
rect 8389 74864 8425 74876
rect 7353 74840 8425 74864
rect 7353 74799 7389 74840
rect 8389 74799 8425 74840
rect 7353 74743 8425 74799
rect 7353 74706 7389 74743
rect 8389 74706 8425 74743
rect 7353 74666 8425 74706
rect 8954 74841 8990 74876
rect 9990 74841 10026 74876
rect 15678 74860 16678 74916
rect 17278 74860 18278 74916
rect 8954 74840 10026 74841
rect 8954 74799 8990 74840
rect 9990 74799 10026 74840
rect 8954 74743 10026 74799
rect 15678 74788 16678 74844
rect 17278 74788 18278 74844
rect 8954 74706 8990 74743
rect 9990 74706 10026 74743
rect 8954 74701 10026 74706
rect 8954 74666 8990 74701
rect 9990 74666 10026 74701
rect 7389 74441 8389 74513
rect 8990 74441 9990 74513
rect 15678 74486 16678 74558
rect 17278 74486 18278 74558
rect 15748 74475 15782 74486
rect 15816 74475 15850 74486
rect 15884 74475 15918 74486
rect 15952 74475 15986 74486
rect 16020 74475 16054 74486
rect 16088 74475 16122 74486
rect 16156 74475 16190 74486
rect 16224 74475 16258 74486
rect 16292 74475 16326 74486
rect 16360 74475 16394 74486
rect 16428 74475 16462 74486
rect 16496 74475 16530 74486
rect 16564 74475 16598 74486
rect 16632 74475 16666 74486
rect 17290 74475 17324 74486
rect 17358 74475 17392 74486
rect 17426 74475 17460 74486
rect 17494 74475 17528 74486
rect 17562 74475 17596 74486
rect 17630 74475 17664 74486
rect 17698 74475 17732 74486
rect 17766 74475 17800 74486
rect 17834 74475 17868 74486
rect 17902 74475 17936 74486
rect 17970 74475 18004 74486
rect 18038 74475 18072 74486
rect 18106 74475 18140 74486
rect 18174 74475 18208 74486
rect 15748 74465 15806 74475
rect 15816 74465 15874 74475
rect 15884 74465 15942 74475
rect 15952 74465 16010 74475
rect 16020 74465 16078 74475
rect 16088 74465 16146 74475
rect 16156 74465 16214 74475
rect 16224 74465 16282 74475
rect 16292 74465 16350 74475
rect 16360 74465 16418 74475
rect 16428 74465 16486 74475
rect 16496 74465 16554 74475
rect 16564 74465 16622 74475
rect 16632 74465 16690 74475
rect 17290 74465 17348 74475
rect 17358 74465 17416 74475
rect 17426 74465 17484 74475
rect 17494 74465 17552 74475
rect 17562 74465 17620 74475
rect 17630 74465 17688 74475
rect 17698 74465 17756 74475
rect 17766 74465 17824 74475
rect 17834 74465 17892 74475
rect 17902 74465 17960 74475
rect 17970 74465 18028 74475
rect 18038 74465 18096 74475
rect 18106 74465 18164 74475
rect 18174 74465 18232 74475
rect 15724 74441 16690 74465
rect 17266 74441 18232 74465
rect 15748 74426 15772 74441
rect 15816 74426 15840 74441
rect 15884 74426 15908 74441
rect 15952 74426 15976 74441
rect 16020 74426 16044 74441
rect 16088 74426 16112 74441
rect 16156 74426 16180 74441
rect 16224 74426 16248 74441
rect 16292 74426 16316 74441
rect 16360 74426 16384 74441
rect 16428 74426 16452 74441
rect 16496 74426 16520 74441
rect 16564 74426 16588 74441
rect 16632 74426 16656 74441
rect 17290 74426 17314 74441
rect 17358 74426 17382 74441
rect 17426 74426 17450 74441
rect 17494 74426 17518 74441
rect 17562 74426 17586 74441
rect 17630 74426 17654 74441
rect 17698 74426 17722 74441
rect 17766 74426 17790 74441
rect 17834 74426 17858 74441
rect 17902 74426 17926 74441
rect 17970 74426 17994 74441
rect 18038 74426 18062 74441
rect 18106 74426 18130 74441
rect 18174 74426 18198 74441
rect 15678 74271 16678 74426
rect 7389 74181 8389 74241
rect 8990 74181 9990 74241
rect 15678 74237 16690 74271
rect 17278 74261 18278 74426
rect 17266 74237 18278 74261
rect 15678 74226 16678 74237
rect 17278 74226 18278 74237
rect 15748 74213 15772 74226
rect 15816 74213 15840 74226
rect 15884 74213 15908 74226
rect 15952 74213 15976 74226
rect 16020 74213 16044 74226
rect 16088 74213 16112 74226
rect 16156 74213 16180 74226
rect 16224 74213 16248 74226
rect 16292 74213 16316 74226
rect 16360 74213 16384 74226
rect 16428 74213 16452 74226
rect 16496 74213 16520 74226
rect 16564 74213 16588 74226
rect 16632 74213 16656 74226
rect 17290 74213 17314 74226
rect 17358 74213 17382 74226
rect 17426 74213 17450 74226
rect 17494 74213 17518 74226
rect 17562 74213 17586 74226
rect 17630 74213 17654 74226
rect 17698 74213 17722 74226
rect 17766 74213 17790 74226
rect 17834 74213 17858 74226
rect 17902 74213 17926 74226
rect 17970 74213 17994 74226
rect 18038 74213 18062 74226
rect 18106 74213 18130 74226
rect 18174 74213 18198 74226
rect 7389 73823 8389 73879
rect 8990 73823 9990 73879
rect 15678 73868 16678 73924
rect 17278 73868 18278 73924
rect 7389 73751 8389 73807
rect 8990 73751 9990 73807
rect 15678 73796 16678 73852
rect 17278 73796 18278 73852
rect 7389 73449 8389 73521
rect 8990 73449 9990 73521
rect 15678 73494 16678 73566
rect 17278 73494 18278 73566
rect 15748 73483 15782 73494
rect 15816 73483 15850 73494
rect 15884 73483 15918 73494
rect 15952 73483 15986 73494
rect 16020 73483 16054 73494
rect 16088 73483 16122 73494
rect 16156 73483 16190 73494
rect 16224 73483 16258 73494
rect 16292 73483 16326 73494
rect 16360 73483 16394 73494
rect 16428 73483 16462 73494
rect 16496 73483 16530 73494
rect 16564 73483 16598 73494
rect 16632 73483 16666 73494
rect 17290 73483 17324 73494
rect 17358 73483 17392 73494
rect 17426 73483 17460 73494
rect 17494 73483 17528 73494
rect 17562 73483 17596 73494
rect 17630 73483 17664 73494
rect 17698 73483 17732 73494
rect 17766 73483 17800 73494
rect 17834 73483 17868 73494
rect 17902 73483 17936 73494
rect 17970 73483 18004 73494
rect 18038 73483 18072 73494
rect 18106 73483 18140 73494
rect 18174 73483 18208 73494
rect 15748 73473 15806 73483
rect 15816 73473 15874 73483
rect 15884 73473 15942 73483
rect 15952 73473 16010 73483
rect 16020 73473 16078 73483
rect 16088 73473 16146 73483
rect 16156 73473 16214 73483
rect 16224 73473 16282 73483
rect 16292 73473 16350 73483
rect 16360 73473 16418 73483
rect 16428 73473 16486 73483
rect 16496 73473 16554 73483
rect 16564 73473 16622 73483
rect 16632 73473 16690 73483
rect 17290 73473 17348 73483
rect 17358 73473 17416 73483
rect 17426 73473 17484 73483
rect 17494 73473 17552 73483
rect 17562 73473 17620 73483
rect 17630 73473 17688 73483
rect 17698 73473 17756 73483
rect 17766 73473 17824 73483
rect 17834 73473 17892 73483
rect 17902 73473 17960 73483
rect 17970 73473 18028 73483
rect 18038 73473 18096 73483
rect 18106 73473 18164 73483
rect 18174 73473 18232 73483
rect 15724 73449 16690 73473
rect 17266 73449 18232 73473
rect 12427 73424 12493 73440
rect 15748 73434 15772 73449
rect 15816 73434 15840 73449
rect 15884 73434 15908 73449
rect 15952 73434 15976 73449
rect 16020 73434 16044 73449
rect 16088 73434 16112 73449
rect 16156 73434 16180 73449
rect 16224 73434 16248 73449
rect 16292 73434 16316 73449
rect 16360 73434 16384 73449
rect 16428 73434 16452 73449
rect 16496 73434 16520 73449
rect 16564 73434 16588 73449
rect 16632 73434 16656 73449
rect 17290 73434 17314 73449
rect 17358 73434 17382 73449
rect 17426 73434 17450 73449
rect 17494 73434 17518 73449
rect 17562 73434 17586 73449
rect 17630 73434 17654 73449
rect 17698 73434 17722 73449
rect 17766 73434 17790 73449
rect 17834 73434 17858 73449
rect 17902 73434 17926 73449
rect 17970 73434 17994 73449
rect 18038 73434 18062 73449
rect 18106 73434 18130 73449
rect 18174 73434 18198 73449
rect 15678 73279 16678 73434
rect 7389 73189 8389 73249
rect 8990 73189 9990 73249
rect 15678 73245 16690 73279
rect 17278 73269 18278 73434
rect 17266 73245 18278 73269
rect 15678 73234 16678 73245
rect 17278 73234 18278 73245
rect 15748 73221 15772 73234
rect 15816 73221 15840 73234
rect 15884 73221 15908 73234
rect 15952 73221 15976 73234
rect 16020 73221 16044 73234
rect 16088 73221 16112 73234
rect 16156 73221 16180 73234
rect 16224 73221 16248 73234
rect 16292 73221 16316 73234
rect 16360 73221 16384 73234
rect 16428 73221 16452 73234
rect 16496 73221 16520 73234
rect 16564 73221 16588 73234
rect 16632 73221 16656 73234
rect 17290 73221 17314 73234
rect 17358 73221 17382 73234
rect 17426 73221 17450 73234
rect 17494 73221 17518 73234
rect 17562 73221 17586 73234
rect 17630 73221 17654 73234
rect 17698 73221 17722 73234
rect 17766 73221 17790 73234
rect 17834 73221 17858 73234
rect 17902 73221 17926 73234
rect 17970 73221 17994 73234
rect 18038 73221 18062 73234
rect 18106 73221 18130 73234
rect 18174 73221 18198 73234
rect 7389 72831 8389 72887
rect 8990 72831 9990 72887
rect 15678 72876 16678 72932
rect 17278 72876 18278 72932
rect 7389 72759 8389 72815
rect 8990 72759 9990 72815
rect 15678 72804 16678 72860
rect 17278 72804 18278 72860
rect 7389 72457 8389 72529
rect 8990 72457 9990 72529
rect 15678 72502 16678 72574
rect 17278 72502 18278 72574
rect 15748 72491 15782 72502
rect 15816 72491 15850 72502
rect 15884 72491 15918 72502
rect 15952 72491 15986 72502
rect 16020 72491 16054 72502
rect 16088 72491 16122 72502
rect 16156 72491 16190 72502
rect 16224 72491 16258 72502
rect 16292 72491 16326 72502
rect 16360 72491 16394 72502
rect 16428 72491 16462 72502
rect 16496 72491 16530 72502
rect 16564 72491 16598 72502
rect 16632 72491 16666 72502
rect 17290 72491 17324 72502
rect 17358 72491 17392 72502
rect 17426 72491 17460 72502
rect 17494 72491 17528 72502
rect 17562 72491 17596 72502
rect 17630 72491 17664 72502
rect 17698 72491 17732 72502
rect 17766 72491 17800 72502
rect 17834 72491 17868 72502
rect 17902 72491 17936 72502
rect 17970 72491 18004 72502
rect 18038 72491 18072 72502
rect 18106 72491 18140 72502
rect 18174 72491 18208 72502
rect 15748 72481 15806 72491
rect 15816 72481 15874 72491
rect 15884 72481 15942 72491
rect 15952 72481 16010 72491
rect 16020 72481 16078 72491
rect 16088 72481 16146 72491
rect 16156 72481 16214 72491
rect 16224 72481 16282 72491
rect 16292 72481 16350 72491
rect 16360 72481 16418 72491
rect 16428 72481 16486 72491
rect 16496 72481 16554 72491
rect 16564 72481 16622 72491
rect 16632 72481 16690 72491
rect 17290 72481 17348 72491
rect 17358 72481 17416 72491
rect 17426 72481 17484 72491
rect 17494 72481 17552 72491
rect 17562 72481 17620 72491
rect 17630 72481 17688 72491
rect 17698 72481 17756 72491
rect 17766 72481 17824 72491
rect 17834 72481 17892 72491
rect 17902 72481 17960 72491
rect 17970 72481 18028 72491
rect 18038 72481 18096 72491
rect 18106 72481 18164 72491
rect 18174 72481 18232 72491
rect 15724 72457 16690 72481
rect 17266 72457 18232 72481
rect 15748 72442 15772 72457
rect 15816 72442 15840 72457
rect 15884 72442 15908 72457
rect 15952 72442 15976 72457
rect 16020 72442 16044 72457
rect 16088 72442 16112 72457
rect 16156 72442 16180 72457
rect 16224 72442 16248 72457
rect 16292 72442 16316 72457
rect 16360 72442 16384 72457
rect 16428 72442 16452 72457
rect 16496 72442 16520 72457
rect 16564 72442 16588 72457
rect 16632 72442 16656 72457
rect 17290 72442 17314 72457
rect 17358 72442 17382 72457
rect 17426 72442 17450 72457
rect 17494 72442 17518 72457
rect 17562 72442 17586 72457
rect 17630 72442 17654 72457
rect 17698 72442 17722 72457
rect 17766 72442 17790 72457
rect 17834 72442 17858 72457
rect 17902 72442 17926 72457
rect 17970 72442 17994 72457
rect 18038 72442 18062 72457
rect 18106 72442 18130 72457
rect 18174 72442 18198 72457
rect 15678 72287 16678 72442
rect 7389 72197 8389 72257
rect 8990 72197 9990 72257
rect 15678 72253 16690 72287
rect 17278 72277 18278 72442
rect 17266 72253 18278 72277
rect 15678 72242 16678 72253
rect 17278 72242 18278 72253
rect 15748 72229 15772 72242
rect 15816 72229 15840 72242
rect 15884 72229 15908 72242
rect 15952 72229 15976 72242
rect 16020 72229 16044 72242
rect 16088 72229 16112 72242
rect 16156 72229 16180 72242
rect 16224 72229 16248 72242
rect 16292 72229 16316 72242
rect 16360 72229 16384 72242
rect 16428 72229 16452 72242
rect 16496 72229 16520 72242
rect 16564 72229 16588 72242
rect 16632 72229 16656 72242
rect 17290 72229 17314 72242
rect 17358 72229 17382 72242
rect 17426 72229 17450 72242
rect 17494 72229 17518 72242
rect 17562 72229 17586 72242
rect 17630 72229 17654 72242
rect 17698 72229 17722 72242
rect 17766 72229 17790 72242
rect 17834 72229 17858 72242
rect 17902 72229 17926 72242
rect 17970 72229 17994 72242
rect 18038 72229 18062 72242
rect 18106 72229 18130 72242
rect 18174 72229 18198 72242
rect 7389 71839 8389 71895
rect 8990 71839 9990 71895
rect 15678 71884 16678 71940
rect 17278 71884 18278 71940
rect 7389 71767 8389 71823
rect 8990 71767 9990 71823
rect 15678 71812 16678 71868
rect 17278 71812 18278 71868
rect 7389 71465 8389 71537
rect 8990 71465 9990 71537
rect 15678 71510 16678 71582
rect 17278 71510 18278 71582
rect 15748 71499 15782 71510
rect 15816 71499 15850 71510
rect 15884 71499 15918 71510
rect 15952 71499 15986 71510
rect 16020 71499 16054 71510
rect 16088 71499 16122 71510
rect 16156 71499 16190 71510
rect 16224 71499 16258 71510
rect 16292 71499 16326 71510
rect 16360 71499 16394 71510
rect 16428 71499 16462 71510
rect 16496 71499 16530 71510
rect 16564 71499 16598 71510
rect 16632 71499 16666 71510
rect 17290 71499 17324 71510
rect 17358 71499 17392 71510
rect 17426 71499 17460 71510
rect 17494 71499 17528 71510
rect 17562 71499 17596 71510
rect 17630 71499 17664 71510
rect 17698 71499 17732 71510
rect 17766 71499 17800 71510
rect 17834 71499 17868 71510
rect 17902 71499 17936 71510
rect 17970 71499 18004 71510
rect 18038 71499 18072 71510
rect 18106 71499 18140 71510
rect 18174 71499 18208 71510
rect 15748 71489 15806 71499
rect 15816 71489 15874 71499
rect 15884 71489 15942 71499
rect 15952 71489 16010 71499
rect 16020 71489 16078 71499
rect 16088 71489 16146 71499
rect 16156 71489 16214 71499
rect 16224 71489 16282 71499
rect 16292 71489 16350 71499
rect 16360 71489 16418 71499
rect 16428 71489 16486 71499
rect 16496 71489 16554 71499
rect 16564 71489 16622 71499
rect 16632 71489 16690 71499
rect 17290 71489 17348 71499
rect 17358 71489 17416 71499
rect 17426 71489 17484 71499
rect 17494 71489 17552 71499
rect 17562 71489 17620 71499
rect 17630 71489 17688 71499
rect 17698 71489 17756 71499
rect 17766 71489 17824 71499
rect 17834 71489 17892 71499
rect 17902 71489 17960 71499
rect 17970 71489 18028 71499
rect 18038 71489 18096 71499
rect 18106 71489 18164 71499
rect 18174 71489 18232 71499
rect 15724 71465 16690 71489
rect 17266 71465 18232 71489
rect 15748 71450 15772 71465
rect 15816 71450 15840 71465
rect 15884 71450 15908 71465
rect 15952 71450 15976 71465
rect 16020 71450 16044 71465
rect 16088 71450 16112 71465
rect 16156 71450 16180 71465
rect 16224 71450 16248 71465
rect 16292 71450 16316 71465
rect 16360 71450 16384 71465
rect 16428 71450 16452 71465
rect 16496 71450 16520 71465
rect 16564 71450 16588 71465
rect 16632 71450 16656 71465
rect 17290 71450 17314 71465
rect 17358 71450 17382 71465
rect 17426 71450 17450 71465
rect 17494 71450 17518 71465
rect 17562 71450 17586 71465
rect 17630 71450 17654 71465
rect 17698 71450 17722 71465
rect 17766 71450 17790 71465
rect 17834 71450 17858 71465
rect 17902 71450 17926 71465
rect 17970 71450 17994 71465
rect 18038 71450 18062 71465
rect 18106 71450 18130 71465
rect 18174 71450 18198 71465
rect 15678 71295 16678 71450
rect 7389 71205 8389 71265
rect 8990 71205 9990 71265
rect 15678 71261 16690 71295
rect 17278 71285 18278 71450
rect 17266 71261 18278 71285
rect 15678 71250 16678 71261
rect 17278 71250 18278 71261
rect 15748 71237 15772 71250
rect 15816 71237 15840 71250
rect 15884 71237 15908 71250
rect 15952 71237 15976 71250
rect 16020 71237 16044 71250
rect 16088 71237 16112 71250
rect 16156 71237 16180 71250
rect 16224 71237 16248 71250
rect 16292 71237 16316 71250
rect 16360 71237 16384 71250
rect 16428 71237 16452 71250
rect 16496 71237 16520 71250
rect 16564 71237 16588 71250
rect 16632 71237 16656 71250
rect 17290 71237 17314 71250
rect 17358 71237 17382 71250
rect 17426 71237 17450 71250
rect 17494 71237 17518 71250
rect 17562 71237 17586 71250
rect 17630 71237 17654 71250
rect 17698 71237 17722 71250
rect 17766 71237 17790 71250
rect 17834 71237 17858 71250
rect 17902 71237 17926 71250
rect 17970 71237 17994 71250
rect 18038 71237 18062 71250
rect 18106 71237 18130 71250
rect 18174 71237 18198 71250
rect 7389 70847 8389 70903
rect 8990 70847 9990 70903
rect 15678 70892 16678 70948
rect 17278 70892 18278 70948
rect 7389 70775 8389 70831
rect 8990 70775 9990 70831
rect 15678 70820 16678 70876
rect 17278 70820 18278 70876
rect 5967 70455 6059 70489
rect 7389 70473 8389 70545
rect 8990 70473 9990 70545
rect 15678 70518 16678 70590
rect 17278 70518 18278 70590
rect 15748 70507 15782 70518
rect 15816 70507 15850 70518
rect 15884 70507 15918 70518
rect 15952 70507 15986 70518
rect 16020 70507 16054 70518
rect 16088 70507 16122 70518
rect 16156 70507 16190 70518
rect 16224 70507 16258 70518
rect 16292 70507 16326 70518
rect 16360 70507 16394 70518
rect 16428 70507 16462 70518
rect 16496 70507 16530 70518
rect 16564 70507 16598 70518
rect 16632 70507 16666 70518
rect 17290 70507 17324 70518
rect 17358 70507 17392 70518
rect 17426 70507 17460 70518
rect 17494 70507 17528 70518
rect 17562 70507 17596 70518
rect 17630 70507 17664 70518
rect 17698 70507 17732 70518
rect 17766 70507 17800 70518
rect 17834 70507 17868 70518
rect 17902 70507 17936 70518
rect 17970 70507 18004 70518
rect 18038 70507 18072 70518
rect 18106 70507 18140 70518
rect 18174 70507 18208 70518
rect 15748 70497 15806 70507
rect 15816 70497 15874 70507
rect 15884 70497 15942 70507
rect 15952 70497 16010 70507
rect 16020 70497 16078 70507
rect 16088 70497 16146 70507
rect 16156 70497 16214 70507
rect 16224 70497 16282 70507
rect 16292 70497 16350 70507
rect 16360 70497 16418 70507
rect 16428 70497 16486 70507
rect 16496 70497 16554 70507
rect 16564 70497 16622 70507
rect 16632 70497 16690 70507
rect 17290 70497 17348 70507
rect 17358 70497 17416 70507
rect 17426 70497 17484 70507
rect 17494 70497 17552 70507
rect 17562 70497 17620 70507
rect 17630 70497 17688 70507
rect 17698 70497 17756 70507
rect 17766 70497 17824 70507
rect 17834 70497 17892 70507
rect 17902 70497 17960 70507
rect 17970 70497 18028 70507
rect 18038 70497 18096 70507
rect 18106 70497 18164 70507
rect 18174 70497 18232 70507
rect 15724 70473 16690 70497
rect 17266 70473 18232 70497
rect 15748 70458 15772 70473
rect 15816 70458 15840 70473
rect 15884 70458 15908 70473
rect 15952 70458 15976 70473
rect 16020 70458 16044 70473
rect 16088 70458 16112 70473
rect 16156 70458 16180 70473
rect 16224 70458 16248 70473
rect 16292 70458 16316 70473
rect 16360 70458 16384 70473
rect 16428 70458 16452 70473
rect 16496 70458 16520 70473
rect 16564 70458 16588 70473
rect 16632 70458 16656 70473
rect 17290 70458 17314 70473
rect 17358 70458 17382 70473
rect 17426 70458 17450 70473
rect 17494 70458 17518 70473
rect 17562 70458 17586 70473
rect 17630 70458 17654 70473
rect 17698 70458 17722 70473
rect 17766 70458 17790 70473
rect 17834 70458 17858 70473
rect 17902 70458 17926 70473
rect 17970 70458 17994 70473
rect 18038 70458 18062 70473
rect 18106 70458 18130 70473
rect 18174 70458 18198 70473
rect 2850 70398 3850 70448
rect 2850 70282 3850 70332
rect 2850 70072 3850 70122
rect 2850 69956 3850 70006
rect 2850 69746 3850 69796
rect 1153 69660 1187 69718
rect 2850 69630 3850 69680
rect 2850 69420 3850 69470
rect 2850 69417 3107 69420
rect 3250 69304 3850 69354
rect 3250 69048 3850 69104
rect 3250 68892 3850 69020
rect 175 68818 1175 68868
rect 175 68662 1175 68790
rect 3250 68736 3850 68792
rect 175 68506 1175 68634
rect 175 68350 1175 68478
rect 175 68194 1175 68322
rect 175 68044 1175 68094
rect 175 67928 1175 67978
rect 175 67772 1175 67828
rect 175 67622 1175 67672
rect 1578 67609 1628 68609
rect 1728 67609 1856 68609
rect 1884 67609 2012 68609
rect 2040 67609 2090 68609
rect 3250 68580 3850 68708
rect 3250 68430 3850 68480
rect 2850 68314 3850 68364
rect 2850 68158 3850 68214
rect 2850 68008 3850 68058
rect 2850 67880 3850 67930
rect 2850 67724 3850 67852
rect 2850 67568 3850 67696
rect 175 67506 1175 67556
rect 175 67350 1175 67478
rect 2850 67412 3850 67468
rect 2850 67256 3850 67384
rect 175 67194 1175 67250
rect 175 67038 1175 67166
rect 175 66888 1175 66938
rect 175 66772 1175 66822
rect 175 66616 1175 66744
rect 1578 66613 1628 67213
rect 1728 66613 1784 67213
rect 1884 66613 1940 67213
rect 2040 66613 2096 67213
rect 2196 66613 2246 67213
rect 2850 67100 3850 67228
rect 2850 66944 3850 67072
rect 2850 66794 3850 66844
rect 2850 66678 3850 66728
rect 2850 66522 3850 66650
rect 175 66460 1175 66516
rect 175 66304 1175 66432
rect 2850 66366 3850 66494
rect 2850 66210 3850 66338
rect 175 66154 1175 66204
rect 803 66151 1175 66154
rect 2850 66054 3850 66110
rect 2850 65898 3850 66026
rect 2850 65742 3850 65870
rect 2850 65586 3850 65642
rect 2850 65436 3850 65486
rect 3926 65455 3960 65491
rect 3967 65339 3989 65455
rect 1638 63869 1688 64869
rect 1848 63869 1976 64869
rect 2064 63869 2114 64869
rect 2850 64275 3050 64287
rect 2850 64162 3850 64212
rect 2850 63946 3850 64074
rect 2850 63730 3850 63786
rect 2850 63514 3850 63642
rect 2850 63304 3850 63354
rect 2850 63188 3850 63238
rect 2850 62978 3850 63028
rect 3926 63015 3960 65339
rect 5169 63315 5191 70429
rect 5488 69194 5538 70194
rect 5658 69194 5708 70194
rect 5488 68073 5538 69073
rect 5658 68073 5708 69073
rect 5488 66952 5538 67952
rect 5658 66952 5708 67952
rect 5488 65842 5538 66842
rect 5658 65842 5708 66842
rect 5488 64721 5538 65721
rect 5658 64721 5708 65721
rect 5488 63600 5538 64600
rect 5658 63600 5708 64600
rect 5971 63386 6059 70455
rect 15678 70303 16678 70458
rect 7389 70213 8389 70273
rect 8990 70213 9990 70273
rect 15678 70269 16690 70303
rect 17278 70293 18278 70458
rect 17266 70269 18278 70293
rect 15678 70258 16678 70269
rect 17278 70258 18278 70269
rect 15748 70245 15772 70258
rect 15816 70245 15840 70258
rect 15884 70245 15908 70258
rect 15952 70245 15976 70258
rect 16020 70245 16044 70258
rect 16088 70245 16112 70258
rect 16156 70245 16180 70258
rect 16224 70245 16248 70258
rect 16292 70245 16316 70258
rect 16360 70245 16384 70258
rect 16428 70245 16452 70258
rect 16496 70245 16520 70258
rect 16564 70245 16588 70258
rect 16632 70245 16656 70258
rect 17290 70245 17314 70258
rect 17358 70245 17382 70258
rect 17426 70245 17450 70258
rect 17494 70245 17518 70258
rect 17562 70245 17586 70258
rect 17630 70245 17654 70258
rect 17698 70245 17722 70258
rect 17766 70245 17790 70258
rect 17834 70245 17858 70258
rect 17902 70245 17926 70258
rect 17970 70245 17994 70258
rect 18038 70245 18062 70258
rect 18106 70245 18130 70258
rect 18174 70245 18198 70258
rect 7389 69855 8389 69911
rect 8990 69855 9990 69911
rect 15678 69900 16678 69956
rect 17278 69900 18278 69956
rect 7389 69783 8389 69839
rect 8990 69783 9990 69839
rect 15678 69828 16678 69884
rect 17278 69828 18278 69884
rect 7389 69481 8389 69553
rect 8990 69481 9990 69553
rect 15678 69526 16678 69598
rect 17278 69526 18278 69598
rect 15748 69515 15782 69526
rect 15816 69515 15850 69526
rect 15884 69515 15918 69526
rect 15952 69515 15986 69526
rect 16020 69515 16054 69526
rect 16088 69515 16122 69526
rect 16156 69515 16190 69526
rect 16224 69515 16258 69526
rect 16292 69515 16326 69526
rect 16360 69515 16394 69526
rect 16428 69515 16462 69526
rect 16496 69515 16530 69526
rect 16564 69515 16598 69526
rect 16632 69515 16666 69526
rect 17290 69515 17324 69526
rect 17358 69515 17392 69526
rect 17426 69515 17460 69526
rect 17494 69515 17528 69526
rect 17562 69515 17596 69526
rect 17630 69515 17664 69526
rect 17698 69515 17732 69526
rect 17766 69515 17800 69526
rect 17834 69515 17868 69526
rect 17902 69515 17936 69526
rect 17970 69515 18004 69526
rect 18038 69515 18072 69526
rect 18106 69515 18140 69526
rect 18174 69515 18208 69526
rect 15748 69505 15806 69515
rect 15816 69505 15874 69515
rect 15884 69505 15942 69515
rect 15952 69505 16010 69515
rect 16020 69505 16078 69515
rect 16088 69505 16146 69515
rect 16156 69505 16214 69515
rect 16224 69505 16282 69515
rect 16292 69505 16350 69515
rect 16360 69505 16418 69515
rect 16428 69505 16486 69515
rect 16496 69505 16554 69515
rect 16564 69505 16622 69515
rect 16632 69505 16690 69515
rect 17290 69505 17348 69515
rect 17358 69505 17416 69515
rect 17426 69505 17484 69515
rect 17494 69505 17552 69515
rect 17562 69505 17620 69515
rect 17630 69505 17688 69515
rect 17698 69505 17756 69515
rect 17766 69505 17824 69515
rect 17834 69505 17892 69515
rect 17902 69505 17960 69515
rect 17970 69505 18028 69515
rect 18038 69505 18096 69515
rect 18106 69505 18164 69515
rect 18174 69505 18232 69515
rect 15724 69481 16690 69505
rect 17266 69481 18232 69505
rect 15748 69466 15772 69481
rect 15816 69466 15840 69481
rect 15884 69466 15908 69481
rect 15952 69466 15976 69481
rect 16020 69466 16044 69481
rect 16088 69466 16112 69481
rect 16156 69466 16180 69481
rect 16224 69466 16248 69481
rect 16292 69466 16316 69481
rect 16360 69466 16384 69481
rect 16428 69466 16452 69481
rect 16496 69466 16520 69481
rect 16564 69466 16588 69481
rect 16632 69466 16656 69481
rect 17290 69466 17314 69481
rect 17358 69466 17382 69481
rect 17426 69466 17450 69481
rect 17494 69466 17518 69481
rect 17562 69466 17586 69481
rect 17630 69466 17654 69481
rect 17698 69466 17722 69481
rect 17766 69466 17790 69481
rect 17834 69466 17858 69481
rect 17902 69466 17926 69481
rect 17970 69466 17994 69481
rect 18038 69466 18062 69481
rect 18106 69466 18130 69481
rect 18174 69466 18198 69481
rect 15678 69311 16678 69466
rect 7389 69221 8389 69281
rect 8990 69221 9990 69281
rect 15678 69277 16690 69311
rect 17278 69301 18278 69466
rect 17266 69277 18278 69301
rect 15678 69266 16678 69277
rect 17278 69266 18278 69277
rect 15748 69253 15772 69266
rect 15816 69253 15840 69266
rect 15884 69253 15908 69266
rect 15952 69253 15976 69266
rect 16020 69253 16044 69266
rect 16088 69253 16112 69266
rect 16156 69253 16180 69266
rect 16224 69253 16248 69266
rect 16292 69253 16316 69266
rect 16360 69253 16384 69266
rect 16428 69253 16452 69266
rect 16496 69253 16520 69266
rect 16564 69253 16588 69266
rect 16632 69253 16656 69266
rect 17290 69253 17314 69266
rect 17358 69253 17382 69266
rect 17426 69253 17450 69266
rect 17494 69253 17518 69266
rect 17562 69253 17586 69266
rect 17630 69253 17654 69266
rect 17698 69253 17722 69266
rect 17766 69253 17790 69266
rect 17834 69253 17858 69266
rect 17902 69253 17926 69266
rect 17970 69253 17994 69266
rect 18038 69253 18062 69266
rect 18106 69253 18130 69266
rect 18174 69253 18198 69266
rect 7389 68863 8389 68919
rect 8990 68863 9990 68919
rect 15678 68908 16678 68964
rect 17278 68908 18278 68964
rect 7389 68791 8389 68847
rect 8990 68791 9990 68847
rect 15678 68836 16678 68892
rect 17278 68836 18278 68892
rect 19480 68867 19516 75817
rect 19547 68867 19583 75817
rect 24572 75738 25172 75866
rect 36785 75864 37385 75920
rect 36785 75688 37385 75744
rect 20809 75650 20833 75684
rect 20809 75582 20833 75616
rect 24572 75588 25172 75638
rect 20809 75514 20833 75548
rect 36785 75518 37385 75568
rect 20809 75446 20833 75480
rect 24572 75458 25172 75508
rect 32930 75457 33530 75507
rect 20809 75378 20833 75412
rect 35287 75391 35887 75441
rect 36785 75402 37385 75452
rect 20809 75310 20833 75344
rect 24572 75308 25172 75358
rect 31463 75307 32063 75357
rect 32930 75301 33530 75357
rect 20809 75242 20833 75276
rect 35287 75215 35887 75343
rect 36785 75226 37385 75282
rect 20809 75174 20833 75208
rect 31463 75151 32063 75207
rect 32930 75151 33530 75201
rect 34079 75157 34679 75207
rect 20809 75106 20833 75140
rect 19844 74051 19894 75051
rect 19994 74051 20122 75051
rect 20150 74051 20278 75051
rect 20306 74051 20434 75051
rect 20462 74051 20512 75051
rect 20809 75038 20833 75072
rect 20809 74970 20833 75004
rect 20973 75000 21007 75024
rect 21041 75000 21075 75024
rect 21109 75000 21143 75024
rect 21177 75000 21211 75024
rect 21245 75000 21279 75024
rect 21313 75000 21347 75024
rect 21381 75000 21415 75024
rect 21449 75000 21483 75024
rect 21517 75000 21551 75024
rect 21585 75000 21619 75024
rect 21653 75000 21687 75024
rect 21721 75000 21755 75024
rect 21789 75000 21823 75024
rect 21857 75000 21891 75024
rect 21925 75000 21959 75024
rect 21993 75000 22027 75024
rect 22061 75000 22095 75024
rect 22129 75000 22163 75024
rect 22197 75000 22210 75024
rect 31463 75001 32063 75051
rect 34079 75001 34679 75057
rect 35287 75039 35887 75095
rect 36785 75050 37385 75106
rect 20809 74902 20833 74936
rect 32596 74929 33596 74979
rect 20809 74834 20833 74868
rect 24573 74820 25173 74870
rect 34079 74851 34679 74901
rect 35287 74869 35887 74919
rect 36785 74880 37385 74930
rect 35287 74866 35559 74869
rect 35716 74866 35887 74869
rect 20809 74766 20833 74800
rect 30171 74795 30771 74845
rect 20809 74698 20833 74732
rect 24573 74664 25173 74792
rect 32596 74773 33596 74829
rect 37993 74704 38593 74754
rect 19844 72521 19894 73921
rect 19994 72521 20122 73921
rect 20150 72521 20278 73921
rect 20306 72521 20434 73921
rect 20462 72521 20512 73921
rect 20809 72219 20833 72253
rect 19844 70759 19894 72159
rect 19994 70759 20122 72159
rect 20150 70759 20278 72159
rect 20306 70759 20434 72159
rect 20462 70759 20512 72159
rect 20809 72151 20833 72185
rect 20809 72083 20833 72117
rect 20809 72015 20833 72049
rect 20809 71947 20833 71981
rect 20809 71879 20833 71913
rect 20809 71811 20833 71845
rect 20809 71743 20833 71777
rect 20809 71675 20833 71709
rect 20809 71607 20833 71641
rect 20809 71539 20833 71573
rect 21263 71518 21313 74518
rect 21413 71518 21541 74518
rect 21569 71518 21697 74518
rect 21725 71518 21853 74518
rect 21881 71518 22009 74518
rect 22037 71518 22165 74518
rect 22193 71518 22321 74518
rect 22349 71518 22399 74518
rect 24573 74508 25173 74636
rect 30171 74619 30771 74675
rect 32596 74623 33596 74673
rect 34110 74589 34710 74639
rect 36785 74620 36797 74624
rect 36785 74609 36800 74620
rect 36970 74609 36985 74624
rect 26348 74530 26372 74564
rect 32596 74507 33596 74557
rect 26348 74461 26372 74495
rect 30171 74449 30771 74499
rect 24573 74352 25173 74408
rect 24573 74196 25173 74324
rect 29993 74310 30993 74360
rect 32596 74351 33596 74479
rect 34110 74433 34710 74561
rect 36785 74429 36985 74609
rect 37993 74534 38593 74584
rect 36785 74418 36800 74429
rect 36785 74414 36797 74418
rect 36970 74414 36985 74429
rect 31347 74317 31362 74332
rect 31535 74328 31547 74332
rect 31532 74317 31547 74328
rect 24573 74040 25173 74168
rect 26490 74122 26690 74172
rect 29993 74160 30993 74210
rect 31347 74137 31547 74317
rect 31347 74122 31362 74137
rect 31532 74126 31547 74137
rect 31535 74122 31547 74126
rect 31607 74317 31622 74332
rect 31795 74328 31807 74332
rect 31792 74317 31807 74328
rect 31607 74137 31807 74317
rect 32596 74195 33596 74323
rect 34110 74277 34710 74405
rect 36785 74384 36797 74388
rect 36785 74373 36800 74384
rect 36970 74373 36985 74388
rect 31607 74122 31622 74137
rect 31792 74126 31807 74137
rect 31795 74122 31807 74126
rect 31347 74081 31362 74096
rect 31535 74092 31547 74096
rect 31532 74081 31547 74092
rect 22906 73855 23212 74025
rect 23406 73855 23712 74025
rect 26490 73966 26690 74022
rect 29993 74001 30993 74051
rect 24573 73890 25173 73940
rect 31347 73901 31547 74081
rect 26490 73816 26690 73866
rect 29993 73851 30993 73901
rect 31347 73886 31362 73901
rect 31532 73890 31547 73901
rect 31535 73886 31547 73890
rect 31607 74081 31622 74096
rect 31795 74092 31807 74096
rect 31792 74081 31807 74092
rect 31607 73901 31807 74081
rect 32596 74039 33596 74167
rect 34110 74121 34710 74249
rect 36785 74193 36985 74373
rect 36785 74182 36800 74193
rect 36785 74178 36797 74182
rect 36970 74178 36985 74193
rect 37083 74373 37098 74388
rect 37083 74193 37120 74373
rect 37083 74178 37098 74193
rect 37998 74108 38598 74158
rect 34110 73971 34710 74021
rect 31607 73886 31622 73901
rect 31792 73890 31807 73901
rect 31795 73886 31807 73890
rect 32596 73883 33596 73939
rect 37998 73932 38598 73988
rect 34110 73855 34710 73905
rect 24573 73760 25173 73810
rect 27691 73682 28291 73732
rect 30253 73721 30268 73736
rect 30441 73732 30453 73736
rect 30438 73721 30453 73732
rect 24573 73610 25173 73660
rect 27691 73532 28291 73582
rect 30253 73541 30453 73721
rect 30253 73526 30268 73541
rect 30438 73530 30453 73541
rect 30441 73526 30453 73530
rect 30513 73721 30528 73736
rect 30701 73732 30713 73736
rect 30698 73721 30713 73732
rect 30513 73541 30713 73721
rect 30513 73526 30528 73541
rect 30698 73530 30713 73541
rect 30701 73526 30713 73530
rect 30773 73721 30788 73736
rect 30961 73732 30973 73736
rect 30958 73721 30973 73732
rect 30773 73541 30973 73721
rect 30773 73526 30788 73541
rect 30958 73530 30973 73541
rect 30961 73526 30973 73530
rect 31087 73721 31102 73736
rect 31275 73732 31287 73736
rect 31272 73721 31287 73732
rect 31087 73541 31287 73721
rect 31087 73526 31102 73541
rect 31272 73530 31287 73541
rect 31275 73526 31287 73530
rect 31347 73721 31362 73736
rect 31535 73732 31547 73736
rect 31532 73721 31547 73732
rect 31347 73541 31547 73721
rect 31347 73526 31362 73541
rect 31532 73530 31547 73541
rect 31535 73526 31547 73530
rect 31607 73721 31622 73736
rect 31795 73732 31807 73736
rect 31792 73721 31807 73732
rect 31607 73541 31807 73721
rect 31607 73526 31622 73541
rect 31792 73530 31807 73541
rect 31795 73526 31807 73530
rect 31867 73721 31882 73736
rect 32055 73732 32067 73736
rect 32052 73721 32067 73732
rect 32596 73727 33596 73855
rect 31867 73541 32067 73721
rect 34110 73699 34710 73827
rect 37998 73762 38598 73812
rect 37998 73759 38220 73762
rect 38245 73759 38539 73762
rect 32596 73571 33596 73699
rect 34110 73543 34710 73671
rect 31867 73526 31882 73541
rect 32052 73530 32067 73541
rect 32055 73526 32067 73530
rect 22619 73446 22647 73474
rect 24573 73438 25173 73488
rect 26490 73416 26690 73466
rect 27691 73402 28291 73452
rect 32596 73415 33596 73543
rect 34110 73387 34710 73515
rect 24573 73288 25173 73338
rect 26490 73260 26690 73316
rect 27691 73246 28291 73374
rect 30253 73361 30268 73376
rect 30441 73372 30453 73376
rect 30438 73361 30453 73372
rect 30253 73331 30453 73361
rect 30253 73316 30268 73331
rect 30438 73320 30453 73331
rect 30441 73316 30453 73320
rect 30513 73361 30528 73376
rect 30701 73372 30713 73376
rect 30698 73361 30713 73372
rect 30513 73331 30713 73361
rect 30513 73316 30528 73331
rect 30698 73320 30713 73331
rect 30701 73316 30713 73320
rect 30773 73361 30788 73376
rect 31347 73361 31362 73376
rect 31535 73372 31547 73376
rect 31532 73361 31547 73372
rect 30773 73331 30793 73361
rect 31347 73331 31547 73361
rect 30773 73316 30788 73331
rect 31347 73316 31362 73331
rect 31532 73320 31547 73331
rect 31535 73316 31547 73320
rect 31607 73361 31622 73376
rect 31795 73372 31807 73376
rect 31792 73361 31807 73372
rect 31607 73331 31807 73361
rect 31607 73316 31622 73331
rect 31792 73320 31807 73331
rect 31795 73316 31807 73320
rect 31867 73361 31882 73376
rect 31867 73331 31921 73361
rect 31867 73316 31882 73331
rect 30253 73275 30268 73290
rect 30441 73286 30453 73290
rect 30438 73275 30453 73286
rect 30253 73245 30453 73275
rect 30253 73230 30268 73245
rect 30438 73234 30453 73245
rect 30441 73230 30453 73234
rect 30513 73275 30528 73290
rect 30701 73286 30713 73290
rect 30698 73275 30713 73286
rect 30513 73245 30713 73275
rect 30513 73230 30528 73245
rect 30698 73234 30713 73245
rect 30701 73230 30713 73234
rect 30773 73275 30788 73290
rect 31347 73275 31362 73290
rect 31535 73286 31547 73290
rect 31532 73275 31547 73286
rect 30773 73245 30793 73275
rect 31347 73245 31547 73275
rect 30773 73230 30788 73245
rect 31347 73230 31362 73245
rect 31532 73234 31547 73245
rect 31535 73230 31547 73234
rect 31607 73275 31622 73290
rect 31795 73286 31807 73290
rect 31792 73275 31807 73286
rect 31607 73245 31807 73275
rect 31607 73230 31622 73245
rect 31792 73234 31807 73245
rect 31795 73230 31807 73234
rect 31867 73275 31882 73290
rect 31867 73245 31921 73275
rect 32596 73265 33596 73315
rect 31867 73230 31882 73245
rect 34110 73231 34710 73287
rect 22906 73055 23212 73225
rect 23406 73055 23712 73225
rect 24573 73158 25173 73208
rect 24573 73002 25173 73130
rect 26490 73107 26690 73160
rect 27691 73090 28291 73218
rect 31823 73084 32061 73118
rect 31481 73080 32061 73084
rect 31481 73068 31797 73080
rect 32596 73063 33596 73113
rect 34110 73075 34710 73203
rect 37998 73133 38148 73145
rect 38317 73133 38467 73145
rect 24573 72846 25173 72974
rect 27691 72934 28291 72990
rect 32596 72907 33596 73035
rect 34110 72919 34710 73047
rect 37998 73020 38598 73070
rect 27691 72778 28291 72906
rect 25286 72758 25310 72762
rect 32596 72751 33596 72879
rect 34110 72763 34710 72891
rect 37998 72844 38598 72900
rect 24573 72690 25173 72746
rect 25286 72687 25310 72721
rect 24573 72534 25173 72662
rect 25286 72615 25310 72649
rect 27691 72622 28291 72750
rect 32596 72595 33596 72723
rect 35287 72695 35487 72707
rect 37998 72674 38598 72724
rect 34110 72607 34710 72663
rect 36785 72650 36797 72654
rect 36785 72639 36800 72650
rect 36970 72639 36985 72654
rect 35134 72582 35734 72632
rect 25286 72543 25310 72577
rect 22906 72255 23212 72425
rect 23406 72255 23712 72425
rect 24573 72378 25173 72506
rect 25286 72471 25310 72505
rect 27691 72472 28291 72522
rect 32596 72439 33596 72567
rect 34110 72451 34710 72507
rect 35134 72432 35734 72482
rect 36785 72459 36985 72639
rect 36785 72448 36800 72459
rect 36785 72444 36797 72448
rect 36970 72444 36985 72459
rect 37083 72639 37098 72654
rect 37083 72459 37120 72639
rect 37083 72444 37098 72459
rect 36785 72414 36797 72418
rect 32596 72283 33596 72411
rect 36785 72403 36800 72414
rect 36970 72403 36985 72418
rect 34110 72295 34710 72351
rect 35134 72316 35734 72366
rect 24573 72228 25173 72278
rect 32596 72127 33596 72255
rect 34110 72145 34710 72195
rect 35134 72160 35734 72288
rect 32596 71971 33596 72099
rect 34110 72029 34710 72079
rect 35134 72004 35734 72132
rect 31481 71862 31797 71880
rect 34110 71873 34710 72001
rect 31823 71828 32061 71860
rect 32596 71821 33596 71871
rect 35134 71848 35734 71976
rect 36071 71805 36098 72295
rect 36785 72223 36985 72403
rect 37993 72248 38593 72298
rect 36785 72212 36800 72223
rect 36785 72208 36797 72212
rect 36970 72208 36985 72223
rect 696597 72200 696600 72320
rect 37993 72078 38593 72128
rect 692376 71983 692396 72017
rect 692463 71993 692532 72017
rect 696191 71993 696239 72017
rect 692487 71983 692532 71993
rect 696204 71983 696239 71993
rect 696340 71983 696360 72017
rect 36785 71902 37385 71952
rect 692487 71915 692502 71939
rect 696200 71915 696215 71939
rect 692454 71891 692478 71915
rect 696224 71891 696248 71915
rect 686755 71800 687355 71850
rect 34110 71717 34710 71773
rect 30253 71701 30268 71716
rect 30441 71712 30453 71716
rect 30438 71701 30453 71712
rect 30253 71671 30453 71701
rect 30253 71656 30268 71671
rect 30438 71660 30453 71671
rect 30441 71656 30453 71660
rect 30513 71701 30528 71716
rect 30701 71712 30713 71716
rect 30698 71701 30713 71712
rect 30513 71671 30713 71701
rect 30513 71656 30528 71671
rect 30698 71660 30713 71671
rect 30701 71656 30713 71660
rect 30773 71701 30788 71716
rect 31347 71701 31362 71716
rect 31535 71712 31547 71716
rect 31532 71701 31547 71712
rect 30773 71671 30793 71701
rect 31347 71671 31547 71701
rect 30773 71656 30788 71671
rect 31347 71656 31362 71671
rect 31532 71660 31547 71671
rect 31535 71656 31547 71660
rect 31607 71701 31622 71716
rect 31795 71712 31807 71716
rect 31792 71701 31807 71712
rect 31607 71671 31807 71701
rect 31607 71656 31622 71671
rect 31792 71660 31807 71671
rect 31795 71656 31807 71660
rect 31867 71701 31882 71716
rect 31867 71671 31921 71701
rect 35134 71698 35734 71770
rect 36785 71726 37385 71782
rect 692487 71748 692505 71752
rect 692479 71718 692505 71748
rect 692487 71698 692505 71718
rect 31867 71656 31882 71671
rect 30253 71615 30268 71630
rect 30441 71626 30453 71630
rect 30438 71615 30453 71626
rect 30253 71585 30453 71615
rect 30253 71570 30268 71585
rect 30438 71574 30453 71585
rect 30441 71570 30453 71574
rect 30513 71615 30528 71630
rect 30701 71626 30713 71630
rect 30698 71615 30713 71626
rect 30513 71585 30713 71615
rect 30513 71570 30528 71585
rect 30698 71574 30713 71585
rect 30701 71570 30713 71574
rect 30773 71615 30788 71630
rect 31347 71615 31362 71630
rect 31535 71626 31547 71630
rect 31532 71615 31547 71626
rect 30773 71585 30793 71615
rect 31347 71585 31547 71615
rect 30773 71570 30788 71585
rect 31347 71570 31362 71585
rect 31532 71574 31547 71585
rect 31535 71570 31547 71574
rect 31607 71615 31622 71630
rect 31795 71626 31807 71630
rect 31792 71615 31807 71626
rect 31607 71585 31807 71615
rect 31607 71570 31622 71585
rect 31792 71574 31807 71585
rect 31795 71570 31807 71574
rect 31867 71615 31882 71630
rect 32546 71619 33546 71669
rect 31867 71585 31921 71615
rect 31867 71570 31882 71585
rect 20809 71471 20833 71505
rect 32546 71463 33546 71591
rect 34110 71561 34710 71689
rect 35134 71645 36134 71695
rect 686755 71624 687355 71680
rect 692485 71674 692505 71698
rect 692509 71674 692517 71718
rect 696215 71698 696223 71748
rect 696203 71674 696223 71698
rect 696227 71674 696245 71752
rect 692485 71640 692521 71674
rect 696203 71640 696249 71674
rect 35134 71489 36134 71617
rect 36785 71550 37385 71606
rect 20809 71403 20833 71437
rect 30253 71405 30268 71420
rect 30441 71416 30453 71420
rect 30438 71405 30453 71416
rect 20809 71335 20833 71369
rect 20809 71267 20833 71301
rect 20809 71199 20833 71233
rect 30253 71225 30453 71405
rect 30253 71210 30268 71225
rect 30438 71214 30453 71225
rect 30441 71210 30453 71214
rect 30513 71405 30528 71420
rect 30701 71416 30713 71420
rect 30698 71405 30713 71416
rect 30513 71225 30713 71405
rect 30513 71210 30528 71225
rect 30698 71214 30713 71225
rect 30701 71210 30713 71214
rect 30773 71405 30788 71420
rect 30961 71416 30973 71420
rect 30958 71405 30973 71416
rect 30773 71225 30973 71405
rect 30773 71210 30788 71225
rect 30958 71214 30973 71225
rect 30961 71210 30973 71214
rect 31087 71405 31102 71420
rect 31275 71416 31287 71420
rect 31272 71405 31287 71416
rect 31087 71225 31287 71405
rect 31087 71210 31102 71225
rect 31272 71214 31287 71225
rect 31275 71210 31287 71214
rect 31347 71405 31362 71420
rect 31535 71416 31547 71420
rect 31532 71405 31547 71416
rect 31347 71225 31547 71405
rect 31347 71210 31362 71225
rect 31532 71214 31547 71225
rect 31535 71210 31547 71214
rect 31607 71405 31622 71420
rect 31795 71416 31807 71420
rect 31792 71405 31807 71416
rect 31607 71225 31807 71405
rect 31607 71210 31622 71225
rect 31792 71214 31807 71225
rect 31795 71210 31807 71214
rect 31867 71405 31882 71420
rect 32055 71416 32067 71420
rect 32052 71405 32067 71416
rect 31867 71225 32067 71405
rect 32546 71307 33546 71435
rect 34110 71411 34710 71461
rect 686755 71448 687355 71504
rect 35134 71339 36134 71389
rect 36785 71380 37385 71430
rect 31867 71210 31882 71225
rect 32052 71214 32067 71225
rect 32055 71210 32067 71214
rect 20809 71131 20833 71165
rect 32546 71151 33546 71279
rect 36785 71248 37385 71298
rect 686755 71278 687355 71328
rect 35285 71162 35319 71172
rect 35353 71162 35387 71172
rect 35421 71162 35455 71172
rect 35489 71162 35523 71172
rect 35564 71162 35598 71172
rect 35632 71162 35666 71172
rect 35700 71162 35734 71172
rect 35768 71162 35802 71172
rect 35836 71162 35870 71172
rect 35904 71162 35938 71172
rect 35972 71162 36006 71172
rect 36040 71162 36074 71172
rect 36108 71162 36142 71172
rect 36176 71162 36210 71172
rect 35255 71126 36255 71138
rect 20809 71063 20833 71097
rect 20940 71085 20983 71103
rect 20940 71069 20949 71085
rect 20974 71069 20983 71085
rect 25113 71069 25349 71093
rect 25383 71069 25417 71093
rect 20974 71051 21008 71069
rect 20809 70995 20833 71029
rect 20974 71028 21003 71051
rect 21361 71045 21409 71069
rect 20949 71027 20983 71028
rect 21385 70991 21409 71045
rect 25113 70991 25137 71069
rect 29993 71045 30993 71095
rect 31347 71045 31362 71060
rect 31535 71056 31547 71060
rect 31532 71045 31547 71056
rect 21361 70967 21409 70991
rect 25089 70967 25137 70991
rect 20809 70927 20833 70961
rect 20809 70859 20833 70893
rect 20809 70791 20833 70825
rect 20809 70723 20833 70757
rect 20809 70655 20833 70689
rect 21413 70638 22813 70681
rect 23685 70638 25085 70681
rect 19844 69229 19894 70629
rect 19994 69229 20122 70629
rect 20150 69229 20278 70629
rect 20306 69229 20434 70629
rect 20462 69229 20512 70629
rect 20809 70587 20833 70621
rect 20809 70519 20833 70553
rect 20809 70451 20833 70485
rect 21413 70475 22813 70603
rect 23685 70475 25085 70603
rect 20809 70383 20833 70417
rect 20809 70315 20833 70349
rect 21413 70312 22813 70440
rect 23685 70312 25085 70440
rect 20809 70247 20833 70281
rect 20809 70179 20833 70213
rect 21413 70149 22813 70277
rect 23685 70149 25085 70277
rect 20809 70111 20833 70145
rect 20809 70043 20833 70077
rect 20809 69975 20833 70009
rect 21413 69986 22813 70114
rect 23685 69986 25085 70114
rect 20809 69907 20833 69941
rect 20809 69839 20833 69873
rect 21413 69823 22813 69951
rect 23685 69823 25085 69951
rect 20809 69771 20833 69805
rect 20809 69703 20833 69737
rect 21413 69673 22813 69716
rect 23685 69673 25085 69716
rect 20809 69635 20833 69669
rect 20809 69567 20833 69601
rect 21361 69552 21419 69586
rect 25089 69552 25147 69586
rect 20809 69499 20833 69533
rect 20809 69431 20833 69465
rect 20809 69363 20833 69397
rect 21361 69373 21419 69397
rect 25089 69373 25147 69397
rect 21385 69363 21419 69373
rect 25113 69363 25147 69373
rect 20809 69295 20833 69329
rect 21385 69291 21419 69325
rect 25113 69291 25147 69325
rect 20809 69227 20833 69261
rect 21385 69219 21419 69253
rect 25113 69219 25147 69253
rect 20809 69159 20833 69193
rect 21385 69171 21419 69181
rect 25113 69171 25147 69181
rect 21361 69147 21419 69171
rect 25089 69147 25147 69171
rect 20809 69091 20833 69125
rect 20809 69023 20833 69057
rect 20809 68955 20833 68989
rect 21361 68969 21409 68993
rect 25089 68969 25137 68993
rect 20809 68887 20833 68921
rect 21385 68915 21409 68969
rect 25113 68915 25137 68969
rect 21361 68891 21409 68915
rect 25089 68891 25137 68915
rect 19480 68831 19583 68867
rect 21413 68754 22813 68804
rect 23685 68754 25085 68804
rect 7389 68489 8389 68561
rect 8990 68489 9990 68561
rect 15678 68534 16678 68606
rect 17278 68534 18278 68606
rect 21413 68591 22813 68719
rect 23685 68591 25085 68719
rect 15748 68523 15782 68534
rect 15816 68523 15850 68534
rect 15884 68523 15918 68534
rect 15952 68523 15986 68534
rect 16020 68523 16054 68534
rect 16088 68523 16122 68534
rect 16156 68523 16190 68534
rect 16224 68523 16258 68534
rect 16292 68523 16326 68534
rect 16360 68523 16394 68534
rect 16428 68523 16462 68534
rect 16496 68523 16530 68534
rect 16564 68523 16598 68534
rect 16632 68523 16666 68534
rect 17290 68523 17324 68534
rect 17358 68523 17392 68534
rect 17426 68523 17460 68534
rect 17494 68523 17528 68534
rect 17562 68523 17596 68534
rect 17630 68523 17664 68534
rect 17698 68523 17732 68534
rect 17766 68523 17800 68534
rect 17834 68523 17868 68534
rect 17902 68523 17936 68534
rect 17970 68523 18004 68534
rect 18038 68523 18072 68534
rect 18106 68523 18140 68534
rect 18174 68523 18208 68534
rect 15748 68513 15806 68523
rect 15816 68513 15874 68523
rect 15884 68513 15942 68523
rect 15952 68513 16010 68523
rect 16020 68513 16078 68523
rect 16088 68513 16146 68523
rect 16156 68513 16214 68523
rect 16224 68513 16282 68523
rect 16292 68513 16350 68523
rect 16360 68513 16418 68523
rect 16428 68513 16486 68523
rect 16496 68513 16554 68523
rect 16564 68513 16622 68523
rect 16632 68513 16690 68523
rect 17290 68513 17348 68523
rect 17358 68513 17416 68523
rect 17426 68513 17484 68523
rect 17494 68513 17552 68523
rect 17562 68513 17620 68523
rect 17630 68513 17688 68523
rect 17698 68513 17756 68523
rect 17766 68513 17824 68523
rect 17834 68513 17892 68523
rect 17902 68513 17960 68523
rect 17970 68513 18028 68523
rect 18038 68513 18096 68523
rect 18106 68513 18164 68523
rect 18174 68513 18232 68523
rect 15724 68489 16690 68513
rect 17266 68489 18232 68513
rect 15748 68474 15772 68489
rect 15816 68474 15840 68489
rect 15884 68474 15908 68489
rect 15952 68474 15976 68489
rect 16020 68474 16044 68489
rect 16088 68474 16112 68489
rect 16156 68474 16180 68489
rect 16224 68474 16248 68489
rect 16292 68474 16316 68489
rect 16360 68474 16384 68489
rect 16428 68474 16452 68489
rect 16496 68474 16520 68489
rect 16564 68474 16588 68489
rect 16632 68474 16656 68489
rect 17290 68474 17314 68489
rect 17358 68474 17382 68489
rect 17426 68474 17450 68489
rect 17494 68474 17518 68489
rect 17562 68474 17586 68489
rect 17630 68474 17654 68489
rect 17698 68474 17722 68489
rect 17766 68474 17790 68489
rect 17834 68474 17858 68489
rect 17902 68474 17926 68489
rect 17970 68474 17994 68489
rect 18038 68474 18062 68489
rect 18106 68474 18130 68489
rect 18174 68474 18198 68489
rect 15678 68319 16678 68474
rect 7389 68229 8389 68289
rect 8990 68229 9990 68289
rect 15678 68285 16690 68319
rect 17278 68309 18278 68474
rect 21413 68428 22813 68556
rect 23685 68428 25085 68556
rect 17266 68285 18278 68309
rect 15678 68274 16678 68285
rect 17278 68274 18278 68285
rect 15748 68261 15772 68274
rect 15816 68261 15840 68274
rect 15884 68261 15908 68274
rect 15952 68261 15976 68274
rect 16020 68261 16044 68274
rect 16088 68261 16112 68274
rect 16156 68261 16180 68274
rect 16224 68261 16248 68274
rect 16292 68261 16316 68274
rect 16360 68261 16384 68274
rect 16428 68261 16452 68274
rect 16496 68261 16520 68274
rect 16564 68261 16588 68274
rect 16632 68261 16656 68274
rect 17290 68261 17314 68274
rect 17358 68261 17382 68274
rect 17426 68261 17450 68274
rect 17494 68261 17518 68274
rect 17562 68261 17586 68274
rect 17630 68261 17654 68274
rect 17698 68261 17722 68274
rect 17766 68261 17790 68274
rect 17834 68261 17858 68274
rect 17902 68261 17926 68274
rect 17970 68261 17994 68274
rect 18038 68261 18062 68274
rect 18106 68261 18130 68274
rect 18174 68261 18198 68274
rect 21413 68265 22813 68393
rect 23685 68265 25085 68393
rect 21413 68102 22813 68230
rect 23685 68102 25085 68230
rect 7389 67871 8389 67927
rect 8990 67871 9990 67927
rect 15678 67916 16678 67972
rect 17278 67916 18278 67972
rect 21413 67952 22813 67995
rect 23685 67952 25085 67995
rect 7389 67799 8389 67855
rect 8990 67799 9990 67855
rect 15678 67844 16678 67900
rect 17278 67844 18278 67900
rect 21406 67865 21430 67889
rect 25068 67865 25092 67889
rect 21382 67841 21385 67865
rect 25113 67841 25116 67865
rect 21382 67763 21396 67787
rect 25102 67763 25116 67787
rect 21348 67739 21372 67763
rect 21406 67739 21430 67763
rect 25068 67739 25092 67763
rect 25126 67739 25150 67763
rect 25524 67703 25548 71001
rect 29993 70895 30993 70945
rect 31347 70865 31547 71045
rect 31347 70850 31362 70865
rect 31532 70854 31547 70865
rect 31535 70850 31547 70854
rect 31607 71045 31622 71060
rect 31795 71056 31807 71060
rect 31792 71045 31807 71056
rect 31607 70865 31807 71045
rect 32546 70995 33546 71123
rect 36785 71072 37385 71128
rect 685547 71102 686147 71152
rect 35255 71019 36255 71069
rect 687155 71007 687170 71022
rect 687343 71018 687355 71022
rect 687340 71007 687355 71018
rect 31607 70850 31622 70865
rect 31792 70854 31807 70865
rect 31795 70850 31807 70854
rect 32546 70839 33546 70967
rect 35255 70843 36255 70971
rect 36785 70896 37385 70952
rect 685547 70932 686147 70982
rect 687155 70827 687355 71007
rect 31347 70809 31362 70824
rect 31535 70820 31547 70824
rect 31532 70809 31547 70820
rect 29993 70736 30993 70786
rect 29993 70586 30993 70636
rect 31347 70629 31547 70809
rect 31347 70614 31362 70629
rect 31532 70618 31547 70629
rect 31535 70614 31547 70618
rect 31607 70809 31622 70824
rect 31795 70820 31807 70824
rect 31792 70809 31807 70820
rect 687155 70812 687170 70827
rect 687340 70816 687355 70827
rect 687343 70812 687355 70816
rect 31607 70629 31807 70809
rect 32546 70683 33546 70811
rect 35255 70667 36255 70795
rect 36785 70726 37385 70776
rect 687042 70771 687057 70786
rect 31607 70614 31622 70629
rect 31792 70618 31807 70629
rect 31795 70614 31807 70618
rect 32546 70527 33546 70655
rect 37993 70550 38593 70600
rect 687020 70591 687057 70771
rect 687155 70771 687170 70786
rect 687343 70782 687355 70786
rect 687340 70771 687355 70782
rect 687155 70591 687355 70771
rect 688210 70630 688260 71630
rect 688360 70740 688488 71630
rect 688516 70740 688644 71630
rect 688672 70740 688800 71630
rect 688828 70740 688956 71630
rect 688984 70740 689112 71630
rect 689140 70740 689268 71630
rect 689296 70740 689424 71630
rect 689452 70740 689580 71630
rect 689608 70740 689736 71630
rect 689764 70740 689892 71630
rect 689920 70740 690048 71630
rect 690076 70740 690204 71630
rect 690232 70740 690360 71630
rect 690388 70630 690438 71630
rect 692485 71606 692505 71640
rect 692509 71606 692517 71640
rect 696203 71606 696223 71640
rect 696227 71606 696245 71640
rect 691275 71523 691875 71573
rect 692485 71572 692521 71606
rect 696203 71572 696249 71606
rect 692485 71538 692505 71572
rect 692509 71538 692517 71572
rect 692485 71504 692521 71538
rect 692583 71528 693983 71571
rect 694719 71528 696119 71571
rect 696203 71538 696223 71572
rect 696227 71538 696245 71572
rect 696203 71504 696249 71538
rect 692485 71470 692505 71504
rect 692509 71470 692517 71504
rect 692485 71436 692521 71470
rect 691275 71373 691875 71423
rect 692485 71402 692505 71436
rect 692509 71402 692517 71436
rect 692485 71368 692521 71402
rect 692485 71334 692505 71368
rect 692509 71334 692517 71368
rect 692583 71365 693983 71493
rect 694719 71365 696119 71493
rect 696203 71470 696223 71504
rect 696227 71470 696245 71504
rect 696203 71436 696249 71470
rect 707624 71441 707658 71475
rect 707695 71441 707729 71475
rect 707769 71441 707803 71475
rect 707840 71441 707874 71475
rect 707914 71441 707948 71475
rect 707985 71441 708019 71475
rect 708059 71441 708093 71475
rect 708130 71441 708164 71475
rect 708204 71441 708238 71475
rect 708275 71441 708309 71475
rect 708369 71441 708403 71475
rect 708446 71441 708480 71475
rect 708520 71441 708554 71465
rect 708588 71441 708610 71465
rect 709211 71441 709234 71465
rect 709270 71441 709304 71475
rect 709364 71441 709398 71475
rect 709435 71441 709469 71475
rect 709509 71441 709543 71475
rect 709580 71441 709614 71475
rect 709654 71441 709688 71475
rect 709725 71441 709759 71475
rect 709799 71441 709833 71475
rect 709870 71441 709904 71475
rect 709944 71441 709978 71475
rect 710015 71441 710049 71475
rect 710089 71441 710123 71475
rect 710160 71441 710194 71475
rect 696203 71402 696223 71436
rect 696227 71402 696245 71436
rect 707610 71431 707624 71441
rect 707658 71431 707695 71441
rect 707729 71431 707769 71441
rect 707803 71431 707840 71441
rect 707874 71431 707914 71441
rect 707948 71431 707985 71441
rect 708019 71431 708059 71441
rect 708093 71431 708130 71441
rect 708164 71431 708204 71441
rect 708238 71431 708275 71441
rect 708309 71431 708369 71441
rect 708403 71431 708446 71441
rect 708480 71431 708520 71441
rect 708554 71431 708588 71441
rect 708610 71431 708634 71441
rect 709211 71431 709270 71441
rect 709304 71431 709364 71441
rect 709398 71431 709435 71441
rect 709469 71431 709509 71441
rect 709543 71431 709580 71441
rect 709614 71431 709654 71441
rect 709688 71431 709725 71441
rect 709759 71431 709799 71441
rect 709833 71431 709870 71441
rect 709904 71431 709944 71441
rect 709978 71431 710015 71441
rect 710049 71431 710089 71441
rect 710123 71431 710160 71441
rect 710194 71431 710211 71441
rect 696203 71368 696249 71402
rect 696203 71334 696223 71368
rect 696227 71334 696245 71368
rect 707610 71337 708610 71431
rect 709211 71337 710211 71431
rect 691275 71251 691875 71301
rect 692485 71300 692521 71334
rect 692485 71266 692505 71300
rect 692509 71266 692517 71300
rect 692485 71232 692521 71266
rect 692485 71198 692505 71232
rect 692509 71198 692517 71232
rect 692583 71202 693983 71330
rect 694719 71202 696119 71330
rect 696203 71300 696249 71334
rect 711579 71317 712463 71331
rect 711579 71307 711619 71317
rect 696203 71266 696223 71300
rect 696227 71266 696245 71300
rect 701730 71290 701747 71292
rect 696203 71232 696249 71266
rect 696203 71198 696223 71232
rect 696227 71198 696245 71232
rect 701692 71220 701722 71254
rect 701730 71220 701760 71290
rect 707610 71241 708610 71301
rect 709211 71241 710211 71301
rect 692485 71164 692521 71198
rect 691275 71101 691875 71151
rect 692485 71130 692505 71164
rect 692509 71130 692517 71164
rect 692485 71096 692521 71130
rect 692485 71062 692505 71096
rect 692509 71062 692517 71096
rect 692485 71028 692521 71062
rect 692583 71039 693983 71167
rect 694719 71039 696119 71167
rect 696203 71164 696249 71198
rect 696203 71130 696223 71164
rect 696227 71130 696245 71164
rect 696203 71096 696249 71130
rect 696203 71062 696223 71096
rect 696227 71062 696245 71096
rect 699322 71064 700322 71097
rect 700922 71064 701922 71097
rect 696203 71028 696249 71062
rect 707610 71044 708610 71048
rect 709211 71044 710211 71048
rect 691275 70975 691875 71025
rect 692485 70994 692505 71028
rect 692509 70994 692517 71028
rect 692485 70960 692521 70994
rect 692485 70926 692505 70960
rect 692509 70926 692517 70960
rect 692485 70892 692521 70926
rect 691275 70825 691875 70875
rect 692485 70858 692505 70892
rect 692509 70858 692517 70892
rect 692583 70876 693983 71004
rect 694719 70876 696119 71004
rect 696203 70994 696223 71028
rect 696227 70994 696245 71028
rect 707574 70994 708646 71030
rect 696203 70960 696249 70994
rect 696203 70926 696223 70960
rect 696227 70926 696245 70960
rect 707574 70953 707610 70994
rect 708610 70953 708646 70994
rect 696203 70892 696249 70926
rect 697284 70894 697350 70910
rect 707574 70897 708646 70953
rect 696203 70858 696223 70892
rect 696227 70858 696245 70892
rect 699322 70877 700322 70894
rect 700922 70877 701922 70894
rect 707574 70881 707610 70897
rect 708610 70881 708646 70897
rect 692485 70824 692521 70858
rect 692485 70790 692505 70824
rect 692509 70790 692517 70824
rect 692485 70756 692521 70790
rect 691275 70703 691875 70753
rect 692485 70740 692505 70756
rect 692509 70740 692517 70756
rect 692583 70740 693983 70841
rect 694719 70740 696119 70841
rect 696203 70824 696249 70858
rect 707574 70825 708646 70881
rect 696203 70790 696223 70824
rect 696227 70790 696245 70824
rect 696203 70756 696249 70790
rect 696203 70740 696223 70756
rect 696227 70740 696245 70756
rect 699322 70740 700322 70811
rect 700922 70740 701922 70811
rect 707574 70788 707610 70825
rect 708610 70788 708646 70825
rect 707574 70748 708646 70788
rect 709175 70994 710247 71030
rect 709175 70953 709211 70994
rect 710211 70953 710247 70994
rect 709175 70897 710247 70953
rect 709175 70881 709211 70897
rect 710211 70881 710247 70897
rect 709175 70825 710247 70881
rect 709175 70788 709211 70825
rect 710211 70788 710247 70825
rect 709175 70748 710247 70788
rect 28647 70450 28671 70477
rect 30171 70447 30771 70497
rect 35255 70491 36255 70547
rect 685542 70506 686142 70556
rect 691275 70553 691875 70603
rect 36785 70466 36797 70470
rect 36785 70455 36800 70466
rect 36970 70455 36985 70470
rect 28683 70397 28717 70431
rect 32546 70377 33546 70427
rect 28683 70328 28717 70362
rect 28683 70259 28717 70293
rect 30171 70271 30771 70327
rect 35255 70321 36255 70371
rect 36785 70275 36985 70455
rect 37993 70380 38593 70430
rect 685542 70330 686142 70386
rect 36785 70264 36800 70275
rect 36785 70260 36797 70264
rect 36970 70260 36985 70275
rect 692583 70237 693983 70280
rect 694719 70237 696119 70280
rect 699322 70278 700322 70418
rect 700922 70278 701922 70418
rect 36785 70230 36797 70234
rect 28683 70190 28717 70224
rect 32596 70175 33596 70225
rect 35359 70156 35375 70222
rect 36143 70156 36159 70222
rect 36785 70219 36800 70230
rect 36970 70219 36985 70234
rect 28683 70121 28717 70155
rect 30171 70101 30771 70151
rect 28683 70052 28717 70086
rect 32596 70019 33596 70147
rect 28683 69983 28717 70017
rect 33959 69994 33975 70060
rect 36143 69994 36159 70060
rect 36785 70039 36985 70219
rect 36785 70028 36800 70039
rect 36785 70024 36797 70028
rect 36970 70024 36985 70039
rect 37083 70219 37098 70234
rect 37083 70039 37120 70219
rect 685542 70160 686142 70210
rect 692583 70101 693983 70144
rect 694719 70101 696119 70144
rect 37083 70024 37098 70039
rect 28683 69914 28717 69948
rect 31463 69895 32063 69945
rect 28683 69845 28717 69879
rect 32596 69863 33596 69991
rect 37998 69954 38598 70004
rect 28683 69776 28717 69810
rect 28683 69707 28717 69741
rect 31463 69739 32063 69795
rect 32596 69707 33596 69835
rect 33959 69832 33975 69898
rect 36143 69832 36159 69898
rect 37998 69778 38598 69834
rect 28683 69638 28717 69672
rect 28683 69569 28717 69603
rect 31463 69589 32063 69639
rect 32596 69551 33596 69679
rect 35359 69670 35375 69736
rect 36143 69670 36159 69736
rect 680215 69678 680815 69728
rect 37998 69608 38598 69658
rect 37998 69605 38220 69608
rect 38245 69605 38539 69608
rect 28683 69500 28717 69534
rect 28683 69431 28717 69465
rect 28683 69362 28717 69396
rect 32596 69395 33596 69523
rect 35255 69521 36255 69571
rect 680215 69502 680815 69558
rect 685551 69516 686551 69566
rect 689154 69480 689204 69897
rect 689304 69480 689360 69897
rect 689460 69480 689516 69897
rect 689616 69480 689672 69897
rect 689772 69480 689828 69897
rect 689928 69480 689978 69897
rect 699322 69860 700322 69916
rect 700922 69860 701922 69916
rect 707610 69905 708610 69961
rect 709211 69905 710211 69961
rect 699322 69788 700322 69844
rect 700922 69788 701922 69844
rect 707610 69833 708610 69889
rect 709211 69833 710211 69889
rect 711579 69525 711605 71307
rect 715956 70297 716006 71297
rect 716106 70740 716234 71297
rect 716262 70297 716312 71297
rect 711579 69480 711595 69495
rect 712409 69480 712431 69485
rect 713640 69480 713641 69785
rect 713750 69772 714750 69822
rect 713750 69562 714750 69612
rect 713750 69480 714750 69496
rect 28683 69293 28717 69327
rect 28683 69224 28717 69258
rect 30015 69256 30718 69272
rect 30015 69246 30721 69256
rect 28683 69155 28717 69189
rect 28683 69086 28717 69120
rect 28683 69017 28717 69051
rect 28683 68948 28717 68982
rect 28683 68879 28717 68913
rect 28683 68810 28717 68844
rect 28683 68741 28717 68775
rect 28683 68672 28717 68706
rect 28683 68603 28717 68637
rect 28683 68534 28717 68568
rect 28683 68465 28717 68499
rect 28683 68396 28717 68430
rect 28682 68361 28683 68366
rect 28682 68332 28717 68361
rect 28647 68303 28671 68332
rect 28647 68234 28671 68268
rect 28647 68165 28671 68199
rect 28647 68096 28671 68130
rect 28647 68027 28671 68061
rect 28647 67958 28671 67992
rect 28647 67889 28671 67923
rect 28647 67820 28671 67854
rect 28647 67751 28671 67785
rect 28647 67682 28671 67716
rect 29778 67695 29802 67719
rect 29802 67671 29826 67683
rect 29880 67681 29914 67715
rect 25524 67635 25548 67669
rect 7389 67497 8389 67569
rect 8990 67497 9990 67569
rect 15678 67542 16678 67614
rect 17278 67542 18278 67614
rect 28647 67613 28671 67647
rect 29778 67635 29802 67659
rect 21361 67586 21409 67610
rect 25089 67586 25137 67610
rect 15748 67531 15782 67542
rect 15816 67531 15850 67542
rect 15884 67531 15918 67542
rect 15952 67531 15986 67542
rect 16020 67531 16054 67542
rect 16088 67531 16122 67542
rect 16156 67531 16190 67542
rect 16224 67531 16258 67542
rect 16292 67531 16326 67542
rect 16360 67531 16394 67542
rect 16428 67531 16462 67542
rect 16496 67531 16530 67542
rect 16564 67531 16598 67542
rect 16632 67531 16666 67542
rect 17290 67531 17324 67542
rect 17358 67531 17392 67542
rect 17426 67531 17460 67542
rect 17494 67531 17528 67542
rect 17562 67531 17596 67542
rect 17630 67531 17664 67542
rect 17698 67531 17732 67542
rect 17766 67531 17800 67542
rect 17834 67531 17868 67542
rect 17902 67531 17936 67542
rect 17970 67531 18004 67542
rect 18038 67531 18072 67542
rect 18106 67531 18140 67542
rect 18174 67531 18208 67542
rect 21385 67532 21409 67586
rect 25113 67532 25137 67586
rect 28647 67544 28671 67578
rect 15748 67521 15806 67531
rect 15816 67521 15874 67531
rect 15884 67521 15942 67531
rect 15952 67521 16010 67531
rect 16020 67521 16078 67531
rect 16088 67521 16146 67531
rect 16156 67521 16214 67531
rect 16224 67521 16282 67531
rect 16292 67521 16350 67531
rect 16360 67521 16418 67531
rect 16428 67521 16486 67531
rect 16496 67521 16554 67531
rect 16564 67521 16622 67531
rect 16632 67521 16690 67531
rect 17290 67521 17348 67531
rect 17358 67521 17416 67531
rect 17426 67521 17484 67531
rect 17494 67521 17552 67531
rect 17562 67521 17620 67531
rect 17630 67521 17688 67531
rect 17698 67521 17756 67531
rect 17766 67521 17824 67531
rect 17834 67521 17892 67531
rect 17902 67521 17960 67531
rect 17970 67521 18028 67531
rect 18038 67521 18096 67531
rect 18106 67521 18164 67531
rect 18174 67521 18232 67531
rect 15724 67497 16690 67521
rect 17266 67497 18232 67521
rect 21361 67508 21409 67532
rect 25089 67508 25137 67532
rect 15748 67482 15772 67497
rect 15816 67482 15840 67497
rect 15884 67482 15908 67497
rect 15952 67482 15976 67497
rect 16020 67482 16044 67497
rect 16088 67482 16112 67497
rect 16156 67482 16180 67497
rect 16224 67482 16248 67497
rect 16292 67482 16316 67497
rect 16360 67482 16384 67497
rect 16428 67482 16452 67497
rect 16496 67482 16520 67497
rect 16564 67482 16588 67497
rect 16632 67482 16656 67497
rect 17290 67482 17314 67497
rect 17358 67482 17382 67497
rect 17426 67482 17450 67497
rect 17494 67482 17518 67497
rect 17562 67482 17586 67497
rect 17630 67482 17654 67497
rect 17698 67482 17722 67497
rect 17766 67482 17790 67497
rect 17834 67482 17858 67497
rect 17902 67482 17926 67497
rect 17970 67482 17994 67497
rect 18038 67482 18062 67497
rect 18106 67482 18130 67497
rect 18174 67482 18198 67497
rect 7389 67237 8389 67297
rect 8990 67237 9990 67297
rect 12559 67273 12865 67375
rect 15678 67327 16678 67482
rect 15678 67293 16690 67327
rect 17278 67317 18278 67482
rect 28647 67475 28671 67509
rect 28647 67406 28671 67440
rect 28647 67337 28671 67371
rect 17266 67293 18278 67317
rect 15678 67282 16678 67293
rect 17278 67282 18278 67293
rect 12543 67257 12881 67273
rect 15748 67269 15772 67282
rect 15816 67269 15840 67282
rect 15884 67269 15908 67282
rect 15952 67269 15976 67282
rect 16020 67269 16044 67282
rect 16088 67269 16112 67282
rect 16156 67269 16180 67282
rect 16224 67269 16248 67282
rect 16292 67269 16316 67282
rect 16360 67269 16384 67282
rect 16428 67269 16452 67282
rect 16496 67269 16520 67282
rect 16564 67269 16588 67282
rect 16632 67269 16656 67282
rect 17290 67269 17314 67282
rect 17358 67269 17382 67282
rect 17426 67269 17450 67282
rect 17494 67269 17518 67282
rect 17562 67269 17586 67282
rect 17630 67269 17654 67282
rect 17698 67269 17722 67282
rect 17766 67269 17790 67282
rect 17834 67269 17858 67282
rect 17902 67269 17926 67282
rect 17970 67269 17994 67282
rect 18038 67269 18062 67282
rect 18106 67269 18130 67282
rect 18174 67269 18198 67282
rect 19980 67048 20286 67218
rect 7389 66879 8389 66935
rect 8990 66879 9990 66935
rect 15678 66924 16678 66980
rect 17278 66924 18278 66980
rect 7389 66807 8389 66863
rect 8990 66807 9990 66863
rect 15678 66852 16678 66908
rect 17278 66852 18278 66908
rect 20945 66796 25553 67332
rect 28647 67268 28671 67302
rect 28647 67199 28671 67233
rect 28647 67154 28671 67164
rect 21413 66706 22813 66796
rect 23685 66706 25085 66796
rect 7389 66505 8389 66577
rect 8990 66505 9990 66577
rect 15678 66550 16678 66622
rect 17278 66550 18278 66622
rect 15748 66539 15782 66550
rect 15816 66539 15850 66550
rect 15884 66539 15918 66550
rect 15952 66539 15986 66550
rect 16020 66539 16054 66550
rect 16088 66539 16122 66550
rect 16156 66539 16190 66550
rect 16224 66539 16258 66550
rect 16292 66539 16326 66550
rect 16360 66539 16394 66550
rect 16428 66539 16462 66550
rect 16496 66539 16530 66550
rect 16564 66539 16598 66550
rect 16632 66539 16666 66550
rect 17290 66539 17324 66550
rect 17358 66539 17392 66550
rect 17426 66539 17460 66550
rect 17494 66539 17528 66550
rect 17562 66539 17596 66550
rect 17630 66539 17664 66550
rect 17698 66539 17732 66550
rect 17766 66539 17800 66550
rect 17834 66539 17868 66550
rect 17902 66539 17936 66550
rect 17970 66539 18004 66550
rect 18038 66539 18072 66550
rect 18106 66539 18140 66550
rect 18174 66539 18208 66550
rect 21413 66543 22813 66671
rect 23685 66543 25085 66671
rect 15748 66529 15806 66539
rect 15816 66529 15874 66539
rect 15884 66529 15942 66539
rect 15952 66529 16010 66539
rect 16020 66529 16078 66539
rect 16088 66529 16146 66539
rect 16156 66529 16214 66539
rect 16224 66529 16282 66539
rect 16292 66529 16350 66539
rect 16360 66529 16418 66539
rect 16428 66529 16486 66539
rect 16496 66529 16554 66539
rect 16564 66529 16622 66539
rect 16632 66529 16690 66539
rect 17290 66529 17348 66539
rect 17358 66529 17416 66539
rect 17426 66529 17484 66539
rect 17494 66529 17552 66539
rect 17562 66529 17620 66539
rect 17630 66529 17688 66539
rect 17698 66529 17756 66539
rect 17766 66529 17824 66539
rect 17834 66529 17892 66539
rect 17902 66529 17960 66539
rect 17970 66529 18028 66539
rect 18038 66529 18096 66539
rect 18106 66529 18164 66539
rect 18174 66529 18232 66539
rect 15724 66505 16690 66529
rect 17266 66505 18232 66529
rect 15748 66490 15772 66505
rect 15816 66490 15840 66505
rect 15884 66490 15908 66505
rect 15952 66490 15976 66505
rect 16020 66490 16044 66505
rect 16088 66490 16112 66505
rect 16156 66490 16180 66505
rect 16224 66490 16248 66505
rect 16292 66490 16316 66505
rect 16360 66490 16384 66505
rect 16428 66490 16452 66505
rect 16496 66490 16520 66505
rect 16564 66490 16588 66505
rect 16632 66490 16656 66505
rect 17290 66490 17314 66505
rect 17358 66490 17382 66505
rect 17426 66490 17450 66505
rect 17494 66490 17518 66505
rect 17562 66490 17586 66505
rect 17630 66490 17654 66505
rect 17698 66490 17722 66505
rect 17766 66490 17790 66505
rect 17834 66490 17858 66505
rect 17902 66490 17926 66505
rect 17970 66490 17994 66505
rect 18038 66490 18062 66505
rect 18106 66490 18130 66505
rect 18174 66490 18198 66505
rect 15678 66335 16678 66490
rect 7389 66245 8389 66305
rect 8990 66245 9990 66305
rect 15678 66301 16690 66335
rect 17278 66325 18278 66490
rect 21413 66380 22813 66508
rect 23685 66380 25085 66508
rect 17266 66301 18278 66325
rect 15678 66290 16678 66301
rect 17278 66290 18278 66301
rect 15748 66277 15772 66290
rect 15816 66277 15840 66290
rect 15884 66277 15908 66290
rect 15952 66277 15976 66290
rect 16020 66277 16044 66290
rect 16088 66277 16112 66290
rect 16156 66277 16180 66290
rect 16224 66277 16248 66290
rect 16292 66277 16316 66290
rect 16360 66277 16384 66290
rect 16428 66277 16452 66290
rect 16496 66277 16520 66290
rect 16564 66277 16588 66290
rect 16632 66277 16656 66290
rect 17290 66277 17314 66290
rect 17358 66277 17382 66290
rect 17426 66277 17450 66290
rect 17494 66277 17518 66290
rect 17562 66277 17586 66290
rect 17630 66277 17654 66290
rect 17698 66277 17722 66290
rect 17766 66277 17790 66290
rect 17834 66277 17858 66290
rect 17902 66277 17926 66290
rect 17970 66277 17994 66290
rect 18038 66277 18062 66290
rect 18106 66277 18130 66290
rect 18174 66277 18198 66290
rect 21413 66217 22813 66345
rect 23685 66217 25085 66345
rect 21413 66054 22813 66182
rect 23685 66054 25085 66182
rect 25936 66132 26936 66182
rect 27274 66033 27358 66036
rect 13899 65998 14059 66002
rect 7389 65887 8389 65943
rect 8990 65887 9990 65943
rect 15678 65932 16678 65988
rect 17278 65932 18278 65988
rect 7389 65815 8389 65871
rect 8990 65815 9990 65871
rect 15678 65860 16678 65916
rect 17278 65860 18278 65916
rect 21413 65891 22813 66019
rect 23685 65891 25085 66019
rect 25936 65976 26936 66032
rect 27158 65983 27358 66033
rect 13899 65852 14059 65856
rect 25936 65820 26936 65876
rect 27158 65807 27358 65935
rect 21413 65741 22813 65784
rect 23685 65741 25085 65784
rect 25936 65664 26936 65720
rect 7389 65513 8389 65585
rect 8990 65513 9990 65585
rect 15678 65558 16678 65630
rect 17278 65558 18278 65630
rect 21413 65605 22813 65648
rect 23685 65605 25085 65648
rect 27158 65631 27358 65687
rect 15748 65547 15782 65558
rect 15816 65547 15850 65558
rect 15884 65547 15918 65558
rect 15952 65547 15986 65558
rect 16020 65547 16054 65558
rect 16088 65547 16122 65558
rect 16156 65547 16190 65558
rect 16224 65547 16258 65558
rect 16292 65547 16326 65558
rect 16360 65547 16394 65558
rect 16428 65547 16462 65558
rect 16496 65547 16530 65558
rect 16564 65547 16598 65558
rect 16632 65547 16666 65558
rect 17290 65547 17324 65558
rect 17358 65547 17392 65558
rect 17426 65547 17460 65558
rect 17494 65547 17528 65558
rect 17562 65547 17596 65558
rect 17630 65547 17664 65558
rect 17698 65547 17732 65558
rect 17766 65547 17800 65558
rect 17834 65547 17868 65558
rect 17902 65547 17936 65558
rect 17970 65547 18004 65558
rect 18038 65547 18072 65558
rect 18106 65547 18140 65558
rect 18174 65547 18208 65558
rect 15748 65537 15806 65547
rect 15816 65537 15874 65547
rect 15884 65537 15942 65547
rect 15952 65537 16010 65547
rect 16020 65537 16078 65547
rect 16088 65537 16146 65547
rect 16156 65537 16214 65547
rect 16224 65537 16282 65547
rect 16292 65537 16350 65547
rect 16360 65537 16418 65547
rect 16428 65537 16486 65547
rect 16496 65537 16554 65547
rect 16564 65537 16622 65547
rect 16632 65537 16690 65547
rect 17290 65537 17348 65547
rect 17358 65537 17416 65547
rect 17426 65537 17484 65547
rect 17494 65537 17552 65547
rect 17562 65537 17620 65547
rect 17630 65537 17688 65547
rect 17698 65537 17756 65547
rect 17766 65537 17824 65547
rect 17834 65537 17892 65547
rect 17902 65537 17960 65547
rect 17970 65537 18028 65547
rect 18038 65537 18096 65547
rect 18106 65537 18164 65547
rect 18174 65537 18232 65547
rect 15724 65513 16690 65537
rect 17266 65513 18232 65537
rect 15748 65498 15772 65513
rect 15816 65498 15840 65513
rect 15884 65498 15908 65513
rect 15952 65498 15976 65513
rect 16020 65498 16044 65513
rect 16088 65498 16112 65513
rect 16156 65498 16180 65513
rect 16224 65498 16248 65513
rect 16292 65498 16316 65513
rect 16360 65498 16384 65513
rect 16428 65498 16452 65513
rect 16496 65498 16520 65513
rect 16564 65498 16588 65513
rect 16632 65498 16656 65513
rect 17290 65498 17314 65513
rect 17358 65498 17382 65513
rect 17426 65498 17450 65513
rect 17494 65498 17518 65513
rect 17562 65498 17586 65513
rect 17630 65498 17654 65513
rect 17698 65498 17722 65513
rect 17766 65498 17790 65513
rect 17834 65498 17858 65513
rect 17902 65498 17926 65513
rect 17970 65498 17994 65513
rect 18038 65498 18062 65513
rect 18106 65498 18130 65513
rect 18174 65498 18198 65513
rect 15678 65343 16678 65498
rect 7389 65253 8389 65313
rect 8990 65253 9990 65313
rect 15678 65309 16690 65343
rect 17278 65333 18278 65498
rect 21413 65442 22813 65570
rect 23685 65442 25085 65570
rect 25936 65514 26936 65564
rect 26393 65511 26477 65514
rect 26726 65511 26810 65514
rect 27158 65455 27358 65583
rect 17266 65309 18278 65333
rect 15678 65298 16678 65309
rect 17278 65298 18278 65309
rect 15748 65285 15772 65298
rect 15816 65285 15840 65298
rect 15884 65285 15908 65298
rect 15952 65285 15976 65298
rect 16020 65285 16044 65298
rect 16088 65285 16112 65298
rect 16156 65285 16180 65298
rect 16224 65285 16248 65298
rect 16292 65285 16316 65298
rect 16360 65285 16384 65298
rect 16428 65285 16452 65298
rect 16496 65285 16520 65298
rect 16564 65285 16588 65298
rect 16632 65285 16656 65298
rect 17290 65285 17314 65298
rect 17358 65285 17382 65298
rect 17426 65285 17450 65298
rect 17494 65285 17518 65298
rect 17562 65285 17586 65298
rect 17630 65285 17654 65298
rect 17698 65285 17722 65298
rect 17766 65285 17790 65298
rect 17834 65285 17858 65298
rect 17902 65285 17926 65298
rect 17970 65285 17994 65298
rect 18038 65285 18062 65298
rect 18106 65285 18130 65298
rect 18174 65285 18198 65298
rect 21413 65279 22813 65407
rect 23685 65279 25085 65407
rect 27158 65279 27358 65335
rect 21413 65116 22813 65244
rect 23685 65116 25085 65244
rect 27158 65103 27358 65231
rect 26393 65100 26477 65103
rect 26726 65100 26810 65103
rect 12543 65069 12881 65085
rect 12559 64967 12865 65069
rect 7389 64895 8389 64951
rect 8990 64895 9990 64951
rect 15678 64940 16678 64996
rect 17278 64940 18278 64996
rect 21413 64953 22813 65081
rect 23685 64953 25085 65081
rect 25936 65050 26936 65100
rect 27622 65095 27672 66095
rect 27772 65095 27828 66095
rect 27928 65095 27984 66095
rect 28084 65095 28140 66095
rect 28240 65095 28296 66095
rect 28396 65637 28446 66095
rect 28396 65553 28449 65637
rect 28396 65305 28446 65553
rect 29778 65320 29802 65344
rect 28396 65221 28449 65305
rect 29802 65296 29826 65309
rect 29880 65299 29914 65333
rect 29778 65261 29802 65285
rect 29890 65275 29914 65299
rect 28396 65095 28446 65221
rect 7389 64823 8389 64879
rect 8990 64823 9990 64879
rect 15678 64868 16678 64924
rect 17278 64868 18278 64924
rect 21413 64790 22813 64918
rect 23685 64790 25085 64918
rect 25936 64894 26936 64950
rect 27158 64927 27358 64983
rect 13899 64656 14059 64660
rect 7389 64521 8389 64593
rect 8990 64521 9990 64593
rect 15678 64566 16678 64638
rect 17278 64566 18278 64638
rect 21413 64627 22813 64755
rect 23685 64627 25085 64755
rect 25936 64738 26936 64794
rect 27158 64751 27358 64879
rect 27912 64757 27962 64873
rect 27909 64673 27962 64757
rect 28082 64673 28210 64873
rect 28258 64673 28314 64873
rect 28434 64673 28562 64873
rect 28610 64673 28660 64873
rect 27917 64669 27951 64673
rect 29880 64672 29914 64706
rect 25936 64582 26936 64638
rect 27158 64581 27358 64631
rect 27274 64578 27358 64581
rect 15748 64555 15782 64566
rect 15816 64555 15850 64566
rect 15884 64555 15918 64566
rect 15952 64555 15986 64566
rect 16020 64555 16054 64566
rect 16088 64555 16122 64566
rect 16156 64555 16190 64566
rect 16224 64555 16258 64566
rect 16292 64555 16326 64566
rect 16360 64555 16394 64566
rect 16428 64555 16462 64566
rect 16496 64555 16530 64566
rect 16564 64555 16598 64566
rect 16632 64555 16666 64566
rect 17290 64555 17324 64566
rect 17358 64555 17392 64566
rect 17426 64555 17460 64566
rect 17494 64555 17528 64566
rect 17562 64555 17596 64566
rect 17630 64555 17664 64566
rect 17698 64555 17732 64566
rect 17766 64555 17800 64566
rect 17834 64555 17868 64566
rect 17902 64555 17936 64566
rect 17970 64555 18004 64566
rect 18038 64555 18072 64566
rect 18106 64555 18140 64566
rect 18174 64555 18208 64566
rect 15748 64545 15806 64555
rect 15816 64545 15874 64555
rect 15884 64545 15942 64555
rect 15952 64545 16010 64555
rect 16020 64545 16078 64555
rect 16088 64545 16146 64555
rect 16156 64545 16214 64555
rect 16224 64545 16282 64555
rect 16292 64545 16350 64555
rect 16360 64545 16418 64555
rect 16428 64545 16486 64555
rect 16496 64545 16554 64555
rect 16564 64545 16622 64555
rect 16632 64545 16690 64555
rect 17290 64545 17348 64555
rect 17358 64545 17416 64555
rect 17426 64545 17484 64555
rect 17494 64545 17552 64555
rect 17562 64545 17620 64555
rect 17630 64545 17688 64555
rect 17698 64545 17756 64555
rect 17766 64545 17824 64555
rect 17834 64545 17892 64555
rect 17902 64545 17960 64555
rect 17970 64545 18028 64555
rect 18038 64545 18096 64555
rect 18106 64545 18164 64555
rect 18174 64545 18232 64555
rect 15724 64521 16690 64545
rect 17266 64521 18232 64545
rect 13901 64510 14061 64514
rect 15748 64506 15772 64521
rect 15816 64506 15840 64521
rect 15884 64506 15908 64521
rect 15952 64506 15976 64521
rect 16020 64506 16044 64521
rect 16088 64506 16112 64521
rect 16156 64506 16180 64521
rect 16224 64506 16248 64521
rect 16292 64506 16316 64521
rect 16360 64506 16384 64521
rect 16428 64506 16452 64521
rect 16496 64506 16520 64521
rect 16564 64506 16588 64521
rect 16632 64506 16656 64521
rect 17290 64506 17314 64521
rect 17358 64506 17382 64521
rect 17426 64506 17450 64521
rect 17494 64506 17518 64521
rect 17562 64506 17586 64521
rect 17630 64506 17654 64521
rect 17698 64506 17722 64521
rect 17766 64506 17790 64521
rect 17834 64506 17858 64521
rect 17902 64506 17926 64521
rect 17970 64506 17994 64521
rect 18038 64506 18062 64521
rect 18106 64506 18130 64521
rect 18174 64506 18198 64521
rect 15678 64351 16678 64506
rect 7389 64261 8389 64321
rect 8990 64261 9990 64321
rect 15678 64317 16690 64351
rect 17278 64341 18278 64506
rect 21413 64470 22813 64520
rect 23685 64470 25085 64520
rect 25936 64432 26936 64482
rect 21349 64390 21373 64414
rect 21407 64390 21431 64414
rect 25067 64390 25091 64414
rect 25125 64390 25149 64414
rect 21383 64356 21397 64390
rect 25101 64356 25115 64390
rect 17266 64317 18278 64341
rect 21349 64332 21373 64356
rect 21407 64332 21431 64356
rect 25067 64332 25091 64356
rect 25125 64332 25149 64356
rect 27917 64325 27951 64329
rect 15678 64306 16678 64317
rect 17278 64306 18278 64317
rect 15748 64293 15772 64306
rect 15816 64293 15840 64306
rect 15884 64293 15908 64306
rect 15952 64293 15976 64306
rect 16020 64293 16044 64306
rect 16088 64293 16112 64306
rect 16156 64293 16180 64306
rect 16224 64293 16248 64306
rect 16292 64293 16316 64306
rect 16360 64293 16384 64306
rect 16428 64293 16452 64306
rect 16496 64293 16520 64306
rect 16564 64293 16588 64306
rect 16632 64293 16656 64306
rect 17290 64293 17314 64306
rect 17358 64293 17382 64306
rect 17426 64293 17450 64306
rect 17494 64293 17518 64306
rect 17562 64293 17586 64306
rect 17630 64293 17654 64306
rect 17698 64293 17722 64306
rect 17766 64293 17790 64306
rect 17834 64293 17858 64306
rect 17902 64293 17926 64306
rect 17970 64293 17994 64306
rect 18038 64293 18062 64306
rect 18106 64293 18130 64306
rect 18174 64293 18198 64306
rect 27909 64241 27962 64325
rect 21634 64101 24864 64203
rect 27912 64125 27962 64241
rect 28082 64125 28210 64325
rect 28258 64125 28314 64325
rect 28434 64125 28562 64325
rect 28610 64125 28660 64325
rect 21186 64047 21210 64071
rect 25288 64047 25312 64071
rect 21162 64023 21186 64037
rect 25312 64023 25336 64037
rect 7389 63903 8389 63959
rect 8990 63903 9990 63959
rect 15678 63948 16678 64004
rect 17278 63948 18278 64004
rect 21072 63989 21084 64013
rect 21186 63989 21210 64013
rect 25288 63989 25312 64013
rect 25414 63989 25426 64013
rect 21385 63944 21403 63948
rect 7389 63831 8389 63887
rect 8990 63831 9990 63887
rect 15678 63876 16678 63932
rect 17278 63876 18278 63932
rect 20250 63914 20316 63930
rect 21377 63914 21403 63944
rect 21385 63904 21403 63914
rect 21383 63880 21403 63904
rect 21407 63880 21415 63914
rect 25113 63904 25121 63944
rect 25101 63880 25121 63904
rect 25125 63880 25143 63948
rect 21383 63846 21419 63880
rect 25101 63846 25147 63880
rect 21383 63812 21403 63846
rect 21407 63812 21415 63846
rect 21383 63778 21419 63812
rect 21481 63784 22881 63834
rect 23617 63784 25017 63834
rect 25101 63812 25121 63846
rect 25125 63812 25143 63846
rect 25101 63778 25147 63812
rect 21383 63744 21403 63778
rect 21407 63744 21415 63778
rect 21383 63710 21419 63744
rect 21383 63676 21403 63710
rect 21407 63676 21415 63710
rect 7389 63529 8389 63601
rect 8990 63529 9990 63601
rect 15678 63574 16678 63646
rect 17278 63574 18278 63646
rect 21383 63642 21419 63676
rect 21383 63608 21403 63642
rect 21407 63608 21415 63642
rect 21481 63621 22881 63749
rect 23617 63621 25017 63749
rect 25101 63744 25121 63778
rect 25125 63744 25143 63778
rect 25101 63710 25147 63744
rect 25101 63676 25121 63710
rect 25125 63676 25143 63710
rect 25101 63642 25147 63676
rect 25101 63608 25121 63642
rect 25125 63608 25143 63642
rect 21383 63574 21419 63608
rect 15748 63563 15782 63574
rect 15816 63563 15850 63574
rect 15884 63563 15918 63574
rect 15952 63563 15986 63574
rect 16020 63563 16054 63574
rect 16088 63563 16122 63574
rect 16156 63563 16190 63574
rect 16224 63563 16258 63574
rect 16292 63563 16326 63574
rect 16360 63563 16394 63574
rect 16428 63563 16462 63574
rect 16496 63563 16530 63574
rect 16564 63563 16598 63574
rect 16632 63563 16666 63574
rect 17290 63563 17324 63574
rect 17358 63563 17392 63574
rect 17426 63563 17460 63574
rect 17494 63563 17528 63574
rect 17562 63563 17596 63574
rect 17630 63563 17664 63574
rect 17698 63563 17732 63574
rect 17766 63563 17800 63574
rect 17834 63563 17868 63574
rect 17902 63563 17936 63574
rect 17970 63563 18004 63574
rect 18038 63563 18072 63574
rect 18106 63563 18140 63574
rect 18174 63563 18208 63574
rect 15748 63553 15806 63563
rect 15816 63553 15874 63563
rect 15884 63553 15942 63563
rect 15952 63553 16010 63563
rect 16020 63553 16078 63563
rect 16088 63553 16146 63563
rect 16156 63553 16214 63563
rect 16224 63553 16282 63563
rect 16292 63553 16350 63563
rect 16360 63553 16418 63563
rect 16428 63553 16486 63563
rect 16496 63553 16554 63563
rect 16564 63553 16622 63563
rect 16632 63553 16690 63563
rect 17290 63553 17348 63563
rect 17358 63553 17416 63563
rect 17426 63553 17484 63563
rect 17494 63553 17552 63563
rect 17562 63553 17620 63563
rect 17630 63553 17688 63563
rect 17698 63553 17756 63563
rect 17766 63553 17824 63563
rect 17834 63553 17892 63563
rect 17902 63553 17960 63563
rect 17970 63553 18028 63563
rect 18038 63553 18096 63563
rect 18106 63553 18164 63563
rect 18174 63553 18232 63563
rect 15724 63529 16690 63553
rect 17266 63529 18232 63553
rect 21383 63540 21403 63574
rect 21407 63540 21415 63574
rect 15748 63514 15772 63529
rect 15816 63514 15840 63529
rect 15884 63514 15908 63529
rect 15952 63514 15976 63529
rect 16020 63514 16044 63529
rect 16088 63514 16112 63529
rect 16156 63514 16180 63529
rect 16224 63514 16248 63529
rect 16292 63514 16316 63529
rect 16360 63514 16384 63529
rect 16428 63514 16452 63529
rect 16496 63514 16520 63529
rect 16564 63514 16588 63529
rect 16632 63514 16656 63529
rect 17290 63514 17314 63529
rect 17358 63514 17382 63529
rect 17426 63514 17450 63529
rect 17494 63514 17518 63529
rect 17562 63514 17586 63529
rect 17630 63514 17654 63529
rect 17698 63514 17722 63529
rect 17766 63514 17790 63529
rect 17834 63514 17858 63529
rect 17902 63514 17926 63529
rect 17970 63514 17994 63529
rect 18038 63514 18062 63529
rect 18106 63514 18130 63529
rect 18174 63514 18198 63529
rect 5937 63318 6089 63386
rect 15678 63359 16678 63514
rect 6005 63315 6089 63318
rect 5967 63305 6059 63315
rect 6005 63275 6021 63305
rect 1288 61503 1338 62503
rect 1438 61503 1566 62503
rect 1594 61503 1644 62503
rect 5995 61493 6021 63275
rect 7389 63269 8389 63329
rect 8990 63269 9990 63329
rect 15678 63325 16690 63359
rect 17278 63349 18278 63514
rect 17266 63325 18278 63349
rect 15678 63314 16678 63325
rect 17278 63314 18278 63325
rect 21383 63506 21419 63540
rect 21383 63472 21403 63506
rect 21407 63472 21415 63506
rect 21383 63438 21419 63472
rect 21481 63458 22881 63586
rect 23617 63458 25017 63586
rect 25101 63574 25147 63608
rect 25101 63540 25121 63574
rect 25125 63540 25143 63574
rect 25101 63506 25147 63540
rect 25101 63472 25121 63506
rect 25125 63472 25143 63506
rect 25101 63438 25147 63472
rect 21383 63404 21403 63438
rect 21407 63404 21415 63438
rect 21383 63370 21419 63404
rect 21383 63336 21403 63370
rect 21407 63336 21415 63370
rect 15748 63301 15772 63314
rect 15816 63301 15840 63314
rect 15884 63301 15908 63314
rect 15952 63301 15976 63314
rect 16020 63301 16044 63314
rect 16088 63301 16112 63314
rect 16156 63301 16180 63314
rect 16224 63301 16248 63314
rect 16292 63301 16316 63314
rect 16360 63301 16384 63314
rect 16428 63301 16452 63314
rect 16496 63301 16520 63314
rect 16564 63301 16588 63314
rect 16632 63301 16656 63314
rect 17290 63301 17314 63314
rect 17358 63301 17382 63314
rect 17426 63301 17450 63314
rect 17494 63301 17518 63314
rect 17562 63301 17586 63314
rect 17630 63301 17654 63314
rect 17698 63301 17722 63314
rect 17766 63301 17790 63314
rect 17834 63301 17858 63314
rect 17902 63301 17926 63314
rect 17970 63301 17994 63314
rect 18038 63301 18062 63314
rect 18106 63301 18130 63314
rect 18174 63301 18198 63314
rect 21383 63302 21419 63336
rect 21383 63268 21403 63302
rect 21407 63268 21415 63302
rect 21481 63295 22881 63423
rect 23617 63295 25017 63423
rect 25101 63404 25121 63438
rect 25125 63404 25143 63438
rect 25101 63370 25147 63404
rect 25101 63336 25121 63370
rect 25125 63336 25143 63370
rect 25101 63302 25147 63336
rect 25101 63268 25121 63302
rect 25125 63268 25143 63302
rect 21383 63234 21419 63268
rect 21383 63200 21403 63234
rect 21407 63200 21415 63234
rect 21383 63166 21419 63200
rect 21383 63132 21403 63166
rect 21407 63132 21415 63166
rect 21481 63132 22881 63260
rect 23617 63132 25017 63260
rect 25101 63234 25147 63268
rect 25101 63200 25121 63234
rect 25125 63200 25143 63234
rect 25101 63166 25147 63200
rect 25101 63132 25121 63166
rect 25125 63132 25143 63166
rect 21383 63098 21419 63132
rect 25101 63098 25147 63132
rect 21383 63064 21403 63098
rect 21407 63064 21415 63098
rect 21383 63030 21419 63064
rect 7389 62911 8389 62967
rect 8990 62911 9990 62967
rect 15678 62956 16678 63012
rect 17278 62956 18278 63012
rect 21383 62996 21403 63030
rect 21407 62996 21415 63030
rect 21383 62962 21419 62996
rect 21481 62969 22881 63097
rect 23617 62969 25017 63097
rect 25101 63064 25121 63098
rect 25125 63064 25143 63098
rect 25101 63030 25147 63064
rect 25101 62996 25121 63030
rect 25125 62996 25143 63030
rect 25101 62962 25147 62996
rect 26478 62985 26648 63291
rect 7389 62839 8389 62895
rect 8990 62839 9990 62895
rect 15678 62884 16678 62940
rect 17278 62884 18278 62940
rect 21383 62928 21403 62962
rect 21407 62928 21415 62962
rect 21383 62894 21419 62928
rect 21383 62860 21403 62894
rect 21407 62860 21415 62894
rect 21383 62826 21419 62860
rect 21383 62792 21403 62826
rect 21407 62792 21415 62826
rect 21481 62806 22881 62934
rect 23617 62806 25017 62934
rect 25101 62928 25121 62962
rect 25125 62928 25143 62962
rect 25101 62894 25147 62928
rect 27622 62903 27672 63903
rect 27772 62903 27828 63903
rect 27928 62903 27984 63903
rect 28084 62903 28140 63903
rect 28240 62903 28296 63903
rect 28396 63777 28446 63903
rect 28396 63693 28449 63777
rect 28396 63445 28446 63693
rect 30015 63523 30027 69246
rect 32596 69239 33596 69367
rect 35255 69345 36255 69401
rect 30135 69062 30735 69112
rect 31049 69042 32049 69092
rect 32596 69083 33596 69211
rect 35255 69169 36255 69297
rect 35255 68993 36255 69121
rect 30135 68886 30735 68942
rect 31049 68886 32049 68942
rect 32596 68927 33596 68983
rect 37998 68979 38148 68991
rect 38317 68979 38467 68991
rect 30135 68716 30735 68766
rect 31049 68736 32049 68786
rect 32596 68777 33596 68827
rect 35255 68823 36255 68873
rect 37998 68866 38598 68916
rect 35255 68754 36255 68766
rect 37998 68690 38598 68746
rect 30135 68600 30735 68650
rect 31049 68600 32049 68650
rect 32596 68575 33196 68625
rect 35255 68621 36255 68671
rect 30135 68424 30735 68480
rect 31049 68444 32049 68500
rect 30135 68248 30735 68376
rect 31049 68288 32049 68344
rect 30135 68072 30735 68200
rect 31049 68132 32049 68188
rect 32596 68141 33196 68191
rect 30135 67896 30735 68024
rect 31049 67982 32049 68032
rect 31049 67866 32049 67916
rect 30135 67726 30735 67776
rect 31049 67710 32049 67838
rect 30135 67610 30735 67660
rect 30135 67434 30735 67562
rect 31049 67554 32049 67682
rect 31049 67398 32049 67526
rect 34152 67490 34202 68478
rect 34322 67490 34372 68478
rect 34492 68465 35092 68515
rect 35255 68445 36255 68573
rect 37998 68520 38598 68570
rect 36785 68496 36797 68500
rect 36785 68485 36800 68496
rect 36970 68485 36985 68500
rect 34492 68289 35092 68345
rect 35255 68269 36255 68325
rect 36785 68305 36985 68485
rect 36785 68294 36800 68305
rect 36785 68290 36797 68294
rect 36970 68290 36985 68305
rect 37083 68485 37098 68500
rect 37083 68305 37120 68485
rect 37083 68290 37098 68305
rect 36785 68260 36797 68264
rect 36785 68249 36800 68260
rect 36970 68249 36985 68264
rect 34492 68119 35092 68169
rect 35255 68099 36255 68149
rect 36785 68069 36985 68249
rect 37993 68094 38593 68144
rect 36785 68058 36800 68069
rect 36785 68054 36797 68058
rect 36970 68054 36985 68069
rect 34491 67849 35091 67899
rect 35255 67883 35855 67933
rect 37993 67924 38593 67974
rect 34491 67673 35091 67729
rect 35255 67707 35855 67763
rect 36785 67748 37385 67798
rect 38920 67761 38946 67787
rect 34491 67503 35091 67553
rect 35255 67531 35855 67659
rect 36785 67572 37385 67628
rect 34019 67418 34029 67490
rect 34152 67478 34372 67490
rect 34091 67415 34101 67418
rect 30135 67258 30735 67314
rect 31049 67242 32049 67370
rect 34091 67365 35091 67415
rect 35255 67361 35855 67411
rect 36785 67396 37385 67452
rect 30135 67082 30735 67210
rect 31049 67086 32049 67214
rect 34091 67195 35091 67245
rect 36785 67226 37385 67276
rect 34091 67192 34101 67195
rect 34202 67192 34302 67195
rect 35255 67159 35855 67209
rect 30135 66912 30735 66962
rect 31049 66930 32049 66986
rect 30135 66796 30735 66846
rect 31049 66774 32049 66902
rect 32481 66898 33081 66948
rect 30135 66620 30735 66748
rect 31049 66618 32049 66746
rect 32481 66742 33081 66870
rect 30135 66444 30735 66572
rect 31049 66462 32049 66590
rect 32481 66586 33081 66714
rect 34152 66532 34202 67132
rect 34302 66532 34352 67132
rect 34491 67066 35091 67116
rect 35255 67003 35855 67131
rect 36785 67094 37385 67144
rect 34491 66890 35091 66946
rect 36785 66918 37385 66974
rect 35255 66847 35855 66903
rect 34491 66720 35091 66770
rect 35255 66691 35855 66819
rect 36785 66742 37385 66798
rect 35255 66541 35855 66591
rect 36785 66572 37385 66622
rect 32481 66436 33081 66486
rect 30135 66268 30735 66396
rect 31049 66306 32049 66434
rect 34491 66379 35091 66429
rect 37993 66396 38593 66446
rect 32481 66306 33081 66356
rect 33261 66287 33861 66323
rect 30135 66092 30735 66220
rect 31049 66150 32049 66278
rect 32481 66150 33081 66278
rect 34491 66203 35091 66331
rect 35255 66287 35855 66337
rect 36785 66312 36797 66316
rect 36785 66301 36800 66312
rect 36970 66301 36985 66316
rect 35255 66131 35855 66259
rect 36785 66121 36985 66301
rect 37993 66226 38593 66276
rect 36785 66110 36800 66121
rect 36785 66106 36797 66110
rect 36970 66106 36985 66121
rect 30135 65916 30735 66044
rect 31049 65994 32049 66050
rect 32481 65994 33081 66050
rect 34491 66027 35091 66083
rect 31049 65818 32049 65946
rect 32481 65838 33081 65966
rect 33261 65907 33861 65963
rect 34491 65851 35091 65979
rect 35255 65975 35855 66103
rect 36785 66076 36797 66080
rect 36785 66065 36800 66076
rect 36970 66065 36985 66080
rect 36785 65885 36985 66065
rect 35255 65819 35855 65875
rect 36785 65874 36800 65885
rect 36785 65870 36797 65874
rect 36970 65870 36985 65885
rect 37083 66065 37098 66080
rect 37083 65885 37120 66065
rect 37083 65870 37098 65885
rect 37998 65800 38598 65850
rect 30135 65740 30735 65796
rect 30135 65564 30735 65692
rect 31049 65642 32049 65770
rect 32481 65688 33081 65738
rect 33261 65723 33861 65773
rect 34491 65681 35091 65731
rect 35255 65669 35855 65719
rect 37998 65624 38598 65680
rect 30135 65388 30735 65516
rect 31049 65466 32049 65594
rect 32481 65558 33081 65608
rect 30135 65212 30735 65340
rect 31049 65290 32049 65418
rect 32481 65402 33081 65458
rect 37998 65454 38598 65504
rect 37998 65451 38220 65454
rect 38245 65451 38539 65454
rect 32481 65252 33081 65302
rect 34427 65259 35027 65309
rect 30135 65036 30735 65164
rect 31049 65114 32049 65242
rect 33672 65183 34272 65233
rect 34427 65083 35027 65211
rect 30135 64860 30735 64988
rect 31049 64938 32049 65066
rect 33672 65007 34272 65063
rect 31049 64762 32049 64890
rect 33672 64831 34272 64959
rect 34427 64907 35027 65035
rect 30135 64684 30735 64740
rect 34427 64731 35027 64859
rect 37998 64825 38148 64837
rect 38317 64825 38467 64837
rect 37998 64712 38598 64762
rect 33672 64655 34272 64711
rect 30135 64508 30735 64636
rect 31049 64592 32049 64642
rect 34427 64555 35027 64683
rect 37998 64536 38598 64592
rect 31049 64476 32049 64526
rect 33672 64479 34272 64535
rect 30135 64332 30735 64388
rect 31049 64320 32049 64448
rect 34427 64379 35027 64435
rect 37998 64366 38598 64416
rect 33672 64303 34272 64359
rect 36785 64342 36797 64346
rect 36785 64331 36800 64342
rect 36970 64331 36985 64346
rect 30135 64156 30735 64284
rect 31049 64164 32049 64292
rect 30135 63980 30735 64036
rect 31049 64008 32049 64136
rect 33672 64127 34272 64255
rect 34427 64203 35027 64331
rect 36785 64151 36985 64331
rect 36785 64140 36800 64151
rect 36785 64136 36797 64140
rect 36970 64136 36985 64151
rect 37083 64331 37098 64346
rect 37083 64151 37120 64331
rect 37083 64136 37098 64151
rect 36785 64106 36797 64110
rect 36785 64095 36800 64106
rect 36970 64095 36985 64110
rect 34427 64033 35027 64083
rect 33672 63957 34272 64007
rect 30135 63804 30735 63932
rect 36785 63915 36985 64095
rect 37993 63940 38593 63990
rect 31049 63852 32049 63908
rect 36785 63904 36800 63915
rect 36785 63900 36797 63904
rect 36970 63900 36985 63915
rect 31049 63696 32049 63824
rect 37993 63770 38593 63820
rect 30135 63634 30735 63684
rect 31049 63540 32049 63668
rect 36785 63594 37385 63644
rect 28396 63361 28449 63445
rect 31049 63384 32049 63512
rect 36785 63418 37385 63474
rect 28396 62903 28446 63361
rect 31049 63234 32049 63284
rect 36785 63242 37385 63298
rect 36785 63072 37385 63122
rect 37939 63039 37963 63063
rect 38085 63039 38109 63063
rect 29925 63003 29931 63032
rect 30271 63003 30305 63027
rect 30342 63003 30376 63027
rect 30413 63003 30447 63027
rect 30484 63003 30518 63027
rect 30555 63003 30589 63027
rect 30626 63003 30660 63027
rect 30697 63003 30731 63027
rect 37963 63015 37987 63038
rect 38061 63015 38085 63038
rect 29931 62962 29939 62986
rect 29955 62962 29961 63003
rect 29891 62938 29915 62962
rect 25101 62860 25121 62894
rect 25125 62860 25143 62894
rect 37759 62867 37783 62891
rect 25101 62826 25147 62860
rect 37792 62843 37807 62867
rect 25101 62792 25121 62826
rect 25125 62792 25143 62826
rect 21383 62758 21419 62792
rect 25101 62758 25147 62792
rect 21383 62724 21403 62758
rect 21407 62724 21415 62758
rect 25101 62724 25121 62758
rect 25125 62724 25143 62758
rect 21383 62690 21419 62724
rect 21383 62656 21403 62690
rect 21407 62656 21415 62690
rect 21481 62656 22881 62699
rect 22892 62675 22920 62703
rect 23617 62656 25017 62699
rect 25101 62690 25147 62724
rect 31458 62703 31608 62715
rect 31777 62703 31927 62715
rect 25101 62656 25121 62690
rect 25125 62656 25143 62690
rect 7389 62628 8389 62632
rect 8990 62628 9990 62632
rect 7353 62578 8425 62614
rect 7353 62537 7389 62578
rect 8389 62537 8425 62578
rect 7353 62501 8425 62537
rect 8954 62578 10026 62614
rect 15678 62582 16678 62654
rect 17278 62582 18278 62654
rect 21383 62622 21419 62656
rect 25101 62622 25147 62656
rect 21383 62588 21403 62622
rect 21407 62588 21415 62622
rect 25101 62588 25121 62622
rect 25125 62588 25143 62622
rect 8954 62537 8990 62578
rect 9990 62537 10026 62578
rect 15748 62571 15782 62582
rect 15816 62571 15850 62582
rect 15884 62571 15918 62582
rect 15952 62571 15986 62582
rect 16020 62571 16054 62582
rect 16088 62571 16122 62582
rect 16156 62571 16190 62582
rect 16224 62571 16258 62582
rect 16292 62571 16326 62582
rect 16360 62571 16394 62582
rect 16428 62571 16462 62582
rect 16496 62571 16530 62582
rect 16564 62571 16598 62582
rect 16632 62571 16666 62582
rect 17290 62571 17324 62582
rect 17358 62571 17392 62582
rect 17426 62571 17460 62582
rect 17494 62571 17528 62582
rect 17562 62571 17596 62582
rect 17630 62571 17664 62582
rect 17698 62571 17732 62582
rect 17766 62571 17800 62582
rect 17834 62571 17868 62582
rect 17902 62571 17936 62582
rect 17970 62571 18004 62582
rect 18038 62571 18072 62582
rect 18106 62571 18140 62582
rect 18174 62571 18208 62582
rect 15748 62561 15806 62571
rect 15816 62561 15874 62571
rect 15884 62561 15942 62571
rect 15952 62561 16010 62571
rect 16020 62561 16078 62571
rect 16088 62561 16146 62571
rect 16156 62561 16214 62571
rect 16224 62561 16282 62571
rect 16292 62561 16350 62571
rect 16360 62561 16418 62571
rect 16428 62561 16486 62571
rect 16496 62561 16554 62571
rect 16564 62561 16622 62571
rect 16632 62561 16690 62571
rect 17290 62561 17348 62571
rect 17358 62561 17416 62571
rect 17426 62561 17484 62571
rect 17494 62561 17552 62571
rect 17562 62561 17620 62571
rect 17630 62561 17688 62571
rect 17698 62561 17756 62571
rect 17766 62561 17824 62571
rect 17834 62561 17892 62571
rect 17902 62561 17960 62571
rect 17970 62561 18028 62571
rect 18038 62561 18096 62571
rect 18106 62561 18164 62571
rect 18174 62561 18232 62571
rect 15724 62537 16690 62561
rect 17266 62537 18232 62561
rect 21383 62554 21419 62588
rect 8954 62501 10026 62537
rect 15748 62522 15772 62537
rect 15816 62522 15840 62537
rect 15884 62522 15908 62537
rect 15952 62522 15976 62537
rect 16020 62522 16044 62537
rect 16088 62522 16112 62537
rect 16156 62522 16180 62537
rect 16224 62522 16248 62537
rect 16292 62522 16316 62537
rect 16360 62522 16384 62537
rect 16428 62522 16452 62537
rect 16496 62522 16520 62537
rect 16564 62522 16588 62537
rect 16632 62522 16656 62537
rect 17290 62522 17314 62537
rect 17358 62522 17382 62537
rect 17426 62522 17450 62537
rect 17494 62522 17518 62537
rect 17562 62522 17586 62537
rect 17630 62522 17654 62537
rect 17698 62522 17722 62537
rect 17766 62522 17790 62537
rect 17834 62522 17858 62537
rect 17902 62522 17926 62537
rect 17970 62522 17994 62537
rect 18038 62522 18062 62537
rect 18106 62522 18130 62537
rect 18174 62522 18198 62537
rect 15678 62367 16678 62522
rect 7389 62277 8389 62337
rect 8990 62277 9990 62337
rect 15678 62333 16690 62367
rect 17278 62357 18278 62522
rect 17266 62333 18278 62357
rect 15678 62322 16678 62333
rect 17278 62322 18278 62333
rect 21383 62520 21403 62554
rect 21407 62520 21415 62554
rect 21481 62520 22881 62563
rect 23617 62520 25017 62563
rect 25101 62554 25147 62588
rect 25414 62573 25438 62607
rect 31458 62590 32058 62640
rect 25101 62520 25121 62554
rect 25125 62520 25143 62554
rect 21383 62486 21419 62520
rect 25101 62486 25147 62520
rect 21383 62452 21403 62486
rect 21407 62452 21415 62486
rect 21383 62418 21419 62452
rect 21383 62384 21403 62418
rect 21407 62384 21415 62418
rect 21383 62350 21419 62384
rect 21481 62357 22881 62485
rect 23617 62357 25017 62485
rect 25101 62452 25121 62486
rect 25125 62452 25143 62486
rect 37792 62470 37807 62494
rect 25101 62418 25147 62452
rect 25101 62384 25121 62418
rect 25125 62384 25143 62418
rect 31458 62414 32058 62470
rect 37759 62446 37783 62470
rect 25101 62350 25147 62384
rect 15748 62309 15772 62322
rect 15816 62309 15840 62322
rect 15884 62309 15908 62322
rect 15952 62309 15976 62322
rect 16020 62309 16044 62322
rect 16088 62309 16112 62322
rect 16156 62309 16180 62322
rect 16224 62309 16248 62322
rect 16292 62309 16316 62322
rect 16360 62309 16384 62322
rect 16428 62309 16452 62322
rect 16496 62309 16520 62322
rect 16564 62309 16588 62322
rect 16632 62309 16656 62322
rect 17290 62309 17314 62322
rect 17358 62309 17382 62322
rect 17426 62309 17450 62322
rect 17494 62309 17518 62322
rect 17562 62309 17586 62322
rect 17630 62309 17654 62322
rect 17698 62309 17722 62322
rect 17766 62309 17790 62322
rect 17834 62309 17858 62322
rect 17902 62309 17926 62322
rect 17970 62309 17994 62322
rect 18038 62309 18062 62322
rect 18106 62309 18130 62322
rect 18174 62309 18198 62322
rect 21383 62316 21403 62350
rect 21407 62316 21415 62350
rect 21383 62282 21419 62316
rect 21383 62248 21403 62282
rect 21407 62248 21415 62282
rect 21383 62214 21419 62248
rect 21383 62180 21403 62214
rect 21407 62180 21415 62214
rect 21481 62194 22881 62322
rect 23617 62194 25017 62322
rect 25101 62316 25121 62350
rect 25125 62316 25143 62350
rect 25101 62282 25147 62316
rect 25101 62248 25121 62282
rect 25125 62248 25143 62282
rect 25101 62214 25147 62248
rect 25101 62180 25121 62214
rect 25125 62180 25143 62214
rect 25725 62197 26325 62247
rect 31458 62244 32058 62294
rect 30245 62220 30257 62224
rect 30245 62209 30260 62220
rect 30430 62209 30445 62224
rect 21383 62146 21419 62180
rect 7389 62066 8389 62070
rect 8990 62066 9990 62070
rect 15678 62061 16678 62133
rect 17278 62061 18278 62133
rect 21383 62112 21403 62146
rect 21407 62112 21415 62146
rect 21383 62078 21419 62112
rect 7353 62016 8425 62052
rect 7353 61975 7389 62016
rect 8389 61975 8425 62016
rect 7353 61919 8425 61975
rect 7353 61903 7389 61919
rect 8389 61903 8425 61919
rect 7353 61847 8425 61903
rect 7353 61810 7389 61847
rect 8389 61810 8425 61847
rect 7353 61770 8425 61810
rect 8954 62016 10026 62052
rect 8954 61975 8990 62016
rect 9990 61975 10026 62016
rect 8954 61919 10026 61975
rect 21383 62044 21403 62078
rect 21407 62044 21415 62078
rect 21383 62010 21419 62044
rect 21481 62031 22881 62159
rect 23617 62031 25017 62159
rect 25101 62146 25147 62180
rect 25101 62112 25121 62146
rect 25125 62112 25143 62146
rect 25101 62078 25147 62112
rect 25101 62044 25121 62078
rect 25125 62044 25143 62078
rect 25725 62047 26325 62097
rect 25101 62010 25147 62044
rect 21383 61976 21403 62010
rect 21407 61976 21415 62010
rect 21383 61942 21419 61976
rect 8954 61903 8990 61919
rect 9990 61903 10026 61919
rect 15678 61906 16678 61923
rect 17278 61906 18278 61923
rect 21383 61908 21403 61942
rect 21407 61908 21415 61942
rect 8954 61847 10026 61903
rect 20250 61890 20316 61906
rect 8954 61810 8990 61847
rect 9990 61810 10026 61847
rect 8954 61770 10026 61810
rect 21383 61874 21419 61908
rect 21383 61840 21403 61874
rect 21407 61840 21415 61874
rect 21481 61868 22881 61996
rect 23617 61868 25017 61996
rect 25101 61976 25121 62010
rect 25125 61976 25143 62010
rect 25101 61942 25147 61976
rect 25101 61908 25121 61942
rect 25125 61908 25143 61942
rect 25725 61925 26325 61975
rect 25101 61874 25147 61908
rect 25101 61840 25121 61874
rect 25125 61840 25143 61874
rect 21383 61806 21419 61840
rect 21383 61772 21403 61806
rect 21407 61772 21415 61806
rect 21383 61738 21419 61772
rect 15678 61703 16678 61736
rect 17278 61703 18278 61736
rect 21383 61704 21403 61738
rect 21407 61704 21415 61738
rect 21481 61705 22881 61833
rect 23617 61705 25017 61833
rect 25101 61806 25147 61840
rect 25101 61772 25121 61806
rect 25125 61772 25143 61806
rect 25725 61775 26325 61825
rect 25101 61738 25147 61772
rect 25101 61704 25121 61738
rect 25125 61704 25143 61738
rect 21383 61670 21419 61704
rect 25101 61670 25147 61704
rect 21383 61636 21403 61670
rect 21407 61636 21415 61670
rect 7389 61559 8389 61631
rect 8990 61559 9990 61631
rect 21383 61602 21419 61636
rect 15840 61510 15870 61580
rect 15878 61546 15908 61580
rect 21383 61568 21403 61602
rect 21407 61568 21415 61602
rect 15853 61508 15870 61510
rect 21383 61534 21419 61568
rect 21481 61542 22881 61670
rect 23617 61542 25017 61670
rect 25101 61636 25121 61670
rect 25125 61636 25143 61670
rect 25725 61649 26325 61699
rect 25101 61602 25147 61636
rect 25101 61568 25121 61602
rect 25125 61568 25143 61602
rect 25101 61534 25147 61568
rect 5981 61483 6021 61493
rect 5137 61469 6021 61483
rect 21383 61500 21403 61534
rect 21407 61500 21415 61534
rect 21383 61466 21419 61500
rect 7389 61369 8389 61463
rect 7389 61359 8413 61369
rect 8990 61359 9990 61463
rect 21383 61432 21403 61466
rect 21407 61432 21415 61466
rect 21383 61398 21419 61432
rect 21383 61364 21403 61398
rect 21407 61364 21415 61398
rect 21481 61379 22881 61507
rect 23617 61379 25017 61507
rect 25101 61500 25121 61534
rect 25125 61500 25143 61534
rect 25101 61466 25147 61500
rect 25725 61499 26325 61549
rect 25101 61432 25121 61466
rect 25125 61432 25143 61466
rect 25101 61398 25147 61432
rect 25101 61364 25121 61398
rect 25125 61364 25143 61398
rect 25725 61377 26325 61427
rect 21383 61330 21419 61364
rect 25101 61330 25147 61364
rect 21383 61296 21403 61330
rect 21407 61296 21415 61330
rect 25101 61296 25121 61330
rect 25125 61296 25143 61330
rect 21383 61262 21419 61296
rect 21383 61228 21403 61262
rect 21407 61228 21415 61262
rect 21481 61229 22881 61272
rect 23617 61229 25017 61272
rect 25101 61262 25147 61296
rect 25101 61228 25121 61262
rect 25125 61228 25143 61262
rect 21383 61194 21419 61228
rect 25101 61194 25147 61228
rect 25725 61227 26325 61277
rect 21383 61160 21403 61194
rect 21407 61160 21415 61194
rect 25101 61160 25121 61194
rect 25125 61160 25143 61194
rect 27162 61170 27212 62170
rect 27312 61170 27440 62170
rect 27468 61170 27596 62170
rect 27624 61170 27752 62170
rect 27780 61170 27908 62170
rect 27936 61170 28064 62170
rect 28092 61170 28220 62170
rect 28248 61170 28376 62170
rect 28404 61170 28532 62170
rect 28560 61170 28688 62170
rect 28716 61170 28844 62170
rect 28872 61170 29000 62170
rect 29028 61170 29156 62170
rect 29184 61170 29312 62170
rect 29340 61170 29390 62170
rect 30245 62029 30445 62209
rect 30245 62018 30260 62029
rect 30245 62014 30257 62018
rect 30430 62014 30445 62029
rect 30543 62209 30558 62224
rect 30543 62029 30580 62209
rect 30543 62014 30558 62029
rect 30245 61984 30257 61988
rect 30245 61973 30260 61984
rect 30430 61973 30445 61988
rect 30245 61793 30445 61973
rect 31453 61818 32053 61868
rect 30245 61782 30260 61793
rect 30245 61778 30257 61782
rect 30430 61778 30445 61793
rect 31453 61648 32053 61698
rect 30245 61472 30845 61522
rect 30245 61296 30845 61352
rect 21383 61126 21419 61160
rect 25101 61126 25147 61160
rect 21383 61102 21403 61126
rect 21385 61048 21403 61102
rect 21407 61082 21415 61126
rect 25101 61102 25121 61126
rect 25113 61082 25121 61102
rect 25125 61048 25143 61126
rect 30245 61120 30845 61176
rect 30245 60950 30845 61000
rect 21000 60800 21003 60920
rect 21352 60885 21376 60909
rect 25122 60885 25146 60909
rect 21385 60861 21400 60885
rect 25098 60861 25113 60885
rect 21274 60783 21294 60851
rect 21410 60817 21430 60851
rect 25068 60817 25088 60851
rect 25204 60817 25224 60851
rect 21385 60807 21430 60817
rect 25102 60807 25137 60817
rect 21361 60783 21430 60807
rect 25089 60783 25137 60807
rect 25238 60783 25258 60817
rect 680480 58427 680517 58520
rect 680615 58427 680815 58520
rect 685793 58483 685993 58520
rect 686053 58483 686253 58520
rect 686607 58440 687607 58490
rect 692427 58392 693027 58448
rect 679007 58216 679607 58266
rect 680615 58191 680815 58371
rect 686829 58301 687429 58351
rect 684004 58243 685004 58293
rect 695201 58282 695251 58520
rect 696287 58282 696337 58520
rect 682890 58161 683490 58211
rect 684004 58127 685004 58177
rect 686829 58125 687429 58181
rect 679007 58046 679607 58096
rect 684004 57971 685004 58027
rect 686829 57955 687429 58005
rect 680215 57870 680815 57920
rect 681713 57881 682313 57931
rect 682921 57899 683521 57949
rect 692427 57930 693027 57980
rect 684004 57821 685004 57871
rect 680215 57694 680815 57750
rect 681713 57705 682313 57761
rect 682921 57743 683521 57799
rect 685537 57749 686137 57799
rect 697088 57749 697138 58520
rect 697706 57749 697756 58520
rect 699322 58374 700322 58514
rect 700922 58374 701922 58514
rect 707610 58098 708610 58099
rect 699322 57956 700322 58012
rect 700922 57956 701922 58012
rect 707610 58001 708610 58057
rect 709211 58001 710211 58057
rect 707610 57959 708610 57960
rect 699322 57884 700322 57940
rect 700922 57884 701922 57940
rect 709211 57936 710211 57960
rect 682921 57593 683521 57643
rect 684070 57599 684670 57649
rect 685537 57593 686137 57649
rect 699322 57623 700322 57673
rect 700922 57623 701922 57673
rect 680215 57518 680815 57574
rect 707610 57523 708610 57617
rect 709211 57523 710211 57591
rect 707610 57513 707624 57523
rect 707658 57513 707695 57523
rect 707729 57513 707769 57523
rect 707803 57513 707840 57523
rect 707874 57513 707914 57523
rect 707948 57513 707985 57523
rect 708019 57513 708059 57523
rect 708093 57513 708130 57523
rect 708164 57513 708204 57523
rect 708238 57513 708275 57523
rect 708309 57513 708369 57523
rect 708403 57513 708446 57523
rect 708480 57513 708522 57523
rect 708556 57513 708604 57523
rect 709219 57513 709270 57523
rect 709304 57513 709364 57523
rect 709398 57513 709435 57523
rect 709469 57513 709509 57523
rect 709543 57513 709580 57523
rect 709614 57513 709654 57523
rect 709688 57513 709725 57523
rect 709759 57513 709799 57523
rect 709833 57513 709870 57523
rect 709904 57513 709944 57523
rect 709978 57513 710015 57523
rect 710049 57513 710089 57523
rect 710123 57513 710160 57523
rect 710194 57513 710211 57523
rect 684070 57443 684670 57499
rect 685537 57443 686137 57493
rect 692428 57442 693028 57492
rect 680215 57348 680815 57398
rect 681713 57359 682313 57409
rect 684070 57293 684670 57343
rect 692428 57292 693028 57342
rect 705107 57336 705173 57352
rect 711579 57301 711595 58520
rect 711892 57697 711942 58520
rect 712062 57697 712112 58520
rect 716071 58357 716074 58358
rect 714645 58323 714752 58357
rect 716071 58356 716072 58357
rect 716073 58356 716074 58357
rect 716071 58355 716074 58356
rect 716208 58357 716211 58358
rect 716208 58356 716209 58357
rect 716210 58356 716211 58357
rect 716208 58355 716211 58356
rect 714964 58247 715998 58329
rect 716284 58247 717318 58329
rect 714175 57398 714225 57998
rect 714425 57398 714475 57998
rect 680215 57232 680815 57282
rect 698017 57232 698053 57260
rect 692428 57162 693028 57212
rect 698030 57198 698077 57232
rect 698017 57164 698053 57198
rect 680215 57056 680815 57112
rect 692428 57006 693028 57134
rect 698030 57130 698077 57164
rect 698017 57096 698053 57130
rect 698030 57062 698077 57096
rect 698017 56983 698053 57062
rect 698084 56983 698120 57260
rect 714781 57191 714863 58226
rect 715134 57955 715828 58037
rect 714686 57123 714863 57191
rect 714645 57089 714863 57123
rect 680215 56880 680815 56936
rect 686719 56893 686739 56917
rect 686743 56893 686753 56917
rect 686719 56859 686757 56893
rect 686719 56822 686739 56859
rect 686743 56822 686753 56859
rect 692428 56850 693028 56978
rect 698017 56947 698210 56983
rect 698084 56935 698210 56947
rect 702756 56959 703645 56983
rect 702756 56935 702853 56959
rect 698084 56828 702853 56935
rect 686719 56788 686757 56822
rect 680215 56704 680815 56760
rect 686719 56751 686739 56788
rect 686743 56751 686753 56788
rect 686719 56741 686757 56751
rect 686699 56717 686767 56741
rect 686719 56704 686739 56717
rect 686743 56704 686753 56717
rect 686719 56695 686753 56704
rect 686719 56693 686743 56695
rect 692428 56694 693028 56750
rect 686685 56656 686709 56680
rect 686743 56656 686767 56680
rect 678799 56503 679399 56553
rect 680215 56534 680815 56584
rect 692428 56538 693028 56666
rect 680593 56531 680815 56534
rect 682009 56501 682069 56516
rect 682024 56465 682054 56501
rect 683708 56387 684308 56437
rect 678799 56327 679399 56383
rect 692428 56382 693028 56510
rect 714781 56308 714863 57089
rect 715063 56609 715145 57915
rect 715289 56777 715339 57719
rect 715633 56777 715683 57719
rect 715382 56672 715422 56756
rect 715542 56672 715582 56756
rect 715342 56632 715382 56672
rect 715582 56632 715622 56672
rect 715815 56609 715897 57915
rect 715134 56387 715828 56469
rect 716100 56308 716182 58226
rect 716454 57955 717148 58037
rect 716385 56609 716467 57915
rect 716599 56777 716649 57719
rect 716943 56777 716993 57719
rect 716700 56672 716740 56756
rect 716860 56672 716900 56756
rect 716660 56632 716700 56672
rect 716900 56632 716940 56672
rect 717137 56609 717219 57915
rect 716454 56387 717148 56469
rect 717419 56308 717501 58226
rect 683708 56237 684308 56287
rect 692428 56232 693028 56282
rect 678799 56157 679399 56207
rect 684565 56160 684790 56168
rect 696597 56000 696600 56120
rect 714964 56095 715998 56177
rect 716284 56095 717318 56177
rect 21000 41000 21003 41120
rect 696597 40200 696600 40320
rect 370961 38920 370987 38946
rect 470961 38920 470987 38946
rect 570961 38920 570987 38946
rect 69734 37993 69784 38593
rect 69904 37993 69954 38593
rect 71447 38201 71497 38801
rect 71617 38201 71673 38801
rect 71793 38201 71843 38801
rect 121734 37993 121784 38593
rect 121904 37993 121954 38593
rect 123447 38201 123497 38801
rect 123617 38201 123673 38801
rect 123793 38201 123843 38801
rect 173734 37993 173784 38593
rect 173904 37993 173954 38593
rect 175447 38201 175497 38801
rect 175617 38201 175673 38801
rect 175793 38201 175843 38801
rect 225734 37993 225784 38593
rect 225904 37993 225954 38593
rect 227447 38201 227497 38801
rect 227617 38201 227673 38801
rect 227793 38201 227843 38801
rect 273734 37993 273784 38593
rect 273904 37993 273954 38593
rect 275447 38201 275497 38801
rect 275617 38201 275673 38801
rect 275793 38201 275843 38801
rect 325734 37993 325784 38593
rect 325904 37993 325954 38593
rect 327447 38201 327497 38801
rect 327617 38201 327673 38801
rect 327793 38201 327843 38801
rect 366239 38085 366263 38109
rect 366215 38061 366238 38085
rect 366970 37993 367020 38593
rect 367140 37993 367190 38593
rect 367566 37998 367616 38598
rect 367736 37998 367792 38598
rect 367912 38539 367962 38598
rect 368654 38539 368704 38598
rect 367912 38467 367965 38539
rect 367912 38220 367962 38467
rect 368025 38317 368037 38467
rect 368651 38317 368704 38539
rect 368654 38220 368704 38317
rect 367912 38148 367965 38220
rect 367912 37998 367962 38148
rect 368025 37998 368037 38148
rect 368651 37998 368704 38220
rect 368824 37998 368880 38598
rect 369000 37998 369050 38598
rect 369426 37993 369476 38593
rect 369596 37993 369646 38593
rect 371124 37993 371174 38593
rect 371294 37993 371344 38593
rect 371720 37998 371770 38598
rect 371890 37998 371946 38598
rect 372066 38539 372116 38598
rect 372808 38539 372858 38598
rect 372066 38467 372119 38539
rect 372066 38220 372116 38467
rect 372179 38317 372191 38467
rect 372805 38317 372858 38539
rect 372808 38220 372858 38317
rect 372066 38148 372119 38220
rect 372066 37998 372116 38148
rect 372179 37998 372191 38148
rect 372805 37998 372858 38220
rect 372978 37998 373034 38598
rect 373154 37998 373204 38598
rect 373580 37993 373630 38593
rect 373750 37993 373800 38593
rect 375278 37993 375328 38593
rect 375448 37993 375498 38593
rect 375874 37998 375924 38598
rect 376044 37998 376100 38598
rect 376220 38539 376270 38598
rect 376962 38539 377012 38598
rect 376220 38467 376273 38539
rect 376220 38220 376270 38467
rect 376333 38317 376345 38467
rect 376959 38317 377012 38539
rect 376962 38220 377012 38317
rect 376220 38148 376273 38220
rect 376220 37998 376270 38148
rect 376333 37998 376345 38148
rect 376959 37998 377012 38220
rect 377132 37998 377188 38598
rect 377308 37998 377358 38598
rect 377734 37993 377784 38593
rect 377904 37993 377954 38593
rect 379447 38201 379497 38801
rect 379617 38201 379673 38801
rect 379793 38201 379843 38801
rect 425734 37993 425784 38593
rect 425904 37993 425954 38593
rect 427447 38201 427497 38801
rect 427617 38201 427673 38801
rect 427793 38201 427843 38801
rect 466239 38085 466263 38109
rect 466215 38061 466238 38085
rect 466970 37993 467020 38593
rect 467140 37993 467190 38593
rect 467566 37998 467616 38598
rect 467736 37998 467792 38598
rect 467912 38539 467962 38598
rect 468654 38539 468704 38598
rect 467912 38467 467965 38539
rect 467912 38220 467962 38467
rect 468025 38317 468037 38467
rect 468651 38317 468704 38539
rect 468654 38220 468704 38317
rect 467912 38148 467965 38220
rect 467912 37998 467962 38148
rect 468025 37998 468037 38148
rect 468651 37998 468704 38220
rect 468824 37998 468880 38598
rect 469000 37998 469050 38598
rect 469426 37993 469476 38593
rect 469596 37993 469646 38593
rect 471124 37993 471174 38593
rect 471294 37993 471344 38593
rect 471720 37998 471770 38598
rect 471890 37998 471946 38598
rect 472066 38539 472116 38598
rect 472808 38539 472858 38598
rect 472066 38467 472119 38539
rect 472066 38220 472116 38467
rect 472179 38317 472191 38467
rect 472805 38317 472858 38539
rect 472808 38220 472858 38317
rect 472066 38148 472119 38220
rect 472066 37998 472116 38148
rect 472179 37998 472191 38148
rect 472805 37998 472858 38220
rect 472978 37998 473034 38598
rect 473154 37998 473204 38598
rect 473580 37993 473630 38593
rect 473750 37993 473800 38593
rect 475278 37993 475328 38593
rect 475448 37993 475498 38593
rect 475874 37998 475924 38598
rect 476044 37998 476100 38598
rect 476220 38539 476270 38598
rect 476962 38539 477012 38598
rect 476220 38467 476273 38539
rect 476220 38220 476270 38467
rect 476333 38317 476345 38467
rect 476959 38317 477012 38539
rect 476962 38220 477012 38317
rect 476220 38148 476273 38220
rect 476220 37998 476270 38148
rect 476333 37998 476345 38148
rect 476959 37998 477012 38220
rect 477132 37998 477188 38598
rect 477308 37998 477358 38598
rect 477734 37993 477784 38593
rect 477904 37993 477954 38593
rect 479447 38201 479497 38801
rect 479617 38201 479673 38801
rect 479793 38201 479843 38801
rect 529734 37993 529784 38593
rect 529904 37993 529954 38593
rect 531447 38201 531497 38801
rect 531617 38201 531673 38801
rect 531793 38201 531843 38801
rect 566239 38085 566263 38109
rect 566215 38061 566238 38085
rect 566970 37993 567020 38593
rect 567140 37993 567190 38593
rect 567566 37998 567616 38598
rect 567736 37998 567792 38598
rect 567912 38539 567962 38598
rect 568654 38539 568704 38598
rect 567912 38467 567965 38539
rect 567912 38220 567962 38467
rect 568025 38317 568037 38467
rect 568651 38317 568704 38539
rect 568654 38220 568704 38317
rect 567912 38148 567965 38220
rect 567912 37998 567962 38148
rect 568025 37998 568037 38148
rect 568651 37998 568704 38220
rect 568824 37998 568880 38598
rect 569000 37998 569050 38598
rect 569426 37993 569476 38593
rect 569596 37993 569646 38593
rect 571124 37993 571174 38593
rect 571294 37993 571344 38593
rect 571720 37998 571770 38598
rect 571890 37998 571946 38598
rect 572066 38539 572116 38598
rect 572808 38539 572858 38598
rect 572066 38467 572119 38539
rect 572066 38220 572116 38467
rect 572179 38317 572191 38467
rect 572805 38317 572858 38539
rect 572808 38220 572858 38317
rect 572066 38148 572119 38220
rect 572066 37998 572116 38148
rect 572179 37998 572191 38148
rect 572805 37998 572858 38220
rect 572978 37998 573034 38598
rect 573154 37998 573204 38598
rect 573580 37993 573630 38593
rect 573750 37993 573800 38593
rect 575278 37993 575328 38593
rect 575448 37993 575498 38593
rect 575874 37998 575924 38598
rect 576044 37998 576100 38598
rect 576220 38539 576270 38598
rect 576962 38539 577012 38598
rect 576220 38467 576273 38539
rect 576220 38220 576270 38467
rect 576333 38317 576345 38467
rect 576959 38317 577012 38539
rect 576962 38220 577012 38317
rect 576220 38148 576273 38220
rect 576220 37998 576270 38148
rect 576333 37998 576345 38148
rect 576959 37998 577012 38220
rect 577132 37998 577188 38598
rect 577308 37998 577358 38598
rect 577734 37993 577784 38593
rect 577904 37993 577954 38593
rect 579447 38201 579497 38801
rect 579617 38201 579673 38801
rect 579793 38201 579843 38801
rect 366215 37963 366238 37987
rect 466215 37963 466238 37987
rect 566215 37963 566238 37987
rect 366239 37939 366263 37963
rect 466239 37939 466263 37963
rect 566239 37939 566263 37963
rect 365670 37792 365694 37807
rect 366043 37792 366067 37807
rect 465670 37792 465694 37807
rect 466043 37792 466067 37807
rect 565670 37792 565694 37807
rect 566043 37792 566067 37807
rect 365646 37759 365670 37783
rect 366067 37759 366091 37783
rect 465646 37759 465670 37783
rect 466067 37759 466091 37783
rect 565646 37759 565670 37783
rect 566067 37759 566091 37783
rect 58272 36785 58322 37385
rect 58442 36785 58498 37385
rect 69480 37083 69573 37120
rect 69480 36785 69573 36985
rect 69629 36785 69809 36985
rect 70080 36785 70130 37385
rect 70250 36785 70306 37385
rect 70426 36785 70482 37385
rect 70602 36785 70652 37385
rect 70718 36785 70768 37385
rect 70888 36785 70944 37385
rect 71064 36785 71120 37385
rect 71240 36785 71296 37385
rect 71416 37007 71466 37385
rect 71416 36935 71469 37007
rect 71416 36785 71466 36935
rect 71529 36785 71541 36935
rect 110272 36785 110322 37385
rect 110442 36785 110498 37385
rect 121480 37083 121573 37120
rect 121480 36785 121573 36985
rect 121629 36785 121809 36985
rect 122080 36785 122130 37385
rect 122250 36785 122306 37385
rect 122426 36785 122482 37385
rect 122602 36785 122652 37385
rect 122718 36785 122768 37385
rect 122888 36785 122944 37385
rect 123064 36785 123120 37385
rect 123240 36785 123296 37385
rect 123416 37007 123466 37385
rect 173480 37083 173573 37120
rect 123416 36935 123469 37007
rect 123416 36785 123466 36935
rect 123529 36785 123541 36935
rect 173480 36785 173573 36985
rect 173629 36785 173809 36985
rect 174080 36785 174130 37385
rect 174250 36785 174306 37385
rect 174426 36785 174482 37385
rect 174602 36785 174652 37385
rect 174718 36785 174768 37385
rect 174888 36785 174944 37385
rect 175064 36785 175120 37385
rect 175240 36785 175296 37385
rect 175416 37007 175466 37385
rect 175416 36935 175469 37007
rect 175416 36785 175466 36935
rect 175529 36785 175541 36935
rect 214272 36785 214322 37385
rect 214442 36785 214498 37385
rect 225480 37083 225573 37120
rect 225480 36785 225573 36985
rect 225629 36785 225809 36985
rect 226080 36785 226130 37385
rect 226250 36785 226306 37385
rect 226426 36785 226482 37385
rect 226602 36785 226652 37385
rect 226718 36785 226768 37385
rect 226888 36785 226944 37385
rect 227064 36785 227120 37385
rect 227240 36785 227296 37385
rect 227416 37007 227466 37385
rect 273480 37083 273573 37120
rect 227416 36935 227469 37007
rect 227416 36785 227466 36935
rect 227529 36785 227541 36935
rect 273480 36785 273573 36985
rect 273629 36785 273809 36985
rect 274080 36785 274130 37385
rect 274250 36785 274306 37385
rect 274426 36785 274482 37385
rect 274602 36785 274652 37385
rect 274718 36785 274768 37385
rect 274888 36785 274944 37385
rect 275064 36785 275120 37385
rect 275240 36785 275296 37385
rect 275416 37007 275466 37385
rect 275416 36935 275469 37007
rect 275416 36785 275466 36935
rect 275529 36785 275541 36935
rect 314272 36785 314322 37385
rect 314442 36785 314498 37385
rect 325480 37083 325573 37120
rect 325480 36785 325573 36985
rect 325629 36785 325809 36985
rect 326080 36785 326130 37385
rect 326250 36785 326306 37385
rect 326426 36785 326482 37385
rect 326602 36785 326652 37385
rect 326718 36785 326768 37385
rect 326888 36785 326944 37385
rect 327064 36785 327120 37385
rect 327240 36785 327296 37385
rect 327416 37007 327466 37385
rect 327416 36935 327469 37007
rect 327416 36785 327466 36935
rect 327529 36785 327541 36935
rect 366272 36785 366322 37385
rect 366442 36785 366498 37385
rect 366618 36785 366674 37385
rect 366794 36785 366844 37385
rect 367351 37098 367531 37120
rect 369085 37098 369265 37120
rect 367336 37083 367546 37098
rect 369070 37083 369280 37098
rect 367100 36970 367310 36985
rect 367336 36970 367546 36985
rect 369070 36970 369280 36985
rect 369306 36970 369516 36985
rect 367115 36800 367295 36970
rect 367351 36800 367531 36970
rect 369085 36800 369265 36970
rect 369321 36800 369501 36970
rect 367104 36797 367306 36800
rect 367340 36797 367542 36800
rect 369074 36797 369276 36800
rect 369310 36797 369512 36800
rect 367100 36785 367310 36797
rect 367336 36785 367546 36797
rect 369070 36785 369280 36797
rect 369306 36785 369516 36797
rect 369772 36785 369822 37385
rect 369942 36785 369998 37385
rect 370118 36785 370174 37385
rect 370294 36785 370344 37385
rect 370426 36785 370476 37385
rect 370596 36785 370652 37385
rect 370772 36785 370828 37385
rect 370948 36785 370998 37385
rect 371505 37098 371685 37120
rect 373239 37098 373419 37120
rect 371490 37083 371700 37098
rect 373224 37083 373434 37098
rect 371254 36970 371464 36985
rect 371490 36970 371700 36985
rect 373224 36970 373434 36985
rect 373460 36970 373670 36985
rect 371269 36800 371449 36970
rect 371505 36800 371685 36970
rect 373239 36800 373419 36970
rect 373475 36800 373655 36970
rect 371258 36797 371460 36800
rect 371494 36797 371696 36800
rect 373228 36797 373430 36800
rect 373464 36797 373666 36800
rect 371254 36785 371464 36797
rect 371490 36785 371700 36797
rect 373224 36785 373434 36797
rect 373460 36785 373670 36797
rect 373926 36785 373976 37385
rect 374096 36785 374152 37385
rect 374272 36785 374328 37385
rect 374448 36785 374498 37385
rect 374580 36785 374630 37385
rect 374750 36785 374806 37385
rect 374926 36785 374982 37385
rect 375102 36785 375152 37385
rect 375659 37098 375839 37120
rect 377393 37098 377573 37120
rect 375644 37083 375854 37098
rect 377378 37083 377588 37098
rect 375408 36970 375618 36985
rect 375644 36970 375854 36985
rect 377378 36970 377588 36985
rect 377614 36970 377824 36985
rect 375423 36800 375603 36970
rect 375659 36800 375839 36970
rect 377393 36800 377573 36970
rect 377629 36800 377809 36970
rect 375412 36797 375614 36800
rect 375648 36797 375850 36800
rect 377382 36797 377584 36800
rect 377618 36797 377820 36800
rect 375408 36785 375618 36797
rect 375644 36785 375854 36797
rect 377378 36785 377588 36797
rect 377614 36785 377824 36797
rect 378080 36785 378130 37385
rect 378250 36785 378306 37385
rect 378426 36785 378482 37385
rect 378602 36785 378652 37385
rect 378718 36785 378768 37385
rect 378888 36785 378944 37385
rect 379064 36785 379120 37385
rect 379240 36785 379296 37385
rect 379416 37007 379466 37385
rect 379416 36935 379469 37007
rect 379416 36785 379466 36935
rect 379529 36785 379541 36935
rect 414272 36785 414322 37385
rect 414442 36785 414498 37385
rect 425480 37083 425573 37120
rect 425480 36785 425573 36985
rect 425629 36785 425809 36985
rect 426080 36785 426130 37385
rect 426250 36785 426306 37385
rect 426426 36785 426482 37385
rect 426602 36785 426652 37385
rect 426718 36785 426768 37385
rect 426888 36785 426944 37385
rect 427064 36785 427120 37385
rect 427240 36785 427296 37385
rect 427416 37007 427466 37385
rect 427416 36935 427469 37007
rect 427416 36785 427466 36935
rect 427529 36785 427541 36935
rect 466272 36785 466322 37385
rect 466442 36785 466498 37385
rect 466618 36785 466674 37385
rect 466794 36785 466844 37385
rect 467351 37098 467531 37120
rect 469085 37098 469265 37120
rect 467336 37083 467546 37098
rect 469070 37083 469280 37098
rect 467100 36970 467310 36985
rect 467336 36970 467546 36985
rect 469070 36970 469280 36985
rect 469306 36970 469516 36985
rect 467115 36800 467295 36970
rect 467351 36800 467531 36970
rect 469085 36800 469265 36970
rect 469321 36800 469501 36970
rect 467104 36797 467306 36800
rect 467340 36797 467542 36800
rect 469074 36797 469276 36800
rect 469310 36797 469512 36800
rect 467100 36785 467310 36797
rect 467336 36785 467546 36797
rect 469070 36785 469280 36797
rect 469306 36785 469516 36797
rect 469772 36785 469822 37385
rect 469942 36785 469998 37385
rect 470118 36785 470174 37385
rect 470294 36785 470344 37385
rect 470426 36785 470476 37385
rect 470596 36785 470652 37385
rect 470772 36785 470828 37385
rect 470948 36785 470998 37385
rect 471505 37098 471685 37120
rect 473239 37098 473419 37120
rect 471490 37083 471700 37098
rect 473224 37083 473434 37098
rect 471254 36970 471464 36985
rect 471490 36970 471700 36985
rect 473224 36970 473434 36985
rect 473460 36970 473670 36985
rect 471269 36800 471449 36970
rect 471505 36800 471685 36970
rect 473239 36800 473419 36970
rect 473475 36800 473655 36970
rect 471258 36797 471460 36800
rect 471494 36797 471696 36800
rect 473228 36797 473430 36800
rect 473464 36797 473666 36800
rect 471254 36785 471464 36797
rect 471490 36785 471700 36797
rect 473224 36785 473434 36797
rect 473460 36785 473670 36797
rect 473926 36785 473976 37385
rect 474096 36785 474152 37385
rect 474272 36785 474328 37385
rect 474448 36785 474498 37385
rect 474580 36785 474630 37385
rect 474750 36785 474806 37385
rect 474926 36785 474982 37385
rect 475102 36785 475152 37385
rect 475659 37098 475839 37120
rect 477393 37098 477573 37120
rect 475644 37083 475854 37098
rect 477378 37083 477588 37098
rect 475408 36970 475618 36985
rect 475644 36970 475854 36985
rect 477378 36970 477588 36985
rect 477614 36970 477824 36985
rect 475423 36800 475603 36970
rect 475659 36800 475839 36970
rect 477393 36800 477573 36970
rect 477629 36800 477809 36970
rect 475412 36797 475614 36800
rect 475648 36797 475850 36800
rect 477382 36797 477584 36800
rect 477618 36797 477820 36800
rect 475408 36785 475618 36797
rect 475644 36785 475854 36797
rect 477378 36785 477588 36797
rect 477614 36785 477824 36797
rect 478080 36785 478130 37385
rect 478250 36785 478306 37385
rect 478426 36785 478482 37385
rect 478602 36785 478652 37385
rect 478718 36785 478768 37385
rect 478888 36785 478944 37385
rect 479064 36785 479120 37385
rect 479240 36785 479296 37385
rect 479416 37007 479466 37385
rect 479416 36935 479469 37007
rect 479416 36785 479466 36935
rect 479529 36785 479541 36935
rect 518272 36785 518322 37385
rect 518442 36785 518498 37385
rect 529480 37083 529573 37120
rect 529480 36785 529573 36985
rect 529629 36785 529809 36985
rect 530080 36785 530130 37385
rect 530250 36785 530306 37385
rect 530426 36785 530482 37385
rect 530602 36785 530652 37385
rect 530718 36785 530768 37385
rect 530888 36785 530944 37385
rect 531064 36785 531120 37385
rect 531240 36785 531296 37385
rect 531416 37007 531466 37385
rect 531416 36935 531469 37007
rect 531416 36785 531466 36935
rect 531529 36785 531541 36935
rect 566272 36785 566322 37385
rect 566442 36785 566498 37385
rect 566618 36785 566674 37385
rect 566794 36785 566844 37385
rect 567351 37098 567531 37120
rect 569085 37098 569265 37120
rect 567336 37083 567546 37098
rect 569070 37083 569280 37098
rect 567100 36970 567310 36985
rect 567336 36970 567546 36985
rect 569070 36970 569280 36985
rect 569306 36970 569516 36985
rect 567115 36800 567295 36970
rect 567351 36800 567531 36970
rect 569085 36800 569265 36970
rect 569321 36800 569501 36970
rect 567104 36797 567306 36800
rect 567340 36797 567542 36800
rect 569074 36797 569276 36800
rect 569310 36797 569512 36800
rect 567100 36785 567310 36797
rect 567336 36785 567546 36797
rect 569070 36785 569280 36797
rect 569306 36785 569516 36797
rect 569772 36785 569822 37385
rect 569942 36785 569998 37385
rect 570118 36785 570174 37385
rect 570294 36785 570344 37385
rect 570426 36785 570476 37385
rect 570596 36785 570652 37385
rect 570772 36785 570828 37385
rect 570948 36785 570998 37385
rect 571505 37098 571685 37120
rect 573239 37098 573419 37120
rect 571490 37083 571700 37098
rect 573224 37083 573434 37098
rect 571254 36970 571464 36985
rect 571490 36970 571700 36985
rect 573224 36970 573434 36985
rect 573460 36970 573670 36985
rect 571269 36800 571449 36970
rect 571505 36800 571685 36970
rect 573239 36800 573419 36970
rect 573475 36800 573655 36970
rect 571258 36797 571460 36800
rect 571494 36797 571696 36800
rect 573228 36797 573430 36800
rect 573464 36797 573666 36800
rect 571254 36785 571464 36797
rect 571490 36785 571700 36797
rect 573224 36785 573434 36797
rect 573460 36785 573670 36797
rect 573926 36785 573976 37385
rect 574096 36785 574152 37385
rect 574272 36785 574328 37385
rect 574448 36785 574498 37385
rect 574580 36785 574630 37385
rect 574750 36785 574806 37385
rect 574926 36785 574982 37385
rect 575102 36785 575152 37385
rect 575659 37098 575839 37120
rect 577393 37098 577573 37120
rect 575644 37083 575854 37098
rect 577378 37083 577588 37098
rect 575408 36970 575618 36985
rect 575644 36970 575854 36985
rect 577378 36970 577588 36985
rect 577614 36970 577824 36985
rect 575423 36800 575603 36970
rect 575659 36800 575839 36970
rect 577393 36800 577573 36970
rect 577629 36800 577809 36970
rect 575412 36797 575614 36800
rect 575648 36797 575850 36800
rect 577382 36797 577584 36800
rect 577618 36797 577820 36800
rect 575408 36785 575618 36797
rect 575644 36785 575854 36797
rect 577378 36785 577588 36797
rect 577614 36785 577824 36797
rect 578080 36785 578130 37385
rect 578250 36785 578306 37385
rect 578426 36785 578482 37385
rect 578602 36785 578652 37385
rect 578718 36785 578768 37385
rect 578888 36785 578944 37385
rect 579064 36785 579120 37385
rect 579240 36785 579296 37385
rect 579416 37007 579466 37385
rect 579416 36935 579469 37007
rect 579416 36785 579466 36935
rect 579529 36785 579541 36935
rect 70069 35287 70119 35887
rect 70239 35287 70295 35887
rect 70591 35287 70641 35887
rect 71484 35576 71499 35591
rect 71484 35546 71535 35576
rect 71484 35531 71499 35546
rect 122069 35287 122119 35887
rect 122239 35287 122295 35887
rect 122591 35287 122641 35887
rect 123484 35576 123499 35591
rect 123484 35546 123535 35576
rect 123484 35531 123499 35546
rect 174069 35287 174119 35887
rect 174239 35287 174295 35887
rect 174591 35287 174641 35887
rect 175484 35576 175499 35591
rect 175484 35546 175535 35576
rect 175484 35531 175499 35546
rect 226069 35287 226119 35887
rect 226239 35287 226295 35887
rect 226591 35287 226641 35887
rect 227484 35576 227499 35591
rect 227484 35546 227535 35576
rect 227484 35531 227499 35546
rect 274069 35287 274119 35887
rect 274239 35287 274295 35887
rect 274591 35287 274641 35887
rect 275484 35576 275499 35591
rect 275484 35546 275535 35576
rect 275484 35531 275499 35546
rect 326069 35287 326119 35887
rect 326239 35287 326295 35887
rect 326591 35287 326641 35887
rect 327484 35576 327499 35591
rect 327484 35546 327535 35576
rect 327484 35531 327499 35546
rect 368869 35255 368919 35855
rect 369019 35255 369075 35855
rect 369175 35255 369303 35855
rect 369331 35255 369459 35855
rect 369487 35255 369537 35855
rect 369741 35255 369791 35855
rect 369891 35255 370019 35855
rect 370047 35255 370103 35855
rect 370203 35255 370331 35855
rect 370359 35255 370409 35855
rect 370561 35255 370611 35855
rect 370731 35255 370859 35855
rect 370907 35255 370963 35855
rect 371083 35255 371133 35855
rect 371299 35255 371349 36255
rect 371469 35255 371525 36255
rect 371645 35255 371773 36255
rect 371821 35255 371871 36255
rect 371954 35255 371966 36255
rect 372023 35255 372073 36255
rect 372193 35255 372321 36255
rect 372369 35255 372497 36255
rect 372545 35255 372601 36255
rect 372721 35255 372771 36255
rect 372870 36143 372936 36159
rect 373032 36143 373098 36159
rect 373194 36143 373260 36159
rect 373356 36143 373422 36159
rect 372870 35359 372936 35375
rect 373356 35359 373422 35375
rect 373521 35255 373571 36255
rect 373691 35255 373747 36255
rect 373867 35255 373995 36255
rect 374043 35255 374171 36255
rect 374219 35255 374269 36255
rect 374326 35255 374338 36255
rect 374362 36176 374372 36210
rect 374362 36108 374372 36142
rect 374362 36040 374372 36074
rect 374362 35972 374372 36006
rect 374362 35904 374372 35938
rect 374362 35836 374372 35870
rect 374362 35768 374372 35802
rect 374362 35700 374372 35734
rect 374362 35632 374372 35666
rect 374362 35564 374372 35598
rect 374362 35489 374372 35523
rect 374362 35421 374372 35455
rect 374362 35353 374372 35387
rect 374362 35285 374372 35319
rect 374539 35134 374589 36134
rect 374689 35134 374817 36134
rect 374845 35806 374895 36134
rect 375005 36071 375495 36098
rect 377994 35887 378006 35936
rect 374845 35794 374898 35806
rect 374838 35734 374898 35794
rect 378066 35788 378119 35887
rect 374845 35134 374895 35734
rect 374898 35134 374970 35734
rect 375048 35134 375176 35734
rect 375204 35134 375332 35734
rect 375360 35134 375488 35734
rect 375516 35134 375566 35734
rect 375632 35134 375682 35734
rect 375782 35559 375832 35734
rect 378069 35559 378119 35788
rect 375782 35487 375835 35559
rect 375782 35134 375832 35487
rect 375895 35287 375907 35487
rect 378066 35287 378119 35559
rect 378239 35287 378295 35887
rect 378415 35287 378543 35887
rect 378591 35287 378641 35887
rect 379484 35576 379499 35591
rect 379484 35546 379535 35576
rect 379484 35531 379499 35546
rect 426069 35287 426119 35887
rect 426239 35287 426295 35887
rect 426591 35287 426641 35887
rect 427484 35576 427499 35591
rect 427484 35546 427535 35576
rect 427484 35531 427499 35546
rect 468869 35255 468919 35855
rect 469019 35255 469075 35855
rect 469175 35255 469303 35855
rect 469331 35255 469459 35855
rect 469487 35255 469537 35855
rect 469741 35255 469791 35855
rect 469891 35255 470019 35855
rect 470047 35255 470103 35855
rect 470203 35255 470331 35855
rect 470359 35255 470409 35855
rect 470561 35255 470611 35855
rect 470731 35255 470859 35855
rect 470907 35255 470963 35855
rect 471083 35255 471133 35855
rect 471299 35255 471349 36255
rect 471469 35255 471525 36255
rect 471645 35255 471773 36255
rect 471821 35255 471871 36255
rect 471954 35255 471966 36255
rect 472023 35255 472073 36255
rect 472193 35255 472321 36255
rect 472369 35255 472497 36255
rect 472545 35255 472601 36255
rect 472721 35255 472771 36255
rect 472870 36143 472936 36159
rect 473032 36143 473098 36159
rect 473194 36143 473260 36159
rect 473356 36143 473422 36159
rect 472870 35359 472936 35375
rect 473356 35359 473422 35375
rect 473521 35255 473571 36255
rect 473691 35255 473747 36255
rect 473867 35255 473995 36255
rect 474043 35255 474171 36255
rect 474219 35255 474269 36255
rect 474326 35255 474338 36255
rect 474362 36176 474372 36210
rect 474362 36108 474372 36142
rect 474362 36040 474372 36074
rect 474362 35972 474372 36006
rect 474362 35904 474372 35938
rect 474362 35836 474372 35870
rect 474362 35768 474372 35802
rect 474362 35700 474372 35734
rect 474362 35632 474372 35666
rect 474362 35564 474372 35598
rect 474362 35489 474372 35523
rect 474362 35421 474372 35455
rect 474362 35353 474372 35387
rect 474362 35285 474372 35319
rect 474539 35134 474589 36134
rect 474689 35134 474817 36134
rect 474845 35806 474895 36134
rect 475005 36071 475495 36098
rect 477994 35887 478006 35936
rect 474845 35794 474898 35806
rect 474838 35734 474898 35794
rect 478066 35788 478119 35887
rect 474845 35134 474895 35734
rect 474898 35134 474970 35734
rect 475048 35134 475176 35734
rect 475204 35134 475332 35734
rect 475360 35134 475488 35734
rect 475516 35134 475566 35734
rect 475632 35134 475682 35734
rect 475782 35559 475832 35734
rect 478069 35559 478119 35788
rect 475782 35487 475835 35559
rect 475782 35134 475832 35487
rect 475895 35287 475907 35487
rect 478066 35287 478119 35559
rect 478239 35287 478295 35887
rect 478415 35287 478543 35887
rect 478591 35287 478641 35887
rect 479484 35576 479499 35591
rect 479484 35546 479535 35576
rect 479484 35531 479499 35546
rect 530069 35287 530119 35887
rect 530239 35287 530295 35887
rect 530591 35287 530641 35887
rect 531484 35576 531499 35591
rect 531484 35546 531535 35576
rect 531484 35531 531499 35546
rect 568869 35255 568919 35855
rect 569019 35255 569075 35855
rect 569175 35255 569303 35855
rect 569331 35255 569459 35855
rect 569487 35255 569537 35855
rect 569741 35255 569791 35855
rect 569891 35255 570019 35855
rect 570047 35255 570103 35855
rect 570203 35255 570331 35855
rect 570359 35255 570409 35855
rect 570561 35255 570611 35855
rect 570731 35255 570859 35855
rect 570907 35255 570963 35855
rect 571083 35255 571133 35855
rect 571299 35255 571349 36255
rect 571469 35255 571525 36255
rect 571645 35255 571773 36255
rect 571821 35255 571871 36255
rect 571954 35255 571966 36255
rect 572023 35255 572073 36255
rect 572193 35255 572321 36255
rect 572369 35255 572497 36255
rect 572545 35255 572601 36255
rect 572721 35255 572771 36255
rect 572870 36143 572936 36159
rect 573032 36143 573098 36159
rect 573194 36143 573260 36159
rect 573356 36143 573422 36159
rect 572870 35359 572936 35375
rect 573356 35359 573422 35375
rect 573521 35255 573571 36255
rect 573691 35255 573747 36255
rect 573867 35255 573995 36255
rect 574043 35255 574171 36255
rect 574219 35255 574269 36255
rect 574326 35255 574338 36255
rect 574362 36176 574372 36210
rect 574362 36108 574372 36142
rect 574362 36040 574372 36074
rect 574362 35972 574372 36006
rect 574362 35904 574372 35938
rect 574362 35836 574372 35870
rect 574362 35768 574372 35802
rect 574362 35700 574372 35734
rect 574362 35632 574372 35666
rect 574362 35564 574372 35598
rect 574362 35489 574372 35523
rect 574362 35421 574372 35455
rect 574362 35353 574372 35387
rect 574362 35285 574372 35319
rect 574539 35134 574589 36134
rect 574689 35134 574817 36134
rect 574845 35806 574895 36134
rect 575005 36071 575495 36098
rect 577994 35887 578006 35936
rect 574845 35794 574898 35806
rect 574838 35734 574898 35794
rect 578066 35788 578119 35887
rect 574845 35134 574895 35734
rect 574898 35134 574970 35734
rect 575048 35134 575176 35734
rect 575204 35134 575332 35734
rect 575360 35134 575488 35734
rect 575516 35134 575566 35734
rect 575632 35134 575682 35734
rect 575782 35559 575832 35734
rect 578069 35559 578119 35788
rect 575782 35487 575835 35559
rect 575782 35134 575832 35487
rect 575895 35287 575907 35487
rect 578066 35287 578119 35559
rect 578239 35287 578295 35887
rect 578415 35287 578543 35887
rect 578591 35287 578641 35887
rect 579484 35576 579499 35591
rect 579484 35546 579535 35576
rect 579484 35531 579499 35546
rect 69789 34110 69839 34710
rect 70051 34079 70101 34679
rect 70201 34079 70257 34679
rect 70357 34079 70407 34679
rect 121789 34110 121839 34710
rect 122051 34079 122101 34679
rect 122201 34079 122257 34679
rect 122357 34079 122407 34679
rect 173789 34110 173839 34710
rect 174051 34079 174101 34679
rect 174201 34079 174257 34679
rect 174357 34079 174407 34679
rect 225789 34110 225839 34710
rect 226051 34079 226101 34679
rect 226201 34079 226257 34679
rect 226357 34079 226407 34679
rect 273789 34110 273839 34710
rect 274051 34079 274101 34679
rect 274201 34079 274257 34679
rect 274357 34079 274407 34679
rect 325789 34110 325839 34710
rect 326051 34079 326101 34679
rect 326201 34079 326257 34679
rect 326357 34079 326407 34679
rect 367233 34427 367283 35027
rect 367403 34427 367531 35027
rect 367579 34427 367635 35027
rect 367755 34427 367883 35027
rect 367931 34427 368059 35027
rect 368107 34427 368235 35027
rect 368283 34427 368411 35027
rect 368459 34427 368509 35027
rect 368881 34491 368931 35091
rect 369051 34491 369179 35091
rect 369227 34491 369283 35091
rect 369403 34491 369531 35091
rect 369579 34491 369629 35091
rect 369920 34491 369970 35091
rect 370090 34491 370146 35091
rect 370266 34491 370316 35091
rect 369732 34302 370332 34352
rect 370395 34302 370445 35091
rect 69707 32596 69757 33596
rect 69823 32596 69873 33596
rect 69973 32596 70029 33596
rect 70129 32596 70179 33596
rect 70351 32930 70401 33530
rect 70501 32930 70557 33530
rect 70657 32930 70707 33530
rect 71563 33292 71613 33892
rect 71713 33292 71763 33892
rect 71862 32810 71870 33035
rect 121707 32596 121757 33596
rect 121823 32596 121873 33596
rect 121973 32596 122029 33596
rect 122129 32596 122179 33596
rect 122351 32930 122401 33530
rect 122501 32930 122557 33530
rect 122657 32930 122707 33530
rect 123563 33292 123613 33892
rect 123713 33292 123763 33892
rect 123862 32810 123870 33035
rect 173707 32596 173757 33596
rect 173823 32596 173873 33596
rect 173973 32596 174029 33596
rect 174129 32596 174179 33596
rect 174351 32930 174401 33530
rect 174501 32930 174557 33530
rect 174657 32930 174707 33530
rect 175563 33292 175613 33892
rect 175713 33292 175763 33892
rect 175862 32810 175870 33035
rect 225707 32596 225757 33596
rect 225823 32596 225873 33596
rect 225973 32596 226029 33596
rect 226129 32596 226179 33596
rect 226351 32930 226401 33530
rect 226501 32930 226557 33530
rect 226657 32930 226707 33530
rect 227563 33292 227613 33892
rect 227713 33292 227763 33892
rect 227862 32810 227870 33035
rect 273707 32596 273757 33596
rect 273823 32596 273873 33596
rect 273973 32596 274029 33596
rect 274129 32596 274179 33596
rect 274351 32930 274401 33530
rect 274501 32930 274557 33530
rect 274657 32930 274707 33530
rect 275563 33292 275613 33892
rect 275713 33292 275763 33892
rect 275862 32810 275870 33035
rect 325707 32596 325757 33596
rect 325823 32596 325873 33596
rect 325973 32596 326029 33596
rect 326129 32596 326179 33596
rect 326351 32930 326401 33530
rect 326501 32930 326557 33530
rect 326657 32930 326707 33530
rect 327563 33292 327613 33892
rect 327713 33292 327763 33892
rect 367157 33672 367207 34272
rect 367327 33672 367455 34272
rect 367503 33672 367559 34272
rect 367679 33672 367735 34272
rect 367855 33672 367911 34272
rect 368031 33672 368159 34272
rect 368207 33672 368263 34272
rect 368383 33672 368433 34272
rect 370392 34202 370445 34302
rect 369732 34152 370332 34202
rect 370395 34101 370445 34202
rect 370392 34091 370445 34101
rect 370565 34101 370615 35091
rect 370703 34491 370753 35091
rect 370873 34491 370929 35091
rect 371049 34491 371099 35091
rect 371319 34492 371369 35092
rect 371489 34492 371545 35092
rect 371665 34492 371715 35092
rect 370678 34322 371678 34372
rect 370678 34202 370690 34322
rect 370678 34152 371678 34202
rect 374611 34110 374661 34710
rect 374761 34110 374889 34710
rect 374917 34110 374973 34710
rect 375073 34110 375201 34710
rect 375229 34110 375279 34710
rect 375345 34110 375395 34710
rect 375495 34110 375551 34710
rect 375651 34110 375707 34710
rect 375807 34110 375863 34710
rect 375963 34110 376091 34710
rect 376119 34110 376247 34710
rect 376275 34110 376403 34710
rect 376431 34110 376487 34710
rect 376587 34110 376715 34710
rect 376743 34110 376871 34710
rect 376899 34110 377027 34710
rect 377055 34110 377105 34710
rect 377171 34110 377221 34710
rect 377321 34110 377449 34710
rect 377477 34110 377605 34710
rect 377633 34110 377761 34710
rect 377789 34110 377839 34710
rect 370565 34091 370618 34101
rect 378051 34079 378101 34679
rect 378201 34079 378257 34679
rect 378357 34079 378407 34679
rect 425789 34110 425839 34710
rect 426051 34079 426101 34679
rect 426201 34079 426257 34679
rect 426357 34079 426407 34679
rect 467233 34427 467283 35027
rect 467403 34427 467531 35027
rect 467579 34427 467635 35027
rect 467755 34427 467883 35027
rect 467931 34427 468059 35027
rect 468107 34427 468235 35027
rect 468283 34427 468411 35027
rect 468459 34427 468509 35027
rect 468881 34491 468931 35091
rect 469051 34491 469179 35091
rect 469227 34491 469283 35091
rect 469403 34491 469531 35091
rect 469579 34491 469629 35091
rect 469920 34491 469970 35091
rect 470090 34491 470146 35091
rect 470266 34491 470316 35091
rect 469732 34302 470332 34352
rect 470395 34302 470445 35091
rect 373032 33959 373098 33975
rect 373194 33959 373260 33975
rect 368923 33261 368973 33861
rect 369107 33261 369163 33861
rect 369487 33261 369523 33861
rect 327862 32810 327870 33035
rect 368452 32481 368502 33081
rect 368602 32481 368658 33081
rect 368758 32481 368808 33081
rect 368888 32481 368938 33081
rect 369038 32481 369166 33081
rect 369194 32481 369250 33081
rect 369350 32481 369478 33081
rect 369506 32481 369556 33081
rect 369636 32481 369686 33081
rect 369786 32481 369914 33081
rect 369942 32481 370070 33081
rect 370098 32481 370148 33081
rect 371341 32596 371391 33196
rect 371775 32596 371825 33196
rect 371977 32596 372027 33596
rect 372127 32596 372183 33596
rect 372283 32596 372411 33596
rect 372439 32596 372567 33596
rect 372595 32596 372723 33596
rect 372751 32596 372879 33596
rect 372907 32596 373035 33596
rect 373063 32596 373191 33596
rect 373219 32596 373347 33596
rect 373375 32596 373425 33596
rect 373577 32546 373627 33546
rect 373727 32546 373855 33546
rect 373883 32546 374011 33546
rect 374039 32546 374167 33546
rect 374195 32546 374323 33546
rect 374351 32546 374479 33546
rect 374507 32546 374635 33546
rect 374663 32546 374791 33546
rect 374819 32546 374869 33546
rect 375021 32596 375071 33596
rect 375171 32596 375299 33596
rect 375327 32596 375455 33596
rect 375483 32596 375611 33596
rect 375639 32596 375767 33596
rect 375795 32596 375923 33596
rect 375951 32596 376079 33596
rect 376107 32596 376235 33596
rect 376263 32596 376313 33596
rect 376465 32596 376515 33596
rect 376615 32596 376743 33596
rect 376771 32596 376899 33596
rect 376927 32596 377055 33596
rect 377083 32596 377139 33596
rect 377239 32596 377367 33596
rect 377395 32596 377523 33596
rect 377551 32596 377679 33596
rect 377707 32596 377757 33596
rect 377823 32596 377873 33596
rect 377973 32596 378029 33596
rect 378129 32596 378179 33596
rect 378351 32930 378401 33530
rect 378501 32930 378557 33530
rect 378657 32930 378707 33530
rect 379563 33292 379613 33892
rect 379713 33292 379763 33892
rect 379862 32810 379870 33035
rect 425707 32596 425757 33596
rect 425823 32596 425873 33596
rect 425973 32596 426029 33596
rect 426129 32596 426179 33596
rect 426351 32930 426401 33530
rect 426501 32930 426557 33530
rect 426657 32930 426707 33530
rect 427563 33292 427613 33892
rect 427713 33292 427763 33892
rect 467157 33672 467207 34272
rect 467327 33672 467455 34272
rect 467503 33672 467559 34272
rect 467679 33672 467735 34272
rect 467855 33672 467911 34272
rect 468031 33672 468159 34272
rect 468207 33672 468263 34272
rect 468383 33672 468433 34272
rect 470392 34202 470445 34302
rect 469732 34152 470332 34202
rect 470395 34101 470445 34202
rect 470392 34091 470445 34101
rect 470565 34101 470615 35091
rect 470703 34491 470753 35091
rect 470873 34491 470929 35091
rect 471049 34491 471099 35091
rect 471319 34492 471369 35092
rect 471489 34492 471545 35092
rect 471665 34492 471715 35092
rect 470678 34322 471678 34372
rect 470678 34202 470690 34322
rect 470678 34152 471678 34202
rect 474611 34110 474661 34710
rect 474761 34110 474889 34710
rect 474917 34110 474973 34710
rect 475073 34110 475201 34710
rect 475229 34110 475279 34710
rect 475345 34110 475395 34710
rect 475495 34110 475551 34710
rect 475651 34110 475707 34710
rect 475807 34110 475863 34710
rect 475963 34110 476091 34710
rect 476119 34110 476247 34710
rect 476275 34110 476403 34710
rect 476431 34110 476487 34710
rect 476587 34110 476715 34710
rect 476743 34110 476871 34710
rect 476899 34110 477027 34710
rect 477055 34110 477105 34710
rect 477171 34110 477221 34710
rect 477321 34110 477449 34710
rect 477477 34110 477605 34710
rect 477633 34110 477761 34710
rect 477789 34110 477839 34710
rect 470565 34091 470618 34101
rect 478051 34079 478101 34679
rect 478201 34079 478257 34679
rect 478357 34079 478407 34679
rect 529789 34110 529839 34710
rect 530051 34079 530101 34679
rect 530201 34079 530257 34679
rect 530357 34079 530407 34679
rect 567233 34427 567283 35027
rect 567403 34427 567531 35027
rect 567579 34427 567635 35027
rect 567755 34427 567883 35027
rect 567931 34427 568059 35027
rect 568107 34427 568235 35027
rect 568283 34427 568411 35027
rect 568459 34427 568509 35027
rect 568881 34491 568931 35091
rect 569051 34491 569179 35091
rect 569227 34491 569283 35091
rect 569403 34491 569531 35091
rect 569579 34491 569629 35091
rect 569920 34491 569970 35091
rect 570090 34491 570146 35091
rect 570266 34491 570316 35091
rect 569732 34302 570332 34352
rect 570395 34302 570445 35091
rect 473032 33959 473098 33975
rect 473194 33959 473260 33975
rect 468923 33261 468973 33861
rect 469107 33261 469163 33861
rect 469487 33261 469523 33861
rect 427862 32810 427870 33035
rect 468452 32481 468502 33081
rect 468602 32481 468658 33081
rect 468758 32481 468808 33081
rect 468888 32481 468938 33081
rect 469038 32481 469166 33081
rect 469194 32481 469250 33081
rect 469350 32481 469478 33081
rect 469506 32481 469556 33081
rect 469636 32481 469686 33081
rect 469786 32481 469914 33081
rect 469942 32481 470070 33081
rect 470098 32481 470148 33081
rect 471341 32596 471391 33196
rect 471775 32596 471825 33196
rect 471977 32596 472027 33596
rect 472127 32596 472183 33596
rect 472283 32596 472411 33596
rect 472439 32596 472567 33596
rect 472595 32596 472723 33596
rect 472751 32596 472879 33596
rect 472907 32596 473035 33596
rect 473063 32596 473191 33596
rect 473219 32596 473347 33596
rect 473375 32596 473425 33596
rect 473577 32546 473627 33546
rect 473727 32546 473855 33546
rect 473883 32546 474011 33546
rect 474039 32546 474167 33546
rect 474195 32546 474323 33546
rect 474351 32546 474479 33546
rect 474507 32546 474635 33546
rect 474663 32546 474791 33546
rect 474819 32546 474869 33546
rect 475021 32596 475071 33596
rect 475171 32596 475299 33596
rect 475327 32596 475455 33596
rect 475483 32596 475611 33596
rect 475639 32596 475767 33596
rect 475795 32596 475923 33596
rect 475951 32596 476079 33596
rect 476107 32596 476235 33596
rect 476263 32596 476313 33596
rect 476465 32596 476515 33596
rect 476615 32596 476743 33596
rect 476771 32596 476899 33596
rect 476927 32596 477055 33596
rect 477083 32596 477139 33596
rect 477239 32596 477367 33596
rect 477395 32596 477523 33596
rect 477551 32596 477679 33596
rect 477707 32596 477757 33596
rect 477823 32596 477873 33596
rect 477973 32596 478029 33596
rect 478129 32596 478179 33596
rect 478351 32930 478401 33530
rect 478501 32930 478557 33530
rect 478657 32930 478707 33530
rect 479563 33292 479613 33892
rect 479713 33292 479763 33892
rect 479862 32810 479870 33035
rect 529707 32596 529757 33596
rect 529823 32596 529873 33596
rect 529973 32596 530029 33596
rect 530129 32596 530179 33596
rect 530351 32930 530401 33530
rect 530501 32930 530557 33530
rect 530657 32930 530707 33530
rect 531563 33292 531613 33892
rect 531713 33292 531763 33892
rect 567157 33672 567207 34272
rect 567327 33672 567455 34272
rect 567503 33672 567559 34272
rect 567679 33672 567735 34272
rect 567855 33672 567911 34272
rect 568031 33672 568159 34272
rect 568207 33672 568263 34272
rect 568383 33672 568433 34272
rect 570392 34202 570445 34302
rect 569732 34152 570332 34202
rect 570395 34101 570445 34202
rect 570392 34091 570445 34101
rect 570565 34101 570615 35091
rect 570703 34491 570753 35091
rect 570873 34491 570929 35091
rect 571049 34491 571099 35091
rect 571319 34492 571369 35092
rect 571489 34492 571545 35092
rect 571665 34492 571715 35092
rect 570678 34322 571678 34372
rect 570678 34202 570690 34322
rect 570678 34152 571678 34202
rect 574611 34110 574661 34710
rect 574761 34110 574889 34710
rect 574917 34110 574973 34710
rect 575073 34110 575201 34710
rect 575229 34110 575279 34710
rect 575345 34110 575395 34710
rect 575495 34110 575551 34710
rect 575651 34110 575707 34710
rect 575807 34110 575863 34710
rect 575963 34110 576091 34710
rect 576119 34110 576247 34710
rect 576275 34110 576403 34710
rect 576431 34110 576487 34710
rect 576587 34110 576715 34710
rect 576743 34110 576871 34710
rect 576899 34110 577027 34710
rect 577055 34110 577105 34710
rect 577171 34110 577221 34710
rect 577321 34110 577449 34710
rect 577477 34110 577605 34710
rect 577633 34110 577761 34710
rect 577789 34110 577839 34710
rect 570565 34091 570618 34101
rect 578051 34079 578101 34679
rect 578201 34079 578257 34679
rect 578357 34079 578407 34679
rect 573032 33959 573098 33975
rect 573194 33959 573260 33975
rect 568923 33261 568973 33861
rect 569107 33261 569163 33861
rect 569487 33261 569523 33861
rect 531862 32810 531870 33035
rect 568452 32481 568502 33081
rect 568602 32481 568658 33081
rect 568758 32481 568808 33081
rect 568888 32481 568938 33081
rect 569038 32481 569166 33081
rect 569194 32481 569250 33081
rect 569350 32481 569478 33081
rect 569506 32481 569556 33081
rect 569636 32481 569686 33081
rect 569786 32481 569914 33081
rect 569942 32481 570070 33081
rect 570098 32481 570148 33081
rect 571341 32596 571391 33196
rect 571775 32596 571825 33196
rect 571977 32596 572027 33596
rect 572127 32596 572183 33596
rect 572283 32596 572411 33596
rect 572439 32596 572567 33596
rect 572595 32596 572723 33596
rect 572751 32596 572879 33596
rect 572907 32596 573035 33596
rect 573063 32596 573191 33596
rect 573219 32596 573347 33596
rect 573375 32596 573425 33596
rect 573577 32546 573627 33546
rect 573727 32546 573855 33546
rect 573883 32546 574011 33546
rect 574039 32546 574167 33546
rect 574195 32546 574323 33546
rect 574351 32546 574479 33546
rect 574507 32546 574635 33546
rect 574663 32546 574791 33546
rect 574819 32546 574869 33546
rect 575021 32596 575071 33596
rect 575171 32596 575299 33596
rect 575327 32596 575455 33596
rect 575483 32596 575611 33596
rect 575639 32596 575767 33596
rect 575795 32596 575923 33596
rect 575951 32596 576079 33596
rect 576107 32596 576235 33596
rect 576263 32596 576313 33596
rect 576465 32596 576515 33596
rect 576615 32596 576743 33596
rect 576771 32596 576899 33596
rect 576927 32596 577055 33596
rect 577083 32596 577139 33596
rect 577239 32596 577367 33596
rect 577395 32596 577523 33596
rect 577551 32596 577679 33596
rect 577707 32596 577757 33596
rect 577823 32596 577873 33596
rect 577973 32596 578029 33596
rect 578129 32596 578179 33596
rect 578351 32930 578401 33530
rect 578501 32930 578557 33530
rect 578657 32930 578707 33530
rect 579563 33292 579613 33892
rect 579713 33292 579763 33892
rect 579862 32810 579870 33035
rect 36262 31387 36264 31512
rect 56848 31453 56898 32053
rect 57018 31453 57068 32053
rect 57444 31458 57494 32058
rect 57614 31458 57670 32058
rect 57790 31458 57840 32058
rect 58434 31049 58484 32049
rect 69480 31607 69517 31807
rect 69480 31347 69517 31547
rect 70201 31463 70251 32063
rect 70351 31463 70407 32063
rect 70507 31463 70557 32063
rect 108848 31453 108898 32053
rect 109018 31453 109068 32053
rect 109444 31458 109494 32058
rect 109614 31458 109670 32058
rect 109790 31458 109840 32058
rect 110434 31049 110484 32049
rect 121480 31607 121517 31807
rect 121480 31347 121517 31547
rect 122201 31463 122251 32063
rect 122351 31463 122407 32063
rect 122507 31463 122557 32063
rect 160848 31453 160898 32053
rect 161018 31453 161068 32053
rect 173480 31607 173517 31807
rect 173480 31347 173517 31547
rect 174201 31463 174251 32063
rect 174351 31463 174407 32063
rect 174507 31463 174557 32063
rect 212848 31453 212898 32053
rect 213018 31453 213068 32053
rect 213444 31458 213494 32058
rect 213614 31458 213670 32058
rect 213790 31458 213840 32058
rect 214434 31049 214484 32049
rect 225480 31607 225517 31807
rect 225480 31347 225517 31547
rect 226201 31463 226251 32063
rect 226351 31463 226407 32063
rect 226507 31463 226557 32063
rect 260848 31453 260898 32053
rect 261018 31453 261068 32053
rect 261444 31458 261494 32058
rect 261614 31458 261670 32058
rect 261790 31458 261840 32058
rect 273480 31607 273517 31807
rect 273480 31347 273517 31547
rect 274201 31463 274251 32063
rect 274351 31463 274407 32063
rect 274507 31463 274557 32063
rect 312848 31453 312898 32053
rect 313018 31453 313068 32053
rect 313444 31458 313494 32058
rect 313614 31458 313670 32058
rect 313790 31458 313840 32058
rect 314434 31049 314484 32049
rect 325480 31607 325517 31807
rect 325480 31347 325517 31547
rect 326201 31463 326251 32063
rect 326351 31463 326407 32063
rect 326507 31463 326557 32063
rect 364848 31453 364898 32053
rect 365018 31453 365068 32053
rect 365444 31458 365494 32058
rect 365614 31458 365670 32058
rect 365790 31999 365840 32058
rect 365790 31927 365843 31999
rect 365790 31680 365840 31927
rect 365903 31777 365915 31927
rect 365790 31608 365843 31680
rect 365790 31458 365840 31608
rect 365903 31458 365915 31608
rect 366434 31049 366484 32049
rect 366584 31049 366712 32049
rect 366740 31049 366868 32049
rect 366896 31049 367024 32049
rect 367052 31049 367108 32049
rect 367208 31049 367336 32049
rect 367364 31049 367492 32049
rect 367520 31049 367648 32049
rect 367676 31049 367726 32049
rect 367792 31049 367842 32049
rect 367962 31049 368090 32049
rect 368138 31049 368266 32049
rect 368314 31049 368442 32049
rect 368490 31049 368618 32049
rect 368666 31049 368794 32049
rect 368842 31049 368970 32049
rect 369018 31049 369146 32049
rect 369194 31049 369250 32049
rect 369350 31049 369478 32049
rect 369506 31049 369634 32049
rect 369662 31049 369790 32049
rect 369818 31049 369946 32049
rect 369974 31049 370102 32049
rect 370130 31049 370186 32049
rect 370286 31049 370414 32049
rect 370442 31049 370570 32049
rect 370598 31049 370726 32049
rect 370754 31049 370882 32049
rect 370910 31049 371038 32049
rect 371066 31049 371116 32049
rect 371182 31049 371232 32049
rect 371332 31049 371388 32049
rect 371488 31049 371544 32049
rect 371644 31049 371700 32049
rect 371800 31049 371850 32049
rect 371936 31049 371986 32049
rect 372086 31049 372142 32049
rect 372242 31049 372292 32049
rect 372789 31463 372839 32063
rect 372939 31463 372995 32063
rect 373095 31463 373145 32063
rect 374410 32055 374620 32067
rect 376284 32061 376318 32087
rect 374414 32052 374616 32055
rect 374425 31882 374605 32052
rect 374785 31882 374815 31921
rect 374871 31882 374901 31921
rect 374410 31867 374620 31882
rect 374770 31867 374830 31882
rect 374856 31867 374916 31882
rect 375028 31823 375060 32061
rect 376280 31823 376318 32061
rect 376726 32055 376936 32067
rect 376730 32052 376932 32055
rect 376445 31882 376475 31921
rect 376531 31882 376561 31921
rect 376741 31882 376921 32052
rect 376430 31867 376490 31882
rect 376516 31867 376576 31882
rect 376726 31867 376936 31882
rect 373814 31795 374024 31807
rect 374050 31795 374260 31807
rect 374410 31795 374620 31807
rect 374770 31795 374830 31807
rect 374856 31795 374916 31807
rect 376280 31797 376284 31823
rect 373818 31792 374020 31795
rect 374054 31792 374256 31795
rect 374414 31792 374616 31795
rect 374774 31792 374826 31795
rect 374860 31792 374912 31795
rect 373829 31622 374009 31792
rect 374065 31622 374245 31792
rect 374425 31622 374605 31792
rect 374785 31622 374815 31792
rect 374871 31622 374901 31792
rect 373814 31607 374024 31622
rect 374050 31607 374260 31622
rect 374410 31607 374620 31622
rect 374770 31607 374830 31622
rect 374856 31607 374916 31622
rect 373814 31535 374024 31547
rect 374050 31535 374260 31547
rect 374410 31535 374620 31547
rect 374770 31535 374830 31547
rect 374856 31535 374916 31547
rect 373818 31532 374020 31535
rect 374054 31532 374256 31535
rect 374414 31532 374616 31535
rect 374774 31532 374826 31535
rect 374860 31532 374912 31535
rect 373829 31362 374009 31532
rect 374065 31362 374245 31532
rect 374425 31362 374605 31532
rect 374785 31362 374815 31532
rect 374871 31362 374901 31532
rect 375062 31481 375080 31797
rect 376268 31481 376284 31797
rect 376430 31795 376490 31807
rect 376516 31795 376576 31807
rect 376726 31795 376936 31807
rect 377086 31795 377296 31807
rect 377322 31795 377532 31807
rect 376434 31792 376486 31795
rect 376520 31792 376572 31795
rect 376730 31792 376932 31795
rect 377090 31792 377292 31795
rect 377326 31792 377528 31795
rect 376445 31622 376475 31792
rect 376531 31622 376561 31792
rect 376741 31622 376921 31792
rect 377101 31622 377281 31792
rect 377337 31622 377517 31792
rect 376430 31607 376490 31622
rect 376516 31607 376576 31622
rect 376726 31607 376936 31622
rect 377086 31607 377296 31622
rect 377322 31607 377532 31622
rect 376430 31535 376490 31547
rect 376516 31535 376576 31547
rect 376726 31535 376936 31547
rect 377086 31535 377296 31547
rect 377322 31535 377532 31547
rect 376434 31532 376486 31535
rect 376520 31532 376572 31535
rect 376730 31532 376932 31535
rect 377090 31532 377292 31535
rect 377326 31532 377528 31535
rect 376445 31362 376475 31532
rect 376531 31362 376561 31532
rect 376741 31362 376921 31532
rect 377101 31362 377281 31532
rect 377337 31362 377517 31532
rect 378201 31463 378251 32063
rect 378351 31463 378407 32063
rect 378507 31463 378557 32063
rect 412848 31453 412898 32053
rect 413018 31453 413068 32053
rect 413444 31458 413494 32058
rect 413614 31458 413670 32058
rect 413790 31458 413840 32058
rect 373814 31347 374024 31362
rect 374050 31347 374260 31362
rect 374410 31347 374620 31362
rect 374770 31347 374830 31362
rect 374856 31347 374916 31362
rect 376430 31347 376490 31362
rect 376516 31347 376576 31362
rect 376726 31347 376936 31362
rect 377086 31347 377296 31362
rect 377322 31347 377532 31362
rect 374410 31275 374620 31287
rect 376726 31275 376936 31287
rect 374414 31272 374616 31275
rect 376730 31272 376932 31275
rect 374425 31102 374605 31272
rect 376741 31102 376921 31272
rect 374410 31087 374620 31102
rect 376726 31087 376936 31102
rect 414434 31049 414484 32049
rect 425480 31607 425517 31807
rect 425480 31347 425517 31547
rect 426201 31463 426251 32063
rect 426351 31463 426407 32063
rect 426507 31463 426557 32063
rect 464848 31453 464898 32053
rect 465018 31453 465068 32053
rect 465444 31458 465494 32058
rect 465614 31458 465670 32058
rect 465790 31999 465840 32058
rect 465790 31927 465843 31999
rect 465790 31680 465840 31927
rect 465903 31777 465915 31927
rect 465790 31608 465843 31680
rect 465790 31458 465840 31608
rect 465903 31458 465915 31608
rect 466434 31049 466484 32049
rect 466584 31049 466712 32049
rect 466740 31049 466868 32049
rect 466896 31049 467024 32049
rect 467052 31049 467108 32049
rect 467208 31049 467336 32049
rect 467364 31049 467492 32049
rect 467520 31049 467648 32049
rect 467676 31049 467726 32049
rect 467792 31049 467842 32049
rect 467962 31049 468090 32049
rect 468138 31049 468266 32049
rect 468314 31049 468442 32049
rect 468490 31049 468618 32049
rect 468666 31049 468794 32049
rect 468842 31049 468970 32049
rect 469018 31049 469146 32049
rect 469194 31049 469250 32049
rect 469350 31049 469478 32049
rect 469506 31049 469634 32049
rect 469662 31049 469790 32049
rect 469818 31049 469946 32049
rect 469974 31049 470102 32049
rect 470130 31049 470186 32049
rect 470286 31049 470414 32049
rect 470442 31049 470570 32049
rect 470598 31049 470726 32049
rect 470754 31049 470882 32049
rect 470910 31049 471038 32049
rect 471066 31049 471116 32049
rect 471182 31049 471232 32049
rect 471332 31049 471388 32049
rect 471488 31049 471544 32049
rect 471644 31049 471700 32049
rect 471800 31049 471850 32049
rect 471936 31049 471986 32049
rect 472086 31049 472142 32049
rect 472242 31049 472292 32049
rect 472789 31463 472839 32063
rect 472939 31463 472995 32063
rect 473095 31463 473145 32063
rect 474410 32055 474620 32067
rect 476284 32061 476318 32087
rect 474414 32052 474616 32055
rect 474425 31882 474605 32052
rect 474785 31882 474815 31921
rect 474871 31882 474901 31921
rect 474410 31867 474620 31882
rect 474770 31867 474830 31882
rect 474856 31867 474916 31882
rect 475028 31823 475060 32061
rect 476280 31823 476318 32061
rect 476726 32055 476936 32067
rect 476730 32052 476932 32055
rect 476445 31882 476475 31921
rect 476531 31882 476561 31921
rect 476741 31882 476921 32052
rect 476430 31867 476490 31882
rect 476516 31867 476576 31882
rect 476726 31867 476936 31882
rect 473814 31795 474024 31807
rect 474050 31795 474260 31807
rect 474410 31795 474620 31807
rect 474770 31795 474830 31807
rect 474856 31795 474916 31807
rect 476280 31797 476284 31823
rect 473818 31792 474020 31795
rect 474054 31792 474256 31795
rect 474414 31792 474616 31795
rect 474774 31792 474826 31795
rect 474860 31792 474912 31795
rect 473829 31622 474009 31792
rect 474065 31622 474245 31792
rect 474425 31622 474605 31792
rect 474785 31622 474815 31792
rect 474871 31622 474901 31792
rect 473814 31607 474024 31622
rect 474050 31607 474260 31622
rect 474410 31607 474620 31622
rect 474770 31607 474830 31622
rect 474856 31607 474916 31622
rect 473814 31535 474024 31547
rect 474050 31535 474260 31547
rect 474410 31535 474620 31547
rect 474770 31535 474830 31547
rect 474856 31535 474916 31547
rect 473818 31532 474020 31535
rect 474054 31532 474256 31535
rect 474414 31532 474616 31535
rect 474774 31532 474826 31535
rect 474860 31532 474912 31535
rect 473829 31362 474009 31532
rect 474065 31362 474245 31532
rect 474425 31362 474605 31532
rect 474785 31362 474815 31532
rect 474871 31362 474901 31532
rect 475062 31481 475080 31797
rect 476268 31481 476284 31797
rect 476430 31795 476490 31807
rect 476516 31795 476576 31807
rect 476726 31795 476936 31807
rect 477086 31795 477296 31807
rect 477322 31795 477532 31807
rect 476434 31792 476486 31795
rect 476520 31792 476572 31795
rect 476730 31792 476932 31795
rect 477090 31792 477292 31795
rect 477326 31792 477528 31795
rect 476445 31622 476475 31792
rect 476531 31622 476561 31792
rect 476741 31622 476921 31792
rect 477101 31622 477281 31792
rect 477337 31622 477517 31792
rect 476430 31607 476490 31622
rect 476516 31607 476576 31622
rect 476726 31607 476936 31622
rect 477086 31607 477296 31622
rect 477322 31607 477532 31622
rect 476430 31535 476490 31547
rect 476516 31535 476576 31547
rect 476726 31535 476936 31547
rect 477086 31535 477296 31547
rect 477322 31535 477532 31547
rect 476434 31532 476486 31535
rect 476520 31532 476572 31535
rect 476730 31532 476932 31535
rect 477090 31532 477292 31535
rect 477326 31532 477528 31535
rect 476445 31362 476475 31532
rect 476531 31362 476561 31532
rect 476741 31362 476921 31532
rect 477101 31362 477281 31532
rect 477337 31362 477517 31532
rect 478201 31463 478251 32063
rect 478351 31463 478407 32063
rect 478507 31463 478557 32063
rect 516848 31453 516898 32053
rect 517018 31453 517068 32053
rect 517444 31458 517494 32058
rect 517614 31458 517670 32058
rect 517790 31458 517840 32058
rect 473814 31347 474024 31362
rect 474050 31347 474260 31362
rect 474410 31347 474620 31362
rect 474770 31347 474830 31362
rect 474856 31347 474916 31362
rect 476430 31347 476490 31362
rect 476516 31347 476576 31362
rect 476726 31347 476936 31362
rect 477086 31347 477296 31362
rect 477322 31347 477532 31362
rect 474410 31275 474620 31287
rect 476726 31275 476936 31287
rect 474414 31272 474616 31275
rect 476730 31272 476932 31275
rect 474425 31102 474605 31272
rect 476741 31102 476921 31272
rect 474410 31087 474620 31102
rect 476726 31087 476936 31102
rect 518434 31049 518484 32049
rect 529480 31607 529517 31807
rect 529480 31347 529517 31547
rect 530201 31463 530251 32063
rect 530351 31463 530407 32063
rect 530507 31463 530557 32063
rect 564848 31453 564898 32053
rect 565018 31453 565068 32053
rect 565444 31458 565494 32058
rect 565614 31458 565670 32058
rect 565790 31999 565840 32058
rect 565790 31927 565843 31999
rect 565790 31680 565840 31927
rect 565903 31777 565915 31927
rect 565790 31608 565843 31680
rect 565790 31458 565840 31608
rect 565903 31458 565915 31608
rect 566434 31049 566484 32049
rect 566584 31049 566712 32049
rect 566740 31049 566868 32049
rect 566896 31049 567024 32049
rect 567052 31049 567108 32049
rect 567208 31049 567336 32049
rect 567364 31049 567492 32049
rect 567520 31049 567648 32049
rect 567676 31049 567726 32049
rect 567792 31049 567842 32049
rect 567962 31049 568090 32049
rect 568138 31049 568266 32049
rect 568314 31049 568442 32049
rect 568490 31049 568618 32049
rect 568666 31049 568794 32049
rect 568842 31049 568970 32049
rect 569018 31049 569146 32049
rect 569194 31049 569250 32049
rect 569350 31049 569478 32049
rect 569506 31049 569634 32049
rect 569662 31049 569790 32049
rect 569818 31049 569946 32049
rect 569974 31049 570102 32049
rect 570130 31049 570186 32049
rect 570286 31049 570414 32049
rect 570442 31049 570570 32049
rect 570598 31049 570726 32049
rect 570754 31049 570882 32049
rect 570910 31049 571038 32049
rect 571066 31049 571116 32049
rect 571182 31049 571232 32049
rect 571332 31049 571388 32049
rect 571488 31049 571544 32049
rect 571644 31049 571700 32049
rect 571800 31049 571850 32049
rect 571936 31049 571986 32049
rect 572086 31049 572142 32049
rect 572242 31049 572292 32049
rect 572789 31463 572839 32063
rect 572939 31463 572995 32063
rect 573095 31463 573145 32063
rect 574410 32055 574620 32067
rect 576284 32061 576318 32087
rect 574414 32052 574616 32055
rect 574425 31882 574605 32052
rect 574785 31882 574815 31921
rect 574871 31882 574901 31921
rect 574410 31867 574620 31882
rect 574770 31867 574830 31882
rect 574856 31867 574916 31882
rect 575028 31823 575060 32061
rect 576280 31823 576318 32061
rect 576726 32055 576936 32067
rect 576730 32052 576932 32055
rect 576445 31882 576475 31921
rect 576531 31882 576561 31921
rect 576741 31882 576921 32052
rect 576430 31867 576490 31882
rect 576516 31867 576576 31882
rect 576726 31867 576936 31882
rect 573814 31795 574024 31807
rect 574050 31795 574260 31807
rect 574410 31795 574620 31807
rect 574770 31795 574830 31807
rect 574856 31795 574916 31807
rect 576280 31797 576284 31823
rect 573818 31792 574020 31795
rect 574054 31792 574256 31795
rect 574414 31792 574616 31795
rect 574774 31792 574826 31795
rect 574860 31792 574912 31795
rect 573829 31622 574009 31792
rect 574065 31622 574245 31792
rect 574425 31622 574605 31792
rect 574785 31622 574815 31792
rect 574871 31622 574901 31792
rect 573814 31607 574024 31622
rect 574050 31607 574260 31622
rect 574410 31607 574620 31622
rect 574770 31607 574830 31622
rect 574856 31607 574916 31622
rect 573814 31535 574024 31547
rect 574050 31535 574260 31547
rect 574410 31535 574620 31547
rect 574770 31535 574830 31547
rect 574856 31535 574916 31547
rect 573818 31532 574020 31535
rect 574054 31532 574256 31535
rect 574414 31532 574616 31535
rect 574774 31532 574826 31535
rect 574860 31532 574912 31535
rect 573829 31362 574009 31532
rect 574065 31362 574245 31532
rect 574425 31362 574605 31532
rect 574785 31362 574815 31532
rect 574871 31362 574901 31532
rect 575062 31481 575080 31797
rect 576268 31481 576284 31797
rect 576430 31795 576490 31807
rect 576516 31795 576576 31807
rect 576726 31795 576936 31807
rect 577086 31795 577296 31807
rect 577322 31795 577532 31807
rect 576434 31792 576486 31795
rect 576520 31792 576572 31795
rect 576730 31792 576932 31795
rect 577090 31792 577292 31795
rect 577326 31792 577528 31795
rect 576445 31622 576475 31792
rect 576531 31622 576561 31792
rect 576741 31622 576921 31792
rect 577101 31622 577281 31792
rect 577337 31622 577517 31792
rect 576430 31607 576490 31622
rect 576516 31607 576576 31622
rect 576726 31607 576936 31622
rect 577086 31607 577296 31622
rect 577322 31607 577532 31622
rect 576430 31535 576490 31547
rect 576516 31535 576576 31547
rect 576726 31535 576936 31547
rect 577086 31535 577296 31547
rect 577322 31535 577532 31547
rect 576434 31532 576486 31535
rect 576520 31532 576572 31535
rect 576730 31532 576932 31535
rect 577090 31532 577292 31535
rect 577326 31532 577528 31535
rect 576445 31362 576475 31532
rect 576531 31362 576561 31532
rect 576741 31362 576921 31532
rect 577101 31362 577281 31532
rect 577337 31362 577517 31532
rect 578201 31463 578251 32063
rect 578351 31463 578407 32063
rect 578507 31463 578557 32063
rect 573814 31347 574024 31362
rect 574050 31347 574260 31362
rect 574410 31347 574620 31362
rect 574770 31347 574830 31362
rect 574856 31347 574916 31362
rect 576430 31347 576490 31362
rect 576516 31347 576576 31362
rect 576726 31347 576936 31362
rect 577086 31347 577296 31362
rect 577322 31347 577532 31362
rect 574410 31275 574620 31287
rect 576726 31275 576936 31287
rect 574414 31272 574616 31275
rect 576730 31272 576932 31275
rect 574425 31102 574605 31272
rect 576741 31102 576921 31272
rect 574410 31087 574620 31102
rect 576726 31087 576936 31102
rect 56150 30245 56200 30845
rect 56320 30245 56376 30845
rect 56496 30245 56552 30845
rect 56672 30245 56722 30845
rect 57229 30558 57409 30580
rect 57214 30543 57409 30558
rect 56978 30430 57188 30445
rect 57214 30430 57409 30445
rect 56993 30260 57173 30430
rect 57229 30260 57409 30430
rect 56982 30257 57184 30260
rect 57218 30257 57409 30260
rect 56978 30245 57188 30257
rect 57214 30245 57409 30257
rect 69510 29993 69560 30993
rect 71107 30907 71141 30911
rect 71178 30907 71212 30911
rect 71249 30907 71283 30911
rect 71083 30891 71335 30907
rect 71107 30887 71141 30891
rect 71178 30887 71212 30891
rect 71249 30887 71283 30891
rect 71083 30881 71305 30887
rect 71083 30867 71307 30881
rect 71296 30857 71307 30867
rect 71259 30833 71283 30857
rect 71320 30833 71344 30857
rect 69649 30171 69699 30771
rect 69819 30171 69875 30771
rect 69995 30171 70045 30771
rect 108150 30245 108200 30845
rect 108320 30245 108376 30845
rect 108496 30245 108552 30845
rect 108672 30245 108722 30845
rect 109229 30558 109409 30580
rect 109214 30543 109409 30558
rect 108978 30430 109188 30445
rect 109214 30430 109409 30445
rect 108993 30260 109173 30430
rect 109229 30260 109409 30430
rect 108982 30257 109184 30260
rect 109218 30257 109409 30260
rect 108978 30245 109188 30257
rect 109214 30245 109409 30257
rect 121510 29993 121560 30993
rect 123107 30907 123141 30911
rect 123178 30907 123212 30911
rect 123249 30907 123283 30911
rect 123083 30891 123335 30907
rect 123107 30887 123141 30891
rect 123178 30887 123212 30891
rect 123249 30887 123283 30891
rect 123083 30881 123305 30887
rect 123083 30867 123307 30881
rect 123296 30857 123307 30867
rect 123259 30833 123283 30857
rect 123320 30833 123344 30857
rect 121649 30171 121699 30771
rect 121819 30171 121875 30771
rect 121995 30171 122045 30771
rect 160150 30245 160200 30845
rect 160320 30245 160376 30845
rect 160496 30245 160552 30845
rect 160672 30245 160722 30845
rect 161229 30558 161280 30580
rect 161214 30543 161280 30558
rect 160978 30430 161188 30445
rect 161214 30430 161280 30445
rect 160993 30260 161173 30430
rect 161229 30260 161280 30430
rect 160982 30257 161184 30260
rect 161218 30257 161280 30260
rect 160978 30245 161188 30257
rect 161214 30245 161280 30257
rect 173510 29993 173560 30993
rect 175107 30907 175141 30911
rect 175178 30907 175212 30911
rect 175249 30907 175283 30911
rect 175083 30891 175335 30907
rect 175107 30887 175141 30891
rect 175178 30887 175212 30891
rect 175249 30887 175283 30891
rect 175083 30881 175305 30887
rect 175083 30867 175307 30881
rect 175296 30857 175307 30867
rect 175259 30833 175283 30857
rect 175320 30833 175344 30857
rect 173649 30171 173699 30771
rect 173819 30171 173875 30771
rect 173995 30171 174045 30771
rect 212150 30245 212200 30845
rect 212320 30245 212376 30845
rect 212496 30245 212552 30845
rect 212672 30245 212722 30845
rect 213229 30558 213409 30580
rect 213214 30543 213409 30558
rect 212978 30430 213188 30445
rect 213214 30430 213409 30445
rect 212993 30260 213173 30430
rect 213229 30260 213409 30430
rect 212982 30257 213184 30260
rect 213218 30257 213409 30260
rect 212978 30245 213188 30257
rect 213214 30245 213409 30257
rect 225510 29993 225560 30993
rect 227107 30907 227141 30911
rect 227178 30907 227212 30911
rect 227249 30907 227283 30911
rect 227083 30891 227335 30907
rect 227107 30887 227141 30891
rect 227178 30887 227212 30891
rect 227249 30887 227283 30891
rect 227083 30881 227305 30887
rect 227083 30867 227307 30881
rect 227296 30857 227307 30867
rect 227259 30833 227283 30857
rect 227320 30833 227344 30857
rect 225649 30171 225699 30771
rect 225819 30171 225875 30771
rect 225995 30171 226045 30771
rect 260150 30245 260200 30845
rect 260320 30245 260376 30845
rect 260496 30245 260552 30845
rect 260672 30245 260722 30845
rect 261229 30558 261409 30580
rect 261214 30543 261409 30558
rect 260978 30430 261188 30445
rect 261214 30430 261409 30445
rect 260993 30260 261173 30430
rect 261229 30260 261409 30430
rect 260982 30257 261184 30260
rect 261218 30257 261409 30260
rect 260978 30245 261188 30257
rect 261214 30245 261409 30257
rect 273510 29993 273560 30993
rect 275107 30907 275141 30911
rect 275178 30907 275212 30911
rect 275249 30907 275283 30911
rect 275083 30891 275335 30907
rect 275107 30887 275141 30891
rect 275178 30887 275212 30891
rect 275249 30887 275283 30891
rect 275083 30881 275305 30887
rect 275083 30867 275307 30881
rect 275296 30857 275307 30867
rect 275259 30833 275283 30857
rect 275320 30833 275344 30857
rect 273649 30171 273699 30771
rect 273819 30171 273875 30771
rect 273995 30171 274045 30771
rect 312150 30245 312200 30845
rect 312320 30245 312376 30845
rect 312496 30245 312552 30845
rect 312672 30245 312722 30845
rect 313229 30558 313409 30580
rect 313214 30543 313409 30558
rect 312978 30430 313188 30445
rect 313214 30430 313409 30445
rect 312993 30260 313173 30430
rect 313229 30260 313409 30430
rect 312982 30257 313184 30260
rect 313218 30257 313409 30260
rect 312978 30245 313188 30257
rect 313214 30245 313409 30257
rect 325510 29993 325560 30993
rect 327107 30907 327141 30911
rect 327178 30907 327212 30911
rect 327249 30907 327283 30911
rect 327083 30891 327335 30907
rect 327107 30887 327141 30891
rect 327178 30887 327212 30891
rect 327249 30887 327283 30891
rect 327083 30881 327305 30887
rect 327083 30867 327307 30881
rect 327296 30857 327307 30867
rect 327259 30833 327283 30857
rect 327320 30833 327344 30857
rect 325649 30171 325699 30771
rect 325819 30171 325875 30771
rect 325995 30171 326045 30771
rect 364150 30245 364200 30845
rect 364320 30245 364376 30845
rect 364496 30245 364552 30845
rect 364672 30245 364722 30845
rect 366203 30697 366227 30731
rect 366203 30626 366227 30660
rect 365229 30558 365409 30580
rect 365214 30543 365424 30558
rect 366203 30555 366227 30589
rect 366203 30484 366227 30518
rect 364978 30430 365188 30445
rect 365214 30430 365424 30445
rect 364993 30260 365173 30430
rect 365229 30260 365409 30430
rect 366203 30413 366227 30447
rect 366203 30342 366227 30376
rect 366203 30271 366227 30305
rect 364982 30257 365184 30260
rect 365218 30257 365420 30260
rect 364978 30245 365188 30257
rect 365214 30245 365424 30257
rect 366834 30135 366884 30735
rect 367004 30135 367132 30735
rect 367180 30135 367236 30735
rect 367356 30135 367484 30735
rect 367532 30135 367588 30735
rect 367708 30135 367836 30735
rect 367884 30135 367940 30735
rect 368060 30135 368188 30735
rect 368236 30135 368364 30735
rect 368412 30135 368540 30735
rect 368588 30135 368716 30735
rect 368764 30135 368892 30735
rect 368940 30135 368996 30735
rect 369116 30135 369244 30735
rect 369292 30135 369420 30735
rect 369468 30135 369596 30735
rect 369644 30135 369772 30735
rect 369820 30135 369948 30735
rect 369996 30135 370046 30735
rect 370112 30135 370162 30735
rect 370282 30135 370410 30735
rect 370458 30135 370514 30735
rect 370634 30135 370762 30735
rect 370810 30135 370860 30735
rect 370926 30135 370976 30735
rect 371096 30135 371224 30735
rect 371272 30135 371400 30735
rect 371448 30135 371576 30735
rect 371624 30135 371680 30735
rect 371800 30135 371850 30735
rect 371916 30135 371966 30735
rect 372086 30135 372142 30735
rect 372262 30135 372312 30735
rect 372446 30718 372456 30721
rect 372446 30027 372472 30718
rect 373301 30171 373351 30771
rect 373471 30171 373527 30771
rect 373647 30171 373697 30771
rect 366723 30015 372472 30027
rect 373786 29993 373836 30993
rect 373936 29993 373986 30993
rect 374095 29993 374145 30993
rect 374245 29993 374295 30993
rect 374410 30961 374620 30973
rect 376726 30961 376936 30973
rect 374414 30958 374616 30961
rect 376730 30958 376932 30961
rect 374425 30788 374605 30958
rect 374785 30788 374815 30793
rect 374871 30788 374901 30793
rect 376445 30788 376475 30793
rect 376531 30788 376561 30793
rect 376741 30788 376921 30958
rect 374410 30773 374620 30788
rect 374770 30773 374830 30788
rect 374856 30773 374916 30788
rect 376430 30773 376490 30788
rect 376516 30773 376576 30788
rect 376726 30773 376936 30788
rect 374410 30701 374620 30713
rect 374770 30701 374830 30713
rect 374856 30701 374916 30713
rect 376430 30701 376490 30713
rect 376516 30701 376576 30713
rect 376726 30701 376936 30713
rect 374414 30698 374616 30701
rect 374774 30698 374826 30701
rect 374860 30698 374912 30701
rect 376434 30698 376486 30701
rect 376520 30698 376572 30701
rect 376730 30698 376932 30701
rect 374425 30528 374605 30698
rect 374785 30528 374815 30698
rect 374871 30528 374901 30698
rect 376445 30528 376475 30698
rect 376531 30528 376561 30698
rect 376741 30528 376921 30698
rect 374410 30513 374620 30528
rect 374770 30513 374830 30528
rect 374856 30513 374916 30528
rect 376430 30513 376490 30528
rect 376516 30513 376576 30528
rect 376726 30513 376936 30528
rect 374410 30441 374620 30453
rect 374770 30441 374830 30453
rect 374856 30441 374916 30453
rect 376430 30441 376490 30453
rect 376516 30441 376576 30453
rect 376726 30441 376936 30453
rect 374414 30438 374616 30441
rect 374774 30438 374826 30441
rect 374860 30438 374912 30441
rect 376434 30438 376486 30441
rect 376520 30438 376572 30441
rect 376730 30438 376932 30441
rect 374425 30268 374605 30438
rect 374785 30268 374815 30438
rect 374871 30268 374901 30438
rect 376445 30268 376475 30438
rect 376531 30268 376561 30438
rect 376741 30268 376921 30438
rect 374410 30253 374620 30268
rect 374770 30253 374830 30268
rect 374856 30253 374916 30268
rect 376430 30253 376490 30268
rect 376516 30253 376576 30268
rect 376726 30253 376936 30268
rect 377051 29993 377101 30993
rect 377201 29993 377251 30993
rect 377360 29993 377410 30993
rect 377510 29993 377560 30993
rect 379107 30907 379141 30911
rect 379178 30907 379212 30911
rect 379249 30907 379283 30911
rect 379083 30891 379335 30907
rect 379107 30887 379141 30891
rect 379178 30887 379212 30891
rect 379249 30887 379283 30891
rect 379083 30881 379305 30887
rect 379083 30867 379307 30881
rect 379296 30857 379307 30867
rect 379259 30833 379283 30857
rect 379320 30833 379344 30857
rect 377649 30171 377699 30771
rect 377819 30171 377875 30771
rect 377995 30171 378045 30771
rect 412150 30245 412200 30845
rect 412320 30245 412376 30845
rect 412496 30245 412552 30845
rect 412672 30245 412722 30845
rect 413229 30558 413409 30580
rect 413214 30543 413409 30558
rect 412978 30430 413188 30445
rect 413214 30430 413409 30445
rect 412993 30260 413173 30430
rect 413229 30260 413409 30430
rect 412982 30257 413184 30260
rect 413218 30257 413409 30260
rect 412978 30245 413188 30257
rect 413214 30245 413409 30257
rect 425510 29993 425560 30993
rect 427107 30907 427141 30911
rect 427178 30907 427212 30911
rect 427249 30907 427283 30911
rect 427083 30891 427335 30907
rect 427107 30887 427141 30891
rect 427178 30887 427212 30891
rect 427249 30887 427283 30891
rect 427083 30881 427305 30887
rect 427083 30867 427307 30881
rect 427296 30857 427307 30867
rect 427259 30833 427283 30857
rect 427320 30833 427344 30857
rect 425649 30171 425699 30771
rect 425819 30171 425875 30771
rect 425995 30171 426045 30771
rect 464150 30245 464200 30845
rect 464320 30245 464376 30845
rect 464496 30245 464552 30845
rect 464672 30245 464722 30845
rect 466203 30697 466227 30731
rect 466203 30626 466227 30660
rect 465229 30558 465409 30580
rect 465214 30543 465424 30558
rect 466203 30555 466227 30589
rect 466203 30484 466227 30518
rect 464978 30430 465188 30445
rect 465214 30430 465424 30445
rect 464993 30260 465173 30430
rect 465229 30260 465409 30430
rect 466203 30413 466227 30447
rect 466203 30342 466227 30376
rect 466203 30271 466227 30305
rect 464982 30257 465184 30260
rect 465218 30257 465420 30260
rect 464978 30245 465188 30257
rect 465214 30245 465424 30257
rect 466834 30135 466884 30735
rect 467004 30135 467132 30735
rect 467180 30135 467236 30735
rect 467356 30135 467484 30735
rect 467532 30135 467588 30735
rect 467708 30135 467836 30735
rect 467884 30135 467940 30735
rect 468060 30135 468188 30735
rect 468236 30135 468364 30735
rect 468412 30135 468540 30735
rect 468588 30135 468716 30735
rect 468764 30135 468892 30735
rect 468940 30135 468996 30735
rect 469116 30135 469244 30735
rect 469292 30135 469420 30735
rect 469468 30135 469596 30735
rect 469644 30135 469772 30735
rect 469820 30135 469948 30735
rect 469996 30135 470046 30735
rect 470112 30135 470162 30735
rect 470282 30135 470410 30735
rect 470458 30135 470514 30735
rect 470634 30135 470762 30735
rect 470810 30135 470860 30735
rect 470926 30135 470976 30735
rect 471096 30135 471224 30735
rect 471272 30135 471400 30735
rect 471448 30135 471576 30735
rect 471624 30135 471680 30735
rect 471800 30135 471850 30735
rect 471916 30135 471966 30735
rect 472086 30135 472142 30735
rect 472262 30135 472312 30735
rect 472446 30718 472456 30721
rect 472446 30027 472472 30718
rect 473301 30171 473351 30771
rect 473471 30171 473527 30771
rect 473647 30171 473697 30771
rect 466723 30015 472472 30027
rect 473786 29993 473836 30993
rect 473936 29993 473986 30993
rect 474095 29993 474145 30993
rect 474245 29993 474295 30993
rect 474410 30961 474620 30973
rect 476726 30961 476936 30973
rect 474414 30958 474616 30961
rect 476730 30958 476932 30961
rect 474425 30788 474605 30958
rect 474785 30788 474815 30793
rect 474871 30788 474901 30793
rect 476445 30788 476475 30793
rect 476531 30788 476561 30793
rect 476741 30788 476921 30958
rect 474410 30773 474620 30788
rect 474770 30773 474830 30788
rect 474856 30773 474916 30788
rect 476430 30773 476490 30788
rect 476516 30773 476576 30788
rect 476726 30773 476936 30788
rect 474410 30701 474620 30713
rect 474770 30701 474830 30713
rect 474856 30701 474916 30713
rect 476430 30701 476490 30713
rect 476516 30701 476576 30713
rect 476726 30701 476936 30713
rect 474414 30698 474616 30701
rect 474774 30698 474826 30701
rect 474860 30698 474912 30701
rect 476434 30698 476486 30701
rect 476520 30698 476572 30701
rect 476730 30698 476932 30701
rect 474425 30528 474605 30698
rect 474785 30528 474815 30698
rect 474871 30528 474901 30698
rect 476445 30528 476475 30698
rect 476531 30528 476561 30698
rect 476741 30528 476921 30698
rect 474410 30513 474620 30528
rect 474770 30513 474830 30528
rect 474856 30513 474916 30528
rect 476430 30513 476490 30528
rect 476516 30513 476576 30528
rect 476726 30513 476936 30528
rect 474410 30441 474620 30453
rect 474770 30441 474830 30453
rect 474856 30441 474916 30453
rect 476430 30441 476490 30453
rect 476516 30441 476576 30453
rect 476726 30441 476936 30453
rect 474414 30438 474616 30441
rect 474774 30438 474826 30441
rect 474860 30438 474912 30441
rect 476434 30438 476486 30441
rect 476520 30438 476572 30441
rect 476730 30438 476932 30441
rect 474425 30268 474605 30438
rect 474785 30268 474815 30438
rect 474871 30268 474901 30438
rect 476445 30268 476475 30438
rect 476531 30268 476561 30438
rect 476741 30268 476921 30438
rect 474410 30253 474620 30268
rect 474770 30253 474830 30268
rect 474856 30253 474916 30268
rect 476430 30253 476490 30268
rect 476516 30253 476576 30268
rect 476726 30253 476936 30268
rect 477051 29993 477101 30993
rect 477201 29993 477251 30993
rect 477360 29993 477410 30993
rect 477510 29993 477560 30993
rect 479107 30907 479141 30911
rect 479178 30907 479212 30911
rect 479249 30907 479283 30911
rect 479083 30891 479335 30907
rect 479107 30887 479141 30891
rect 479178 30887 479212 30891
rect 479249 30887 479283 30891
rect 479083 30881 479305 30887
rect 479083 30867 479307 30881
rect 479296 30857 479307 30867
rect 479259 30833 479283 30857
rect 479320 30833 479344 30857
rect 477649 30171 477699 30771
rect 477819 30171 477875 30771
rect 477995 30171 478045 30771
rect 516150 30245 516200 30845
rect 516320 30245 516376 30845
rect 516496 30245 516552 30845
rect 516672 30245 516722 30845
rect 517229 30558 517409 30580
rect 517214 30543 517409 30558
rect 516978 30430 517188 30445
rect 517214 30430 517409 30445
rect 516993 30260 517173 30430
rect 517229 30260 517409 30430
rect 516982 30257 517184 30260
rect 517218 30257 517409 30260
rect 516978 30245 517188 30257
rect 517214 30245 517409 30257
rect 529510 29993 529560 30993
rect 531107 30907 531141 30911
rect 531178 30907 531212 30911
rect 531249 30907 531283 30911
rect 531083 30891 531335 30907
rect 531107 30887 531141 30891
rect 531178 30887 531212 30891
rect 531249 30887 531283 30891
rect 531083 30881 531305 30887
rect 531083 30867 531307 30881
rect 531296 30857 531307 30867
rect 531259 30833 531283 30857
rect 531320 30833 531344 30857
rect 529649 30171 529699 30771
rect 529819 30171 529875 30771
rect 529995 30171 530045 30771
rect 564150 30245 564200 30845
rect 564320 30245 564376 30845
rect 564496 30245 564552 30845
rect 564672 30245 564722 30845
rect 566203 30697 566227 30731
rect 566203 30626 566227 30660
rect 565229 30558 565409 30580
rect 565214 30543 565424 30558
rect 566203 30555 566227 30589
rect 566203 30484 566227 30518
rect 564978 30430 565188 30445
rect 565214 30430 565424 30445
rect 564993 30260 565173 30430
rect 565229 30260 565409 30430
rect 566203 30413 566227 30447
rect 566203 30342 566227 30376
rect 566203 30271 566227 30305
rect 564982 30257 565184 30260
rect 565218 30257 565420 30260
rect 564978 30245 565188 30257
rect 565214 30245 565424 30257
rect 566834 30135 566884 30735
rect 567004 30135 567132 30735
rect 567180 30135 567236 30735
rect 567356 30135 567484 30735
rect 567532 30135 567588 30735
rect 567708 30135 567836 30735
rect 567884 30135 567940 30735
rect 568060 30135 568188 30735
rect 568236 30135 568364 30735
rect 568412 30135 568540 30735
rect 568588 30135 568716 30735
rect 568764 30135 568892 30735
rect 568940 30135 568996 30735
rect 569116 30135 569244 30735
rect 569292 30135 569420 30735
rect 569468 30135 569596 30735
rect 569644 30135 569772 30735
rect 569820 30135 569948 30735
rect 569996 30135 570046 30735
rect 570112 30135 570162 30735
rect 570282 30135 570410 30735
rect 570458 30135 570514 30735
rect 570634 30135 570762 30735
rect 570810 30135 570860 30735
rect 570926 30135 570976 30735
rect 571096 30135 571224 30735
rect 571272 30135 571400 30735
rect 571448 30135 571576 30735
rect 571624 30135 571680 30735
rect 571800 30135 571850 30735
rect 571916 30135 571966 30735
rect 572086 30135 572142 30735
rect 572262 30135 572312 30735
rect 572446 30718 572456 30721
rect 572446 30027 572472 30718
rect 573301 30171 573351 30771
rect 573471 30171 573527 30771
rect 573647 30171 573697 30771
rect 566723 30015 572472 30027
rect 573786 29993 573836 30993
rect 573936 29993 573986 30993
rect 574095 29993 574145 30993
rect 574245 29993 574295 30993
rect 574410 30961 574620 30973
rect 576726 30961 576936 30973
rect 574414 30958 574616 30961
rect 576730 30958 576932 30961
rect 574425 30788 574605 30958
rect 574785 30788 574815 30793
rect 574871 30788 574901 30793
rect 576445 30788 576475 30793
rect 576531 30788 576561 30793
rect 576741 30788 576921 30958
rect 574410 30773 574620 30788
rect 574770 30773 574830 30788
rect 574856 30773 574916 30788
rect 576430 30773 576490 30788
rect 576516 30773 576576 30788
rect 576726 30773 576936 30788
rect 574410 30701 574620 30713
rect 574770 30701 574830 30713
rect 574856 30701 574916 30713
rect 576430 30701 576490 30713
rect 576516 30701 576576 30713
rect 576726 30701 576936 30713
rect 574414 30698 574616 30701
rect 574774 30698 574826 30701
rect 574860 30698 574912 30701
rect 576434 30698 576486 30701
rect 576520 30698 576572 30701
rect 576730 30698 576932 30701
rect 574425 30528 574605 30698
rect 574785 30528 574815 30698
rect 574871 30528 574901 30698
rect 576445 30528 576475 30698
rect 576531 30528 576561 30698
rect 576741 30528 576921 30698
rect 574410 30513 574620 30528
rect 574770 30513 574830 30528
rect 574856 30513 574916 30528
rect 576430 30513 576490 30528
rect 576516 30513 576576 30528
rect 576726 30513 576936 30528
rect 574410 30441 574620 30453
rect 574770 30441 574830 30453
rect 574856 30441 574916 30453
rect 576430 30441 576490 30453
rect 576516 30441 576576 30453
rect 576726 30441 576936 30453
rect 574414 30438 574616 30441
rect 574774 30438 574826 30441
rect 574860 30438 574912 30441
rect 576434 30438 576486 30441
rect 576520 30438 576572 30441
rect 576730 30438 576932 30441
rect 574425 30268 574605 30438
rect 574785 30268 574815 30438
rect 574871 30268 574901 30438
rect 576445 30268 576475 30438
rect 576531 30268 576561 30438
rect 576741 30268 576921 30438
rect 574410 30253 574620 30268
rect 574770 30253 574830 30268
rect 574856 30253 574916 30268
rect 576430 30253 576490 30268
rect 576516 30253 576576 30268
rect 576726 30253 576936 30268
rect 577051 29993 577101 30993
rect 577201 29993 577251 30993
rect 577360 29993 577410 30993
rect 577510 29993 577560 30993
rect 579107 30907 579141 30911
rect 579178 30907 579212 30911
rect 579249 30907 579283 30911
rect 579083 30891 579335 30907
rect 579107 30887 579141 30891
rect 579178 30887 579212 30891
rect 579249 30887 579283 30891
rect 579083 30881 579305 30887
rect 579083 30867 579307 30881
rect 579296 30857 579307 30867
rect 579259 30833 579283 30857
rect 579320 30833 579344 30857
rect 577649 30171 577699 30771
rect 577819 30171 577875 30771
rect 577995 30171 578045 30771
rect 366162 29955 366203 29961
rect 466162 29955 466203 29961
rect 566162 29955 566203 29961
rect 366162 29931 366186 29939
rect 466162 29931 466186 29939
rect 566162 29931 566186 29939
rect 366138 29891 366162 29915
rect 367872 29880 367906 29914
rect 368475 29890 368533 29914
rect 368499 29880 368533 29890
rect 370881 29880 370915 29914
rect 466138 29891 466162 29915
rect 467872 29880 467906 29914
rect 468475 29890 468533 29914
rect 468499 29880 468533 29890
rect 470881 29880 470915 29914
rect 566138 29891 566162 29915
rect 567872 29880 567906 29914
rect 568475 29890 568533 29914
rect 568499 29880 568533 29890
rect 570881 29880 570915 29914
rect 368496 29802 368509 29826
rect 370871 29802 370883 29826
rect 468496 29802 468509 29826
rect 470871 29802 470883 29826
rect 568496 29802 568509 29826
rect 570871 29802 570883 29826
rect 368461 29778 368485 29802
rect 368520 29778 368544 29802
rect 370835 29778 370859 29802
rect 370895 29778 370919 29802
rect 468461 29778 468485 29802
rect 468520 29778 468544 29802
rect 470835 29778 470859 29802
rect 470895 29778 470919 29802
rect 568461 29778 568485 29802
rect 568520 29778 568544 29802
rect 570835 29778 570859 29802
rect 570895 29778 570919 29802
rect 56370 29340 57370 29390
rect 108370 29340 109370 29390
rect 160370 29340 161280 29390
rect 212370 29340 213370 29390
rect 260370 29340 261370 29390
rect 312370 29340 313370 29390
rect 364370 29340 365370 29390
rect 412370 29340 413370 29390
rect 464370 29340 465370 29390
rect 516370 29340 517370 29390
rect 564370 29340 565370 29390
rect 56370 29184 57260 29312
rect 108370 29184 109260 29312
rect 160370 29184 161260 29312
rect 212370 29184 213260 29312
rect 260370 29184 261260 29312
rect 312370 29184 313260 29312
rect 364370 29184 365370 29312
rect 412370 29184 413260 29312
rect 464370 29184 465370 29312
rect 516370 29184 517260 29312
rect 564370 29184 565370 29312
rect 56370 29028 57260 29156
rect 108370 29028 109260 29156
rect 160370 29028 161260 29156
rect 212370 29028 213260 29156
rect 260370 29028 261260 29156
rect 312370 29028 313260 29156
rect 364370 29028 365370 29156
rect 412370 29028 413260 29156
rect 464370 29028 465370 29156
rect 516370 29028 517260 29156
rect 564370 29028 565370 29156
rect 56370 28872 57260 29000
rect 108370 28872 109260 29000
rect 160370 28872 161260 29000
rect 212370 28872 213260 29000
rect 260370 28872 261260 29000
rect 312370 28872 313260 29000
rect 364370 28872 365370 29000
rect 412370 28872 413260 29000
rect 464370 28872 465370 29000
rect 516370 28872 517260 29000
rect 564370 28872 565370 29000
rect 56370 28716 57260 28844
rect 108370 28716 109260 28844
rect 160370 28716 161260 28844
rect 212370 28716 213260 28844
rect 260370 28716 261260 28844
rect 312370 28716 313260 28844
rect 364370 28716 365370 28844
rect 371498 28716 371561 28717
rect 56370 28560 57260 28688
rect 108370 28560 109260 28688
rect 160370 28560 161260 28688
rect 212370 28560 213260 28688
rect 260370 28560 261260 28688
rect 312370 28560 313260 28688
rect 364370 28560 365370 28688
rect 371498 28683 371527 28716
rect 371532 28683 371561 28716
rect 371596 28683 371630 28717
rect 371665 28683 371699 28717
rect 371734 28683 371768 28717
rect 371803 28683 371837 28717
rect 371872 28683 371906 28717
rect 371941 28683 371975 28717
rect 372010 28683 372044 28717
rect 372079 28683 372113 28717
rect 372148 28683 372182 28717
rect 372217 28683 372251 28717
rect 372286 28683 372320 28717
rect 372355 28683 372389 28717
rect 372424 28683 372458 28717
rect 372493 28683 372527 28717
rect 372562 28683 372596 28717
rect 372631 28683 372665 28717
rect 372700 28683 372734 28717
rect 372769 28683 372803 28717
rect 372838 28683 372872 28717
rect 372907 28683 372941 28717
rect 372976 28683 373010 28717
rect 373045 28683 373079 28717
rect 373114 28683 373148 28717
rect 373183 28683 373217 28717
rect 373252 28683 373286 28717
rect 373321 28683 373355 28717
rect 373390 28683 373424 28717
rect 373459 28683 373493 28717
rect 373528 28683 373562 28717
rect 373597 28683 373631 28717
rect 412370 28716 413260 28844
rect 464370 28716 465370 28844
rect 471498 28716 471561 28717
rect 371532 28682 371566 28683
rect 367325 28610 367525 28660
rect 367873 28610 368073 28660
rect 370354 28647 370364 28671
rect 370399 28647 370433 28671
rect 370468 28647 370502 28671
rect 370537 28647 370571 28671
rect 370606 28647 370640 28671
rect 370675 28647 370709 28671
rect 370744 28647 370778 28671
rect 370813 28647 370847 28671
rect 370882 28647 370916 28671
rect 370951 28647 370985 28671
rect 371020 28647 371054 28671
rect 371089 28647 371123 28671
rect 371158 28647 371192 28671
rect 371227 28647 371261 28671
rect 371296 28647 371330 28671
rect 371365 28647 371399 28671
rect 371434 28647 371468 28671
rect 371503 28647 371532 28671
rect 373650 28647 373677 28671
rect 56370 28404 57260 28532
rect 58103 28396 58520 28446
rect 108370 28404 109260 28532
rect 110103 28396 110520 28446
rect 160370 28404 161260 28532
rect 212370 28404 213260 28532
rect 214103 28396 214520 28446
rect 260370 28404 261260 28532
rect 312370 28404 313260 28532
rect 314103 28396 314520 28446
rect 364370 28404 365370 28532
rect 366561 28446 366645 28449
rect 366893 28446 366977 28449
rect 366103 28396 367103 28446
rect 367325 28434 367525 28562
rect 367873 28434 368073 28562
rect 412370 28560 413260 28688
rect 464370 28560 465370 28688
rect 471498 28683 471527 28716
rect 471532 28683 471561 28716
rect 471596 28683 471630 28717
rect 471665 28683 471699 28717
rect 471734 28683 471768 28717
rect 471803 28683 471837 28717
rect 471872 28683 471906 28717
rect 471941 28683 471975 28717
rect 472010 28683 472044 28717
rect 472079 28683 472113 28717
rect 472148 28683 472182 28717
rect 472217 28683 472251 28717
rect 472286 28683 472320 28717
rect 472355 28683 472389 28717
rect 472424 28683 472458 28717
rect 472493 28683 472527 28717
rect 472562 28683 472596 28717
rect 472631 28683 472665 28717
rect 472700 28683 472734 28717
rect 472769 28683 472803 28717
rect 472838 28683 472872 28717
rect 472907 28683 472941 28717
rect 472976 28683 473010 28717
rect 473045 28683 473079 28717
rect 473114 28683 473148 28717
rect 473183 28683 473217 28717
rect 473252 28683 473286 28717
rect 473321 28683 473355 28717
rect 473390 28683 473424 28717
rect 473459 28683 473493 28717
rect 473528 28683 473562 28717
rect 473597 28683 473631 28717
rect 516370 28716 517260 28844
rect 564370 28716 565370 28844
rect 571498 28716 571561 28717
rect 471532 28682 471566 28683
rect 467325 28610 467525 28660
rect 467873 28610 468073 28660
rect 470354 28647 470364 28671
rect 470399 28647 470433 28671
rect 470468 28647 470502 28671
rect 470537 28647 470571 28671
rect 470606 28647 470640 28671
rect 470675 28647 470709 28671
rect 470744 28647 470778 28671
rect 470813 28647 470847 28671
rect 470882 28647 470916 28671
rect 470951 28647 470985 28671
rect 471020 28647 471054 28671
rect 471089 28647 471123 28671
rect 471158 28647 471192 28671
rect 471227 28647 471261 28671
rect 471296 28647 471330 28671
rect 471365 28647 471399 28671
rect 471434 28647 471468 28671
rect 471503 28647 471532 28671
rect 473650 28647 473677 28671
rect 368421 28446 368505 28449
rect 368753 28446 368837 28449
rect 368295 28396 369295 28446
rect 412370 28404 413260 28532
rect 414103 28396 414520 28446
rect 464370 28404 465370 28532
rect 466561 28446 466645 28449
rect 466893 28446 466977 28449
rect 466103 28396 467103 28446
rect 467325 28434 467525 28562
rect 467873 28434 468073 28562
rect 516370 28560 517260 28688
rect 564370 28560 565370 28688
rect 571498 28683 571527 28716
rect 571532 28683 571561 28716
rect 571596 28683 571630 28717
rect 571665 28683 571699 28717
rect 571734 28683 571768 28717
rect 571803 28683 571837 28717
rect 571872 28683 571906 28717
rect 571941 28683 571975 28717
rect 572010 28683 572044 28717
rect 572079 28683 572113 28717
rect 572148 28683 572182 28717
rect 572217 28683 572251 28717
rect 572286 28683 572320 28717
rect 572355 28683 572389 28717
rect 572424 28683 572458 28717
rect 572493 28683 572527 28717
rect 572562 28683 572596 28717
rect 572631 28683 572665 28717
rect 572700 28683 572734 28717
rect 572769 28683 572803 28717
rect 572838 28683 572872 28717
rect 572907 28683 572941 28717
rect 572976 28683 573010 28717
rect 573045 28683 573079 28717
rect 573114 28683 573148 28717
rect 573183 28683 573217 28717
rect 573252 28683 573286 28717
rect 573321 28683 573355 28717
rect 573390 28683 573424 28717
rect 573459 28683 573493 28717
rect 573528 28683 573562 28717
rect 573597 28683 573631 28717
rect 571532 28682 571566 28683
rect 567325 28610 567525 28660
rect 567873 28610 568073 28660
rect 570354 28647 570364 28671
rect 570399 28647 570433 28671
rect 570468 28647 570502 28671
rect 570537 28647 570571 28671
rect 570606 28647 570640 28671
rect 570675 28647 570709 28671
rect 570744 28647 570778 28671
rect 570813 28647 570847 28671
rect 570882 28647 570916 28671
rect 570951 28647 570985 28671
rect 571020 28647 571054 28671
rect 571089 28647 571123 28671
rect 571158 28647 571192 28671
rect 571227 28647 571261 28671
rect 571296 28647 571330 28671
rect 571365 28647 571399 28671
rect 571434 28647 571468 28671
rect 571503 28647 571532 28671
rect 573650 28647 573677 28671
rect 468421 28446 468505 28449
rect 468753 28446 468837 28449
rect 468295 28396 469295 28446
rect 516370 28404 517260 28532
rect 518103 28396 518520 28446
rect 564370 28404 565370 28532
rect 566561 28446 566645 28449
rect 566893 28446 566977 28449
rect 566103 28396 567103 28446
rect 567325 28434 567525 28562
rect 567873 28434 568073 28562
rect 568421 28446 568505 28449
rect 568753 28446 568837 28449
rect 568295 28396 569295 28446
rect 56370 28248 57260 28376
rect 58103 28240 58520 28296
rect 108370 28248 109260 28376
rect 110103 28240 110520 28296
rect 160370 28248 161260 28376
rect 212370 28248 213260 28376
rect 214103 28240 214520 28296
rect 260370 28248 261260 28376
rect 312370 28248 313260 28376
rect 314103 28240 314520 28296
rect 364370 28248 365370 28376
rect 366103 28240 367103 28296
rect 367325 28258 367525 28314
rect 367873 28258 368073 28314
rect 368295 28240 369295 28296
rect 56370 28092 57260 28220
rect 58103 28084 58520 28140
rect 108370 28092 109260 28220
rect 110103 28084 110520 28140
rect 160370 28092 161260 28220
rect 212370 28092 213260 28220
rect 214103 28084 214520 28140
rect 260370 28092 261260 28220
rect 312370 28092 313260 28220
rect 314103 28084 314520 28140
rect 364370 28092 365370 28220
rect 366103 28084 367103 28140
rect 367325 28082 367525 28210
rect 367873 28082 368073 28210
rect 368295 28084 369295 28140
rect 56370 27936 57260 28064
rect 58103 27928 58520 27984
rect 108370 27936 109260 28064
rect 110103 27928 110520 27984
rect 160370 27936 161260 28064
rect 212370 27936 213260 28064
rect 214103 27928 214520 27984
rect 260370 27936 261260 28064
rect 312370 27936 313260 28064
rect 314103 27928 314520 27984
rect 364370 27936 365370 28064
rect 366103 27928 367103 27984
rect 367325 27912 367525 27962
rect 367873 27951 368073 27962
rect 367869 27917 368073 27951
rect 368295 27928 369295 27984
rect 367441 27909 367525 27912
rect 367873 27912 368073 27917
rect 367873 27909 367957 27912
rect 56370 27780 57260 27908
rect 58103 27772 58520 27828
rect 108370 27780 109260 27908
rect 110103 27772 110520 27828
rect 160370 27780 161260 27908
rect 212370 27780 213260 27908
rect 214103 27772 214520 27828
rect 260370 27780 261260 27908
rect 312370 27780 313260 27908
rect 314103 27772 314520 27828
rect 364370 27780 365370 27908
rect 366103 27772 367103 27828
rect 368295 27772 369295 27828
rect 56370 27624 57260 27752
rect 58103 27622 58520 27672
rect 108370 27624 109260 27752
rect 110103 27622 110520 27672
rect 160370 27624 161260 27752
rect 212370 27624 213260 27752
rect 214103 27622 214520 27672
rect 260370 27624 261260 27752
rect 312370 27624 313260 27752
rect 314103 27622 314520 27672
rect 364370 27624 365370 27752
rect 375672 27691 375722 28291
rect 375822 27691 375950 28291
rect 375978 27691 376106 28291
rect 376134 27691 376190 28291
rect 376290 27691 376418 28291
rect 376446 27691 376574 28291
rect 376602 27691 376652 28291
rect 376732 27691 376782 28291
rect 376882 27691 376932 28291
rect 412370 28248 413260 28376
rect 414103 28240 414520 28296
rect 464370 28248 465370 28376
rect 466103 28240 467103 28296
rect 467325 28258 467525 28314
rect 467873 28258 468073 28314
rect 468295 28240 469295 28296
rect 412370 28092 413260 28220
rect 414103 28084 414520 28140
rect 464370 28092 465370 28220
rect 466103 28084 467103 28140
rect 467325 28082 467525 28210
rect 467873 28082 468073 28210
rect 468295 28084 469295 28140
rect 412370 27936 413260 28064
rect 414103 27928 414520 27984
rect 464370 27936 465370 28064
rect 466103 27928 467103 27984
rect 467325 27912 467525 27962
rect 467873 27951 468073 27962
rect 467869 27917 468073 27951
rect 468295 27928 469295 27984
rect 467441 27909 467525 27912
rect 467873 27912 468073 27917
rect 467873 27909 467957 27912
rect 412370 27780 413260 27908
rect 414103 27772 414520 27828
rect 464370 27780 465370 27908
rect 466103 27772 467103 27828
rect 468295 27772 469295 27828
rect 366103 27622 367103 27672
rect 368295 27622 369295 27672
rect 412370 27624 413260 27752
rect 414103 27622 414520 27672
rect 464370 27624 465370 27752
rect 475672 27691 475722 28291
rect 475822 27691 475950 28291
rect 475978 27691 476106 28291
rect 476134 27691 476190 28291
rect 476290 27691 476418 28291
rect 476446 27691 476574 28291
rect 476602 27691 476652 28291
rect 476732 27691 476782 28291
rect 476882 27691 476932 28291
rect 516370 28248 517260 28376
rect 518103 28240 518520 28296
rect 564370 28248 565370 28376
rect 566103 28240 567103 28296
rect 567325 28258 567525 28314
rect 567873 28258 568073 28314
rect 568295 28240 569295 28296
rect 516370 28092 517260 28220
rect 518103 28084 518520 28140
rect 564370 28092 565370 28220
rect 566103 28084 567103 28140
rect 567325 28082 567525 28210
rect 567873 28082 568073 28210
rect 568295 28084 569295 28140
rect 516370 27936 517260 28064
rect 518103 27928 518520 27984
rect 564370 27936 565370 28064
rect 566103 27928 567103 27984
rect 567325 27912 567525 27962
rect 567873 27951 568073 27962
rect 567869 27917 568073 27951
rect 568295 27928 569295 27984
rect 567441 27909 567525 27912
rect 567873 27912 568073 27917
rect 567873 27909 567957 27912
rect 516370 27780 517260 27908
rect 518103 27772 518520 27828
rect 564370 27780 565370 27908
rect 566103 27772 567103 27828
rect 568295 27772 569295 27828
rect 466103 27622 467103 27672
rect 468295 27622 469295 27672
rect 516370 27624 517260 27752
rect 518103 27622 518520 27672
rect 564370 27624 565370 27752
rect 575672 27691 575722 28291
rect 575822 27691 575950 28291
rect 575978 27691 576106 28291
rect 576134 27691 576190 28291
rect 576290 27691 576418 28291
rect 576446 27691 576574 28291
rect 576602 27691 576652 28291
rect 576732 27691 576782 28291
rect 576882 27691 576932 28291
rect 566103 27622 567103 27672
rect 568295 27622 569295 27672
rect 56370 27468 57260 27596
rect 108370 27468 109260 27596
rect 160370 27468 161260 27596
rect 212370 27468 213260 27596
rect 260370 27468 261260 27596
rect 312370 27468 313260 27596
rect 364370 27468 365370 27596
rect 412370 27468 413260 27596
rect 464370 27468 465370 27596
rect 516370 27468 517260 27596
rect 564370 27468 565370 27596
rect 56370 27312 57260 27440
rect 108370 27312 109260 27440
rect 160370 27312 161260 27440
rect 212370 27312 213260 27440
rect 260370 27312 261260 27440
rect 312370 27312 313260 27440
rect 364370 27312 365370 27440
rect 367786 27358 367820 27362
rect 369194 27358 369228 27362
rect 367778 27274 367831 27358
rect 56370 27162 57370 27212
rect 108370 27162 109370 27212
rect 160370 27162 161280 27212
rect 212370 27162 213370 27212
rect 260370 27162 261370 27212
rect 312370 27162 313370 27212
rect 364370 27162 365370 27212
rect 367781 27158 367831 27274
rect 367951 27158 368079 27358
rect 368127 27158 368183 27358
rect 368303 27158 368431 27358
rect 368479 27158 368535 27358
rect 368655 27158 368783 27358
rect 368831 27158 368887 27358
rect 369007 27158 369135 27358
rect 369183 27274 369236 27358
rect 412370 27312 413260 27440
rect 464370 27312 465370 27440
rect 467786 27358 467820 27362
rect 469194 27358 469228 27362
rect 467778 27274 467831 27358
rect 369183 27158 369233 27274
rect 412370 27162 413370 27212
rect 464370 27162 465370 27212
rect 467781 27158 467831 27274
rect 467951 27158 468079 27358
rect 468127 27158 468183 27358
rect 468303 27158 468431 27358
rect 468479 27158 468535 27358
rect 468655 27158 468783 27358
rect 468831 27158 468887 27358
rect 469007 27158 469135 27358
rect 469183 27274 469236 27358
rect 516370 27312 517260 27440
rect 564370 27312 565370 27440
rect 567786 27358 567820 27362
rect 569194 27358 569228 27362
rect 567778 27274 567831 27358
rect 469183 27158 469233 27274
rect 516370 27162 517370 27212
rect 564370 27162 565370 27212
rect 567781 27158 567831 27274
rect 567951 27158 568079 27358
rect 568127 27158 568183 27358
rect 568303 27158 568431 27358
rect 568479 27158 568535 27358
rect 568655 27158 568783 27358
rect 568831 27158 568887 27358
rect 569007 27158 569135 27358
rect 569183 27274 569236 27358
rect 569183 27158 569233 27274
rect 366185 26478 366491 26648
rect 56427 25725 56477 26325
rect 56577 25725 56627 26325
rect 56699 25725 56749 26325
rect 56849 25725 56899 26325
rect 56975 25725 57025 26325
rect 57125 25725 57175 26325
rect 57247 25725 57297 26325
rect 57397 25725 57447 26325
rect 108427 25725 108477 26325
rect 108577 25725 108627 26325
rect 108699 25725 108749 26325
rect 108849 25725 108899 26325
rect 108975 25725 109025 26325
rect 109125 25725 109175 26325
rect 109247 25725 109297 26325
rect 109397 25725 109447 26325
rect 160427 25725 160477 26325
rect 160577 25725 160627 26325
rect 160699 25725 160749 26325
rect 160849 25725 160899 26325
rect 160975 25725 161025 26325
rect 161125 25725 161175 26325
rect 161247 25725 161280 26325
rect 212427 25725 212477 26325
rect 212577 25725 212627 26325
rect 212699 25725 212749 26325
rect 212849 25725 212899 26325
rect 212975 25725 213025 26325
rect 213125 25725 213175 26325
rect 213247 25725 213297 26325
rect 213397 25725 213447 26325
rect 260427 25725 260477 26325
rect 260577 25725 260627 26325
rect 260699 25725 260749 26325
rect 260849 25725 260899 26325
rect 260975 25725 261025 26325
rect 261125 25725 261175 26325
rect 261247 25725 261297 26325
rect 261397 25725 261447 26325
rect 312427 25725 312477 26325
rect 312577 25725 312627 26325
rect 312699 25725 312749 26325
rect 312849 25725 312899 26325
rect 312975 25725 313025 26325
rect 313125 25725 313175 26325
rect 313247 25725 313297 26325
rect 313397 25725 313447 26325
rect 364427 25725 364477 26325
rect 364577 25725 364627 26325
rect 364699 25725 364749 26325
rect 364849 25725 364899 26325
rect 364975 25725 365025 26325
rect 365125 25725 365175 26325
rect 365247 25725 365297 26325
rect 365397 25725 365447 26325
rect 367632 25936 367682 26936
rect 367782 25936 367838 26936
rect 367938 25936 367994 26936
rect 368094 25936 368150 26936
rect 368250 26810 368300 26936
rect 368714 26810 368764 26936
rect 368250 26726 368303 26810
rect 368711 26726 368764 26810
rect 368250 26477 368300 26726
rect 368714 26477 368764 26726
rect 368250 26393 368303 26477
rect 368711 26393 368764 26477
rect 368250 25936 368300 26393
rect 368714 25936 368764 26393
rect 368864 25936 368920 26936
rect 369020 25936 369076 26936
rect 369176 25936 369232 26936
rect 369332 25936 369382 26936
rect 376307 26490 376360 26690
rect 376460 26490 376516 26690
rect 376616 26490 376666 26690
rect 377016 26490 377066 26690
rect 377166 26490 377222 26690
rect 377322 26490 377372 26690
rect 466185 26478 466491 26648
rect 377661 26348 377695 26372
rect 377730 26348 377764 26372
rect 412427 25725 412477 26325
rect 412577 25725 412627 26325
rect 412699 25725 412749 26325
rect 412849 25725 412899 26325
rect 412975 25725 413025 26325
rect 413125 25725 413175 26325
rect 413247 25725 413297 26325
rect 413397 25725 413447 26325
rect 464427 25725 464477 26325
rect 464577 25725 464627 26325
rect 464699 25725 464749 26325
rect 464849 25725 464899 26325
rect 464975 25725 465025 26325
rect 465125 25725 465175 26325
rect 465247 25725 465297 26325
rect 465397 25725 465447 26325
rect 467632 25936 467682 26936
rect 467782 25936 467838 26936
rect 467938 25936 467994 26936
rect 468094 25936 468150 26936
rect 468250 26810 468300 26936
rect 468714 26810 468764 26936
rect 468250 26726 468303 26810
rect 468711 26726 468764 26810
rect 468250 26477 468300 26726
rect 468714 26477 468764 26726
rect 468250 26393 468303 26477
rect 468711 26393 468764 26477
rect 468250 25936 468300 26393
rect 468714 25936 468764 26393
rect 468864 25936 468920 26936
rect 469020 25936 469076 26936
rect 469176 25936 469232 26936
rect 469332 25936 469382 26936
rect 476307 26490 476360 26690
rect 476460 26490 476516 26690
rect 476616 26490 476666 26690
rect 477016 26490 477066 26690
rect 477166 26490 477222 26690
rect 477322 26490 477372 26690
rect 566185 26478 566491 26648
rect 477661 26348 477695 26372
rect 477730 26348 477764 26372
rect 516427 25725 516477 26325
rect 516577 25725 516627 26325
rect 516699 25725 516749 26325
rect 516849 25725 516899 26325
rect 516975 25725 517025 26325
rect 517125 25725 517175 26325
rect 517247 25725 517297 26325
rect 517397 25725 517447 26325
rect 564427 25725 564477 26325
rect 564577 25725 564627 26325
rect 564699 25725 564749 26325
rect 564849 25725 564899 26325
rect 564975 25725 565025 26325
rect 565125 25725 565175 26325
rect 565247 25725 565297 26325
rect 565397 25725 565447 26325
rect 567632 25936 567682 26936
rect 567782 25936 567838 26936
rect 567938 25936 567994 26936
rect 568094 25936 568150 26936
rect 568250 26810 568300 26936
rect 568714 26810 568764 26936
rect 568250 26726 568303 26810
rect 568711 26726 568764 26810
rect 568250 26477 568300 26726
rect 568714 26477 568764 26726
rect 568250 26393 568303 26477
rect 568711 26393 568764 26477
rect 568250 25936 568300 26393
rect 568714 25936 568764 26393
rect 568864 25936 568920 26936
rect 569020 25936 569076 26936
rect 569176 25936 569232 26936
rect 569332 25936 569382 26936
rect 576307 26490 576360 26690
rect 576460 26490 576516 26690
rect 576616 26490 576666 26690
rect 577016 26490 577066 26690
rect 577166 26490 577222 26690
rect 577322 26490 577372 26690
rect 577661 26348 577695 26372
rect 577730 26348 577764 26372
rect 365773 25414 365807 25438
rect 367223 25312 367237 25336
rect 367189 25288 367213 25312
rect 367247 25288 367271 25312
rect 55983 25238 56017 25258
rect 107983 25238 108017 25258
rect 159983 25238 160017 25258
rect 211983 25238 212017 25258
rect 259983 25238 260017 25258
rect 311983 25238 312017 25258
rect 363983 25238 364017 25258
rect 55983 25102 56017 25137
rect 56085 25122 56109 25146
rect 56326 25143 56360 25147
rect 56394 25143 56428 25147
rect 56462 25143 56496 25147
rect 56530 25143 56564 25147
rect 56598 25143 56632 25147
rect 56666 25143 56700 25147
rect 56734 25143 56768 25147
rect 56802 25143 56836 25147
rect 56870 25143 56904 25147
rect 56938 25143 56972 25147
rect 57006 25143 57040 25147
rect 57074 25143 57108 25147
rect 57142 25143 57176 25147
rect 57210 25143 57244 25147
rect 56248 25125 57260 25143
rect 56326 25121 56360 25125
rect 56394 25121 56428 25125
rect 56462 25121 56496 25125
rect 56530 25121 56564 25125
rect 56598 25121 56632 25125
rect 56666 25121 56700 25125
rect 56734 25121 56768 25125
rect 56802 25121 56836 25125
rect 56870 25121 56904 25125
rect 56938 25121 56972 25125
rect 57006 25121 57040 25125
rect 57074 25121 57108 25125
rect 57142 25121 57176 25125
rect 57210 25121 57244 25125
rect 56252 25113 57260 25121
rect 55983 25089 56007 25102
rect 56061 25098 56085 25113
rect 56302 25101 57260 25113
rect 56429 23617 56472 25017
rect 56579 23617 56707 25017
rect 56742 23617 56870 25017
rect 56905 23617 57033 25017
rect 57068 23617 57196 25017
rect 57231 23617 57260 25017
rect 57720 23617 57763 25017
rect 57856 23617 57899 25017
rect 69552 24573 69608 25173
rect 70020 24573 70070 25173
rect 70508 24572 70558 25172
rect 70658 24572 70708 25172
rect 70788 24572 70838 25172
rect 70938 24572 71066 25172
rect 71094 24572 71222 25172
rect 71250 24572 71306 25172
rect 71406 24572 71534 25172
rect 71562 24572 71690 25172
rect 71718 24572 71768 25172
rect 107983 25102 108017 25137
rect 108085 25122 108109 25146
rect 108326 25143 108360 25147
rect 108394 25143 108428 25147
rect 108462 25143 108496 25147
rect 108530 25143 108564 25147
rect 108598 25143 108632 25147
rect 108666 25143 108700 25147
rect 108734 25143 108768 25147
rect 108802 25143 108836 25147
rect 108870 25143 108904 25147
rect 108938 25143 108972 25147
rect 109006 25143 109040 25147
rect 109074 25143 109108 25147
rect 109142 25143 109176 25147
rect 109210 25143 109244 25147
rect 108248 25125 109260 25143
rect 108326 25121 108360 25125
rect 108394 25121 108428 25125
rect 108462 25121 108496 25125
rect 108530 25121 108564 25125
rect 108598 25121 108632 25125
rect 108666 25121 108700 25125
rect 108734 25121 108768 25125
rect 108802 25121 108836 25125
rect 108870 25121 108904 25125
rect 108938 25121 108972 25125
rect 109006 25121 109040 25125
rect 109074 25121 109108 25125
rect 109142 25121 109176 25125
rect 109210 25121 109244 25125
rect 108252 25113 109260 25121
rect 107983 25089 108007 25102
rect 108061 25098 108085 25113
rect 108302 25101 109260 25113
rect 108429 23617 108472 25017
rect 108579 23617 108707 25017
rect 108742 23617 108870 25017
rect 108905 23617 109033 25017
rect 109068 23617 109196 25017
rect 109231 23617 109260 25017
rect 109720 23617 109763 25017
rect 109856 23617 109899 25017
rect 121552 24573 121608 25173
rect 122020 24573 122070 25173
rect 122508 24572 122558 25172
rect 122658 24572 122708 25172
rect 122788 24572 122838 25172
rect 122938 24572 123066 25172
rect 123094 24572 123222 25172
rect 123250 24572 123306 25172
rect 123406 24572 123534 25172
rect 123562 24572 123690 25172
rect 123718 24572 123768 25172
rect 159983 25102 160017 25137
rect 160085 25122 160109 25146
rect 160326 25143 160360 25147
rect 160394 25143 160428 25147
rect 160462 25143 160496 25147
rect 160530 25143 160564 25147
rect 160598 25143 160632 25147
rect 160666 25143 160700 25147
rect 160734 25143 160768 25147
rect 160802 25143 160836 25147
rect 160870 25143 160904 25147
rect 160938 25143 160972 25147
rect 161006 25143 161040 25147
rect 161074 25143 161108 25147
rect 161142 25143 161176 25147
rect 161210 25143 161244 25147
rect 160248 25125 161260 25143
rect 160326 25121 160360 25125
rect 160394 25121 160428 25125
rect 160462 25121 160496 25125
rect 160530 25121 160564 25125
rect 160598 25121 160632 25125
rect 160666 25121 160700 25125
rect 160734 25121 160768 25125
rect 160802 25121 160836 25125
rect 160870 25121 160904 25125
rect 160938 25121 160972 25125
rect 161006 25121 161040 25125
rect 161074 25121 161108 25125
rect 161142 25121 161176 25125
rect 161210 25121 161244 25125
rect 160252 25113 161260 25121
rect 159983 25089 160007 25102
rect 160061 25098 160085 25113
rect 160302 25101 161260 25113
rect 160429 23617 160472 25017
rect 160579 23617 160707 25017
rect 160742 23617 160870 25017
rect 160905 23617 161033 25017
rect 161068 23617 161196 25017
rect 161231 23617 161260 25017
rect 173552 24573 173608 25173
rect 174020 24573 174070 25173
rect 174508 24572 174558 25172
rect 174658 24572 174708 25172
rect 174788 24572 174838 25172
rect 174938 24572 175066 25172
rect 175094 24572 175222 25172
rect 175250 24572 175306 25172
rect 175406 24572 175534 25172
rect 175562 24572 175690 25172
rect 175718 24572 175768 25172
rect 211983 25102 212017 25137
rect 212085 25122 212109 25146
rect 212326 25143 212360 25147
rect 212394 25143 212428 25147
rect 212462 25143 212496 25147
rect 212530 25143 212564 25147
rect 212598 25143 212632 25147
rect 212666 25143 212700 25147
rect 212734 25143 212768 25147
rect 212802 25143 212836 25147
rect 212870 25143 212904 25147
rect 212938 25143 212972 25147
rect 213006 25143 213040 25147
rect 213074 25143 213108 25147
rect 213142 25143 213176 25147
rect 213210 25143 213244 25147
rect 212248 25125 213260 25143
rect 212326 25121 212360 25125
rect 212394 25121 212428 25125
rect 212462 25121 212496 25125
rect 212530 25121 212564 25125
rect 212598 25121 212632 25125
rect 212666 25121 212700 25125
rect 212734 25121 212768 25125
rect 212802 25121 212836 25125
rect 212870 25121 212904 25125
rect 212938 25121 212972 25125
rect 213006 25121 213040 25125
rect 213074 25121 213108 25125
rect 213142 25121 213176 25125
rect 213210 25121 213244 25125
rect 212252 25113 213260 25121
rect 211983 25089 212007 25102
rect 212061 25098 212085 25113
rect 212302 25101 213260 25113
rect 212429 23617 212472 25017
rect 212579 23617 212707 25017
rect 212742 23617 212870 25017
rect 212905 23617 213033 25017
rect 213068 23617 213196 25017
rect 213231 23617 213260 25017
rect 213720 23617 213763 25017
rect 213856 23617 213899 25017
rect 225552 24573 225608 25173
rect 226020 24573 226070 25173
rect 226508 24572 226558 25172
rect 226658 24572 226708 25172
rect 226788 24572 226838 25172
rect 226938 24572 227066 25172
rect 227094 24572 227222 25172
rect 227250 24572 227306 25172
rect 227406 24572 227534 25172
rect 227562 24572 227690 25172
rect 227718 24572 227768 25172
rect 259983 25102 260017 25137
rect 260085 25122 260109 25146
rect 260326 25143 260360 25147
rect 260394 25143 260428 25147
rect 260462 25143 260496 25147
rect 260530 25143 260564 25147
rect 260598 25143 260632 25147
rect 260666 25143 260700 25147
rect 260734 25143 260768 25147
rect 260802 25143 260836 25147
rect 260870 25143 260904 25147
rect 260938 25143 260972 25147
rect 261006 25143 261040 25147
rect 261074 25143 261108 25147
rect 261142 25143 261176 25147
rect 261210 25143 261244 25147
rect 260248 25125 261260 25143
rect 260326 25121 260360 25125
rect 260394 25121 260428 25125
rect 260462 25121 260496 25125
rect 260530 25121 260564 25125
rect 260598 25121 260632 25125
rect 260666 25121 260700 25125
rect 260734 25121 260768 25125
rect 260802 25121 260836 25125
rect 260870 25121 260904 25125
rect 260938 25121 260972 25125
rect 261006 25121 261040 25125
rect 261074 25121 261108 25125
rect 261142 25121 261176 25125
rect 261210 25121 261244 25125
rect 260252 25113 261260 25121
rect 259983 25089 260007 25102
rect 260061 25098 260085 25113
rect 260302 25101 261260 25113
rect 260429 23617 260472 25017
rect 260579 23617 260707 25017
rect 260742 23617 260870 25017
rect 260905 23617 261033 25017
rect 261068 23617 261196 25017
rect 261231 23617 261260 25017
rect 261720 23617 261763 25017
rect 261856 23617 261899 25017
rect 273552 24573 273608 25173
rect 274020 24573 274070 25173
rect 274508 24572 274558 25172
rect 274658 24572 274708 25172
rect 274788 24572 274838 25172
rect 274938 24572 275066 25172
rect 275094 24572 275222 25172
rect 275250 24572 275306 25172
rect 275406 24572 275534 25172
rect 275562 24572 275690 25172
rect 275718 24572 275768 25172
rect 311983 25102 312017 25137
rect 312085 25122 312109 25146
rect 312326 25143 312360 25147
rect 312394 25143 312428 25147
rect 312462 25143 312496 25147
rect 312530 25143 312564 25147
rect 312598 25143 312632 25147
rect 312666 25143 312700 25147
rect 312734 25143 312768 25147
rect 312802 25143 312836 25147
rect 312870 25143 312904 25147
rect 312938 25143 312972 25147
rect 313006 25143 313040 25147
rect 313074 25143 313108 25147
rect 313142 25143 313176 25147
rect 313210 25143 313244 25147
rect 312248 25125 313260 25143
rect 312326 25121 312360 25125
rect 312394 25121 312428 25125
rect 312462 25121 312496 25125
rect 312530 25121 312564 25125
rect 312598 25121 312632 25125
rect 312666 25121 312700 25125
rect 312734 25121 312768 25125
rect 312802 25121 312836 25125
rect 312870 25121 312904 25125
rect 312938 25121 312972 25125
rect 313006 25121 313040 25125
rect 313074 25121 313108 25125
rect 313142 25121 313176 25125
rect 313210 25121 313244 25125
rect 312252 25113 313260 25121
rect 311983 25089 312007 25102
rect 312061 25098 312085 25113
rect 312302 25101 313260 25113
rect 312429 23617 312472 25017
rect 312579 23617 312707 25017
rect 312742 23617 312870 25017
rect 312905 23617 313033 25017
rect 313068 23617 313196 25017
rect 313231 23617 313260 25017
rect 313720 23617 313763 25017
rect 313856 23617 313899 25017
rect 325552 24573 325608 25173
rect 326020 24573 326070 25173
rect 326508 24572 326558 25172
rect 326658 24572 326708 25172
rect 326788 24572 326838 25172
rect 326938 24572 327066 25172
rect 327094 24572 327222 25172
rect 327250 24572 327306 25172
rect 327406 24572 327534 25172
rect 327562 24572 327690 25172
rect 327718 24572 327768 25172
rect 363983 25102 364017 25137
rect 364085 25122 364109 25146
rect 364326 25143 364360 25147
rect 364394 25143 364428 25147
rect 364462 25143 364496 25147
rect 364530 25143 364564 25147
rect 364598 25143 364632 25147
rect 364666 25143 364700 25147
rect 364734 25143 364768 25147
rect 364802 25143 364836 25147
rect 364870 25143 364904 25147
rect 364938 25143 364972 25147
rect 365006 25143 365040 25147
rect 365074 25143 365108 25147
rect 365142 25143 365176 25147
rect 365210 25143 365244 25147
rect 365278 25143 365312 25147
rect 365346 25143 365380 25147
rect 365414 25143 365448 25147
rect 365482 25143 365516 25147
rect 365550 25143 365584 25147
rect 365618 25143 365652 25147
rect 365686 25143 365720 25147
rect 365754 25143 365788 25147
rect 365822 25143 365856 25147
rect 365890 25143 365924 25147
rect 365958 25143 365992 25147
rect 366026 25143 366060 25147
rect 366094 25143 366128 25147
rect 366162 25143 366196 25147
rect 366230 25143 366264 25147
rect 366298 25143 366332 25147
rect 366366 25143 366400 25147
rect 366434 25143 366468 25147
rect 366502 25143 366536 25147
rect 366570 25143 366604 25147
rect 366638 25143 366672 25147
rect 366706 25143 366740 25147
rect 366774 25143 366808 25147
rect 366842 25143 366876 25147
rect 366910 25143 366944 25147
rect 366978 25143 367012 25147
rect 367046 25143 367080 25147
rect 364248 25125 367148 25143
rect 367532 25125 367556 25149
rect 367590 25125 367614 25149
rect 364326 25121 364360 25125
rect 364394 25121 364428 25125
rect 364462 25121 364496 25125
rect 364530 25121 364564 25125
rect 364598 25121 364632 25125
rect 364666 25121 364700 25125
rect 364734 25121 364768 25125
rect 364802 25121 364836 25125
rect 364870 25121 364904 25125
rect 364938 25121 364972 25125
rect 365006 25121 365040 25125
rect 365074 25121 365108 25125
rect 365142 25121 365176 25125
rect 365210 25121 365244 25125
rect 365278 25121 365312 25125
rect 365346 25121 365380 25125
rect 365414 25121 365448 25125
rect 365482 25121 365516 25125
rect 365550 25121 365584 25125
rect 365618 25121 365652 25125
rect 365686 25121 365720 25125
rect 365754 25121 365788 25125
rect 365822 25121 365856 25125
rect 365890 25121 365924 25125
rect 365958 25121 365992 25125
rect 366026 25121 366060 25125
rect 366094 25121 366128 25125
rect 366162 25121 366196 25125
rect 366230 25121 366264 25125
rect 366298 25121 366332 25125
rect 366366 25121 366400 25125
rect 366434 25121 366468 25125
rect 366502 25121 366536 25125
rect 366570 25121 366604 25125
rect 366638 25121 366672 25125
rect 366706 25121 366740 25125
rect 366774 25121 366808 25125
rect 366842 25121 366876 25125
rect 366910 25121 366944 25125
rect 366978 25121 367012 25125
rect 367046 25121 367080 25125
rect 364252 25113 367144 25121
rect 363983 25089 364007 25102
rect 364061 25098 364085 25113
rect 364302 25101 367104 25113
rect 367556 25101 367590 25115
rect 367532 25067 367556 25091
rect 367590 25067 367614 25091
rect 369996 25085 370532 25553
rect 370835 25524 370869 25548
rect 370903 25524 374201 25548
rect 374269 25383 374293 25417
rect 465773 25414 465807 25438
rect 370708 25113 370810 25137
rect 370939 25126 370963 25150
rect 370708 25089 370732 25113
rect 370786 25089 370810 25113
rect 370963 25102 370987 25116
rect 371041 25113 371065 25116
rect 372091 25113 372193 25137
rect 364429 23617 364472 25017
rect 364579 23617 364707 25017
rect 364742 23617 364870 25017
rect 364905 23617 365033 25017
rect 365068 23617 365196 25017
rect 365231 23617 365359 25017
rect 365394 23617 365522 25017
rect 365557 23617 365685 25017
rect 365720 23617 365763 25017
rect 365856 23617 365899 25017
rect 366006 23617 366134 25017
rect 366169 23617 366297 25017
rect 366332 23617 366460 25017
rect 366495 23617 366623 25017
rect 366658 23617 366786 25017
rect 366821 23617 366949 25017
rect 366984 23617 367034 25017
rect 367301 23300 367403 24864
rect 367670 23685 367720 25085
rect 367827 23685 367955 25085
rect 367990 23685 368118 25085
rect 368153 23685 368281 25085
rect 368316 23685 368444 25085
rect 368479 23685 368607 25085
rect 368642 23685 368770 25085
rect 368805 23685 368848 25085
rect 368941 23685 368984 25085
rect 369091 23685 369219 25085
rect 369254 23685 369382 25085
rect 369417 23685 369545 25085
rect 369580 23685 369708 25085
rect 369743 23685 369871 25085
rect 369906 23685 370532 25085
rect 370939 25068 370963 25092
rect 371065 25068 371089 25092
rect 372091 25089 372115 25113
rect 372169 25089 372193 25113
rect 372347 25113 372381 25147
rect 372419 25113 372453 25147
rect 372491 25113 372525 25147
rect 372563 25113 372597 25147
rect 372347 25089 372371 25113
rect 372573 25089 372597 25113
rect 372752 25089 372786 25147
rect 374269 25137 374293 25349
rect 467223 25312 467237 25336
rect 375671 25286 375705 25310
rect 375743 25286 375777 25310
rect 375815 25286 375849 25310
rect 375887 25286 375921 25310
rect 375958 25286 375962 25310
rect 467189 25288 467213 25312
rect 467247 25288 467271 25312
rect 411983 25238 412017 25258
rect 463983 25238 464017 25258
rect 374167 25113 374293 25137
rect 374167 25089 374191 25113
rect 371152 23685 371195 25085
rect 371302 23685 371430 25085
rect 371465 23685 371593 25085
rect 371628 23685 371756 25085
rect 371791 23685 371919 25085
rect 371954 23685 372004 25085
rect 372873 23685 372916 25085
rect 373023 23685 373151 25085
rect 373186 23685 373314 25085
rect 373349 23685 373477 25085
rect 373512 23685 373640 25085
rect 373675 23685 373803 25085
rect 373838 23685 373881 25085
rect 375428 24573 375478 25173
rect 375578 24573 375706 25173
rect 375734 24573 375862 25173
rect 375890 24573 375946 25173
rect 376046 24573 376174 25173
rect 376202 24573 376330 25173
rect 376358 24573 376408 25173
rect 376488 24573 376538 25173
rect 376638 24573 376688 25173
rect 376810 24573 376860 25173
rect 376960 24573 377010 25173
rect 377090 24573 377140 25173
rect 377240 24573 377368 25173
rect 377396 24573 377524 25173
rect 377552 24573 377608 25173
rect 377708 24573 377836 25173
rect 377864 24573 377992 25173
rect 378020 24573 378070 25173
rect 378508 24572 378558 25172
rect 378658 24572 378708 25172
rect 378788 24572 378838 25172
rect 378938 24572 379066 25172
rect 379094 24572 379222 25172
rect 379250 24572 379306 25172
rect 379406 24572 379534 25172
rect 379562 24572 379690 25172
rect 379718 24572 379768 25172
rect 411983 25102 412017 25137
rect 412085 25122 412109 25146
rect 412326 25143 412360 25147
rect 412394 25143 412428 25147
rect 412462 25143 412496 25147
rect 412530 25143 412564 25147
rect 412598 25143 412632 25147
rect 412666 25143 412700 25147
rect 412734 25143 412768 25147
rect 412802 25143 412836 25147
rect 412870 25143 412904 25147
rect 412938 25143 412972 25147
rect 413006 25143 413040 25147
rect 413074 25143 413108 25147
rect 413142 25143 413176 25147
rect 413210 25143 413244 25147
rect 412248 25125 413260 25143
rect 412326 25121 412360 25125
rect 412394 25121 412428 25125
rect 412462 25121 412496 25125
rect 412530 25121 412564 25125
rect 412598 25121 412632 25125
rect 412666 25121 412700 25125
rect 412734 25121 412768 25125
rect 412802 25121 412836 25125
rect 412870 25121 412904 25125
rect 412938 25121 412972 25125
rect 413006 25121 413040 25125
rect 413074 25121 413108 25125
rect 413142 25121 413176 25125
rect 413210 25121 413244 25125
rect 412252 25113 413260 25121
rect 411983 25089 412007 25102
rect 412061 25098 412085 25113
rect 412302 25101 413260 25113
rect 367335 23276 367369 23300
rect 367335 23198 367369 23222
rect 56429 21481 56472 22881
rect 56579 21481 56707 22881
rect 56742 21481 56870 22881
rect 56905 21481 57033 22881
rect 57068 21481 57196 22881
rect 57231 21481 57260 22881
rect 57720 21481 57763 22881
rect 57856 21481 57899 22881
rect 69480 22349 69718 22399
rect 108429 21481 108472 22881
rect 108579 21481 108707 22881
rect 108742 21481 108870 22881
rect 108905 21481 109033 22881
rect 109068 21481 109196 22881
rect 109231 21481 109260 22881
rect 109720 21481 109763 22881
rect 109856 21481 109899 22881
rect 121480 22349 121718 22399
rect 160429 21481 160472 22881
rect 160579 21481 160707 22881
rect 160742 21481 160870 22881
rect 160905 21481 161033 22881
rect 161068 21481 161196 22881
rect 161231 21481 161260 22881
rect 173480 22349 173718 22399
rect 212429 21481 212472 22881
rect 212579 21481 212707 22881
rect 212742 21481 212870 22881
rect 212905 21481 213033 22881
rect 213068 21481 213196 22881
rect 213231 21481 213260 22881
rect 213720 21481 213763 22881
rect 213856 21481 213899 22881
rect 225480 22349 225718 22399
rect 260429 21481 260472 22881
rect 260579 21481 260707 22881
rect 260742 21481 260870 22881
rect 260905 21481 261033 22881
rect 261068 21481 261196 22881
rect 261231 21481 261260 22881
rect 261720 21481 261763 22881
rect 261856 21481 261899 22881
rect 273480 22349 273718 22399
rect 312429 21481 312472 22881
rect 312579 21481 312707 22881
rect 312742 21481 312870 22881
rect 312905 21481 313033 22881
rect 313068 21481 313196 22881
rect 313231 21481 313260 22881
rect 313720 21481 313763 22881
rect 313856 21481 313899 22881
rect 325480 22349 325718 22399
rect 364429 21481 364472 22881
rect 364579 21481 364707 22881
rect 364742 21481 364870 22881
rect 364905 21481 365033 22881
rect 365068 21481 365196 22881
rect 365231 21481 365359 22881
rect 365394 21481 365522 22881
rect 365557 21481 365685 22881
rect 365720 21481 365763 22881
rect 365856 21481 365899 22881
rect 366006 21481 366134 22881
rect 366169 21481 366297 22881
rect 366332 21481 366460 22881
rect 366495 21481 366623 22881
rect 366658 21481 366786 22881
rect 366821 21481 366949 22881
rect 366984 21481 367034 22881
rect 367301 21634 367403 23198
rect 369996 22813 370532 23685
rect 375455 23406 375625 23712
rect 376255 23406 376425 23712
rect 377055 23406 377225 23712
rect 412429 23617 412472 25017
rect 412579 23617 412707 25017
rect 412742 23617 412870 25017
rect 412905 23617 413033 25017
rect 413068 23617 413196 25017
rect 413231 23617 413260 25017
rect 413720 23617 413763 25017
rect 413856 23617 413899 25017
rect 425552 24573 425608 25173
rect 426020 24573 426070 25173
rect 426508 24572 426558 25172
rect 426658 24572 426708 25172
rect 426788 24572 426838 25172
rect 426938 24572 427066 25172
rect 427094 24572 427222 25172
rect 427250 24572 427306 25172
rect 427406 24572 427534 25172
rect 427562 24572 427690 25172
rect 427718 24572 427768 25172
rect 463983 25102 464017 25137
rect 464085 25122 464109 25146
rect 464326 25143 464360 25147
rect 464394 25143 464428 25147
rect 464462 25143 464496 25147
rect 464530 25143 464564 25147
rect 464598 25143 464632 25147
rect 464666 25143 464700 25147
rect 464734 25143 464768 25147
rect 464802 25143 464836 25147
rect 464870 25143 464904 25147
rect 464938 25143 464972 25147
rect 465006 25143 465040 25147
rect 465074 25143 465108 25147
rect 465142 25143 465176 25147
rect 465210 25143 465244 25147
rect 465278 25143 465312 25147
rect 465346 25143 465380 25147
rect 465414 25143 465448 25147
rect 465482 25143 465516 25147
rect 465550 25143 465584 25147
rect 465618 25143 465652 25147
rect 465686 25143 465720 25147
rect 465754 25143 465788 25147
rect 465822 25143 465856 25147
rect 465890 25143 465924 25147
rect 465958 25143 465992 25147
rect 466026 25143 466060 25147
rect 466094 25143 466128 25147
rect 466162 25143 466196 25147
rect 466230 25143 466264 25147
rect 466298 25143 466332 25147
rect 466366 25143 466400 25147
rect 466434 25143 466468 25147
rect 466502 25143 466536 25147
rect 466570 25143 466604 25147
rect 466638 25143 466672 25147
rect 466706 25143 466740 25147
rect 466774 25143 466808 25147
rect 466842 25143 466876 25147
rect 466910 25143 466944 25147
rect 466978 25143 467012 25147
rect 467046 25143 467080 25147
rect 464248 25125 467148 25143
rect 467532 25125 467556 25149
rect 467590 25125 467614 25149
rect 464326 25121 464360 25125
rect 464394 25121 464428 25125
rect 464462 25121 464496 25125
rect 464530 25121 464564 25125
rect 464598 25121 464632 25125
rect 464666 25121 464700 25125
rect 464734 25121 464768 25125
rect 464802 25121 464836 25125
rect 464870 25121 464904 25125
rect 464938 25121 464972 25125
rect 465006 25121 465040 25125
rect 465074 25121 465108 25125
rect 465142 25121 465176 25125
rect 465210 25121 465244 25125
rect 465278 25121 465312 25125
rect 465346 25121 465380 25125
rect 465414 25121 465448 25125
rect 465482 25121 465516 25125
rect 465550 25121 465584 25125
rect 465618 25121 465652 25125
rect 465686 25121 465720 25125
rect 465754 25121 465788 25125
rect 465822 25121 465856 25125
rect 465890 25121 465924 25125
rect 465958 25121 465992 25125
rect 466026 25121 466060 25125
rect 466094 25121 466128 25125
rect 466162 25121 466196 25125
rect 466230 25121 466264 25125
rect 466298 25121 466332 25125
rect 466366 25121 466400 25125
rect 466434 25121 466468 25125
rect 466502 25121 466536 25125
rect 466570 25121 466604 25125
rect 466638 25121 466672 25125
rect 466706 25121 466740 25125
rect 466774 25121 466808 25125
rect 466842 25121 466876 25125
rect 466910 25121 466944 25125
rect 466978 25121 467012 25125
rect 467046 25121 467080 25125
rect 464252 25113 467144 25121
rect 463983 25089 464007 25102
rect 464061 25098 464085 25113
rect 464302 25101 467104 25113
rect 467556 25101 467590 25115
rect 467532 25067 467556 25091
rect 467590 25067 467614 25091
rect 469996 25085 470532 25553
rect 470835 25524 470869 25548
rect 470903 25524 474201 25548
rect 474269 25383 474293 25417
rect 565773 25414 565807 25438
rect 470708 25113 470810 25137
rect 470939 25126 470963 25150
rect 470708 25089 470732 25113
rect 470786 25089 470810 25113
rect 470963 25102 470987 25116
rect 471041 25113 471065 25116
rect 472091 25113 472193 25137
rect 464429 23617 464472 25017
rect 464579 23617 464707 25017
rect 464742 23617 464870 25017
rect 464905 23617 465033 25017
rect 465068 23617 465196 25017
rect 465231 23617 465359 25017
rect 465394 23617 465522 25017
rect 465557 23617 465685 25017
rect 465720 23617 465763 25017
rect 465856 23617 465899 25017
rect 466006 23617 466134 25017
rect 466169 23617 466297 25017
rect 466332 23617 466460 25017
rect 466495 23617 466623 25017
rect 466658 23617 466786 25017
rect 466821 23617 466949 25017
rect 466984 23617 467034 25017
rect 467301 23300 467403 24864
rect 467670 23685 467720 25085
rect 467827 23685 467955 25085
rect 467990 23685 468118 25085
rect 468153 23685 468281 25085
rect 468316 23685 468444 25085
rect 468479 23685 468607 25085
rect 468642 23685 468770 25085
rect 468805 23685 468848 25085
rect 468941 23685 468984 25085
rect 469091 23685 469219 25085
rect 469254 23685 469382 25085
rect 469417 23685 469545 25085
rect 469580 23685 469708 25085
rect 469743 23685 469871 25085
rect 469906 23685 470532 25085
rect 470939 25068 470963 25092
rect 471065 25068 471089 25092
rect 472091 25089 472115 25113
rect 472169 25089 472193 25113
rect 472347 25113 472381 25147
rect 472419 25113 472453 25147
rect 472491 25113 472525 25147
rect 472563 25113 472597 25147
rect 472347 25089 472371 25113
rect 472573 25089 472597 25113
rect 472752 25089 472786 25147
rect 474269 25137 474293 25349
rect 567223 25312 567237 25336
rect 475671 25286 475705 25310
rect 475743 25286 475777 25310
rect 475815 25286 475849 25310
rect 475887 25286 475921 25310
rect 475958 25286 475962 25310
rect 567189 25288 567213 25312
rect 567247 25288 567271 25312
rect 515983 25238 516017 25258
rect 563983 25238 564017 25258
rect 474167 25113 474293 25137
rect 474167 25089 474191 25113
rect 471152 23685 471195 25085
rect 471302 23685 471430 25085
rect 471465 23685 471593 25085
rect 471628 23685 471756 25085
rect 471791 23685 471919 25085
rect 471954 23685 472004 25085
rect 472873 23685 472916 25085
rect 473023 23685 473151 25085
rect 473186 23685 473314 25085
rect 473349 23685 473477 25085
rect 473512 23685 473640 25085
rect 473675 23685 473803 25085
rect 473838 23685 473881 25085
rect 475428 24573 475478 25173
rect 475578 24573 475706 25173
rect 475734 24573 475862 25173
rect 475890 24573 475946 25173
rect 476046 24573 476174 25173
rect 476202 24573 476330 25173
rect 476358 24573 476408 25173
rect 476488 24573 476538 25173
rect 476638 24573 476688 25173
rect 476810 24573 476860 25173
rect 476960 24573 477010 25173
rect 477090 24573 477140 25173
rect 477240 24573 477368 25173
rect 477396 24573 477524 25173
rect 477552 24573 477608 25173
rect 477708 24573 477836 25173
rect 477864 24573 477992 25173
rect 478020 24573 478070 25173
rect 478508 24572 478558 25172
rect 478658 24572 478708 25172
rect 478788 24572 478838 25172
rect 478938 24572 479066 25172
rect 479094 24572 479222 25172
rect 479250 24572 479306 25172
rect 479406 24572 479534 25172
rect 479562 24572 479690 25172
rect 479718 24572 479768 25172
rect 515983 25102 516017 25137
rect 516085 25122 516109 25146
rect 516326 25143 516360 25147
rect 516394 25143 516428 25147
rect 516462 25143 516496 25147
rect 516530 25143 516564 25147
rect 516598 25143 516632 25147
rect 516666 25143 516700 25147
rect 516734 25143 516768 25147
rect 516802 25143 516836 25147
rect 516870 25143 516904 25147
rect 516938 25143 516972 25147
rect 517006 25143 517040 25147
rect 517074 25143 517108 25147
rect 517142 25143 517176 25147
rect 517210 25143 517244 25147
rect 516248 25125 517260 25143
rect 516326 25121 516360 25125
rect 516394 25121 516428 25125
rect 516462 25121 516496 25125
rect 516530 25121 516564 25125
rect 516598 25121 516632 25125
rect 516666 25121 516700 25125
rect 516734 25121 516768 25125
rect 516802 25121 516836 25125
rect 516870 25121 516904 25125
rect 516938 25121 516972 25125
rect 517006 25121 517040 25125
rect 517074 25121 517108 25125
rect 517142 25121 517176 25125
rect 517210 25121 517244 25125
rect 516252 25113 517260 25121
rect 515983 25089 516007 25102
rect 516061 25098 516085 25113
rect 516302 25101 517260 25113
rect 467335 23276 467369 23300
rect 375455 22906 375625 23212
rect 376255 22906 376425 23212
rect 377055 22906 377225 23212
rect 467335 23198 467369 23222
rect 55983 21410 56051 21430
rect 56326 21415 56360 21419
rect 56394 21415 56428 21419
rect 56462 21415 56496 21419
rect 56530 21415 56564 21419
rect 56598 21415 56632 21419
rect 56666 21415 56700 21419
rect 56734 21415 56768 21419
rect 56802 21415 56836 21419
rect 56870 21415 56904 21419
rect 56938 21415 56972 21419
rect 57006 21415 57040 21419
rect 57074 21415 57108 21419
rect 57142 21415 57176 21419
rect 57210 21415 57244 21419
rect 55983 21385 56017 21410
rect 56282 21407 57260 21415
rect 107983 21410 108051 21430
rect 108326 21415 108360 21419
rect 108394 21415 108428 21419
rect 108462 21415 108496 21419
rect 108530 21415 108564 21419
rect 108598 21415 108632 21419
rect 108666 21415 108700 21419
rect 108734 21415 108768 21419
rect 108802 21415 108836 21419
rect 108870 21415 108904 21419
rect 108938 21415 108972 21419
rect 109006 21415 109040 21419
rect 109074 21415 109108 21419
rect 109142 21415 109176 21419
rect 109210 21415 109244 21419
rect 56326 21403 56360 21407
rect 56394 21403 56428 21407
rect 56462 21403 56496 21407
rect 56530 21403 56564 21407
rect 56598 21403 56632 21407
rect 56666 21403 56700 21407
rect 56734 21403 56768 21407
rect 56802 21403 56836 21407
rect 56870 21403 56904 21407
rect 56938 21403 56972 21407
rect 57006 21403 57040 21407
rect 57074 21403 57108 21407
rect 57142 21403 57176 21407
rect 57210 21403 57244 21407
rect 56061 21385 56085 21400
rect 56248 21385 57260 21403
rect 55983 21361 56007 21385
rect 56302 21383 57260 21385
rect 107983 21385 108017 21410
rect 108282 21407 109260 21415
rect 159983 21410 160051 21430
rect 160326 21415 160360 21419
rect 160394 21415 160428 21419
rect 160462 21415 160496 21419
rect 160530 21415 160564 21419
rect 160598 21415 160632 21419
rect 160666 21415 160700 21419
rect 160734 21415 160768 21419
rect 160802 21415 160836 21419
rect 160870 21415 160904 21419
rect 160938 21415 160972 21419
rect 161006 21415 161040 21419
rect 161074 21415 161108 21419
rect 161142 21415 161176 21419
rect 161210 21415 161244 21419
rect 108326 21403 108360 21407
rect 108394 21403 108428 21407
rect 108462 21403 108496 21407
rect 108530 21403 108564 21407
rect 108598 21403 108632 21407
rect 108666 21403 108700 21407
rect 108734 21403 108768 21407
rect 108802 21403 108836 21407
rect 108870 21403 108904 21407
rect 108938 21403 108972 21407
rect 109006 21403 109040 21407
rect 109074 21403 109108 21407
rect 109142 21403 109176 21407
rect 109210 21403 109244 21407
rect 108061 21385 108085 21400
rect 108248 21385 109260 21403
rect 56085 21352 56109 21376
rect 107983 21361 108007 21385
rect 108302 21383 109260 21385
rect 159983 21385 160017 21410
rect 160282 21407 161260 21415
rect 211983 21410 212051 21430
rect 212326 21415 212360 21419
rect 212394 21415 212428 21419
rect 212462 21415 212496 21419
rect 212530 21415 212564 21419
rect 212598 21415 212632 21419
rect 212666 21415 212700 21419
rect 212734 21415 212768 21419
rect 212802 21415 212836 21419
rect 212870 21415 212904 21419
rect 212938 21415 212972 21419
rect 213006 21415 213040 21419
rect 213074 21415 213108 21419
rect 213142 21415 213176 21419
rect 213210 21415 213244 21419
rect 160326 21403 160360 21407
rect 160394 21403 160428 21407
rect 160462 21403 160496 21407
rect 160530 21403 160564 21407
rect 160598 21403 160632 21407
rect 160666 21403 160700 21407
rect 160734 21403 160768 21407
rect 160802 21403 160836 21407
rect 160870 21403 160904 21407
rect 160938 21403 160972 21407
rect 161006 21403 161040 21407
rect 161074 21403 161108 21407
rect 161142 21403 161176 21407
rect 161210 21403 161244 21407
rect 160061 21385 160085 21400
rect 160248 21385 161260 21403
rect 108085 21352 108109 21376
rect 159983 21361 160007 21385
rect 160302 21383 161260 21385
rect 211983 21385 212017 21410
rect 212282 21407 213260 21415
rect 259983 21410 260051 21430
rect 260326 21415 260360 21419
rect 260394 21415 260428 21419
rect 260462 21415 260496 21419
rect 260530 21415 260564 21419
rect 260598 21415 260632 21419
rect 260666 21415 260700 21419
rect 260734 21415 260768 21419
rect 260802 21415 260836 21419
rect 260870 21415 260904 21419
rect 260938 21415 260972 21419
rect 261006 21415 261040 21419
rect 261074 21415 261108 21419
rect 261142 21415 261176 21419
rect 261210 21415 261244 21419
rect 212326 21403 212360 21407
rect 212394 21403 212428 21407
rect 212462 21403 212496 21407
rect 212530 21403 212564 21407
rect 212598 21403 212632 21407
rect 212666 21403 212700 21407
rect 212734 21403 212768 21407
rect 212802 21403 212836 21407
rect 212870 21403 212904 21407
rect 212938 21403 212972 21407
rect 213006 21403 213040 21407
rect 213074 21403 213108 21407
rect 213142 21403 213176 21407
rect 213210 21403 213244 21407
rect 212061 21385 212085 21400
rect 212248 21385 213260 21403
rect 160085 21352 160109 21376
rect 211983 21361 212007 21385
rect 212302 21383 213260 21385
rect 259983 21385 260017 21410
rect 260282 21407 261260 21415
rect 311983 21410 312051 21430
rect 312326 21415 312360 21419
rect 312394 21415 312428 21419
rect 312462 21415 312496 21419
rect 312530 21415 312564 21419
rect 312598 21415 312632 21419
rect 312666 21415 312700 21419
rect 312734 21415 312768 21419
rect 312802 21415 312836 21419
rect 312870 21415 312904 21419
rect 312938 21415 312972 21419
rect 313006 21415 313040 21419
rect 313074 21415 313108 21419
rect 313142 21415 313176 21419
rect 313210 21415 313244 21419
rect 260326 21403 260360 21407
rect 260394 21403 260428 21407
rect 260462 21403 260496 21407
rect 260530 21403 260564 21407
rect 260598 21403 260632 21407
rect 260666 21403 260700 21407
rect 260734 21403 260768 21407
rect 260802 21403 260836 21407
rect 260870 21403 260904 21407
rect 260938 21403 260972 21407
rect 261006 21403 261040 21407
rect 261074 21403 261108 21407
rect 261142 21403 261176 21407
rect 261210 21403 261244 21407
rect 260061 21385 260085 21400
rect 260248 21385 261260 21403
rect 212085 21352 212109 21376
rect 259983 21361 260007 21385
rect 260302 21383 261260 21385
rect 311983 21385 312017 21410
rect 312282 21407 313260 21415
rect 363983 21410 364051 21430
rect 364326 21415 364360 21419
rect 364394 21415 364428 21419
rect 364462 21415 364496 21419
rect 364530 21415 364564 21419
rect 364598 21415 364632 21419
rect 364666 21415 364700 21419
rect 364734 21415 364768 21419
rect 364802 21415 364836 21419
rect 364870 21415 364904 21419
rect 364938 21415 364972 21419
rect 365006 21415 365040 21419
rect 365074 21415 365108 21419
rect 365142 21415 365176 21419
rect 365210 21415 365244 21419
rect 365278 21415 365312 21419
rect 365346 21415 365380 21419
rect 365414 21415 365448 21419
rect 365482 21415 365516 21419
rect 365550 21415 365584 21419
rect 365618 21415 365652 21419
rect 365686 21415 365720 21419
rect 365754 21415 365788 21419
rect 365822 21415 365856 21419
rect 365890 21415 365924 21419
rect 365958 21415 365992 21419
rect 366026 21415 366060 21419
rect 366094 21415 366128 21419
rect 366162 21415 366196 21419
rect 366230 21415 366264 21419
rect 366298 21415 366332 21419
rect 366366 21415 366400 21419
rect 366434 21415 366468 21419
rect 366502 21415 366536 21419
rect 366570 21415 366604 21419
rect 366638 21415 366672 21419
rect 366706 21415 366740 21419
rect 366774 21415 366808 21419
rect 366842 21415 366876 21419
rect 366910 21415 366944 21419
rect 366978 21415 367012 21419
rect 367046 21415 367080 21419
rect 312326 21403 312360 21407
rect 312394 21403 312428 21407
rect 312462 21403 312496 21407
rect 312530 21403 312564 21407
rect 312598 21403 312632 21407
rect 312666 21403 312700 21407
rect 312734 21403 312768 21407
rect 312802 21403 312836 21407
rect 312870 21403 312904 21407
rect 312938 21403 312972 21407
rect 313006 21403 313040 21407
rect 313074 21403 313108 21407
rect 313142 21403 313176 21407
rect 313210 21403 313244 21407
rect 312061 21385 312085 21400
rect 312248 21385 313260 21403
rect 260085 21352 260109 21376
rect 311983 21361 312007 21385
rect 312302 21383 313260 21385
rect 363983 21385 364017 21410
rect 364282 21407 367114 21415
rect 367532 21407 367556 21431
rect 367590 21407 367614 21431
rect 367670 21413 367720 22813
rect 367827 21413 367955 22813
rect 367990 21413 368118 22813
rect 368153 21413 368281 22813
rect 368316 21413 368444 22813
rect 368479 21413 368607 22813
rect 368642 21413 368770 22813
rect 368805 21413 368848 22813
rect 368941 21413 368984 22813
rect 369091 21413 369219 22813
rect 369254 21413 369382 22813
rect 369417 21413 369545 22813
rect 369580 21413 369708 22813
rect 369743 21413 369871 22813
rect 369906 21413 370532 22813
rect 364326 21403 364360 21407
rect 364394 21403 364428 21407
rect 364462 21403 364496 21407
rect 364530 21403 364564 21407
rect 364598 21403 364632 21407
rect 364666 21403 364700 21407
rect 364734 21403 364768 21407
rect 364802 21403 364836 21407
rect 364870 21403 364904 21407
rect 364938 21403 364972 21407
rect 365006 21403 365040 21407
rect 365074 21403 365108 21407
rect 365142 21403 365176 21407
rect 365210 21403 365244 21407
rect 365278 21403 365312 21407
rect 365346 21403 365380 21407
rect 365414 21403 365448 21407
rect 365482 21403 365516 21407
rect 365550 21403 365584 21407
rect 365618 21403 365652 21407
rect 365686 21403 365720 21407
rect 365754 21403 365788 21407
rect 365822 21403 365856 21407
rect 365890 21403 365924 21407
rect 365958 21403 365992 21407
rect 366026 21403 366060 21407
rect 366094 21403 366128 21407
rect 366162 21403 366196 21407
rect 366230 21403 366264 21407
rect 366298 21403 366332 21407
rect 366366 21403 366400 21407
rect 366434 21403 366468 21407
rect 366502 21403 366536 21407
rect 366570 21403 366604 21407
rect 366638 21403 366672 21407
rect 366706 21403 366740 21407
rect 366774 21403 366808 21407
rect 366842 21403 366876 21407
rect 366910 21403 366944 21407
rect 366978 21403 367012 21407
rect 367046 21403 367080 21407
rect 364061 21385 364085 21400
rect 364248 21385 367148 21403
rect 312085 21352 312109 21376
rect 363983 21361 364007 21385
rect 364302 21383 367104 21385
rect 367556 21383 367590 21397
rect 364085 21352 364109 21376
rect 367532 21349 367556 21373
rect 367590 21349 367614 21373
rect 55983 21274 56051 21294
rect 69480 21263 69718 21313
rect 107983 21274 108051 21294
rect 121480 21263 121718 21313
rect 159983 21274 160051 21294
rect 173480 21263 173718 21313
rect 211983 21274 212051 21294
rect 225480 21263 225718 21313
rect 259983 21274 260051 21294
rect 273480 21263 273718 21313
rect 311983 21274 312051 21294
rect 325480 21263 325718 21313
rect 363983 21274 364051 21294
rect 367189 21186 367213 21210
rect 367247 21186 367271 21210
rect 367223 21162 367237 21186
rect 40200 21000 40320 21003
rect 56000 21000 56120 21003
rect 72200 21000 72320 21003
rect 108000 21000 108120 21003
rect 124200 21000 124320 21003
rect 160000 21000 160120 21003
rect 176200 21000 176320 21003
rect 212000 21000 212120 21003
rect 228200 21000 228320 21003
rect 260000 21000 260120 21003
rect 276200 21000 276320 21003
rect 312000 21000 312120 21003
rect 328200 21000 328320 21003
rect 364000 21000 364120 21003
rect 369996 20945 370532 21413
rect 370708 21385 370810 21409
rect 370939 21406 370963 21430
rect 371065 21406 371089 21430
rect 371152 21413 371195 22813
rect 371302 21413 371430 22813
rect 371465 21413 371593 22813
rect 371628 21413 371756 22813
rect 371791 21413 371919 22813
rect 371954 21413 372004 22813
rect 370708 21361 370732 21385
rect 370786 21361 370810 21385
rect 370963 21382 370987 21396
rect 372091 21385 372193 21409
rect 371041 21382 371065 21385
rect 370939 21348 370963 21372
rect 372091 21361 372115 21385
rect 372169 21361 372193 21385
rect 372347 21385 372381 21419
rect 372419 21385 372453 21419
rect 372491 21385 372525 21419
rect 372563 21385 372597 21419
rect 372347 21361 372371 21385
rect 372573 21361 372597 21385
rect 372752 21361 372786 21419
rect 372873 21413 372916 22813
rect 373023 21413 373151 22813
rect 373186 21413 373314 22813
rect 373349 21413 373477 22813
rect 373512 21413 373640 22813
rect 373675 21413 373803 22813
rect 373838 21413 373881 22813
rect 374718 22349 377718 22399
rect 374718 22193 377718 22321
rect 378200 22197 378224 22210
rect 374718 22037 377718 22165
rect 378200 22129 378224 22163
rect 378200 22061 378224 22095
rect 374718 21881 377718 22009
rect 378200 21993 378224 22027
rect 378200 21925 378224 21959
rect 378200 21857 378224 21891
rect 374718 21725 377718 21853
rect 378200 21789 378224 21823
rect 378200 21721 378224 21755
rect 374718 21569 377718 21697
rect 378200 21653 378224 21687
rect 378200 21585 378224 21619
rect 374599 21471 374627 21499
rect 374718 21413 377718 21541
rect 378200 21517 378224 21551
rect 378200 21449 378224 21483
rect 412429 21481 412472 22881
rect 412579 21481 412707 22881
rect 412742 21481 412870 22881
rect 412905 21481 413033 22881
rect 413068 21481 413196 22881
rect 413231 21481 413260 22881
rect 413720 21481 413763 22881
rect 413856 21481 413899 22881
rect 425480 22349 425718 22399
rect 464429 21481 464472 22881
rect 464579 21481 464707 22881
rect 464742 21481 464870 22881
rect 464905 21481 465033 22881
rect 465068 21481 465196 22881
rect 465231 21481 465359 22881
rect 465394 21481 465522 22881
rect 465557 21481 465685 22881
rect 465720 21481 465763 22881
rect 465856 21481 465899 22881
rect 466006 21481 466134 22881
rect 466169 21481 466297 22881
rect 466332 21481 466460 22881
rect 466495 21481 466623 22881
rect 466658 21481 466786 22881
rect 466821 21481 466949 22881
rect 466984 21481 467034 22881
rect 467301 21634 467403 23198
rect 469996 22813 470532 23685
rect 475455 23406 475625 23712
rect 476255 23406 476425 23712
rect 477055 23406 477225 23712
rect 516429 23617 516472 25017
rect 516579 23617 516707 25017
rect 516742 23617 516870 25017
rect 516905 23617 517033 25017
rect 517068 23617 517196 25017
rect 517231 23617 517260 25017
rect 517720 23617 517763 25017
rect 517856 23617 517899 25017
rect 529552 24573 529608 25173
rect 530020 24573 530070 25173
rect 530508 24572 530558 25172
rect 530658 24572 530708 25172
rect 530788 24572 530838 25172
rect 530938 24572 531066 25172
rect 531094 24572 531222 25172
rect 531250 24572 531306 25172
rect 531406 24572 531534 25172
rect 531562 24572 531690 25172
rect 531718 24572 531768 25172
rect 563983 25102 564017 25137
rect 564085 25122 564109 25146
rect 564326 25143 564360 25147
rect 564394 25143 564428 25147
rect 564462 25143 564496 25147
rect 564530 25143 564564 25147
rect 564598 25143 564632 25147
rect 564666 25143 564700 25147
rect 564734 25143 564768 25147
rect 564802 25143 564836 25147
rect 564870 25143 564904 25147
rect 564938 25143 564972 25147
rect 565006 25143 565040 25147
rect 565074 25143 565108 25147
rect 565142 25143 565176 25147
rect 565210 25143 565244 25147
rect 565278 25143 565312 25147
rect 565346 25143 565380 25147
rect 565414 25143 565448 25147
rect 565482 25143 565516 25147
rect 565550 25143 565584 25147
rect 565618 25143 565652 25147
rect 565686 25143 565720 25147
rect 565754 25143 565788 25147
rect 565822 25143 565856 25147
rect 565890 25143 565924 25147
rect 565958 25143 565992 25147
rect 566026 25143 566060 25147
rect 566094 25143 566128 25147
rect 566162 25143 566196 25147
rect 566230 25143 566264 25147
rect 566298 25143 566332 25147
rect 566366 25143 566400 25147
rect 566434 25143 566468 25147
rect 566502 25143 566536 25147
rect 566570 25143 566604 25147
rect 566638 25143 566672 25147
rect 566706 25143 566740 25147
rect 566774 25143 566808 25147
rect 566842 25143 566876 25147
rect 566910 25143 566944 25147
rect 566978 25143 567012 25147
rect 567046 25143 567080 25147
rect 564248 25125 567148 25143
rect 567532 25125 567556 25149
rect 567590 25125 567614 25149
rect 564326 25121 564360 25125
rect 564394 25121 564428 25125
rect 564462 25121 564496 25125
rect 564530 25121 564564 25125
rect 564598 25121 564632 25125
rect 564666 25121 564700 25125
rect 564734 25121 564768 25125
rect 564802 25121 564836 25125
rect 564870 25121 564904 25125
rect 564938 25121 564972 25125
rect 565006 25121 565040 25125
rect 565074 25121 565108 25125
rect 565142 25121 565176 25125
rect 565210 25121 565244 25125
rect 565278 25121 565312 25125
rect 565346 25121 565380 25125
rect 565414 25121 565448 25125
rect 565482 25121 565516 25125
rect 565550 25121 565584 25125
rect 565618 25121 565652 25125
rect 565686 25121 565720 25125
rect 565754 25121 565788 25125
rect 565822 25121 565856 25125
rect 565890 25121 565924 25125
rect 565958 25121 565992 25125
rect 566026 25121 566060 25125
rect 566094 25121 566128 25125
rect 566162 25121 566196 25125
rect 566230 25121 566264 25125
rect 566298 25121 566332 25125
rect 566366 25121 566400 25125
rect 566434 25121 566468 25125
rect 566502 25121 566536 25125
rect 566570 25121 566604 25125
rect 566638 25121 566672 25125
rect 566706 25121 566740 25125
rect 566774 25121 566808 25125
rect 566842 25121 566876 25125
rect 566910 25121 566944 25125
rect 566978 25121 567012 25125
rect 567046 25121 567080 25125
rect 564252 25113 567144 25121
rect 563983 25089 564007 25102
rect 564061 25098 564085 25113
rect 564302 25101 567104 25113
rect 567556 25101 567590 25115
rect 567532 25067 567556 25091
rect 567590 25067 567614 25091
rect 569996 25085 570532 25553
rect 570835 25524 570869 25548
rect 570903 25524 574201 25548
rect 574269 25383 574293 25417
rect 570708 25113 570810 25137
rect 570939 25126 570963 25150
rect 570708 25089 570732 25113
rect 570786 25089 570810 25113
rect 570963 25102 570987 25116
rect 571041 25113 571065 25116
rect 572091 25113 572193 25137
rect 564429 23617 564472 25017
rect 564579 23617 564707 25017
rect 564742 23617 564870 25017
rect 564905 23617 565033 25017
rect 565068 23617 565196 25017
rect 565231 23617 565359 25017
rect 565394 23617 565522 25017
rect 565557 23617 565685 25017
rect 565720 23617 565763 25017
rect 565856 23617 565899 25017
rect 566006 23617 566134 25017
rect 566169 23617 566297 25017
rect 566332 23617 566460 25017
rect 566495 23617 566623 25017
rect 566658 23617 566786 25017
rect 566821 23617 566949 25017
rect 566984 23617 567034 25017
rect 567301 23300 567403 24864
rect 567670 23685 567720 25085
rect 567827 23685 567955 25085
rect 567990 23685 568118 25085
rect 568153 23685 568281 25085
rect 568316 23685 568444 25085
rect 568479 23685 568607 25085
rect 568642 23685 568770 25085
rect 568805 23685 568848 25085
rect 568941 23685 568984 25085
rect 569091 23685 569219 25085
rect 569254 23685 569382 25085
rect 569417 23685 569545 25085
rect 569580 23685 569708 25085
rect 569743 23685 569871 25085
rect 569906 23685 570532 25085
rect 570939 25068 570963 25092
rect 571065 25068 571089 25092
rect 572091 25089 572115 25113
rect 572169 25089 572193 25113
rect 572347 25113 572381 25147
rect 572419 25113 572453 25147
rect 572491 25113 572525 25147
rect 572563 25113 572597 25147
rect 572347 25089 572371 25113
rect 572573 25089 572597 25113
rect 572752 25089 572786 25147
rect 574269 25137 574293 25349
rect 575671 25286 575705 25310
rect 575743 25286 575777 25310
rect 575815 25286 575849 25310
rect 575887 25286 575921 25310
rect 575958 25286 575962 25310
rect 574167 25113 574293 25137
rect 574167 25089 574191 25113
rect 571152 23685 571195 25085
rect 571302 23685 571430 25085
rect 571465 23685 571593 25085
rect 571628 23685 571756 25085
rect 571791 23685 571919 25085
rect 571954 23685 572004 25085
rect 572873 23685 572916 25085
rect 573023 23685 573151 25085
rect 573186 23685 573314 25085
rect 573349 23685 573477 25085
rect 573512 23685 573640 25085
rect 573675 23685 573803 25085
rect 573838 23685 573881 25085
rect 575428 24573 575478 25173
rect 575578 24573 575706 25173
rect 575734 24573 575862 25173
rect 575890 24573 575946 25173
rect 576046 24573 576174 25173
rect 576202 24573 576330 25173
rect 576358 24573 576408 25173
rect 576488 24573 576538 25173
rect 576638 24573 576688 25173
rect 576810 24573 576860 25173
rect 576960 24573 577010 25173
rect 577090 24573 577140 25173
rect 577240 24573 577368 25173
rect 577396 24573 577524 25173
rect 577552 24573 577608 25173
rect 577708 24573 577836 25173
rect 577864 24573 577992 25173
rect 578020 24573 578070 25173
rect 578508 24572 578558 25172
rect 578658 24572 578708 25172
rect 578788 24572 578838 25172
rect 578938 24572 579066 25172
rect 579094 24572 579222 25172
rect 579250 24572 579306 25172
rect 579406 24572 579534 25172
rect 579562 24572 579690 25172
rect 579718 24572 579768 25172
rect 567335 23276 567369 23300
rect 475455 22906 475625 23212
rect 476255 22906 476425 23212
rect 477055 22906 477225 23212
rect 567335 23198 567369 23222
rect 374167 21385 374269 21409
rect 374167 21361 374191 21385
rect 374245 21361 374269 21385
rect 378200 21381 378224 21415
rect 411983 21410 412051 21430
rect 412326 21415 412360 21419
rect 412394 21415 412428 21419
rect 412462 21415 412496 21419
rect 412530 21415 412564 21419
rect 412598 21415 412632 21419
rect 412666 21415 412700 21419
rect 412734 21415 412768 21419
rect 412802 21415 412836 21419
rect 412870 21415 412904 21419
rect 412938 21415 412972 21419
rect 413006 21415 413040 21419
rect 413074 21415 413108 21419
rect 413142 21415 413176 21419
rect 413210 21415 413244 21419
rect 411983 21385 412017 21410
rect 412282 21407 413260 21415
rect 463983 21410 464051 21430
rect 464326 21415 464360 21419
rect 464394 21415 464428 21419
rect 464462 21415 464496 21419
rect 464530 21415 464564 21419
rect 464598 21415 464632 21419
rect 464666 21415 464700 21419
rect 464734 21415 464768 21419
rect 464802 21415 464836 21419
rect 464870 21415 464904 21419
rect 464938 21415 464972 21419
rect 465006 21415 465040 21419
rect 465074 21415 465108 21419
rect 465142 21415 465176 21419
rect 465210 21415 465244 21419
rect 465278 21415 465312 21419
rect 465346 21415 465380 21419
rect 465414 21415 465448 21419
rect 465482 21415 465516 21419
rect 465550 21415 465584 21419
rect 465618 21415 465652 21419
rect 465686 21415 465720 21419
rect 465754 21415 465788 21419
rect 465822 21415 465856 21419
rect 465890 21415 465924 21419
rect 465958 21415 465992 21419
rect 466026 21415 466060 21419
rect 466094 21415 466128 21419
rect 466162 21415 466196 21419
rect 466230 21415 466264 21419
rect 466298 21415 466332 21419
rect 466366 21415 466400 21419
rect 466434 21415 466468 21419
rect 466502 21415 466536 21419
rect 466570 21415 466604 21419
rect 466638 21415 466672 21419
rect 466706 21415 466740 21419
rect 466774 21415 466808 21419
rect 466842 21415 466876 21419
rect 466910 21415 466944 21419
rect 466978 21415 467012 21419
rect 467046 21415 467080 21419
rect 412326 21403 412360 21407
rect 412394 21403 412428 21407
rect 412462 21403 412496 21407
rect 412530 21403 412564 21407
rect 412598 21403 412632 21407
rect 412666 21403 412700 21407
rect 412734 21403 412768 21407
rect 412802 21403 412836 21407
rect 412870 21403 412904 21407
rect 412938 21403 412972 21407
rect 413006 21403 413040 21407
rect 413074 21403 413108 21407
rect 413142 21403 413176 21407
rect 413210 21403 413244 21407
rect 412061 21385 412085 21400
rect 412248 21385 413260 21403
rect 411983 21361 412007 21385
rect 412302 21383 413260 21385
rect 463983 21385 464017 21410
rect 464282 21407 467114 21415
rect 467532 21407 467556 21431
rect 467590 21407 467614 21431
rect 467670 21413 467720 22813
rect 467827 21413 467955 22813
rect 467990 21413 468118 22813
rect 468153 21413 468281 22813
rect 468316 21413 468444 22813
rect 468479 21413 468607 22813
rect 468642 21413 468770 22813
rect 468805 21413 468848 22813
rect 468941 21413 468984 22813
rect 469091 21413 469219 22813
rect 469254 21413 469382 22813
rect 469417 21413 469545 22813
rect 469580 21413 469708 22813
rect 469743 21413 469871 22813
rect 469906 21413 470532 22813
rect 464326 21403 464360 21407
rect 464394 21403 464428 21407
rect 464462 21403 464496 21407
rect 464530 21403 464564 21407
rect 464598 21403 464632 21407
rect 464666 21403 464700 21407
rect 464734 21403 464768 21407
rect 464802 21403 464836 21407
rect 464870 21403 464904 21407
rect 464938 21403 464972 21407
rect 465006 21403 465040 21407
rect 465074 21403 465108 21407
rect 465142 21403 465176 21407
rect 465210 21403 465244 21407
rect 465278 21403 465312 21407
rect 465346 21403 465380 21407
rect 465414 21403 465448 21407
rect 465482 21403 465516 21407
rect 465550 21403 465584 21407
rect 465618 21403 465652 21407
rect 465686 21403 465720 21407
rect 465754 21403 465788 21407
rect 465822 21403 465856 21407
rect 465890 21403 465924 21407
rect 465958 21403 465992 21407
rect 466026 21403 466060 21407
rect 466094 21403 466128 21407
rect 466162 21403 466196 21407
rect 466230 21403 466264 21407
rect 466298 21403 466332 21407
rect 466366 21403 466400 21407
rect 466434 21403 466468 21407
rect 466502 21403 466536 21407
rect 466570 21403 466604 21407
rect 466638 21403 466672 21407
rect 466706 21403 466740 21407
rect 466774 21403 466808 21407
rect 466842 21403 466876 21407
rect 466910 21403 466944 21407
rect 466978 21403 467012 21407
rect 467046 21403 467080 21407
rect 464061 21385 464085 21400
rect 464248 21385 467148 21403
rect 412085 21352 412109 21376
rect 463983 21361 464007 21385
rect 464302 21383 467104 21385
rect 467556 21383 467590 21397
rect 464085 21352 464109 21376
rect 467532 21349 467556 21373
rect 467590 21349 467614 21373
rect 378200 21313 378224 21347
rect 374718 21263 377718 21313
rect 378200 21245 378224 21279
rect 411983 21274 412051 21294
rect 425480 21263 425718 21313
rect 463983 21274 464051 21294
rect 378200 21177 378224 21211
rect 467189 21186 467213 21210
rect 467247 21186 467271 21210
rect 467223 21162 467237 21186
rect 378200 21109 378224 21143
rect 378200 21041 378224 21075
rect 374251 21003 374269 21008
rect 374228 20983 374269 21003
rect 374227 20974 374303 20983
rect 374227 20949 374228 20974
rect 378200 20973 378224 21007
rect 380200 21000 380320 21003
rect 412000 21000 412120 21003
rect 428200 21000 428320 21003
rect 464000 21000 464120 21003
rect 469996 20945 470532 21413
rect 470708 21385 470810 21409
rect 470939 21406 470963 21430
rect 471065 21406 471089 21430
rect 471152 21413 471195 22813
rect 471302 21413 471430 22813
rect 471465 21413 471593 22813
rect 471628 21413 471756 22813
rect 471791 21413 471919 22813
rect 471954 21413 472004 22813
rect 470708 21361 470732 21385
rect 470786 21361 470810 21385
rect 470963 21382 470987 21396
rect 472091 21385 472193 21409
rect 471041 21382 471065 21385
rect 470939 21348 470963 21372
rect 472091 21361 472115 21385
rect 472169 21361 472193 21385
rect 472347 21385 472381 21419
rect 472419 21385 472453 21419
rect 472491 21385 472525 21419
rect 472563 21385 472597 21419
rect 472347 21361 472371 21385
rect 472573 21361 472597 21385
rect 472752 21361 472786 21419
rect 472873 21413 472916 22813
rect 473023 21413 473151 22813
rect 473186 21413 473314 22813
rect 473349 21413 473477 22813
rect 473512 21413 473640 22813
rect 473675 21413 473803 22813
rect 473838 21413 473881 22813
rect 474718 22349 477718 22399
rect 474718 22193 477718 22321
rect 478200 22197 478224 22210
rect 474718 22037 477718 22165
rect 478200 22129 478224 22163
rect 478200 22061 478224 22095
rect 474718 21881 477718 22009
rect 478200 21993 478224 22027
rect 478200 21925 478224 21959
rect 478200 21857 478224 21891
rect 474718 21725 477718 21853
rect 478200 21789 478224 21823
rect 478200 21721 478224 21755
rect 474718 21569 477718 21697
rect 478200 21653 478224 21687
rect 478200 21585 478224 21619
rect 474599 21471 474627 21499
rect 474718 21413 477718 21541
rect 478200 21517 478224 21551
rect 478200 21449 478224 21483
rect 516429 21481 516472 22881
rect 516579 21481 516707 22881
rect 516742 21481 516870 22881
rect 516905 21481 517033 22881
rect 517068 21481 517196 22881
rect 517231 21481 517260 22881
rect 517720 21481 517763 22881
rect 517856 21481 517899 22881
rect 529480 22349 529718 22399
rect 564429 21481 564472 22881
rect 564579 21481 564707 22881
rect 564742 21481 564870 22881
rect 564905 21481 565033 22881
rect 565068 21481 565196 22881
rect 565231 21481 565359 22881
rect 565394 21481 565522 22881
rect 565557 21481 565685 22881
rect 565720 21481 565763 22881
rect 565856 21481 565899 22881
rect 566006 21481 566134 22881
rect 566169 21481 566297 22881
rect 566332 21481 566460 22881
rect 566495 21481 566623 22881
rect 566658 21481 566786 22881
rect 566821 21481 566949 22881
rect 566984 21481 567034 22881
rect 567301 21634 567403 23198
rect 569996 22813 570532 23685
rect 575455 23406 575625 23712
rect 576255 23406 576425 23712
rect 577055 23406 577225 23712
rect 575455 22906 575625 23212
rect 576255 22906 576425 23212
rect 577055 22906 577225 23212
rect 474167 21385 474269 21409
rect 474167 21361 474191 21385
rect 474245 21361 474269 21385
rect 478200 21381 478224 21415
rect 515983 21410 516051 21430
rect 516326 21415 516360 21419
rect 516394 21415 516428 21419
rect 516462 21415 516496 21419
rect 516530 21415 516564 21419
rect 516598 21415 516632 21419
rect 516666 21415 516700 21419
rect 516734 21415 516768 21419
rect 516802 21415 516836 21419
rect 516870 21415 516904 21419
rect 516938 21415 516972 21419
rect 517006 21415 517040 21419
rect 517074 21415 517108 21419
rect 517142 21415 517176 21419
rect 517210 21415 517244 21419
rect 515983 21385 516017 21410
rect 516282 21407 517260 21415
rect 563983 21410 564051 21430
rect 564326 21415 564360 21419
rect 564394 21415 564428 21419
rect 564462 21415 564496 21419
rect 564530 21415 564564 21419
rect 564598 21415 564632 21419
rect 564666 21415 564700 21419
rect 564734 21415 564768 21419
rect 564802 21415 564836 21419
rect 564870 21415 564904 21419
rect 564938 21415 564972 21419
rect 565006 21415 565040 21419
rect 565074 21415 565108 21419
rect 565142 21415 565176 21419
rect 565210 21415 565244 21419
rect 565278 21415 565312 21419
rect 565346 21415 565380 21419
rect 565414 21415 565448 21419
rect 565482 21415 565516 21419
rect 565550 21415 565584 21419
rect 565618 21415 565652 21419
rect 565686 21415 565720 21419
rect 565754 21415 565788 21419
rect 565822 21415 565856 21419
rect 565890 21415 565924 21419
rect 565958 21415 565992 21419
rect 566026 21415 566060 21419
rect 566094 21415 566128 21419
rect 566162 21415 566196 21419
rect 566230 21415 566264 21419
rect 566298 21415 566332 21419
rect 566366 21415 566400 21419
rect 566434 21415 566468 21419
rect 566502 21415 566536 21419
rect 566570 21415 566604 21419
rect 566638 21415 566672 21419
rect 566706 21415 566740 21419
rect 566774 21415 566808 21419
rect 566842 21415 566876 21419
rect 566910 21415 566944 21419
rect 566978 21415 567012 21419
rect 567046 21415 567080 21419
rect 516326 21403 516360 21407
rect 516394 21403 516428 21407
rect 516462 21403 516496 21407
rect 516530 21403 516564 21407
rect 516598 21403 516632 21407
rect 516666 21403 516700 21407
rect 516734 21403 516768 21407
rect 516802 21403 516836 21407
rect 516870 21403 516904 21407
rect 516938 21403 516972 21407
rect 517006 21403 517040 21407
rect 517074 21403 517108 21407
rect 517142 21403 517176 21407
rect 517210 21403 517244 21407
rect 516061 21385 516085 21400
rect 516248 21385 517260 21403
rect 515983 21361 516007 21385
rect 516302 21383 517260 21385
rect 563983 21385 564017 21410
rect 564282 21407 567114 21415
rect 567532 21407 567556 21431
rect 567590 21407 567614 21431
rect 567670 21413 567720 22813
rect 567827 21413 567955 22813
rect 567990 21413 568118 22813
rect 568153 21413 568281 22813
rect 568316 21413 568444 22813
rect 568479 21413 568607 22813
rect 568642 21413 568770 22813
rect 568805 21413 568848 22813
rect 568941 21413 568984 22813
rect 569091 21413 569219 22813
rect 569254 21413 569382 22813
rect 569417 21413 569545 22813
rect 569580 21413 569708 22813
rect 569743 21413 569871 22813
rect 569906 21413 570532 22813
rect 564326 21403 564360 21407
rect 564394 21403 564428 21407
rect 564462 21403 564496 21407
rect 564530 21403 564564 21407
rect 564598 21403 564632 21407
rect 564666 21403 564700 21407
rect 564734 21403 564768 21407
rect 564802 21403 564836 21407
rect 564870 21403 564904 21407
rect 564938 21403 564972 21407
rect 565006 21403 565040 21407
rect 565074 21403 565108 21407
rect 565142 21403 565176 21407
rect 565210 21403 565244 21407
rect 565278 21403 565312 21407
rect 565346 21403 565380 21407
rect 565414 21403 565448 21407
rect 565482 21403 565516 21407
rect 565550 21403 565584 21407
rect 565618 21403 565652 21407
rect 565686 21403 565720 21407
rect 565754 21403 565788 21407
rect 565822 21403 565856 21407
rect 565890 21403 565924 21407
rect 565958 21403 565992 21407
rect 566026 21403 566060 21407
rect 566094 21403 566128 21407
rect 566162 21403 566196 21407
rect 566230 21403 566264 21407
rect 566298 21403 566332 21407
rect 566366 21403 566400 21407
rect 566434 21403 566468 21407
rect 566502 21403 566536 21407
rect 566570 21403 566604 21407
rect 566638 21403 566672 21407
rect 566706 21403 566740 21407
rect 566774 21403 566808 21407
rect 566842 21403 566876 21407
rect 566910 21403 566944 21407
rect 566978 21403 567012 21407
rect 567046 21403 567080 21407
rect 564061 21385 564085 21400
rect 564248 21385 567148 21403
rect 516085 21352 516109 21376
rect 563983 21361 564007 21385
rect 564302 21383 567104 21385
rect 567556 21383 567590 21397
rect 564085 21352 564109 21376
rect 567532 21349 567556 21373
rect 567590 21349 567614 21373
rect 478200 21313 478224 21347
rect 474718 21263 477718 21313
rect 478200 21245 478224 21279
rect 515983 21274 516051 21294
rect 529480 21263 529718 21313
rect 563983 21274 564051 21294
rect 478200 21177 478224 21211
rect 567189 21186 567213 21210
rect 567247 21186 567271 21210
rect 567223 21162 567237 21186
rect 478200 21109 478224 21143
rect 478200 21041 478224 21075
rect 474251 21003 474269 21008
rect 474228 20983 474269 21003
rect 474227 20974 474303 20983
rect 474227 20949 474228 20974
rect 478200 20973 478224 21007
rect 480200 21000 480320 21003
rect 516000 21000 516120 21003
rect 532200 21000 532320 21003
rect 564000 21000 564120 21003
rect 569996 20945 570532 21413
rect 570708 21385 570810 21409
rect 570939 21406 570963 21430
rect 571065 21406 571089 21430
rect 571152 21413 571195 22813
rect 571302 21413 571430 22813
rect 571465 21413 571593 22813
rect 571628 21413 571756 22813
rect 571791 21413 571919 22813
rect 571954 21413 572004 22813
rect 570708 21361 570732 21385
rect 570786 21361 570810 21385
rect 570963 21382 570987 21396
rect 572091 21385 572193 21409
rect 571041 21382 571065 21385
rect 570939 21348 570963 21372
rect 572091 21361 572115 21385
rect 572169 21361 572193 21385
rect 572347 21385 572381 21419
rect 572419 21385 572453 21419
rect 572491 21385 572525 21419
rect 572563 21385 572597 21419
rect 572347 21361 572371 21385
rect 572573 21361 572597 21385
rect 572752 21361 572786 21419
rect 572873 21413 572916 22813
rect 573023 21413 573151 22813
rect 573186 21413 573314 22813
rect 573349 21413 573477 22813
rect 573512 21413 573640 22813
rect 573675 21413 573803 22813
rect 573838 21413 573881 22813
rect 574718 22349 577718 22399
rect 574718 22193 577718 22321
rect 578200 22197 578224 22210
rect 574718 22037 577718 22165
rect 578200 22129 578224 22163
rect 578200 22061 578224 22095
rect 574718 21881 577718 22009
rect 578200 21993 578224 22027
rect 578200 21925 578224 21959
rect 578200 21857 578224 21891
rect 574718 21725 577718 21853
rect 578200 21789 578224 21823
rect 578200 21721 578224 21755
rect 574718 21569 577718 21697
rect 578200 21653 578224 21687
rect 578200 21585 578224 21619
rect 574599 21471 574627 21499
rect 574718 21413 577718 21541
rect 578200 21517 578224 21551
rect 578200 21449 578224 21483
rect 574167 21385 574269 21409
rect 574167 21361 574191 21385
rect 574245 21361 574269 21385
rect 578200 21381 578224 21415
rect 578200 21313 578224 21347
rect 574718 21263 577718 21313
rect 578200 21245 578224 21279
rect 578200 21177 578224 21211
rect 578200 21109 578224 21143
rect 578200 21041 578224 21075
rect 574251 21003 574269 21008
rect 574228 20983 574269 21003
rect 574227 20974 574303 20983
rect 574227 20949 574228 20974
rect 578200 20973 578224 21007
rect 580200 21000 580320 21003
rect 70740 20809 70748 20833
rect 70782 20809 70816 20833
rect 70850 20809 70884 20833
rect 122740 20809 122748 20833
rect 122782 20809 122816 20833
rect 122850 20809 122884 20833
rect 174740 20809 174748 20833
rect 174782 20809 174816 20833
rect 174850 20809 174884 20833
rect 226740 20809 226748 20833
rect 226782 20809 226816 20833
rect 226850 20809 226884 20833
rect 274740 20809 274748 20833
rect 274782 20809 274816 20833
rect 274850 20809 274884 20833
rect 326740 20809 326748 20833
rect 326782 20809 326816 20833
rect 326850 20809 326884 20833
rect 372087 20809 372121 20833
rect 372155 20809 372189 20833
rect 372223 20809 372257 20833
rect 372291 20809 372325 20833
rect 372359 20809 372393 20833
rect 372427 20809 372461 20833
rect 372495 20809 372529 20833
rect 372563 20809 372597 20833
rect 372631 20809 372665 20833
rect 372699 20809 372733 20833
rect 372767 20809 372801 20833
rect 372835 20809 372869 20833
rect 372903 20809 372937 20833
rect 372971 20809 373005 20833
rect 373039 20809 373073 20833
rect 373107 20809 373141 20833
rect 373175 20809 373209 20833
rect 373243 20809 373277 20833
rect 373311 20809 373345 20833
rect 373379 20809 373413 20833
rect 373447 20809 373481 20833
rect 373515 20809 373549 20833
rect 373583 20809 373617 20833
rect 373651 20809 373685 20833
rect 373719 20809 373753 20833
rect 373787 20809 373821 20833
rect 373855 20809 373889 20833
rect 373923 20809 373957 20833
rect 373991 20809 374025 20833
rect 374059 20809 374093 20833
rect 374127 20809 374161 20833
rect 374195 20809 374229 20833
rect 374263 20809 374297 20833
rect 374331 20809 374365 20833
rect 374399 20809 374433 20833
rect 374467 20809 374501 20833
rect 374535 20809 374569 20833
rect 374603 20809 374637 20833
rect 374671 20809 374705 20833
rect 374739 20809 374773 20833
rect 374807 20809 374841 20833
rect 374875 20809 374909 20833
rect 374943 20809 374977 20833
rect 375011 20809 375045 20833
rect 375079 20809 375113 20833
rect 375147 20809 375181 20833
rect 375215 20809 375249 20833
rect 375283 20809 375317 20833
rect 375351 20809 375385 20833
rect 375419 20809 375453 20833
rect 377898 20809 377932 20833
rect 377966 20809 378000 20833
rect 378034 20809 378068 20833
rect 378102 20809 378136 20833
rect 378170 20809 378204 20833
rect 378238 20809 378272 20833
rect 378306 20809 378340 20833
rect 378374 20809 378408 20833
rect 378442 20809 378476 20833
rect 378510 20809 378544 20833
rect 378578 20809 378612 20833
rect 378646 20809 378680 20833
rect 378714 20809 378748 20833
rect 378782 20809 378816 20833
rect 378850 20809 378884 20833
rect 426740 20809 426748 20833
rect 426782 20809 426816 20833
rect 426850 20809 426884 20833
rect 472087 20809 472121 20833
rect 472155 20809 472189 20833
rect 472223 20809 472257 20833
rect 472291 20809 472325 20833
rect 472359 20809 472393 20833
rect 472427 20809 472461 20833
rect 472495 20809 472529 20833
rect 472563 20809 472597 20833
rect 472631 20809 472665 20833
rect 472699 20809 472733 20833
rect 472767 20809 472801 20833
rect 472835 20809 472869 20833
rect 472903 20809 472937 20833
rect 472971 20809 473005 20833
rect 473039 20809 473073 20833
rect 473107 20809 473141 20833
rect 473175 20809 473209 20833
rect 473243 20809 473277 20833
rect 473311 20809 473345 20833
rect 473379 20809 473413 20833
rect 473447 20809 473481 20833
rect 473515 20809 473549 20833
rect 473583 20809 473617 20833
rect 473651 20809 473685 20833
rect 473719 20809 473753 20833
rect 473787 20809 473821 20833
rect 473855 20809 473889 20833
rect 473923 20809 473957 20833
rect 473991 20809 474025 20833
rect 474059 20809 474093 20833
rect 474127 20809 474161 20833
rect 474195 20809 474229 20833
rect 474263 20809 474297 20833
rect 474331 20809 474365 20833
rect 474399 20809 474433 20833
rect 474467 20809 474501 20833
rect 474535 20809 474569 20833
rect 474603 20809 474637 20833
rect 474671 20809 474705 20833
rect 474739 20809 474773 20833
rect 474807 20809 474841 20833
rect 474875 20809 474909 20833
rect 474943 20809 474977 20833
rect 475011 20809 475045 20833
rect 475079 20809 475113 20833
rect 475147 20809 475181 20833
rect 475215 20809 475249 20833
rect 475283 20809 475317 20833
rect 475351 20809 475385 20833
rect 475419 20809 475453 20833
rect 477898 20809 477932 20833
rect 477966 20809 478000 20833
rect 478034 20809 478068 20833
rect 478102 20809 478136 20833
rect 478170 20809 478204 20833
rect 478238 20809 478272 20833
rect 478306 20809 478340 20833
rect 478374 20809 478408 20833
rect 478442 20809 478476 20833
rect 478510 20809 478544 20833
rect 478578 20809 478612 20833
rect 478646 20809 478680 20833
rect 478714 20809 478748 20833
rect 478782 20809 478816 20833
rect 478850 20809 478884 20833
rect 530740 20809 530748 20833
rect 530782 20809 530816 20833
rect 530850 20809 530884 20833
rect 572087 20809 572121 20833
rect 572155 20809 572189 20833
rect 572223 20809 572257 20833
rect 572291 20809 572325 20833
rect 572359 20809 572393 20833
rect 572427 20809 572461 20833
rect 572495 20809 572529 20833
rect 572563 20809 572597 20833
rect 572631 20809 572665 20833
rect 572699 20809 572733 20833
rect 572767 20809 572801 20833
rect 572835 20809 572869 20833
rect 572903 20809 572937 20833
rect 572971 20809 573005 20833
rect 573039 20809 573073 20833
rect 573107 20809 573141 20833
rect 573175 20809 573209 20833
rect 573243 20809 573277 20833
rect 573311 20809 573345 20833
rect 573379 20809 573413 20833
rect 573447 20809 573481 20833
rect 573515 20809 573549 20833
rect 573583 20809 573617 20833
rect 573651 20809 573685 20833
rect 573719 20809 573753 20833
rect 573787 20809 573821 20833
rect 573855 20809 573889 20833
rect 573923 20809 573957 20833
rect 573991 20809 574025 20833
rect 574059 20809 574093 20833
rect 574127 20809 574161 20833
rect 574195 20809 574229 20833
rect 574263 20809 574297 20833
rect 574331 20809 574365 20833
rect 574399 20809 574433 20833
rect 574467 20809 574501 20833
rect 574535 20809 574569 20833
rect 574603 20809 574637 20833
rect 574671 20809 574705 20833
rect 574739 20809 574773 20833
rect 574807 20809 574841 20833
rect 574875 20809 574909 20833
rect 574943 20809 574977 20833
rect 575011 20809 575045 20833
rect 575079 20809 575113 20833
rect 575147 20809 575181 20833
rect 575215 20809 575249 20833
rect 575283 20809 575317 20833
rect 575351 20809 575385 20833
rect 575419 20809 575453 20833
rect 577898 20809 577932 20833
rect 577966 20809 578000 20833
rect 578034 20809 578068 20833
rect 578102 20809 578136 20833
rect 578170 20809 578204 20833
rect 578238 20809 578272 20833
rect 578306 20809 578340 20833
rect 578374 20809 578408 20833
rect 578442 20809 578476 20833
rect 578510 20809 578544 20833
rect 578578 20809 578612 20833
rect 578646 20809 578680 20833
rect 578714 20809 578748 20833
rect 578782 20809 578816 20833
rect 578850 20809 578884 20833
rect 71017 20659 71041 20693
rect 123017 20659 123041 20693
rect 175017 20659 175041 20693
rect 227017 20659 227041 20693
rect 275017 20659 275041 20693
rect 327017 20659 327041 20693
rect 379017 20659 379041 20693
rect 427017 20659 427041 20693
rect 479017 20659 479041 20693
rect 531017 20659 531041 20693
rect 579017 20659 579041 20693
rect 71017 20591 71041 20625
rect 123017 20591 123041 20625
rect 175017 20591 175041 20625
rect 227017 20591 227041 20625
rect 275017 20591 275041 20625
rect 327017 20591 327041 20625
rect 379017 20591 379041 20625
rect 427017 20591 427041 20625
rect 479017 20591 479041 20625
rect 531017 20591 531041 20625
rect 579017 20591 579041 20625
rect 71017 20523 71041 20557
rect 123017 20523 123041 20557
rect 175017 20523 175041 20557
rect 227017 20523 227041 20557
rect 275017 20523 275041 20557
rect 327017 20523 327041 20557
rect 379017 20523 379041 20557
rect 427017 20523 427041 20557
rect 479017 20523 479041 20557
rect 531017 20523 531041 20557
rect 579017 20523 579041 20557
rect 69480 20462 70251 20512
rect 71017 20455 71041 20489
rect 121480 20462 122251 20512
rect 123017 20455 123041 20489
rect 173480 20462 174251 20512
rect 175017 20455 175041 20489
rect 225480 20462 226251 20512
rect 227017 20455 227041 20489
rect 273480 20462 274251 20512
rect 275017 20455 275041 20489
rect 325480 20462 326251 20512
rect 327017 20455 327041 20489
rect 372429 20462 373829 20512
rect 373959 20462 375359 20512
rect 375721 20462 377121 20512
rect 377251 20462 378251 20512
rect 379017 20455 379041 20489
rect 425480 20462 426251 20512
rect 427017 20455 427041 20489
rect 472429 20462 473829 20512
rect 473959 20462 475359 20512
rect 475721 20462 477121 20512
rect 477251 20462 478251 20512
rect 479017 20455 479041 20489
rect 529480 20462 530251 20512
rect 531017 20455 531041 20489
rect 572429 20462 573829 20512
rect 573959 20462 575359 20512
rect 575721 20462 577121 20512
rect 577251 20462 578251 20512
rect 579017 20455 579041 20489
rect 71017 20387 71041 20421
rect 123017 20387 123041 20421
rect 175017 20387 175041 20421
rect 227017 20387 227041 20421
rect 275017 20387 275041 20421
rect 327017 20387 327041 20421
rect 71017 20319 71041 20353
rect 123017 20319 123041 20353
rect 175017 20319 175041 20353
rect 227017 20319 227041 20353
rect 275017 20319 275041 20353
rect 327017 20319 327041 20353
rect 57090 20250 57106 20316
rect 71017 20251 71041 20285
rect 109090 20250 109106 20316
rect 123017 20251 123041 20285
rect 161090 20250 161106 20316
rect 175017 20251 175041 20285
rect 213090 20250 213106 20316
rect 227017 20251 227041 20285
rect 261090 20250 261106 20316
rect 275017 20251 275041 20285
rect 313090 20250 313106 20316
rect 327017 20251 327041 20285
rect 365090 20250 365106 20316
rect 367114 20250 367130 20316
rect 372429 20306 373829 20434
rect 373959 20306 375359 20434
rect 375721 20306 377121 20434
rect 377251 20306 378251 20434
rect 379017 20387 379041 20421
rect 427017 20387 427041 20421
rect 379017 20319 379041 20353
rect 427017 20319 427041 20353
rect 71017 20183 71041 20217
rect 123017 20183 123041 20217
rect 175017 20183 175041 20217
rect 227017 20183 227041 20217
rect 275017 20183 275041 20217
rect 327017 20183 327041 20217
rect 71017 20115 71041 20149
rect 123017 20115 123041 20149
rect 175017 20115 175041 20149
rect 227017 20115 227041 20149
rect 275017 20115 275041 20149
rect 327017 20115 327041 20149
rect 71017 20047 71041 20081
rect 123017 20047 123041 20081
rect 175017 20047 175041 20081
rect 227017 20047 227041 20081
rect 275017 20047 275041 20081
rect 327017 20047 327041 20081
rect 71017 19979 71041 20013
rect 123017 19979 123041 20013
rect 175017 19979 175041 20013
rect 227017 19979 227041 20013
rect 275017 19979 275041 20013
rect 327017 19979 327041 20013
rect 370248 19980 370418 20286
rect 372429 20150 373829 20278
rect 373959 20150 375359 20278
rect 375721 20150 377121 20278
rect 377251 20150 378251 20278
rect 379017 20251 379041 20285
rect 413090 20250 413106 20316
rect 427017 20251 427041 20285
rect 465090 20250 465106 20316
rect 467114 20250 467130 20316
rect 472429 20306 473829 20434
rect 473959 20306 475359 20434
rect 475721 20306 477121 20434
rect 477251 20306 478251 20434
rect 479017 20387 479041 20421
rect 531017 20387 531041 20421
rect 479017 20319 479041 20353
rect 531017 20319 531041 20353
rect 379017 20183 379041 20217
rect 427017 20183 427041 20217
rect 372429 19994 373829 20122
rect 373959 19994 375359 20122
rect 375721 19994 377121 20122
rect 377251 19994 378251 20122
rect 379017 20115 379041 20149
rect 427017 20115 427041 20149
rect 379017 20047 379041 20081
rect 427017 20047 427041 20081
rect 379017 19979 379041 20013
rect 427017 19979 427041 20013
rect 470248 19980 470418 20286
rect 472429 20150 473829 20278
rect 473959 20150 475359 20278
rect 475721 20150 477121 20278
rect 477251 20150 478251 20278
rect 479017 20251 479041 20285
rect 517090 20250 517106 20316
rect 531017 20251 531041 20285
rect 565090 20250 565106 20316
rect 567114 20250 567130 20316
rect 572429 20306 573829 20434
rect 573959 20306 575359 20434
rect 575721 20306 577121 20434
rect 577251 20306 578251 20434
rect 579017 20387 579041 20421
rect 579017 20319 579041 20353
rect 479017 20183 479041 20217
rect 531017 20183 531041 20217
rect 472429 19994 473829 20122
rect 473959 19994 475359 20122
rect 475721 19994 477121 20122
rect 477251 19994 478251 20122
rect 479017 20115 479041 20149
rect 531017 20115 531041 20149
rect 479017 20047 479041 20081
rect 531017 20047 531041 20081
rect 479017 19979 479041 20013
rect 531017 19979 531041 20013
rect 570248 19980 570418 20286
rect 572429 20150 573829 20278
rect 573959 20150 575359 20278
rect 575721 20150 577121 20278
rect 577251 20150 578251 20278
rect 579017 20251 579041 20285
rect 579017 20183 579041 20217
rect 572429 19994 573829 20122
rect 573959 19994 575359 20122
rect 575721 19994 577121 20122
rect 577251 19994 578251 20122
rect 579017 20115 579041 20149
rect 579017 20047 579041 20081
rect 579017 19979 579041 20013
rect 71017 19911 71041 19945
rect 123017 19911 123041 19945
rect 175017 19911 175041 19945
rect 227017 19911 227041 19945
rect 275017 19911 275041 19945
rect 327017 19911 327041 19945
rect 379017 19911 379041 19945
rect 427017 19911 427041 19945
rect 479017 19911 479041 19945
rect 531017 19911 531041 19945
rect 579017 19911 579041 19945
rect 69480 19844 70251 19894
rect 71017 19843 71041 19877
rect 121480 19844 122251 19894
rect 123017 19843 123041 19877
rect 173480 19844 174251 19894
rect 175017 19843 175041 19877
rect 225480 19844 226251 19894
rect 227017 19843 227041 19877
rect 273480 19844 274251 19894
rect 275017 19843 275041 19877
rect 325480 19844 326251 19894
rect 327017 19843 327041 19877
rect 372429 19844 373829 19894
rect 373959 19844 375359 19894
rect 375721 19844 377121 19894
rect 377251 19844 378251 19894
rect 379017 19843 379041 19877
rect 425480 19844 426251 19894
rect 427017 19843 427041 19877
rect 472429 19844 473829 19894
rect 473959 19844 475359 19894
rect 475721 19844 477121 19894
rect 477251 19844 478251 19894
rect 479017 19843 479041 19877
rect 529480 19844 530251 19894
rect 531017 19843 531041 19877
rect 572429 19844 573829 19894
rect 573959 19844 575359 19894
rect 575721 19844 577121 19894
rect 577251 19844 578251 19894
rect 579017 19843 579041 19877
rect 71017 19775 71041 19809
rect 123017 19775 123041 19809
rect 175017 19775 175041 19809
rect 227017 19775 227041 19809
rect 275017 19775 275041 19809
rect 327017 19775 327041 19809
rect 379017 19775 379041 19809
rect 427017 19775 427041 19809
rect 479017 19775 479041 19809
rect 531017 19775 531041 19809
rect 579017 19775 579041 19809
rect 71017 19707 71041 19741
rect 123017 19707 123041 19741
rect 175017 19707 175041 19741
rect 227017 19707 227041 19741
rect 275017 19707 275041 19741
rect 327017 19707 327041 19741
rect 379017 19707 379041 19741
rect 427017 19707 427041 19741
rect 479017 19707 479041 19741
rect 531017 19707 531041 19741
rect 579017 19707 579041 19741
rect 71017 19639 71041 19673
rect 123017 19639 123041 19673
rect 175017 19639 175041 19673
rect 227017 19639 227041 19673
rect 275017 19639 275041 19673
rect 327017 19639 327041 19673
rect 379017 19639 379041 19673
rect 427017 19639 427041 19673
rect 479017 19639 479041 19673
rect 531017 19639 531041 19673
rect 579017 19639 579041 19673
rect 71017 19583 71041 19605
rect 123017 19583 123041 19605
rect 175017 19583 175041 19605
rect 227017 19583 227041 19605
rect 275017 19583 275041 19605
rect 327017 19583 327041 19605
rect 379017 19583 379041 19605
rect 427017 19583 427041 19605
rect 479017 19583 479041 19605
rect 531017 19583 531041 19605
rect 579017 19583 579041 19605
rect 70740 19547 71053 19583
rect 122740 19547 123053 19583
rect 174740 19547 175053 19583
rect 226740 19547 227053 19583
rect 274740 19547 275053 19583
rect 326740 19547 327053 19583
rect 71017 19516 71053 19547
rect 123017 19516 123053 19547
rect 175017 19516 175053 19547
rect 227017 19516 227053 19547
rect 275017 19516 275053 19547
rect 327017 19516 327053 19547
rect 372031 19547 379053 19583
rect 426740 19547 427053 19583
rect 372031 19516 372067 19547
rect 379017 19516 379053 19547
rect 427017 19516 427053 19547
rect 472031 19547 479053 19583
rect 530740 19547 531053 19583
rect 472031 19516 472067 19547
rect 479017 19516 479053 19547
rect 531017 19516 531053 19547
rect 572031 19547 579053 19583
rect 572031 19516 572067 19547
rect 579017 19516 579053 19547
rect 70740 19480 71172 19516
rect 122740 19480 123172 19516
rect 174740 19480 175172 19516
rect 226740 19480 227172 19516
rect 274740 19480 275172 19516
rect 326740 19480 327172 19516
rect 372031 19480 379172 19516
rect 426740 19480 427172 19516
rect 472031 19480 479172 19516
rect 530740 19480 531172 19516
rect 572031 19480 579172 19516
rect 71017 19390 71172 19480
rect 123017 19390 123172 19480
rect 175017 19390 175172 19480
rect 227017 19390 227172 19480
rect 275017 19390 275172 19480
rect 327017 19390 327172 19480
rect 379017 19390 379172 19480
rect 427017 19390 427172 19480
rect 479017 19390 479172 19480
rect 531017 19390 531172 19480
rect 579017 19390 579172 19480
rect 56903 17278 56936 18278
rect 57106 17278 57123 18278
rect 57582 17278 57722 18278
rect 58084 17278 58140 18278
rect 58156 17278 58212 18278
rect 69486 17278 69626 18278
rect 69988 17278 70044 18278
rect 70060 17278 70116 18278
rect 70327 17278 70377 18278
rect 56746 15878 56780 15908
rect 56708 15840 56780 15870
rect 56903 15678 56936 16678
rect 57106 15678 57123 16678
rect 57582 15678 57722 16678
rect 58084 15678 58140 16678
rect 58156 15678 58212 16678
rect 69486 15678 69626 16678
rect 69988 15678 70044 16678
rect 70060 15678 70116 16678
rect 70327 15678 70377 16678
rect 71065 14844 71172 19390
rect 108903 17278 108936 18278
rect 109106 17278 109123 18278
rect 109582 17278 109722 18278
rect 110084 17278 110140 18278
rect 110156 17278 110212 18278
rect 121486 17278 121626 18278
rect 121988 17278 122044 18278
rect 122060 17278 122116 18278
rect 122327 17278 122377 18278
rect 108746 15878 108780 15908
rect 108708 15840 108780 15870
rect 108903 15678 108936 16678
rect 109106 15678 109123 16678
rect 109582 15678 109722 16678
rect 110084 15678 110140 16678
rect 110156 15678 110212 16678
rect 121486 15678 121626 16678
rect 121988 15678 122044 16678
rect 122060 15678 122116 16678
rect 122327 15678 122377 16678
rect 123065 14844 123172 19390
rect 160903 17278 160936 18278
rect 161106 17278 161123 18278
rect 173486 17278 173626 18278
rect 173988 17278 174044 18278
rect 174060 17278 174116 18278
rect 174327 17278 174377 18278
rect 160746 15878 160780 15908
rect 160708 15840 160780 15870
rect 160903 15678 160936 16678
rect 161106 15678 161123 16678
rect 173486 15678 173626 16678
rect 173988 15678 174044 16678
rect 174060 15678 174116 16678
rect 174327 15678 174377 16678
rect 175065 14844 175172 19390
rect 212903 17278 212936 18278
rect 213106 17278 213123 18278
rect 213582 17278 213722 18278
rect 214084 17278 214140 18278
rect 214156 17278 214212 18278
rect 225486 17278 225626 18278
rect 225988 17278 226044 18278
rect 226060 17278 226116 18278
rect 226327 17278 226377 18278
rect 212746 15878 212780 15908
rect 212708 15840 212780 15870
rect 212903 15678 212936 16678
rect 213106 15678 213123 16678
rect 213582 15678 213722 16678
rect 214084 15678 214140 16678
rect 214156 15678 214212 16678
rect 225486 15678 225626 16678
rect 225988 15678 226044 16678
rect 226060 15678 226116 16678
rect 226327 15678 226377 16678
rect 227065 14844 227172 19390
rect 260903 17278 260936 18278
rect 261106 17278 261123 18278
rect 261582 17278 261722 18278
rect 273486 17278 273626 18278
rect 273988 17278 274044 18278
rect 274060 17278 274116 18278
rect 274327 17278 274377 18278
rect 260746 15878 260780 15908
rect 260708 15840 260780 15870
rect 260903 15678 260936 16678
rect 261106 15678 261123 16678
rect 261582 15678 261722 16678
rect 273486 15678 273626 16678
rect 273988 15678 274044 16678
rect 274060 15678 274116 16678
rect 274327 15678 274377 16678
rect 275065 14844 275172 19390
rect 312903 17278 312936 18278
rect 313106 17278 313123 18278
rect 313582 17278 313722 18278
rect 314084 17278 314140 18278
rect 314156 17278 314212 18278
rect 325486 17278 325626 18278
rect 325988 17278 326044 18278
rect 326060 17278 326116 18278
rect 326327 17278 326377 18278
rect 312746 15878 312780 15908
rect 312708 15840 312780 15870
rect 312903 15678 312936 16678
rect 313106 15678 313123 16678
rect 313582 15678 313722 16678
rect 314084 15678 314140 16678
rect 314156 15678 314212 16678
rect 325486 15678 325626 16678
rect 325988 15678 326044 16678
rect 326060 15678 326116 16678
rect 326327 15678 326377 16678
rect 327065 14844 327172 19390
rect 364903 17278 364936 18278
rect 365106 17278 365123 18278
rect 365261 17278 365333 18278
rect 365522 18198 365722 18278
rect 365737 18208 365771 18232
rect 365782 18208 365854 18278
rect 365737 18198 365854 18208
rect 365509 18174 365854 18198
rect 365522 18130 365722 18174
rect 365737 18164 365761 18174
rect 365737 18140 365771 18164
rect 365782 18140 365854 18174
rect 365737 18130 365854 18140
rect 365509 18106 365854 18130
rect 365522 18062 365722 18106
rect 365737 18096 365761 18106
rect 365737 18072 365771 18096
rect 365782 18072 365854 18106
rect 365737 18062 365854 18072
rect 365509 18038 365854 18062
rect 365522 17994 365722 18038
rect 365737 18028 365761 18038
rect 365737 18004 365771 18028
rect 365782 18004 365854 18038
rect 365737 17994 365854 18004
rect 365509 17970 365854 17994
rect 365522 17926 365722 17970
rect 365737 17960 365761 17970
rect 365737 17936 365771 17960
rect 365782 17936 365854 17970
rect 365737 17926 365854 17936
rect 365509 17902 365854 17926
rect 365522 17858 365722 17902
rect 365737 17892 365761 17902
rect 365737 17868 365771 17892
rect 365782 17868 365854 17902
rect 365737 17858 365854 17868
rect 365509 17834 365854 17858
rect 365522 17790 365722 17834
rect 365737 17824 365761 17834
rect 365737 17800 365771 17824
rect 365782 17800 365854 17834
rect 365737 17790 365854 17800
rect 365509 17766 365854 17790
rect 365522 17722 365722 17766
rect 365737 17756 365761 17766
rect 365737 17732 365771 17756
rect 365782 17732 365854 17766
rect 365737 17722 365854 17732
rect 365509 17698 365854 17722
rect 365522 17654 365722 17698
rect 365737 17688 365761 17698
rect 365737 17664 365771 17688
rect 365782 17664 365854 17698
rect 365737 17654 365854 17664
rect 365509 17630 365854 17654
rect 365522 17586 365722 17630
rect 365737 17620 365761 17630
rect 365737 17596 365771 17620
rect 365782 17596 365854 17630
rect 365737 17586 365854 17596
rect 365509 17562 365854 17586
rect 365522 17518 365722 17562
rect 365737 17552 365761 17562
rect 365737 17528 365771 17552
rect 365782 17528 365854 17562
rect 365737 17518 365854 17528
rect 365509 17494 365854 17518
rect 365522 17450 365722 17494
rect 365737 17484 365761 17494
rect 365737 17460 365771 17484
rect 365782 17460 365854 17494
rect 365737 17450 365854 17460
rect 365509 17426 365854 17450
rect 365522 17382 365722 17426
rect 365737 17416 365761 17426
rect 365737 17392 365771 17416
rect 365782 17392 365854 17426
rect 365737 17382 365854 17392
rect 365509 17358 365854 17382
rect 365522 17314 365722 17358
rect 365737 17348 365761 17358
rect 365737 17324 365771 17348
rect 365782 17324 365854 17358
rect 365737 17314 365854 17324
rect 365509 17290 365854 17314
rect 365522 17278 365722 17290
rect 365533 17266 365557 17278
rect 365737 17266 365761 17290
rect 365782 17278 365854 17290
rect 366084 17278 366140 18278
rect 366156 17278 366212 18278
rect 366514 18198 366714 18278
rect 366729 18208 366763 18232
rect 366774 18208 366846 18278
rect 366729 18198 366846 18208
rect 366501 18174 366846 18198
rect 366514 18130 366714 18174
rect 366729 18164 366753 18174
rect 366729 18140 366763 18164
rect 366774 18140 366846 18174
rect 366729 18130 366846 18140
rect 366501 18106 366846 18130
rect 366514 18062 366714 18106
rect 366729 18096 366753 18106
rect 366729 18072 366763 18096
rect 366774 18072 366846 18106
rect 366729 18062 366846 18072
rect 366501 18038 366846 18062
rect 366514 17994 366714 18038
rect 366729 18028 366753 18038
rect 366729 18004 366763 18028
rect 366774 18004 366846 18038
rect 366729 17994 366846 18004
rect 366501 17970 366846 17994
rect 366514 17926 366714 17970
rect 366729 17960 366753 17970
rect 366729 17936 366763 17960
rect 366774 17936 366846 17970
rect 366729 17926 366846 17936
rect 366501 17902 366846 17926
rect 366514 17858 366714 17902
rect 366729 17892 366753 17902
rect 366729 17868 366763 17892
rect 366774 17868 366846 17902
rect 366729 17858 366846 17868
rect 366501 17834 366846 17858
rect 366514 17790 366714 17834
rect 366729 17824 366753 17834
rect 366729 17800 366763 17824
rect 366774 17800 366846 17834
rect 366729 17790 366846 17800
rect 366501 17766 366846 17790
rect 366514 17722 366714 17766
rect 366729 17756 366753 17766
rect 366729 17732 366763 17756
rect 366774 17732 366846 17766
rect 366729 17722 366846 17732
rect 366501 17698 366846 17722
rect 366514 17654 366714 17698
rect 366729 17688 366753 17698
rect 366729 17664 366763 17688
rect 366774 17664 366846 17698
rect 366729 17654 366846 17664
rect 366501 17630 366846 17654
rect 366514 17586 366714 17630
rect 366729 17620 366753 17630
rect 366729 17596 366763 17620
rect 366774 17596 366846 17630
rect 366729 17586 366846 17596
rect 366501 17562 366846 17586
rect 366514 17518 366714 17562
rect 366729 17552 366753 17562
rect 366729 17528 366763 17552
rect 366774 17528 366846 17562
rect 366729 17518 366846 17528
rect 366501 17494 366846 17518
rect 366514 17450 366714 17494
rect 366729 17484 366753 17494
rect 366729 17460 366763 17484
rect 366774 17460 366846 17494
rect 366729 17450 366846 17460
rect 366501 17426 366846 17450
rect 366514 17382 366714 17426
rect 366729 17416 366753 17426
rect 366729 17392 366763 17416
rect 366774 17392 366846 17426
rect 366729 17382 366846 17392
rect 366501 17358 366846 17382
rect 366514 17314 366714 17358
rect 366729 17348 366753 17358
rect 366729 17324 366763 17348
rect 366774 17324 366846 17358
rect 366729 17314 366846 17324
rect 366501 17290 366846 17314
rect 366514 17278 366714 17290
rect 366525 17266 366549 17278
rect 366729 17266 366753 17290
rect 366774 17278 366846 17290
rect 367076 17278 367132 18278
rect 367148 17278 367204 18278
rect 367506 18198 367706 18278
rect 367721 18208 367755 18232
rect 367766 18208 367838 18278
rect 367721 18198 367838 18208
rect 367493 18174 367838 18198
rect 367506 18130 367706 18174
rect 367721 18164 367745 18174
rect 367721 18140 367755 18164
rect 367766 18140 367838 18174
rect 367721 18130 367838 18140
rect 367493 18106 367838 18130
rect 367506 18062 367706 18106
rect 367721 18096 367745 18106
rect 367721 18072 367755 18096
rect 367766 18072 367838 18106
rect 367721 18062 367838 18072
rect 367493 18038 367838 18062
rect 367506 17994 367706 18038
rect 367721 18028 367745 18038
rect 367721 18004 367755 18028
rect 367766 18004 367838 18038
rect 367721 17994 367838 18004
rect 367493 17970 367838 17994
rect 367506 17926 367706 17970
rect 367721 17960 367745 17970
rect 367721 17936 367755 17960
rect 367766 17936 367838 17970
rect 367721 17926 367838 17936
rect 367493 17902 367838 17926
rect 367506 17858 367706 17902
rect 367721 17892 367745 17902
rect 367721 17868 367755 17892
rect 367766 17868 367838 17902
rect 367721 17858 367838 17868
rect 367493 17834 367838 17858
rect 367506 17790 367706 17834
rect 367721 17824 367745 17834
rect 367721 17800 367755 17824
rect 367766 17800 367838 17834
rect 367721 17790 367838 17800
rect 367493 17766 367838 17790
rect 367506 17722 367706 17766
rect 367721 17756 367745 17766
rect 367721 17732 367755 17756
rect 367766 17732 367838 17766
rect 367721 17722 367838 17732
rect 367493 17698 367838 17722
rect 367506 17654 367706 17698
rect 367721 17688 367745 17698
rect 367721 17664 367755 17688
rect 367766 17664 367838 17698
rect 367721 17654 367838 17664
rect 367493 17630 367838 17654
rect 367506 17586 367706 17630
rect 367721 17620 367745 17630
rect 367721 17596 367755 17620
rect 367766 17596 367838 17630
rect 367721 17586 367838 17596
rect 367493 17562 367838 17586
rect 367506 17518 367706 17562
rect 367721 17552 367745 17562
rect 367721 17528 367755 17552
rect 367766 17528 367838 17562
rect 367721 17518 367838 17528
rect 367493 17494 367838 17518
rect 367506 17450 367706 17494
rect 367721 17484 367745 17494
rect 367721 17460 367755 17484
rect 367766 17460 367838 17494
rect 367721 17450 367838 17460
rect 367493 17426 367838 17450
rect 367506 17382 367706 17426
rect 367721 17416 367745 17426
rect 367721 17392 367755 17416
rect 367766 17392 367838 17426
rect 367721 17382 367838 17392
rect 367493 17358 367838 17382
rect 367506 17314 367706 17358
rect 367721 17348 367745 17358
rect 367721 17324 367755 17348
rect 367766 17324 367838 17358
rect 367721 17314 367838 17324
rect 367493 17290 367838 17314
rect 367506 17278 367706 17290
rect 367517 17266 367541 17278
rect 367721 17266 367745 17290
rect 367766 17278 367838 17290
rect 368068 17278 368124 18278
rect 368140 17278 368196 18278
rect 368498 18198 368698 18278
rect 368713 18208 368747 18232
rect 368758 18208 368830 18278
rect 368713 18198 368830 18208
rect 368485 18174 368830 18198
rect 368498 18130 368698 18174
rect 368713 18164 368737 18174
rect 368713 18140 368747 18164
rect 368758 18140 368830 18174
rect 368713 18130 368830 18140
rect 368485 18106 368830 18130
rect 368498 18062 368698 18106
rect 368713 18096 368737 18106
rect 368713 18072 368747 18096
rect 368758 18072 368830 18106
rect 368713 18062 368830 18072
rect 368485 18038 368830 18062
rect 368498 17994 368698 18038
rect 368713 18028 368737 18038
rect 368713 18004 368747 18028
rect 368758 18004 368830 18038
rect 368713 17994 368830 18004
rect 368485 17970 368830 17994
rect 368498 17926 368698 17970
rect 368713 17960 368737 17970
rect 368713 17936 368747 17960
rect 368758 17936 368830 17970
rect 368713 17926 368830 17936
rect 368485 17902 368830 17926
rect 368498 17858 368698 17902
rect 368713 17892 368737 17902
rect 368713 17868 368747 17892
rect 368758 17868 368830 17902
rect 368713 17858 368830 17868
rect 368485 17834 368830 17858
rect 368498 17790 368698 17834
rect 368713 17824 368737 17834
rect 368713 17800 368747 17824
rect 368758 17800 368830 17834
rect 368713 17790 368830 17800
rect 368485 17766 368830 17790
rect 368498 17722 368698 17766
rect 368713 17756 368737 17766
rect 368713 17732 368747 17756
rect 368758 17732 368830 17766
rect 368713 17722 368830 17732
rect 368485 17698 368830 17722
rect 368498 17654 368698 17698
rect 368713 17688 368737 17698
rect 368713 17664 368747 17688
rect 368758 17664 368830 17698
rect 368713 17654 368830 17664
rect 368485 17630 368830 17654
rect 368498 17586 368698 17630
rect 368713 17620 368737 17630
rect 368713 17596 368747 17620
rect 368758 17596 368830 17630
rect 368713 17586 368830 17596
rect 368485 17562 368830 17586
rect 368498 17518 368698 17562
rect 368713 17552 368737 17562
rect 368713 17528 368747 17552
rect 368758 17528 368830 17562
rect 368713 17518 368830 17528
rect 368485 17494 368830 17518
rect 368498 17450 368698 17494
rect 368713 17484 368737 17494
rect 368713 17460 368747 17484
rect 368758 17460 368830 17494
rect 368713 17450 368830 17460
rect 368485 17426 368830 17450
rect 368498 17382 368698 17426
rect 368713 17416 368737 17426
rect 368713 17392 368747 17416
rect 368758 17392 368830 17426
rect 368713 17382 368830 17392
rect 368485 17358 368830 17382
rect 368498 17314 368698 17358
rect 368713 17348 368737 17358
rect 368713 17324 368747 17348
rect 368758 17324 368830 17358
rect 368713 17314 368830 17324
rect 368485 17290 368830 17314
rect 368498 17278 368698 17290
rect 368509 17266 368533 17278
rect 368713 17266 368737 17290
rect 368758 17278 368830 17290
rect 369060 17278 369116 18278
rect 369132 17278 369188 18278
rect 369490 18198 369690 18278
rect 369705 18208 369739 18232
rect 369750 18208 369822 18278
rect 369705 18198 369822 18208
rect 369477 18174 369822 18198
rect 369490 18130 369690 18174
rect 369705 18164 369729 18174
rect 369705 18140 369739 18164
rect 369750 18140 369822 18174
rect 369705 18130 369822 18140
rect 369477 18106 369822 18130
rect 369490 18062 369690 18106
rect 369705 18096 369729 18106
rect 369705 18072 369739 18096
rect 369750 18072 369822 18106
rect 369705 18062 369822 18072
rect 369477 18038 369822 18062
rect 369490 17994 369690 18038
rect 369705 18028 369729 18038
rect 369705 18004 369739 18028
rect 369750 18004 369822 18038
rect 369705 17994 369822 18004
rect 369477 17970 369822 17994
rect 369490 17926 369690 17970
rect 369705 17960 369729 17970
rect 369705 17936 369739 17960
rect 369750 17936 369822 17970
rect 369705 17926 369822 17936
rect 369477 17902 369822 17926
rect 369490 17858 369690 17902
rect 369705 17892 369729 17902
rect 369705 17868 369739 17892
rect 369750 17868 369822 17902
rect 369705 17858 369822 17868
rect 369477 17834 369822 17858
rect 369490 17790 369690 17834
rect 369705 17824 369729 17834
rect 369705 17800 369739 17824
rect 369750 17800 369822 17834
rect 369705 17790 369822 17800
rect 369477 17766 369822 17790
rect 369490 17722 369690 17766
rect 369705 17756 369729 17766
rect 369705 17732 369739 17756
rect 369750 17732 369822 17766
rect 369705 17722 369822 17732
rect 369477 17698 369822 17722
rect 369490 17654 369690 17698
rect 369705 17688 369729 17698
rect 369705 17664 369739 17688
rect 369750 17664 369822 17698
rect 369705 17654 369822 17664
rect 369477 17630 369822 17654
rect 369490 17586 369690 17630
rect 369705 17620 369729 17630
rect 369705 17596 369739 17620
rect 369750 17596 369822 17630
rect 369705 17586 369822 17596
rect 369477 17562 369822 17586
rect 369490 17518 369690 17562
rect 369705 17552 369729 17562
rect 369705 17528 369739 17552
rect 369750 17528 369822 17562
rect 369705 17518 369822 17528
rect 369477 17494 369822 17518
rect 369490 17450 369690 17494
rect 369705 17484 369729 17494
rect 369705 17460 369739 17484
rect 369750 17460 369822 17494
rect 369705 17450 369822 17460
rect 369477 17426 369822 17450
rect 369490 17382 369690 17426
rect 369705 17416 369729 17426
rect 369705 17392 369739 17416
rect 369750 17392 369822 17426
rect 369705 17382 369822 17392
rect 369477 17358 369822 17382
rect 369490 17314 369690 17358
rect 369705 17348 369729 17358
rect 369705 17324 369739 17348
rect 369750 17324 369822 17358
rect 369705 17314 369822 17324
rect 369477 17290 369822 17314
rect 369490 17278 369690 17290
rect 369501 17266 369525 17278
rect 369705 17266 369729 17290
rect 369750 17278 369822 17290
rect 370052 17278 370108 18278
rect 370124 17278 370180 18278
rect 370482 18198 370682 18278
rect 370697 18208 370731 18232
rect 370742 18208 370814 18278
rect 370697 18198 370814 18208
rect 370469 18174 370814 18198
rect 370482 18130 370682 18174
rect 370697 18164 370721 18174
rect 370697 18140 370731 18164
rect 370742 18140 370814 18174
rect 370697 18130 370814 18140
rect 370469 18106 370814 18130
rect 370482 18062 370682 18106
rect 370697 18096 370721 18106
rect 370697 18072 370731 18096
rect 370742 18072 370814 18106
rect 370697 18062 370814 18072
rect 370469 18038 370814 18062
rect 370482 17994 370682 18038
rect 370697 18028 370721 18038
rect 370697 18004 370731 18028
rect 370742 18004 370814 18038
rect 370697 17994 370814 18004
rect 370469 17970 370814 17994
rect 370482 17926 370682 17970
rect 370697 17960 370721 17970
rect 370697 17936 370731 17960
rect 370742 17936 370814 17970
rect 370697 17926 370814 17936
rect 370469 17902 370814 17926
rect 370482 17858 370682 17902
rect 370697 17892 370721 17902
rect 370697 17868 370731 17892
rect 370742 17868 370814 17902
rect 370697 17858 370814 17868
rect 370469 17834 370814 17858
rect 370482 17790 370682 17834
rect 370697 17824 370721 17834
rect 370697 17800 370731 17824
rect 370742 17800 370814 17834
rect 370697 17790 370814 17800
rect 370469 17766 370814 17790
rect 370482 17722 370682 17766
rect 370697 17756 370721 17766
rect 370697 17732 370731 17756
rect 370742 17732 370814 17766
rect 370697 17722 370814 17732
rect 370469 17698 370814 17722
rect 370482 17654 370682 17698
rect 370697 17688 370721 17698
rect 370697 17664 370731 17688
rect 370742 17664 370814 17698
rect 370697 17654 370814 17664
rect 370469 17630 370814 17654
rect 370482 17586 370682 17630
rect 370697 17620 370721 17630
rect 370697 17596 370731 17620
rect 370742 17596 370814 17630
rect 370697 17586 370814 17596
rect 370469 17562 370814 17586
rect 370482 17518 370682 17562
rect 370697 17552 370721 17562
rect 370697 17528 370731 17552
rect 370742 17528 370814 17562
rect 370697 17518 370814 17528
rect 370469 17494 370814 17518
rect 370482 17450 370682 17494
rect 370697 17484 370721 17494
rect 370697 17460 370731 17484
rect 370742 17460 370814 17494
rect 370697 17450 370814 17460
rect 370469 17426 370814 17450
rect 370482 17382 370682 17426
rect 370697 17416 370721 17426
rect 370697 17392 370731 17416
rect 370742 17392 370814 17426
rect 370697 17382 370814 17392
rect 370469 17358 370814 17382
rect 370482 17314 370682 17358
rect 370697 17348 370721 17358
rect 370697 17324 370731 17348
rect 370742 17324 370814 17358
rect 370697 17314 370814 17324
rect 370469 17290 370814 17314
rect 370482 17278 370682 17290
rect 370493 17266 370517 17278
rect 370697 17266 370721 17290
rect 370742 17278 370814 17290
rect 371044 17278 371100 18278
rect 371116 17278 371172 18278
rect 371474 18198 371674 18278
rect 371689 18208 371723 18232
rect 371734 18208 371806 18278
rect 371689 18198 371806 18208
rect 371461 18174 371806 18198
rect 371474 18130 371674 18174
rect 371689 18164 371713 18174
rect 371689 18140 371723 18164
rect 371734 18140 371806 18174
rect 371689 18130 371806 18140
rect 371461 18106 371806 18130
rect 371474 18062 371674 18106
rect 371689 18096 371713 18106
rect 371689 18072 371723 18096
rect 371734 18072 371806 18106
rect 371689 18062 371806 18072
rect 371461 18038 371806 18062
rect 371474 17994 371674 18038
rect 371689 18028 371713 18038
rect 371689 18004 371723 18028
rect 371734 18004 371806 18038
rect 371689 17994 371806 18004
rect 371461 17970 371806 17994
rect 371474 17926 371674 17970
rect 371689 17960 371713 17970
rect 371689 17936 371723 17960
rect 371734 17936 371806 17970
rect 371689 17926 371806 17936
rect 371461 17902 371806 17926
rect 371474 17858 371674 17902
rect 371689 17892 371713 17902
rect 371689 17868 371723 17892
rect 371734 17868 371806 17902
rect 371689 17858 371806 17868
rect 371461 17834 371806 17858
rect 371474 17790 371674 17834
rect 371689 17824 371713 17834
rect 371689 17800 371723 17824
rect 371734 17800 371806 17834
rect 371689 17790 371806 17800
rect 371461 17766 371806 17790
rect 371474 17722 371674 17766
rect 371689 17756 371713 17766
rect 371689 17732 371723 17756
rect 371734 17732 371806 17766
rect 371689 17722 371806 17732
rect 371461 17698 371806 17722
rect 371474 17654 371674 17698
rect 371689 17688 371713 17698
rect 371689 17664 371723 17688
rect 371734 17664 371806 17698
rect 371689 17654 371806 17664
rect 371461 17630 371806 17654
rect 371474 17586 371674 17630
rect 371689 17620 371713 17630
rect 371689 17596 371723 17620
rect 371734 17596 371806 17630
rect 371689 17586 371806 17596
rect 371461 17562 371806 17586
rect 371474 17518 371674 17562
rect 371689 17552 371713 17562
rect 371689 17528 371723 17552
rect 371734 17528 371806 17562
rect 371689 17518 371806 17528
rect 371461 17494 371806 17518
rect 371474 17450 371674 17494
rect 371689 17484 371713 17494
rect 371689 17460 371723 17484
rect 371734 17460 371806 17494
rect 371689 17450 371806 17460
rect 371461 17426 371806 17450
rect 371474 17382 371674 17426
rect 371689 17416 371713 17426
rect 371689 17392 371723 17416
rect 371734 17392 371806 17426
rect 371689 17382 371806 17392
rect 371461 17358 371806 17382
rect 371474 17314 371674 17358
rect 371689 17348 371713 17358
rect 371689 17324 371723 17348
rect 371734 17324 371806 17358
rect 371689 17314 371806 17324
rect 371461 17290 371806 17314
rect 371474 17278 371674 17290
rect 371485 17266 371509 17278
rect 371689 17266 371713 17290
rect 371734 17278 371806 17290
rect 372036 17278 372092 18278
rect 372108 17278 372164 18278
rect 372466 18198 372666 18278
rect 372681 18208 372715 18232
rect 372726 18208 372798 18278
rect 372681 18198 372798 18208
rect 372453 18174 372798 18198
rect 372466 18130 372666 18174
rect 372681 18164 372705 18174
rect 372681 18140 372715 18164
rect 372726 18140 372798 18174
rect 372681 18130 372798 18140
rect 372453 18106 372798 18130
rect 372466 18062 372666 18106
rect 372681 18096 372705 18106
rect 372681 18072 372715 18096
rect 372726 18072 372798 18106
rect 372681 18062 372798 18072
rect 372453 18038 372798 18062
rect 372466 17994 372666 18038
rect 372681 18028 372705 18038
rect 372681 18004 372715 18028
rect 372726 18004 372798 18038
rect 372681 17994 372798 18004
rect 372453 17970 372798 17994
rect 372466 17926 372666 17970
rect 372681 17960 372705 17970
rect 372681 17936 372715 17960
rect 372726 17936 372798 17970
rect 372681 17926 372798 17936
rect 372453 17902 372798 17926
rect 372466 17858 372666 17902
rect 372681 17892 372705 17902
rect 372681 17868 372715 17892
rect 372726 17868 372798 17902
rect 372681 17858 372798 17868
rect 372453 17834 372798 17858
rect 372466 17790 372666 17834
rect 372681 17824 372705 17834
rect 372681 17800 372715 17824
rect 372726 17800 372798 17834
rect 372681 17790 372798 17800
rect 372453 17766 372798 17790
rect 372466 17722 372666 17766
rect 372681 17756 372705 17766
rect 372681 17732 372715 17756
rect 372726 17732 372798 17766
rect 372681 17722 372798 17732
rect 372453 17698 372798 17722
rect 372466 17654 372666 17698
rect 372681 17688 372705 17698
rect 372681 17664 372715 17688
rect 372726 17664 372798 17698
rect 372681 17654 372798 17664
rect 372453 17630 372798 17654
rect 372466 17586 372666 17630
rect 372681 17620 372705 17630
rect 372681 17596 372715 17620
rect 372726 17596 372798 17630
rect 372681 17586 372798 17596
rect 372453 17562 372798 17586
rect 372466 17518 372666 17562
rect 372681 17552 372705 17562
rect 372681 17528 372715 17552
rect 372726 17528 372798 17562
rect 372681 17518 372798 17528
rect 372453 17494 372798 17518
rect 372466 17450 372666 17494
rect 372681 17484 372705 17494
rect 372681 17460 372715 17484
rect 372726 17460 372798 17494
rect 372681 17450 372798 17460
rect 372453 17426 372798 17450
rect 372466 17382 372666 17426
rect 372681 17416 372705 17426
rect 372681 17392 372715 17416
rect 372726 17392 372798 17426
rect 372681 17382 372798 17392
rect 372453 17358 372798 17382
rect 372466 17314 372666 17358
rect 372681 17348 372705 17358
rect 372681 17324 372715 17348
rect 372726 17324 372798 17358
rect 372681 17314 372798 17324
rect 372453 17290 372798 17314
rect 372466 17278 372666 17290
rect 372477 17266 372501 17278
rect 372681 17266 372705 17290
rect 372726 17278 372798 17290
rect 373028 17278 373084 18278
rect 373100 17278 373156 18278
rect 373458 18198 373658 18278
rect 373673 18208 373707 18232
rect 373718 18208 373790 18278
rect 373673 18198 373790 18208
rect 373445 18174 373790 18198
rect 373458 18130 373658 18174
rect 373673 18164 373697 18174
rect 373673 18140 373707 18164
rect 373718 18140 373790 18174
rect 373673 18130 373790 18140
rect 373445 18106 373790 18130
rect 373458 18062 373658 18106
rect 373673 18096 373697 18106
rect 373673 18072 373707 18096
rect 373718 18072 373790 18106
rect 373673 18062 373790 18072
rect 373445 18038 373790 18062
rect 373458 17994 373658 18038
rect 373673 18028 373697 18038
rect 373673 18004 373707 18028
rect 373718 18004 373790 18038
rect 373673 17994 373790 18004
rect 373445 17970 373790 17994
rect 373458 17926 373658 17970
rect 373673 17960 373697 17970
rect 373673 17936 373707 17960
rect 373718 17936 373790 17970
rect 373673 17926 373790 17936
rect 373445 17902 373790 17926
rect 373458 17858 373658 17902
rect 373673 17892 373697 17902
rect 373673 17868 373707 17892
rect 373718 17868 373790 17902
rect 373673 17858 373790 17868
rect 373445 17834 373790 17858
rect 373458 17790 373658 17834
rect 373673 17824 373697 17834
rect 373673 17800 373707 17824
rect 373718 17800 373790 17834
rect 373673 17790 373790 17800
rect 373445 17766 373790 17790
rect 373458 17722 373658 17766
rect 373673 17756 373697 17766
rect 373673 17732 373707 17756
rect 373718 17732 373790 17766
rect 373673 17722 373790 17732
rect 373445 17698 373790 17722
rect 373458 17654 373658 17698
rect 373673 17688 373697 17698
rect 373673 17664 373707 17688
rect 373718 17664 373790 17698
rect 373673 17654 373790 17664
rect 373445 17630 373790 17654
rect 373458 17586 373658 17630
rect 373673 17620 373697 17630
rect 373673 17596 373707 17620
rect 373718 17596 373790 17630
rect 373673 17586 373790 17596
rect 373445 17562 373790 17586
rect 373458 17518 373658 17562
rect 373673 17552 373697 17562
rect 373673 17528 373707 17552
rect 373718 17528 373790 17562
rect 373673 17518 373790 17528
rect 373445 17494 373790 17518
rect 373458 17450 373658 17494
rect 373673 17484 373697 17494
rect 373673 17460 373707 17484
rect 373718 17460 373790 17494
rect 373673 17450 373790 17460
rect 373445 17426 373790 17450
rect 373458 17382 373658 17426
rect 373673 17416 373697 17426
rect 373673 17392 373707 17416
rect 373718 17392 373790 17426
rect 373673 17382 373790 17392
rect 373445 17358 373790 17382
rect 373458 17314 373658 17358
rect 373673 17348 373697 17358
rect 373673 17324 373707 17348
rect 373718 17324 373790 17358
rect 373673 17314 373790 17324
rect 373445 17290 373790 17314
rect 373458 17278 373658 17290
rect 373469 17266 373493 17278
rect 373673 17266 373697 17290
rect 373718 17278 373790 17290
rect 374020 17278 374076 18278
rect 374092 17278 374148 18278
rect 374450 18198 374650 18278
rect 374665 18208 374699 18232
rect 374710 18208 374782 18278
rect 374665 18198 374782 18208
rect 374437 18174 374782 18198
rect 374450 18130 374650 18174
rect 374665 18164 374689 18174
rect 374665 18140 374699 18164
rect 374710 18140 374782 18174
rect 374665 18130 374782 18140
rect 374437 18106 374782 18130
rect 374450 18062 374650 18106
rect 374665 18096 374689 18106
rect 374665 18072 374699 18096
rect 374710 18072 374782 18106
rect 374665 18062 374782 18072
rect 374437 18038 374782 18062
rect 374450 17994 374650 18038
rect 374665 18028 374689 18038
rect 374665 18004 374699 18028
rect 374710 18004 374782 18038
rect 374665 17994 374782 18004
rect 374437 17970 374782 17994
rect 374450 17926 374650 17970
rect 374665 17960 374689 17970
rect 374665 17936 374699 17960
rect 374710 17936 374782 17970
rect 374665 17926 374782 17936
rect 374437 17902 374782 17926
rect 374450 17858 374650 17902
rect 374665 17892 374689 17902
rect 374665 17868 374699 17892
rect 374710 17868 374782 17902
rect 374665 17858 374782 17868
rect 374437 17834 374782 17858
rect 374450 17790 374650 17834
rect 374665 17824 374689 17834
rect 374665 17800 374699 17824
rect 374710 17800 374782 17834
rect 374665 17790 374782 17800
rect 374437 17766 374782 17790
rect 374450 17722 374650 17766
rect 374665 17756 374689 17766
rect 374665 17732 374699 17756
rect 374710 17732 374782 17766
rect 374665 17722 374782 17732
rect 374437 17698 374782 17722
rect 374450 17654 374650 17698
rect 374665 17688 374689 17698
rect 374665 17664 374699 17688
rect 374710 17664 374782 17698
rect 374665 17654 374782 17664
rect 374437 17630 374782 17654
rect 374450 17586 374650 17630
rect 374665 17620 374689 17630
rect 374665 17596 374699 17620
rect 374710 17596 374782 17630
rect 374665 17586 374782 17596
rect 374437 17562 374782 17586
rect 374450 17518 374650 17562
rect 374665 17552 374689 17562
rect 374665 17528 374699 17552
rect 374710 17528 374782 17562
rect 374665 17518 374782 17528
rect 374437 17494 374782 17518
rect 374450 17450 374650 17494
rect 374665 17484 374689 17494
rect 374665 17460 374699 17484
rect 374710 17460 374782 17494
rect 374665 17450 374782 17460
rect 374437 17426 374782 17450
rect 374450 17382 374650 17426
rect 374665 17416 374689 17426
rect 374665 17392 374699 17416
rect 374710 17392 374782 17426
rect 374665 17382 374782 17392
rect 374437 17358 374782 17382
rect 374450 17314 374650 17358
rect 374665 17348 374689 17358
rect 374665 17324 374699 17348
rect 374710 17324 374782 17358
rect 374665 17314 374782 17324
rect 374437 17290 374782 17314
rect 374450 17278 374650 17290
rect 374461 17266 374485 17278
rect 374665 17266 374689 17290
rect 374710 17278 374782 17290
rect 375012 17278 375068 18278
rect 375084 17278 375140 18278
rect 375442 18198 375642 18278
rect 375657 18208 375691 18232
rect 375702 18208 375774 18278
rect 375657 18198 375774 18208
rect 375429 18174 375774 18198
rect 375442 18130 375642 18174
rect 375657 18164 375681 18174
rect 375657 18140 375691 18164
rect 375702 18140 375774 18174
rect 375657 18130 375774 18140
rect 375429 18106 375774 18130
rect 375442 18062 375642 18106
rect 375657 18096 375681 18106
rect 375657 18072 375691 18096
rect 375702 18072 375774 18106
rect 375657 18062 375774 18072
rect 375429 18038 375774 18062
rect 375442 17994 375642 18038
rect 375657 18028 375681 18038
rect 375657 18004 375691 18028
rect 375702 18004 375774 18038
rect 375657 17994 375774 18004
rect 375429 17970 375774 17994
rect 375442 17926 375642 17970
rect 375657 17960 375681 17970
rect 375657 17936 375691 17960
rect 375702 17936 375774 17970
rect 375657 17926 375774 17936
rect 375429 17902 375774 17926
rect 375442 17858 375642 17902
rect 375657 17892 375681 17902
rect 375657 17868 375691 17892
rect 375702 17868 375774 17902
rect 375657 17858 375774 17868
rect 375429 17834 375774 17858
rect 375442 17790 375642 17834
rect 375657 17824 375681 17834
rect 375657 17800 375691 17824
rect 375702 17800 375774 17834
rect 375657 17790 375774 17800
rect 375429 17766 375774 17790
rect 375442 17722 375642 17766
rect 375657 17756 375681 17766
rect 375657 17732 375691 17756
rect 375702 17732 375774 17766
rect 375657 17722 375774 17732
rect 375429 17698 375774 17722
rect 375442 17654 375642 17698
rect 375657 17688 375681 17698
rect 375657 17664 375691 17688
rect 375702 17664 375774 17698
rect 375657 17654 375774 17664
rect 375429 17630 375774 17654
rect 375442 17586 375642 17630
rect 375657 17620 375681 17630
rect 375657 17596 375691 17620
rect 375702 17596 375774 17630
rect 375657 17586 375774 17596
rect 375429 17562 375774 17586
rect 375442 17518 375642 17562
rect 375657 17552 375681 17562
rect 375657 17528 375691 17552
rect 375702 17528 375774 17562
rect 375657 17518 375774 17528
rect 375429 17494 375774 17518
rect 375442 17450 375642 17494
rect 375657 17484 375681 17494
rect 375657 17460 375691 17484
rect 375702 17460 375774 17494
rect 375657 17450 375774 17460
rect 375429 17426 375774 17450
rect 375442 17382 375642 17426
rect 375657 17416 375681 17426
rect 375657 17392 375691 17416
rect 375702 17392 375774 17426
rect 375657 17382 375774 17392
rect 375429 17358 375774 17382
rect 375442 17314 375642 17358
rect 375657 17348 375681 17358
rect 375657 17324 375691 17348
rect 375702 17324 375774 17358
rect 375657 17314 375774 17324
rect 375429 17290 375774 17314
rect 375442 17278 375642 17290
rect 375453 17266 375477 17278
rect 375657 17266 375681 17290
rect 375702 17278 375774 17290
rect 376004 17278 376060 18278
rect 376076 17278 376132 18278
rect 376434 18198 376634 18278
rect 376649 18208 376683 18232
rect 376694 18208 376766 18278
rect 376649 18198 376766 18208
rect 376421 18174 376766 18198
rect 376434 18130 376634 18174
rect 376649 18164 376673 18174
rect 376649 18140 376683 18164
rect 376694 18140 376766 18174
rect 376649 18130 376766 18140
rect 376421 18106 376766 18130
rect 376434 18062 376634 18106
rect 376649 18096 376673 18106
rect 376649 18072 376683 18096
rect 376694 18072 376766 18106
rect 376649 18062 376766 18072
rect 376421 18038 376766 18062
rect 376434 17994 376634 18038
rect 376649 18028 376673 18038
rect 376649 18004 376683 18028
rect 376694 18004 376766 18038
rect 376649 17994 376766 18004
rect 376421 17970 376766 17994
rect 376434 17926 376634 17970
rect 376649 17960 376673 17970
rect 376649 17936 376683 17960
rect 376694 17936 376766 17970
rect 376649 17926 376766 17936
rect 376421 17902 376766 17926
rect 376434 17858 376634 17902
rect 376649 17892 376673 17902
rect 376649 17868 376683 17892
rect 376694 17868 376766 17902
rect 376649 17858 376766 17868
rect 376421 17834 376766 17858
rect 376434 17790 376634 17834
rect 376649 17824 376673 17834
rect 376649 17800 376683 17824
rect 376694 17800 376766 17834
rect 376649 17790 376766 17800
rect 376421 17766 376766 17790
rect 376434 17722 376634 17766
rect 376649 17756 376673 17766
rect 376649 17732 376683 17756
rect 376694 17732 376766 17766
rect 376649 17722 376766 17732
rect 376421 17698 376766 17722
rect 376434 17654 376634 17698
rect 376649 17688 376673 17698
rect 376649 17664 376683 17688
rect 376694 17664 376766 17698
rect 376649 17654 376766 17664
rect 376421 17630 376766 17654
rect 376434 17586 376634 17630
rect 376649 17620 376673 17630
rect 376649 17596 376683 17620
rect 376694 17596 376766 17630
rect 376649 17586 376766 17596
rect 376421 17562 376766 17586
rect 376434 17518 376634 17562
rect 376649 17552 376673 17562
rect 376649 17528 376683 17552
rect 376694 17528 376766 17562
rect 376649 17518 376766 17528
rect 376421 17494 376766 17518
rect 376434 17450 376634 17494
rect 376649 17484 376673 17494
rect 376649 17460 376683 17484
rect 376694 17460 376766 17494
rect 376649 17450 376766 17460
rect 376421 17426 376766 17450
rect 376434 17382 376634 17426
rect 376649 17416 376673 17426
rect 376649 17392 376683 17416
rect 376694 17392 376766 17426
rect 376649 17382 376766 17392
rect 376421 17358 376766 17382
rect 376434 17314 376634 17358
rect 376649 17348 376673 17358
rect 376649 17324 376683 17348
rect 376694 17324 376766 17358
rect 376649 17314 376766 17324
rect 376421 17290 376766 17314
rect 376434 17278 376634 17290
rect 376445 17266 376469 17278
rect 376649 17266 376673 17290
rect 376694 17278 376766 17290
rect 376996 17278 377052 18278
rect 377068 17278 377124 18278
rect 377426 18198 377626 18278
rect 377641 18208 377675 18232
rect 377686 18208 377758 18278
rect 377641 18198 377758 18208
rect 377413 18174 377758 18198
rect 377426 18130 377626 18174
rect 377641 18164 377665 18174
rect 377641 18140 377675 18164
rect 377686 18140 377758 18174
rect 377641 18130 377758 18140
rect 377413 18106 377758 18130
rect 377426 18062 377626 18106
rect 377641 18096 377665 18106
rect 377641 18072 377675 18096
rect 377686 18072 377758 18106
rect 377641 18062 377758 18072
rect 377413 18038 377758 18062
rect 377426 17994 377626 18038
rect 377641 18028 377665 18038
rect 377641 18004 377675 18028
rect 377686 18004 377758 18038
rect 377641 17994 377758 18004
rect 377413 17970 377758 17994
rect 377426 17926 377626 17970
rect 377641 17960 377665 17970
rect 377641 17936 377675 17960
rect 377686 17936 377758 17970
rect 377641 17926 377758 17936
rect 377413 17902 377758 17926
rect 377426 17858 377626 17902
rect 377641 17892 377665 17902
rect 377641 17868 377675 17892
rect 377686 17868 377758 17902
rect 377641 17858 377758 17868
rect 377413 17834 377758 17858
rect 377426 17790 377626 17834
rect 377641 17824 377665 17834
rect 377641 17800 377675 17824
rect 377686 17800 377758 17834
rect 377641 17790 377758 17800
rect 377413 17766 377758 17790
rect 377426 17722 377626 17766
rect 377641 17756 377665 17766
rect 377641 17732 377675 17756
rect 377686 17732 377758 17766
rect 377641 17722 377758 17732
rect 377413 17698 377758 17722
rect 377426 17654 377626 17698
rect 377641 17688 377665 17698
rect 377641 17664 377675 17688
rect 377686 17664 377758 17698
rect 377641 17654 377758 17664
rect 377413 17630 377758 17654
rect 377426 17586 377626 17630
rect 377641 17620 377665 17630
rect 377641 17596 377675 17620
rect 377686 17596 377758 17630
rect 377641 17586 377758 17596
rect 377413 17562 377758 17586
rect 377426 17518 377626 17562
rect 377641 17552 377665 17562
rect 377641 17528 377675 17552
rect 377686 17528 377758 17562
rect 377641 17518 377758 17528
rect 377413 17494 377758 17518
rect 377426 17450 377626 17494
rect 377641 17484 377665 17494
rect 377641 17460 377675 17484
rect 377686 17460 377758 17494
rect 377641 17450 377758 17460
rect 377413 17426 377758 17450
rect 377426 17382 377626 17426
rect 377641 17416 377665 17426
rect 377641 17392 377675 17416
rect 377686 17392 377758 17426
rect 377641 17382 377758 17392
rect 377413 17358 377758 17382
rect 377426 17314 377626 17358
rect 377641 17348 377665 17358
rect 377641 17324 377675 17348
rect 377686 17324 377758 17358
rect 377641 17314 377758 17324
rect 377413 17290 377758 17314
rect 377426 17278 377626 17290
rect 377437 17266 377461 17278
rect 377641 17266 377665 17290
rect 377686 17278 377758 17290
rect 377988 17278 378044 18278
rect 378060 17278 378116 18278
rect 378327 17278 378377 18278
rect 365533 16678 365567 16690
rect 364746 15878 364780 15908
rect 364708 15840 364780 15870
rect 364903 15678 364936 16678
rect 365106 15678 365123 16678
rect 365261 15678 365333 16678
rect 365522 16656 365722 16678
rect 365737 16666 365771 16690
rect 366525 16678 366559 16690
rect 365782 16666 365854 16678
rect 365737 16656 365854 16666
rect 365509 16632 365854 16656
rect 365522 16588 365722 16632
rect 365737 16622 365761 16632
rect 365737 16598 365771 16622
rect 365782 16598 365854 16632
rect 365737 16588 365854 16598
rect 365509 16564 365854 16588
rect 365522 16520 365722 16564
rect 365737 16554 365761 16564
rect 365737 16530 365771 16554
rect 365782 16530 365854 16564
rect 365737 16520 365854 16530
rect 365509 16496 365854 16520
rect 365522 16452 365722 16496
rect 365737 16486 365761 16496
rect 365737 16462 365771 16486
rect 365782 16462 365854 16496
rect 365737 16452 365854 16462
rect 365509 16428 365854 16452
rect 365522 16384 365722 16428
rect 365737 16418 365761 16428
rect 365737 16394 365771 16418
rect 365782 16394 365854 16428
rect 365737 16384 365854 16394
rect 365509 16360 365854 16384
rect 365522 16316 365722 16360
rect 365737 16350 365761 16360
rect 365737 16326 365771 16350
rect 365782 16326 365854 16360
rect 365737 16316 365854 16326
rect 365509 16292 365854 16316
rect 365522 16248 365722 16292
rect 365737 16282 365761 16292
rect 365737 16258 365771 16282
rect 365782 16258 365854 16292
rect 365737 16248 365854 16258
rect 365509 16224 365854 16248
rect 365522 16180 365722 16224
rect 365737 16214 365761 16224
rect 365737 16190 365771 16214
rect 365782 16190 365854 16224
rect 365737 16180 365854 16190
rect 365509 16156 365854 16180
rect 365522 16112 365722 16156
rect 365737 16146 365761 16156
rect 365737 16122 365771 16146
rect 365782 16122 365854 16156
rect 365737 16112 365854 16122
rect 365509 16088 365854 16112
rect 365522 16044 365722 16088
rect 365737 16078 365761 16088
rect 365737 16054 365771 16078
rect 365782 16054 365854 16088
rect 365737 16044 365854 16054
rect 365509 16020 365854 16044
rect 365522 15976 365722 16020
rect 365737 16010 365761 16020
rect 365737 15986 365771 16010
rect 365782 15986 365854 16020
rect 365737 15976 365854 15986
rect 365509 15952 365854 15976
rect 365522 15908 365722 15952
rect 365737 15942 365761 15952
rect 365737 15918 365771 15942
rect 365782 15918 365854 15952
rect 365737 15908 365854 15918
rect 365509 15884 365854 15908
rect 365522 15840 365722 15884
rect 365737 15874 365761 15884
rect 365737 15850 365771 15874
rect 365782 15850 365854 15884
rect 365737 15840 365854 15850
rect 365509 15816 365854 15840
rect 365522 15772 365722 15816
rect 365737 15806 365761 15816
rect 365737 15782 365771 15806
rect 365782 15782 365854 15816
rect 365737 15772 365854 15782
rect 365509 15748 365854 15772
rect 365522 15678 365722 15748
rect 365737 15724 365761 15748
rect 365782 15678 365854 15748
rect 366084 15678 366140 16678
rect 366156 15678 366212 16678
rect 366514 16656 366714 16678
rect 366729 16666 366763 16690
rect 367517 16678 367551 16690
rect 366774 16666 366846 16678
rect 366729 16656 366846 16666
rect 366501 16632 366846 16656
rect 366514 16588 366714 16632
rect 366729 16622 366753 16632
rect 366729 16598 366763 16622
rect 366774 16598 366846 16632
rect 366729 16588 366846 16598
rect 366501 16564 366846 16588
rect 366514 16520 366714 16564
rect 366729 16554 366753 16564
rect 366729 16530 366763 16554
rect 366774 16530 366846 16564
rect 366729 16520 366846 16530
rect 366501 16496 366846 16520
rect 366514 16452 366714 16496
rect 366729 16486 366753 16496
rect 366729 16462 366763 16486
rect 366774 16462 366846 16496
rect 366729 16452 366846 16462
rect 366501 16428 366846 16452
rect 366514 16384 366714 16428
rect 366729 16418 366753 16428
rect 366729 16394 366763 16418
rect 366774 16394 366846 16428
rect 366729 16384 366846 16394
rect 366501 16360 366846 16384
rect 366514 16316 366714 16360
rect 366729 16350 366753 16360
rect 366729 16326 366763 16350
rect 366774 16326 366846 16360
rect 366729 16316 366846 16326
rect 366501 16292 366846 16316
rect 366514 16248 366714 16292
rect 366729 16282 366753 16292
rect 366729 16258 366763 16282
rect 366774 16258 366846 16292
rect 366729 16248 366846 16258
rect 366501 16224 366846 16248
rect 366514 16180 366714 16224
rect 366729 16214 366753 16224
rect 366729 16190 366763 16214
rect 366774 16190 366846 16224
rect 366729 16180 366846 16190
rect 366501 16156 366846 16180
rect 366514 16112 366714 16156
rect 366729 16146 366753 16156
rect 366729 16122 366763 16146
rect 366774 16122 366846 16156
rect 366729 16112 366846 16122
rect 366501 16088 366846 16112
rect 366514 16044 366714 16088
rect 366729 16078 366753 16088
rect 366729 16054 366763 16078
rect 366774 16054 366846 16088
rect 366729 16044 366846 16054
rect 366501 16020 366846 16044
rect 366514 15976 366714 16020
rect 366729 16010 366753 16020
rect 366729 15986 366763 16010
rect 366774 15986 366846 16020
rect 366729 15976 366846 15986
rect 366501 15952 366846 15976
rect 366514 15908 366714 15952
rect 366729 15942 366753 15952
rect 366729 15918 366763 15942
rect 366774 15918 366846 15952
rect 366729 15908 366846 15918
rect 366501 15884 366846 15908
rect 366514 15840 366714 15884
rect 366729 15874 366753 15884
rect 366729 15850 366763 15874
rect 366774 15850 366846 15884
rect 366729 15840 366846 15850
rect 366501 15816 366846 15840
rect 366514 15772 366714 15816
rect 366729 15806 366753 15816
rect 366729 15782 366763 15806
rect 366774 15782 366846 15816
rect 366729 15772 366846 15782
rect 366501 15748 366846 15772
rect 366514 15678 366714 15748
rect 366729 15724 366753 15748
rect 366774 15678 366846 15748
rect 367076 15678 367132 16678
rect 367148 15678 367204 16678
rect 367506 16656 367706 16678
rect 367721 16666 367755 16690
rect 368509 16678 368543 16690
rect 367766 16666 367838 16678
rect 367721 16656 367838 16666
rect 367493 16632 367838 16656
rect 367506 16588 367706 16632
rect 367721 16622 367745 16632
rect 367721 16598 367755 16622
rect 367766 16598 367838 16632
rect 367721 16588 367838 16598
rect 367493 16564 367838 16588
rect 367506 16520 367706 16564
rect 367721 16554 367745 16564
rect 367721 16530 367755 16554
rect 367766 16530 367838 16564
rect 367721 16520 367838 16530
rect 367493 16496 367838 16520
rect 367506 16452 367706 16496
rect 367721 16486 367745 16496
rect 367721 16462 367755 16486
rect 367766 16462 367838 16496
rect 367721 16452 367838 16462
rect 367493 16428 367838 16452
rect 367506 16384 367706 16428
rect 367721 16418 367745 16428
rect 367721 16394 367755 16418
rect 367766 16394 367838 16428
rect 367721 16384 367838 16394
rect 367493 16360 367838 16384
rect 367506 16316 367706 16360
rect 367721 16350 367745 16360
rect 367721 16326 367755 16350
rect 367766 16326 367838 16360
rect 367721 16316 367838 16326
rect 367493 16292 367838 16316
rect 367506 16248 367706 16292
rect 367721 16282 367745 16292
rect 367721 16258 367755 16282
rect 367766 16258 367838 16292
rect 367721 16248 367838 16258
rect 367493 16224 367838 16248
rect 367506 16180 367706 16224
rect 367721 16214 367745 16224
rect 367721 16190 367755 16214
rect 367766 16190 367838 16224
rect 367721 16180 367838 16190
rect 367493 16156 367838 16180
rect 367506 16112 367706 16156
rect 367721 16146 367745 16156
rect 367721 16122 367755 16146
rect 367766 16122 367838 16156
rect 367721 16112 367838 16122
rect 367493 16088 367838 16112
rect 367506 16044 367706 16088
rect 367721 16078 367745 16088
rect 367721 16054 367755 16078
rect 367766 16054 367838 16088
rect 367721 16044 367838 16054
rect 367493 16020 367838 16044
rect 367506 15976 367706 16020
rect 367721 16010 367745 16020
rect 367721 15986 367755 16010
rect 367766 15986 367838 16020
rect 367721 15976 367838 15986
rect 367493 15952 367838 15976
rect 367506 15908 367706 15952
rect 367721 15942 367745 15952
rect 367721 15918 367755 15942
rect 367766 15918 367838 15952
rect 367721 15908 367838 15918
rect 367493 15884 367838 15908
rect 367506 15840 367706 15884
rect 367721 15874 367745 15884
rect 367721 15850 367755 15874
rect 367766 15850 367838 15884
rect 367721 15840 367838 15850
rect 367493 15816 367838 15840
rect 367506 15772 367706 15816
rect 367721 15806 367745 15816
rect 367721 15782 367755 15806
rect 367766 15782 367838 15816
rect 367721 15772 367838 15782
rect 367493 15748 367838 15772
rect 367506 15678 367706 15748
rect 367721 15724 367745 15748
rect 367766 15678 367838 15748
rect 368068 15678 368124 16678
rect 368140 15678 368196 16678
rect 368498 16656 368698 16678
rect 368713 16666 368747 16690
rect 369501 16678 369535 16690
rect 368758 16666 368830 16678
rect 368713 16656 368830 16666
rect 368485 16632 368830 16656
rect 368498 16588 368698 16632
rect 368713 16622 368737 16632
rect 368713 16598 368747 16622
rect 368758 16598 368830 16632
rect 368713 16588 368830 16598
rect 368485 16564 368830 16588
rect 368498 16520 368698 16564
rect 368713 16554 368737 16564
rect 368713 16530 368747 16554
rect 368758 16530 368830 16564
rect 368713 16520 368830 16530
rect 368485 16496 368830 16520
rect 368498 16452 368698 16496
rect 368713 16486 368737 16496
rect 368713 16462 368747 16486
rect 368758 16462 368830 16496
rect 368713 16452 368830 16462
rect 368485 16428 368830 16452
rect 368498 16384 368698 16428
rect 368713 16418 368737 16428
rect 368713 16394 368747 16418
rect 368758 16394 368830 16428
rect 368713 16384 368830 16394
rect 368485 16360 368830 16384
rect 368498 16316 368698 16360
rect 368713 16350 368737 16360
rect 368713 16326 368747 16350
rect 368758 16326 368830 16360
rect 368713 16316 368830 16326
rect 368485 16292 368830 16316
rect 368498 16248 368698 16292
rect 368713 16282 368737 16292
rect 368713 16258 368747 16282
rect 368758 16258 368830 16292
rect 368713 16248 368830 16258
rect 368485 16224 368830 16248
rect 368498 16180 368698 16224
rect 368713 16214 368737 16224
rect 368713 16190 368747 16214
rect 368758 16190 368830 16224
rect 368713 16180 368830 16190
rect 368485 16156 368830 16180
rect 368498 16112 368698 16156
rect 368713 16146 368737 16156
rect 368713 16122 368747 16146
rect 368758 16122 368830 16156
rect 368713 16112 368830 16122
rect 368485 16088 368830 16112
rect 368498 16044 368698 16088
rect 368713 16078 368737 16088
rect 368713 16054 368747 16078
rect 368758 16054 368830 16088
rect 368713 16044 368830 16054
rect 368485 16020 368830 16044
rect 368498 15976 368698 16020
rect 368713 16010 368737 16020
rect 368713 15986 368747 16010
rect 368758 15986 368830 16020
rect 368713 15976 368830 15986
rect 368485 15952 368830 15976
rect 368498 15908 368698 15952
rect 368713 15942 368737 15952
rect 368713 15918 368747 15942
rect 368758 15918 368830 15952
rect 368713 15908 368830 15918
rect 368485 15884 368830 15908
rect 368498 15840 368698 15884
rect 368713 15874 368737 15884
rect 368713 15850 368747 15874
rect 368758 15850 368830 15884
rect 368713 15840 368830 15850
rect 368485 15816 368830 15840
rect 368498 15772 368698 15816
rect 368713 15806 368737 15816
rect 368713 15782 368747 15806
rect 368758 15782 368830 15816
rect 368713 15772 368830 15782
rect 368485 15748 368830 15772
rect 368498 15678 368698 15748
rect 368713 15724 368737 15748
rect 368758 15678 368830 15748
rect 369060 15678 369116 16678
rect 369132 15678 369188 16678
rect 369490 16656 369690 16678
rect 369705 16666 369739 16690
rect 370493 16678 370527 16690
rect 369750 16666 369822 16678
rect 369705 16656 369822 16666
rect 369477 16632 369822 16656
rect 369490 16588 369690 16632
rect 369705 16622 369729 16632
rect 369705 16598 369739 16622
rect 369750 16598 369822 16632
rect 369705 16588 369822 16598
rect 369477 16564 369822 16588
rect 369490 16520 369690 16564
rect 369705 16554 369729 16564
rect 369705 16530 369739 16554
rect 369750 16530 369822 16564
rect 369705 16520 369822 16530
rect 369477 16496 369822 16520
rect 369490 16452 369690 16496
rect 369705 16486 369729 16496
rect 369705 16462 369739 16486
rect 369750 16462 369822 16496
rect 369705 16452 369822 16462
rect 369477 16428 369822 16452
rect 369490 16384 369690 16428
rect 369705 16418 369729 16428
rect 369705 16394 369739 16418
rect 369750 16394 369822 16428
rect 369705 16384 369822 16394
rect 369477 16360 369822 16384
rect 369490 16316 369690 16360
rect 369705 16350 369729 16360
rect 369705 16326 369739 16350
rect 369750 16326 369822 16360
rect 369705 16316 369822 16326
rect 369477 16292 369822 16316
rect 369490 16248 369690 16292
rect 369705 16282 369729 16292
rect 369705 16258 369739 16282
rect 369750 16258 369822 16292
rect 369705 16248 369822 16258
rect 369477 16224 369822 16248
rect 369490 16180 369690 16224
rect 369705 16214 369729 16224
rect 369705 16190 369739 16214
rect 369750 16190 369822 16224
rect 369705 16180 369822 16190
rect 369477 16156 369822 16180
rect 369490 16112 369690 16156
rect 369705 16146 369729 16156
rect 369705 16122 369739 16146
rect 369750 16122 369822 16156
rect 369705 16112 369822 16122
rect 369477 16088 369822 16112
rect 369490 16044 369690 16088
rect 369705 16078 369729 16088
rect 369705 16054 369739 16078
rect 369750 16054 369822 16088
rect 369705 16044 369822 16054
rect 369477 16020 369822 16044
rect 369490 15976 369690 16020
rect 369705 16010 369729 16020
rect 369705 15986 369739 16010
rect 369750 15986 369822 16020
rect 369705 15976 369822 15986
rect 369477 15952 369822 15976
rect 369490 15908 369690 15952
rect 369705 15942 369729 15952
rect 369705 15918 369739 15942
rect 369750 15918 369822 15952
rect 369705 15908 369822 15918
rect 369477 15884 369822 15908
rect 369490 15840 369690 15884
rect 369705 15874 369729 15884
rect 369705 15850 369739 15874
rect 369750 15850 369822 15884
rect 369705 15840 369822 15850
rect 369477 15816 369822 15840
rect 369490 15772 369690 15816
rect 369705 15806 369729 15816
rect 369705 15782 369739 15806
rect 369750 15782 369822 15816
rect 369705 15772 369822 15782
rect 369477 15748 369822 15772
rect 369490 15678 369690 15748
rect 369705 15724 369729 15748
rect 369750 15678 369822 15748
rect 370052 15678 370108 16678
rect 370124 15678 370180 16678
rect 370482 16656 370682 16678
rect 370697 16666 370731 16690
rect 371485 16678 371519 16690
rect 370742 16666 370814 16678
rect 370697 16656 370814 16666
rect 370469 16632 370814 16656
rect 370482 16588 370682 16632
rect 370697 16622 370721 16632
rect 370697 16598 370731 16622
rect 370742 16598 370814 16632
rect 370697 16588 370814 16598
rect 370469 16564 370814 16588
rect 370482 16520 370682 16564
rect 370697 16554 370721 16564
rect 370697 16530 370731 16554
rect 370742 16530 370814 16564
rect 370697 16520 370814 16530
rect 370469 16496 370814 16520
rect 370482 16452 370682 16496
rect 370697 16486 370721 16496
rect 370697 16462 370731 16486
rect 370742 16462 370814 16496
rect 370697 16452 370814 16462
rect 370469 16428 370814 16452
rect 370482 16384 370682 16428
rect 370697 16418 370721 16428
rect 370697 16394 370731 16418
rect 370742 16394 370814 16428
rect 370697 16384 370814 16394
rect 370469 16360 370814 16384
rect 370482 16316 370682 16360
rect 370697 16350 370721 16360
rect 370697 16326 370731 16350
rect 370742 16326 370814 16360
rect 370697 16316 370814 16326
rect 370469 16292 370814 16316
rect 370482 16248 370682 16292
rect 370697 16282 370721 16292
rect 370697 16258 370731 16282
rect 370742 16258 370814 16292
rect 370697 16248 370814 16258
rect 370469 16224 370814 16248
rect 370482 16180 370682 16224
rect 370697 16214 370721 16224
rect 370697 16190 370731 16214
rect 370742 16190 370814 16224
rect 370697 16180 370814 16190
rect 370469 16156 370814 16180
rect 370482 16112 370682 16156
rect 370697 16146 370721 16156
rect 370697 16122 370731 16146
rect 370742 16122 370814 16156
rect 370697 16112 370814 16122
rect 370469 16088 370814 16112
rect 370482 16044 370682 16088
rect 370697 16078 370721 16088
rect 370697 16054 370731 16078
rect 370742 16054 370814 16088
rect 370697 16044 370814 16054
rect 370469 16020 370814 16044
rect 370482 15976 370682 16020
rect 370697 16010 370721 16020
rect 370697 15986 370731 16010
rect 370742 15986 370814 16020
rect 370697 15976 370814 15986
rect 370469 15952 370814 15976
rect 370482 15908 370682 15952
rect 370697 15942 370721 15952
rect 370697 15918 370731 15942
rect 370742 15918 370814 15952
rect 370697 15908 370814 15918
rect 370469 15884 370814 15908
rect 370482 15840 370682 15884
rect 370697 15874 370721 15884
rect 370697 15850 370731 15874
rect 370742 15850 370814 15884
rect 370697 15840 370814 15850
rect 370469 15816 370814 15840
rect 370482 15772 370682 15816
rect 370697 15806 370721 15816
rect 370697 15782 370731 15806
rect 370742 15782 370814 15816
rect 370697 15772 370814 15782
rect 370469 15748 370814 15772
rect 370482 15678 370682 15748
rect 370697 15724 370721 15748
rect 370742 15678 370814 15748
rect 371044 15678 371100 16678
rect 371116 15678 371172 16678
rect 371474 16656 371674 16678
rect 371689 16666 371723 16690
rect 372477 16678 372511 16690
rect 371734 16666 371806 16678
rect 371689 16656 371806 16666
rect 371461 16632 371806 16656
rect 371474 16588 371674 16632
rect 371689 16622 371713 16632
rect 371689 16598 371723 16622
rect 371734 16598 371806 16632
rect 371689 16588 371806 16598
rect 371461 16564 371806 16588
rect 371474 16520 371674 16564
rect 371689 16554 371713 16564
rect 371689 16530 371723 16554
rect 371734 16530 371806 16564
rect 371689 16520 371806 16530
rect 371461 16496 371806 16520
rect 371474 16452 371674 16496
rect 371689 16486 371713 16496
rect 371689 16462 371723 16486
rect 371734 16462 371806 16496
rect 371689 16452 371806 16462
rect 371461 16428 371806 16452
rect 371474 16384 371674 16428
rect 371689 16418 371713 16428
rect 371689 16394 371723 16418
rect 371734 16394 371806 16428
rect 371689 16384 371806 16394
rect 371461 16360 371806 16384
rect 371474 16316 371674 16360
rect 371689 16350 371713 16360
rect 371689 16326 371723 16350
rect 371734 16326 371806 16360
rect 371689 16316 371806 16326
rect 371461 16292 371806 16316
rect 371474 16248 371674 16292
rect 371689 16282 371713 16292
rect 371689 16258 371723 16282
rect 371734 16258 371806 16292
rect 371689 16248 371806 16258
rect 371461 16224 371806 16248
rect 371474 16180 371674 16224
rect 371689 16214 371713 16224
rect 371689 16190 371723 16214
rect 371734 16190 371806 16224
rect 371689 16180 371806 16190
rect 371461 16156 371806 16180
rect 371474 16112 371674 16156
rect 371689 16146 371713 16156
rect 371689 16122 371723 16146
rect 371734 16122 371806 16156
rect 371689 16112 371806 16122
rect 371461 16088 371806 16112
rect 371474 16044 371674 16088
rect 371689 16078 371713 16088
rect 371689 16054 371723 16078
rect 371734 16054 371806 16088
rect 371689 16044 371806 16054
rect 371461 16020 371806 16044
rect 371474 15976 371674 16020
rect 371689 16010 371713 16020
rect 371689 15986 371723 16010
rect 371734 15986 371806 16020
rect 371689 15976 371806 15986
rect 371461 15952 371806 15976
rect 371474 15908 371674 15952
rect 371689 15942 371713 15952
rect 371689 15918 371723 15942
rect 371734 15918 371806 15952
rect 371689 15908 371806 15918
rect 371461 15884 371806 15908
rect 371474 15840 371674 15884
rect 371689 15874 371713 15884
rect 371689 15850 371723 15874
rect 371734 15850 371806 15884
rect 371689 15840 371806 15850
rect 371461 15816 371806 15840
rect 371474 15772 371674 15816
rect 371689 15806 371713 15816
rect 371689 15782 371723 15806
rect 371734 15782 371806 15816
rect 371689 15772 371806 15782
rect 371461 15748 371806 15772
rect 371474 15678 371674 15748
rect 371689 15724 371713 15748
rect 371734 15678 371806 15748
rect 372036 15678 372092 16678
rect 372108 15678 372164 16678
rect 372466 16656 372666 16678
rect 372681 16666 372715 16690
rect 373469 16678 373503 16690
rect 372726 16666 372798 16678
rect 372681 16656 372798 16666
rect 372453 16632 372798 16656
rect 372466 16588 372666 16632
rect 372681 16622 372705 16632
rect 372681 16598 372715 16622
rect 372726 16598 372798 16632
rect 372681 16588 372798 16598
rect 372453 16564 372798 16588
rect 372466 16520 372666 16564
rect 372681 16554 372705 16564
rect 372681 16530 372715 16554
rect 372726 16530 372798 16564
rect 372681 16520 372798 16530
rect 372453 16496 372798 16520
rect 372466 16452 372666 16496
rect 372681 16486 372705 16496
rect 372681 16462 372715 16486
rect 372726 16462 372798 16496
rect 372681 16452 372798 16462
rect 372453 16428 372798 16452
rect 372466 16384 372666 16428
rect 372681 16418 372705 16428
rect 372681 16394 372715 16418
rect 372726 16394 372798 16428
rect 372681 16384 372798 16394
rect 372453 16360 372798 16384
rect 372466 16316 372666 16360
rect 372681 16350 372705 16360
rect 372681 16326 372715 16350
rect 372726 16326 372798 16360
rect 372681 16316 372798 16326
rect 372453 16292 372798 16316
rect 372466 16248 372666 16292
rect 372681 16282 372705 16292
rect 372681 16258 372715 16282
rect 372726 16258 372798 16292
rect 372681 16248 372798 16258
rect 372453 16224 372798 16248
rect 372466 16180 372666 16224
rect 372681 16214 372705 16224
rect 372681 16190 372715 16214
rect 372726 16190 372798 16224
rect 372681 16180 372798 16190
rect 372453 16156 372798 16180
rect 372466 16112 372666 16156
rect 372681 16146 372705 16156
rect 372681 16122 372715 16146
rect 372726 16122 372798 16156
rect 372681 16112 372798 16122
rect 372453 16088 372798 16112
rect 372466 16044 372666 16088
rect 372681 16078 372705 16088
rect 372681 16054 372715 16078
rect 372726 16054 372798 16088
rect 372681 16044 372798 16054
rect 372453 16020 372798 16044
rect 372466 15976 372666 16020
rect 372681 16010 372705 16020
rect 372681 15986 372715 16010
rect 372726 15986 372798 16020
rect 372681 15976 372798 15986
rect 372453 15952 372798 15976
rect 372466 15908 372666 15952
rect 372681 15942 372705 15952
rect 372681 15918 372715 15942
rect 372726 15918 372798 15952
rect 372681 15908 372798 15918
rect 372453 15884 372798 15908
rect 372466 15840 372666 15884
rect 372681 15874 372705 15884
rect 372681 15850 372715 15874
rect 372726 15850 372798 15884
rect 372681 15840 372798 15850
rect 372453 15816 372798 15840
rect 372466 15772 372666 15816
rect 372681 15806 372705 15816
rect 372681 15782 372715 15806
rect 372726 15782 372798 15816
rect 372681 15772 372798 15782
rect 372453 15748 372798 15772
rect 372466 15678 372666 15748
rect 372681 15724 372705 15748
rect 372726 15678 372798 15748
rect 373028 15678 373084 16678
rect 373100 15678 373156 16678
rect 373458 16656 373658 16678
rect 373673 16666 373707 16690
rect 374461 16678 374495 16690
rect 373718 16666 373790 16678
rect 373673 16656 373790 16666
rect 373445 16632 373790 16656
rect 373458 16588 373658 16632
rect 373673 16622 373697 16632
rect 373673 16598 373707 16622
rect 373718 16598 373790 16632
rect 373673 16588 373790 16598
rect 373445 16564 373790 16588
rect 373458 16520 373658 16564
rect 373673 16554 373697 16564
rect 373673 16530 373707 16554
rect 373718 16530 373790 16564
rect 373673 16520 373790 16530
rect 373445 16496 373790 16520
rect 373458 16452 373658 16496
rect 373673 16486 373697 16496
rect 373673 16462 373707 16486
rect 373718 16462 373790 16496
rect 373673 16452 373790 16462
rect 373445 16428 373790 16452
rect 373458 16384 373658 16428
rect 373673 16418 373697 16428
rect 373673 16394 373707 16418
rect 373718 16394 373790 16428
rect 373673 16384 373790 16394
rect 373445 16360 373790 16384
rect 373458 16316 373658 16360
rect 373673 16350 373697 16360
rect 373673 16326 373707 16350
rect 373718 16326 373790 16360
rect 373673 16316 373790 16326
rect 373445 16292 373790 16316
rect 373458 16248 373658 16292
rect 373673 16282 373697 16292
rect 373673 16258 373707 16282
rect 373718 16258 373790 16292
rect 373673 16248 373790 16258
rect 373445 16224 373790 16248
rect 373458 16180 373658 16224
rect 373673 16214 373697 16224
rect 373673 16190 373707 16214
rect 373718 16190 373790 16224
rect 373673 16180 373790 16190
rect 373445 16156 373790 16180
rect 373458 16112 373658 16156
rect 373673 16146 373697 16156
rect 373673 16122 373707 16146
rect 373718 16122 373790 16156
rect 373673 16112 373790 16122
rect 373445 16088 373790 16112
rect 373458 16044 373658 16088
rect 373673 16078 373697 16088
rect 373673 16054 373707 16078
rect 373718 16054 373790 16088
rect 373673 16044 373790 16054
rect 373445 16020 373790 16044
rect 373458 15976 373658 16020
rect 373673 16010 373697 16020
rect 373673 15986 373707 16010
rect 373718 15986 373790 16020
rect 373673 15976 373790 15986
rect 373445 15952 373790 15976
rect 373458 15908 373658 15952
rect 373673 15942 373697 15952
rect 373673 15918 373707 15942
rect 373718 15918 373790 15952
rect 373673 15908 373790 15918
rect 373445 15884 373790 15908
rect 373458 15840 373658 15884
rect 373673 15874 373697 15884
rect 373673 15850 373707 15874
rect 373718 15850 373790 15884
rect 373673 15840 373790 15850
rect 373445 15816 373790 15840
rect 373458 15772 373658 15816
rect 373673 15806 373697 15816
rect 373673 15782 373707 15806
rect 373718 15782 373790 15816
rect 373673 15772 373790 15782
rect 373445 15748 373790 15772
rect 373458 15678 373658 15748
rect 373673 15724 373697 15748
rect 373718 15678 373790 15748
rect 374020 15678 374076 16678
rect 374092 15678 374148 16678
rect 374450 16656 374650 16678
rect 374665 16666 374699 16690
rect 375453 16678 375487 16690
rect 374710 16666 374782 16678
rect 374665 16656 374782 16666
rect 374437 16632 374782 16656
rect 374450 16588 374650 16632
rect 374665 16622 374689 16632
rect 374665 16598 374699 16622
rect 374710 16598 374782 16632
rect 374665 16588 374782 16598
rect 374437 16564 374782 16588
rect 374450 16520 374650 16564
rect 374665 16554 374689 16564
rect 374665 16530 374699 16554
rect 374710 16530 374782 16564
rect 374665 16520 374782 16530
rect 374437 16496 374782 16520
rect 374450 16452 374650 16496
rect 374665 16486 374689 16496
rect 374665 16462 374699 16486
rect 374710 16462 374782 16496
rect 374665 16452 374782 16462
rect 374437 16428 374782 16452
rect 374450 16384 374650 16428
rect 374665 16418 374689 16428
rect 374665 16394 374699 16418
rect 374710 16394 374782 16428
rect 374665 16384 374782 16394
rect 374437 16360 374782 16384
rect 374450 16316 374650 16360
rect 374665 16350 374689 16360
rect 374665 16326 374699 16350
rect 374710 16326 374782 16360
rect 374665 16316 374782 16326
rect 374437 16292 374782 16316
rect 374450 16248 374650 16292
rect 374665 16282 374689 16292
rect 374665 16258 374699 16282
rect 374710 16258 374782 16292
rect 374665 16248 374782 16258
rect 374437 16224 374782 16248
rect 374450 16180 374650 16224
rect 374665 16214 374689 16224
rect 374665 16190 374699 16214
rect 374710 16190 374782 16224
rect 374665 16180 374782 16190
rect 374437 16156 374782 16180
rect 374450 16112 374650 16156
rect 374665 16146 374689 16156
rect 374665 16122 374699 16146
rect 374710 16122 374782 16156
rect 374665 16112 374782 16122
rect 374437 16088 374782 16112
rect 374450 16044 374650 16088
rect 374665 16078 374689 16088
rect 374665 16054 374699 16078
rect 374710 16054 374782 16088
rect 374665 16044 374782 16054
rect 374437 16020 374782 16044
rect 374450 15976 374650 16020
rect 374665 16010 374689 16020
rect 374665 15986 374699 16010
rect 374710 15986 374782 16020
rect 374665 15976 374782 15986
rect 374437 15952 374782 15976
rect 374450 15908 374650 15952
rect 374665 15942 374689 15952
rect 374665 15918 374699 15942
rect 374710 15918 374782 15952
rect 374665 15908 374782 15918
rect 374437 15884 374782 15908
rect 374450 15840 374650 15884
rect 374665 15874 374689 15884
rect 374665 15850 374699 15874
rect 374710 15850 374782 15884
rect 374665 15840 374782 15850
rect 374437 15816 374782 15840
rect 374450 15772 374650 15816
rect 374665 15806 374689 15816
rect 374665 15782 374699 15806
rect 374710 15782 374782 15816
rect 374665 15772 374782 15782
rect 374437 15748 374782 15772
rect 374450 15678 374650 15748
rect 374665 15724 374689 15748
rect 374710 15678 374782 15748
rect 375012 15678 375068 16678
rect 375084 15678 375140 16678
rect 375442 16656 375642 16678
rect 375657 16666 375691 16690
rect 376445 16678 376479 16690
rect 375702 16666 375774 16678
rect 375657 16656 375774 16666
rect 375429 16632 375774 16656
rect 375442 16588 375642 16632
rect 375657 16622 375681 16632
rect 375657 16598 375691 16622
rect 375702 16598 375774 16632
rect 375657 16588 375774 16598
rect 375429 16564 375774 16588
rect 375442 16520 375642 16564
rect 375657 16554 375681 16564
rect 375657 16530 375691 16554
rect 375702 16530 375774 16564
rect 375657 16520 375774 16530
rect 375429 16496 375774 16520
rect 375442 16452 375642 16496
rect 375657 16486 375681 16496
rect 375657 16462 375691 16486
rect 375702 16462 375774 16496
rect 375657 16452 375774 16462
rect 375429 16428 375774 16452
rect 375442 16384 375642 16428
rect 375657 16418 375681 16428
rect 375657 16394 375691 16418
rect 375702 16394 375774 16428
rect 375657 16384 375774 16394
rect 375429 16360 375774 16384
rect 375442 16316 375642 16360
rect 375657 16350 375681 16360
rect 375657 16326 375691 16350
rect 375702 16326 375774 16360
rect 375657 16316 375774 16326
rect 375429 16292 375774 16316
rect 375442 16248 375642 16292
rect 375657 16282 375681 16292
rect 375657 16258 375691 16282
rect 375702 16258 375774 16292
rect 375657 16248 375774 16258
rect 375429 16224 375774 16248
rect 375442 16180 375642 16224
rect 375657 16214 375681 16224
rect 375657 16190 375691 16214
rect 375702 16190 375774 16224
rect 375657 16180 375774 16190
rect 375429 16156 375774 16180
rect 375442 16112 375642 16156
rect 375657 16146 375681 16156
rect 375657 16122 375691 16146
rect 375702 16122 375774 16156
rect 375657 16112 375774 16122
rect 375429 16088 375774 16112
rect 375442 16044 375642 16088
rect 375657 16078 375681 16088
rect 375657 16054 375691 16078
rect 375702 16054 375774 16088
rect 375657 16044 375774 16054
rect 375429 16020 375774 16044
rect 375442 15976 375642 16020
rect 375657 16010 375681 16020
rect 375657 15986 375691 16010
rect 375702 15986 375774 16020
rect 375657 15976 375774 15986
rect 375429 15952 375774 15976
rect 375442 15908 375642 15952
rect 375657 15942 375681 15952
rect 375657 15918 375691 15942
rect 375702 15918 375774 15952
rect 375657 15908 375774 15918
rect 375429 15884 375774 15908
rect 375442 15840 375642 15884
rect 375657 15874 375681 15884
rect 375657 15850 375691 15874
rect 375702 15850 375774 15884
rect 375657 15840 375774 15850
rect 375429 15816 375774 15840
rect 375442 15772 375642 15816
rect 375657 15806 375681 15816
rect 375657 15782 375691 15806
rect 375702 15782 375774 15816
rect 375657 15772 375774 15782
rect 375429 15748 375774 15772
rect 375442 15678 375642 15748
rect 375657 15724 375681 15748
rect 375702 15678 375774 15748
rect 376004 15678 376060 16678
rect 376076 15678 376132 16678
rect 376434 16656 376634 16678
rect 376649 16666 376683 16690
rect 377437 16678 377471 16690
rect 376694 16666 376766 16678
rect 376649 16656 376766 16666
rect 376421 16632 376766 16656
rect 376434 16588 376634 16632
rect 376649 16622 376673 16632
rect 376649 16598 376683 16622
rect 376694 16598 376766 16632
rect 376649 16588 376766 16598
rect 376421 16564 376766 16588
rect 376434 16520 376634 16564
rect 376649 16554 376673 16564
rect 376649 16530 376683 16554
rect 376694 16530 376766 16564
rect 376649 16520 376766 16530
rect 376421 16496 376766 16520
rect 376434 16452 376634 16496
rect 376649 16486 376673 16496
rect 376649 16462 376683 16486
rect 376694 16462 376766 16496
rect 376649 16452 376766 16462
rect 376421 16428 376766 16452
rect 376434 16384 376634 16428
rect 376649 16418 376673 16428
rect 376649 16394 376683 16418
rect 376694 16394 376766 16428
rect 376649 16384 376766 16394
rect 376421 16360 376766 16384
rect 376434 16316 376634 16360
rect 376649 16350 376673 16360
rect 376649 16326 376683 16350
rect 376694 16326 376766 16360
rect 376649 16316 376766 16326
rect 376421 16292 376766 16316
rect 376434 16248 376634 16292
rect 376649 16282 376673 16292
rect 376649 16258 376683 16282
rect 376694 16258 376766 16292
rect 376649 16248 376766 16258
rect 376421 16224 376766 16248
rect 376434 16180 376634 16224
rect 376649 16214 376673 16224
rect 376649 16190 376683 16214
rect 376694 16190 376766 16224
rect 376649 16180 376766 16190
rect 376421 16156 376766 16180
rect 376434 16112 376634 16156
rect 376649 16146 376673 16156
rect 376649 16122 376683 16146
rect 376694 16122 376766 16156
rect 376649 16112 376766 16122
rect 376421 16088 376766 16112
rect 376434 16044 376634 16088
rect 376649 16078 376673 16088
rect 376649 16054 376683 16078
rect 376694 16054 376766 16088
rect 376649 16044 376766 16054
rect 376421 16020 376766 16044
rect 376434 15976 376634 16020
rect 376649 16010 376673 16020
rect 376649 15986 376683 16010
rect 376694 15986 376766 16020
rect 376649 15976 376766 15986
rect 376421 15952 376766 15976
rect 376434 15908 376634 15952
rect 376649 15942 376673 15952
rect 376649 15918 376683 15942
rect 376694 15918 376766 15952
rect 376649 15908 376766 15918
rect 376421 15884 376766 15908
rect 376434 15840 376634 15884
rect 376649 15874 376673 15884
rect 376649 15850 376683 15874
rect 376694 15850 376766 15884
rect 376649 15840 376766 15850
rect 376421 15816 376766 15840
rect 376434 15772 376634 15816
rect 376649 15806 376673 15816
rect 376649 15782 376683 15806
rect 376694 15782 376766 15816
rect 376649 15772 376766 15782
rect 376421 15748 376766 15772
rect 376434 15678 376634 15748
rect 376649 15724 376673 15748
rect 376694 15678 376766 15748
rect 376996 15678 377052 16678
rect 377068 15678 377124 16678
rect 377426 16656 377626 16678
rect 377641 16666 377675 16690
rect 377686 16666 377758 16678
rect 377641 16656 377758 16666
rect 377413 16632 377758 16656
rect 377426 16588 377626 16632
rect 377641 16622 377665 16632
rect 377641 16598 377675 16622
rect 377686 16598 377758 16632
rect 377641 16588 377758 16598
rect 377413 16564 377758 16588
rect 377426 16520 377626 16564
rect 377641 16554 377665 16564
rect 377641 16530 377675 16554
rect 377686 16530 377758 16564
rect 377641 16520 377758 16530
rect 377413 16496 377758 16520
rect 377426 16452 377626 16496
rect 377641 16486 377665 16496
rect 377641 16462 377675 16486
rect 377686 16462 377758 16496
rect 377641 16452 377758 16462
rect 377413 16428 377758 16452
rect 377426 16384 377626 16428
rect 377641 16418 377665 16428
rect 377641 16394 377675 16418
rect 377686 16394 377758 16428
rect 377641 16384 377758 16394
rect 377413 16360 377758 16384
rect 377426 16316 377626 16360
rect 377641 16350 377665 16360
rect 377641 16326 377675 16350
rect 377686 16326 377758 16360
rect 377641 16316 377758 16326
rect 377413 16292 377758 16316
rect 377426 16248 377626 16292
rect 377641 16282 377665 16292
rect 377641 16258 377675 16282
rect 377686 16258 377758 16292
rect 377641 16248 377758 16258
rect 377413 16224 377758 16248
rect 377426 16180 377626 16224
rect 377641 16214 377665 16224
rect 377641 16190 377675 16214
rect 377686 16190 377758 16224
rect 377641 16180 377758 16190
rect 377413 16156 377758 16180
rect 377426 16112 377626 16156
rect 377641 16146 377665 16156
rect 377641 16122 377675 16146
rect 377686 16122 377758 16156
rect 377641 16112 377758 16122
rect 377413 16088 377758 16112
rect 377426 16044 377626 16088
rect 377641 16078 377665 16088
rect 377641 16054 377675 16078
rect 377686 16054 377758 16088
rect 377641 16044 377758 16054
rect 377413 16020 377758 16044
rect 377426 15976 377626 16020
rect 377641 16010 377665 16020
rect 377641 15986 377675 16010
rect 377686 15986 377758 16020
rect 377641 15976 377758 15986
rect 377413 15952 377758 15976
rect 377426 15908 377626 15952
rect 377641 15942 377665 15952
rect 377641 15918 377675 15942
rect 377686 15918 377758 15952
rect 377641 15908 377758 15918
rect 377413 15884 377758 15908
rect 377426 15840 377626 15884
rect 377641 15874 377665 15884
rect 377641 15850 377675 15874
rect 377686 15850 377758 15884
rect 377641 15840 377758 15850
rect 377413 15816 377758 15840
rect 377426 15772 377626 15816
rect 377641 15806 377665 15816
rect 377641 15782 377675 15806
rect 377686 15782 377758 15816
rect 377641 15772 377758 15782
rect 377413 15748 377758 15772
rect 377426 15678 377626 15748
rect 377641 15724 377665 15748
rect 377686 15678 377758 15748
rect 377988 15678 378044 16678
rect 378060 15678 378116 16678
rect 378327 15678 378377 16678
rect 379065 14844 379172 19390
rect 412903 17278 412936 18278
rect 413106 17278 413123 18278
rect 413582 17278 413722 18278
rect 414084 17278 414140 18278
rect 414156 17278 414212 18278
rect 425486 17278 425626 18278
rect 425988 17278 426044 18278
rect 426060 17278 426116 18278
rect 426327 17278 426377 18278
rect 412746 15878 412780 15908
rect 412708 15840 412780 15870
rect 412903 15678 412936 16678
rect 413106 15678 413123 16678
rect 413582 15678 413722 16678
rect 414084 15678 414140 16678
rect 414156 15678 414212 16678
rect 425486 15678 425626 16678
rect 425988 15678 426044 16678
rect 426060 15678 426116 16678
rect 426327 15678 426377 16678
rect 427065 14844 427172 19390
rect 464903 17278 464936 18278
rect 465106 17278 465123 18278
rect 465261 17278 465333 18278
rect 465522 18198 465722 18278
rect 465737 18208 465771 18232
rect 465782 18208 465854 18278
rect 465737 18198 465854 18208
rect 465509 18174 465854 18198
rect 465522 18130 465722 18174
rect 465737 18164 465761 18174
rect 465737 18140 465771 18164
rect 465782 18140 465854 18174
rect 465737 18130 465854 18140
rect 465509 18106 465854 18130
rect 465522 18062 465722 18106
rect 465737 18096 465761 18106
rect 465737 18072 465771 18096
rect 465782 18072 465854 18106
rect 465737 18062 465854 18072
rect 465509 18038 465854 18062
rect 465522 17994 465722 18038
rect 465737 18028 465761 18038
rect 465737 18004 465771 18028
rect 465782 18004 465854 18038
rect 465737 17994 465854 18004
rect 465509 17970 465854 17994
rect 465522 17926 465722 17970
rect 465737 17960 465761 17970
rect 465737 17936 465771 17960
rect 465782 17936 465854 17970
rect 465737 17926 465854 17936
rect 465509 17902 465854 17926
rect 465522 17858 465722 17902
rect 465737 17892 465761 17902
rect 465737 17868 465771 17892
rect 465782 17868 465854 17902
rect 465737 17858 465854 17868
rect 465509 17834 465854 17858
rect 465522 17790 465722 17834
rect 465737 17824 465761 17834
rect 465737 17800 465771 17824
rect 465782 17800 465854 17834
rect 465737 17790 465854 17800
rect 465509 17766 465854 17790
rect 465522 17722 465722 17766
rect 465737 17756 465761 17766
rect 465737 17732 465771 17756
rect 465782 17732 465854 17766
rect 465737 17722 465854 17732
rect 465509 17698 465854 17722
rect 465522 17654 465722 17698
rect 465737 17688 465761 17698
rect 465737 17664 465771 17688
rect 465782 17664 465854 17698
rect 465737 17654 465854 17664
rect 465509 17630 465854 17654
rect 465522 17586 465722 17630
rect 465737 17620 465761 17630
rect 465737 17596 465771 17620
rect 465782 17596 465854 17630
rect 465737 17586 465854 17596
rect 465509 17562 465854 17586
rect 465522 17518 465722 17562
rect 465737 17552 465761 17562
rect 465737 17528 465771 17552
rect 465782 17528 465854 17562
rect 465737 17518 465854 17528
rect 465509 17494 465854 17518
rect 465522 17450 465722 17494
rect 465737 17484 465761 17494
rect 465737 17460 465771 17484
rect 465782 17460 465854 17494
rect 465737 17450 465854 17460
rect 465509 17426 465854 17450
rect 465522 17382 465722 17426
rect 465737 17416 465761 17426
rect 465737 17392 465771 17416
rect 465782 17392 465854 17426
rect 465737 17382 465854 17392
rect 465509 17358 465854 17382
rect 465522 17314 465722 17358
rect 465737 17348 465761 17358
rect 465737 17324 465771 17348
rect 465782 17324 465854 17358
rect 465737 17314 465854 17324
rect 465509 17290 465854 17314
rect 465522 17278 465722 17290
rect 465533 17266 465557 17278
rect 465737 17266 465761 17290
rect 465782 17278 465854 17290
rect 466084 17278 466140 18278
rect 466156 17278 466212 18278
rect 466514 18198 466714 18278
rect 466729 18208 466763 18232
rect 466774 18208 466846 18278
rect 466729 18198 466846 18208
rect 466501 18174 466846 18198
rect 466514 18130 466714 18174
rect 466729 18164 466753 18174
rect 466729 18140 466763 18164
rect 466774 18140 466846 18174
rect 466729 18130 466846 18140
rect 466501 18106 466846 18130
rect 466514 18062 466714 18106
rect 466729 18096 466753 18106
rect 466729 18072 466763 18096
rect 466774 18072 466846 18106
rect 466729 18062 466846 18072
rect 466501 18038 466846 18062
rect 466514 17994 466714 18038
rect 466729 18028 466753 18038
rect 466729 18004 466763 18028
rect 466774 18004 466846 18038
rect 466729 17994 466846 18004
rect 466501 17970 466846 17994
rect 466514 17926 466714 17970
rect 466729 17960 466753 17970
rect 466729 17936 466763 17960
rect 466774 17936 466846 17970
rect 466729 17926 466846 17936
rect 466501 17902 466846 17926
rect 466514 17858 466714 17902
rect 466729 17892 466753 17902
rect 466729 17868 466763 17892
rect 466774 17868 466846 17902
rect 466729 17858 466846 17868
rect 466501 17834 466846 17858
rect 466514 17790 466714 17834
rect 466729 17824 466753 17834
rect 466729 17800 466763 17824
rect 466774 17800 466846 17834
rect 466729 17790 466846 17800
rect 466501 17766 466846 17790
rect 466514 17722 466714 17766
rect 466729 17756 466753 17766
rect 466729 17732 466763 17756
rect 466774 17732 466846 17766
rect 466729 17722 466846 17732
rect 466501 17698 466846 17722
rect 466514 17654 466714 17698
rect 466729 17688 466753 17698
rect 466729 17664 466763 17688
rect 466774 17664 466846 17698
rect 466729 17654 466846 17664
rect 466501 17630 466846 17654
rect 466514 17586 466714 17630
rect 466729 17620 466753 17630
rect 466729 17596 466763 17620
rect 466774 17596 466846 17630
rect 466729 17586 466846 17596
rect 466501 17562 466846 17586
rect 466514 17518 466714 17562
rect 466729 17552 466753 17562
rect 466729 17528 466763 17552
rect 466774 17528 466846 17562
rect 466729 17518 466846 17528
rect 466501 17494 466846 17518
rect 466514 17450 466714 17494
rect 466729 17484 466753 17494
rect 466729 17460 466763 17484
rect 466774 17460 466846 17494
rect 466729 17450 466846 17460
rect 466501 17426 466846 17450
rect 466514 17382 466714 17426
rect 466729 17416 466753 17426
rect 466729 17392 466763 17416
rect 466774 17392 466846 17426
rect 466729 17382 466846 17392
rect 466501 17358 466846 17382
rect 466514 17314 466714 17358
rect 466729 17348 466753 17358
rect 466729 17324 466763 17348
rect 466774 17324 466846 17358
rect 466729 17314 466846 17324
rect 466501 17290 466846 17314
rect 466514 17278 466714 17290
rect 466525 17266 466549 17278
rect 466729 17266 466753 17290
rect 466774 17278 466846 17290
rect 467076 17278 467132 18278
rect 467148 17278 467204 18278
rect 467506 18198 467706 18278
rect 467721 18208 467755 18232
rect 467766 18208 467838 18278
rect 467721 18198 467838 18208
rect 467493 18174 467838 18198
rect 467506 18130 467706 18174
rect 467721 18164 467745 18174
rect 467721 18140 467755 18164
rect 467766 18140 467838 18174
rect 467721 18130 467838 18140
rect 467493 18106 467838 18130
rect 467506 18062 467706 18106
rect 467721 18096 467745 18106
rect 467721 18072 467755 18096
rect 467766 18072 467838 18106
rect 467721 18062 467838 18072
rect 467493 18038 467838 18062
rect 467506 17994 467706 18038
rect 467721 18028 467745 18038
rect 467721 18004 467755 18028
rect 467766 18004 467838 18038
rect 467721 17994 467838 18004
rect 467493 17970 467838 17994
rect 467506 17926 467706 17970
rect 467721 17960 467745 17970
rect 467721 17936 467755 17960
rect 467766 17936 467838 17970
rect 467721 17926 467838 17936
rect 467493 17902 467838 17926
rect 467506 17858 467706 17902
rect 467721 17892 467745 17902
rect 467721 17868 467755 17892
rect 467766 17868 467838 17902
rect 467721 17858 467838 17868
rect 467493 17834 467838 17858
rect 467506 17790 467706 17834
rect 467721 17824 467745 17834
rect 467721 17800 467755 17824
rect 467766 17800 467838 17834
rect 467721 17790 467838 17800
rect 467493 17766 467838 17790
rect 467506 17722 467706 17766
rect 467721 17756 467745 17766
rect 467721 17732 467755 17756
rect 467766 17732 467838 17766
rect 467721 17722 467838 17732
rect 467493 17698 467838 17722
rect 467506 17654 467706 17698
rect 467721 17688 467745 17698
rect 467721 17664 467755 17688
rect 467766 17664 467838 17698
rect 467721 17654 467838 17664
rect 467493 17630 467838 17654
rect 467506 17586 467706 17630
rect 467721 17620 467745 17630
rect 467721 17596 467755 17620
rect 467766 17596 467838 17630
rect 467721 17586 467838 17596
rect 467493 17562 467838 17586
rect 467506 17518 467706 17562
rect 467721 17552 467745 17562
rect 467721 17528 467755 17552
rect 467766 17528 467838 17562
rect 467721 17518 467838 17528
rect 467493 17494 467838 17518
rect 467506 17450 467706 17494
rect 467721 17484 467745 17494
rect 467721 17460 467755 17484
rect 467766 17460 467838 17494
rect 467721 17450 467838 17460
rect 467493 17426 467838 17450
rect 467506 17382 467706 17426
rect 467721 17416 467745 17426
rect 467721 17392 467755 17416
rect 467766 17392 467838 17426
rect 467721 17382 467838 17392
rect 467493 17358 467838 17382
rect 467506 17314 467706 17358
rect 467721 17348 467745 17358
rect 467721 17324 467755 17348
rect 467766 17324 467838 17358
rect 467721 17314 467838 17324
rect 467493 17290 467838 17314
rect 467506 17278 467706 17290
rect 467517 17266 467541 17278
rect 467721 17266 467745 17290
rect 467766 17278 467838 17290
rect 468068 17278 468124 18278
rect 468140 17278 468196 18278
rect 468498 18198 468698 18278
rect 468713 18208 468747 18232
rect 468758 18208 468830 18278
rect 468713 18198 468830 18208
rect 468485 18174 468830 18198
rect 468498 18130 468698 18174
rect 468713 18164 468737 18174
rect 468713 18140 468747 18164
rect 468758 18140 468830 18174
rect 468713 18130 468830 18140
rect 468485 18106 468830 18130
rect 468498 18062 468698 18106
rect 468713 18096 468737 18106
rect 468713 18072 468747 18096
rect 468758 18072 468830 18106
rect 468713 18062 468830 18072
rect 468485 18038 468830 18062
rect 468498 17994 468698 18038
rect 468713 18028 468737 18038
rect 468713 18004 468747 18028
rect 468758 18004 468830 18038
rect 468713 17994 468830 18004
rect 468485 17970 468830 17994
rect 468498 17926 468698 17970
rect 468713 17960 468737 17970
rect 468713 17936 468747 17960
rect 468758 17936 468830 17970
rect 468713 17926 468830 17936
rect 468485 17902 468830 17926
rect 468498 17858 468698 17902
rect 468713 17892 468737 17902
rect 468713 17868 468747 17892
rect 468758 17868 468830 17902
rect 468713 17858 468830 17868
rect 468485 17834 468830 17858
rect 468498 17790 468698 17834
rect 468713 17824 468737 17834
rect 468713 17800 468747 17824
rect 468758 17800 468830 17834
rect 468713 17790 468830 17800
rect 468485 17766 468830 17790
rect 468498 17722 468698 17766
rect 468713 17756 468737 17766
rect 468713 17732 468747 17756
rect 468758 17732 468830 17766
rect 468713 17722 468830 17732
rect 468485 17698 468830 17722
rect 468498 17654 468698 17698
rect 468713 17688 468737 17698
rect 468713 17664 468747 17688
rect 468758 17664 468830 17698
rect 468713 17654 468830 17664
rect 468485 17630 468830 17654
rect 468498 17586 468698 17630
rect 468713 17620 468737 17630
rect 468713 17596 468747 17620
rect 468758 17596 468830 17630
rect 468713 17586 468830 17596
rect 468485 17562 468830 17586
rect 468498 17518 468698 17562
rect 468713 17552 468737 17562
rect 468713 17528 468747 17552
rect 468758 17528 468830 17562
rect 468713 17518 468830 17528
rect 468485 17494 468830 17518
rect 468498 17450 468698 17494
rect 468713 17484 468737 17494
rect 468713 17460 468747 17484
rect 468758 17460 468830 17494
rect 468713 17450 468830 17460
rect 468485 17426 468830 17450
rect 468498 17382 468698 17426
rect 468713 17416 468737 17426
rect 468713 17392 468747 17416
rect 468758 17392 468830 17426
rect 468713 17382 468830 17392
rect 468485 17358 468830 17382
rect 468498 17314 468698 17358
rect 468713 17348 468737 17358
rect 468713 17324 468747 17348
rect 468758 17324 468830 17358
rect 468713 17314 468830 17324
rect 468485 17290 468830 17314
rect 468498 17278 468698 17290
rect 468509 17266 468533 17278
rect 468713 17266 468737 17290
rect 468758 17278 468830 17290
rect 469060 17278 469116 18278
rect 469132 17278 469188 18278
rect 469490 18198 469690 18278
rect 469705 18208 469739 18232
rect 469750 18208 469822 18278
rect 469705 18198 469822 18208
rect 469477 18174 469822 18198
rect 469490 18130 469690 18174
rect 469705 18164 469729 18174
rect 469705 18140 469739 18164
rect 469750 18140 469822 18174
rect 469705 18130 469822 18140
rect 469477 18106 469822 18130
rect 469490 18062 469690 18106
rect 469705 18096 469729 18106
rect 469705 18072 469739 18096
rect 469750 18072 469822 18106
rect 469705 18062 469822 18072
rect 469477 18038 469822 18062
rect 469490 17994 469690 18038
rect 469705 18028 469729 18038
rect 469705 18004 469739 18028
rect 469750 18004 469822 18038
rect 469705 17994 469822 18004
rect 469477 17970 469822 17994
rect 469490 17926 469690 17970
rect 469705 17960 469729 17970
rect 469705 17936 469739 17960
rect 469750 17936 469822 17970
rect 469705 17926 469822 17936
rect 469477 17902 469822 17926
rect 469490 17858 469690 17902
rect 469705 17892 469729 17902
rect 469705 17868 469739 17892
rect 469750 17868 469822 17902
rect 469705 17858 469822 17868
rect 469477 17834 469822 17858
rect 469490 17790 469690 17834
rect 469705 17824 469729 17834
rect 469705 17800 469739 17824
rect 469750 17800 469822 17834
rect 469705 17790 469822 17800
rect 469477 17766 469822 17790
rect 469490 17722 469690 17766
rect 469705 17756 469729 17766
rect 469705 17732 469739 17756
rect 469750 17732 469822 17766
rect 469705 17722 469822 17732
rect 469477 17698 469822 17722
rect 469490 17654 469690 17698
rect 469705 17688 469729 17698
rect 469705 17664 469739 17688
rect 469750 17664 469822 17698
rect 469705 17654 469822 17664
rect 469477 17630 469822 17654
rect 469490 17586 469690 17630
rect 469705 17620 469729 17630
rect 469705 17596 469739 17620
rect 469750 17596 469822 17630
rect 469705 17586 469822 17596
rect 469477 17562 469822 17586
rect 469490 17518 469690 17562
rect 469705 17552 469729 17562
rect 469705 17528 469739 17552
rect 469750 17528 469822 17562
rect 469705 17518 469822 17528
rect 469477 17494 469822 17518
rect 469490 17450 469690 17494
rect 469705 17484 469729 17494
rect 469705 17460 469739 17484
rect 469750 17460 469822 17494
rect 469705 17450 469822 17460
rect 469477 17426 469822 17450
rect 469490 17382 469690 17426
rect 469705 17416 469729 17426
rect 469705 17392 469739 17416
rect 469750 17392 469822 17426
rect 469705 17382 469822 17392
rect 469477 17358 469822 17382
rect 469490 17314 469690 17358
rect 469705 17348 469729 17358
rect 469705 17324 469739 17348
rect 469750 17324 469822 17358
rect 469705 17314 469822 17324
rect 469477 17290 469822 17314
rect 469490 17278 469690 17290
rect 469501 17266 469525 17278
rect 469705 17266 469729 17290
rect 469750 17278 469822 17290
rect 470052 17278 470108 18278
rect 470124 17278 470180 18278
rect 470482 18198 470682 18278
rect 470697 18208 470731 18232
rect 470742 18208 470814 18278
rect 470697 18198 470814 18208
rect 470469 18174 470814 18198
rect 470482 18130 470682 18174
rect 470697 18164 470721 18174
rect 470697 18140 470731 18164
rect 470742 18140 470814 18174
rect 470697 18130 470814 18140
rect 470469 18106 470814 18130
rect 470482 18062 470682 18106
rect 470697 18096 470721 18106
rect 470697 18072 470731 18096
rect 470742 18072 470814 18106
rect 470697 18062 470814 18072
rect 470469 18038 470814 18062
rect 470482 17994 470682 18038
rect 470697 18028 470721 18038
rect 470697 18004 470731 18028
rect 470742 18004 470814 18038
rect 470697 17994 470814 18004
rect 470469 17970 470814 17994
rect 470482 17926 470682 17970
rect 470697 17960 470721 17970
rect 470697 17936 470731 17960
rect 470742 17936 470814 17970
rect 470697 17926 470814 17936
rect 470469 17902 470814 17926
rect 470482 17858 470682 17902
rect 470697 17892 470721 17902
rect 470697 17868 470731 17892
rect 470742 17868 470814 17902
rect 470697 17858 470814 17868
rect 470469 17834 470814 17858
rect 470482 17790 470682 17834
rect 470697 17824 470721 17834
rect 470697 17800 470731 17824
rect 470742 17800 470814 17834
rect 470697 17790 470814 17800
rect 470469 17766 470814 17790
rect 470482 17722 470682 17766
rect 470697 17756 470721 17766
rect 470697 17732 470731 17756
rect 470742 17732 470814 17766
rect 470697 17722 470814 17732
rect 470469 17698 470814 17722
rect 470482 17654 470682 17698
rect 470697 17688 470721 17698
rect 470697 17664 470731 17688
rect 470742 17664 470814 17698
rect 470697 17654 470814 17664
rect 470469 17630 470814 17654
rect 470482 17586 470682 17630
rect 470697 17620 470721 17630
rect 470697 17596 470731 17620
rect 470742 17596 470814 17630
rect 470697 17586 470814 17596
rect 470469 17562 470814 17586
rect 470482 17518 470682 17562
rect 470697 17552 470721 17562
rect 470697 17528 470731 17552
rect 470742 17528 470814 17562
rect 470697 17518 470814 17528
rect 470469 17494 470814 17518
rect 470482 17450 470682 17494
rect 470697 17484 470721 17494
rect 470697 17460 470731 17484
rect 470742 17460 470814 17494
rect 470697 17450 470814 17460
rect 470469 17426 470814 17450
rect 470482 17382 470682 17426
rect 470697 17416 470721 17426
rect 470697 17392 470731 17416
rect 470742 17392 470814 17426
rect 470697 17382 470814 17392
rect 470469 17358 470814 17382
rect 470482 17314 470682 17358
rect 470697 17348 470721 17358
rect 470697 17324 470731 17348
rect 470742 17324 470814 17358
rect 470697 17314 470814 17324
rect 470469 17290 470814 17314
rect 470482 17278 470682 17290
rect 470493 17266 470517 17278
rect 470697 17266 470721 17290
rect 470742 17278 470814 17290
rect 471044 17278 471100 18278
rect 471116 17278 471172 18278
rect 471474 18198 471674 18278
rect 471689 18208 471723 18232
rect 471734 18208 471806 18278
rect 471689 18198 471806 18208
rect 471461 18174 471806 18198
rect 471474 18130 471674 18174
rect 471689 18164 471713 18174
rect 471689 18140 471723 18164
rect 471734 18140 471806 18174
rect 471689 18130 471806 18140
rect 471461 18106 471806 18130
rect 471474 18062 471674 18106
rect 471689 18096 471713 18106
rect 471689 18072 471723 18096
rect 471734 18072 471806 18106
rect 471689 18062 471806 18072
rect 471461 18038 471806 18062
rect 471474 17994 471674 18038
rect 471689 18028 471713 18038
rect 471689 18004 471723 18028
rect 471734 18004 471806 18038
rect 471689 17994 471806 18004
rect 471461 17970 471806 17994
rect 471474 17926 471674 17970
rect 471689 17960 471713 17970
rect 471689 17936 471723 17960
rect 471734 17936 471806 17970
rect 471689 17926 471806 17936
rect 471461 17902 471806 17926
rect 471474 17858 471674 17902
rect 471689 17892 471713 17902
rect 471689 17868 471723 17892
rect 471734 17868 471806 17902
rect 471689 17858 471806 17868
rect 471461 17834 471806 17858
rect 471474 17790 471674 17834
rect 471689 17824 471713 17834
rect 471689 17800 471723 17824
rect 471734 17800 471806 17834
rect 471689 17790 471806 17800
rect 471461 17766 471806 17790
rect 471474 17722 471674 17766
rect 471689 17756 471713 17766
rect 471689 17732 471723 17756
rect 471734 17732 471806 17766
rect 471689 17722 471806 17732
rect 471461 17698 471806 17722
rect 471474 17654 471674 17698
rect 471689 17688 471713 17698
rect 471689 17664 471723 17688
rect 471734 17664 471806 17698
rect 471689 17654 471806 17664
rect 471461 17630 471806 17654
rect 471474 17586 471674 17630
rect 471689 17620 471713 17630
rect 471689 17596 471723 17620
rect 471734 17596 471806 17630
rect 471689 17586 471806 17596
rect 471461 17562 471806 17586
rect 471474 17518 471674 17562
rect 471689 17552 471713 17562
rect 471689 17528 471723 17552
rect 471734 17528 471806 17562
rect 471689 17518 471806 17528
rect 471461 17494 471806 17518
rect 471474 17450 471674 17494
rect 471689 17484 471713 17494
rect 471689 17460 471723 17484
rect 471734 17460 471806 17494
rect 471689 17450 471806 17460
rect 471461 17426 471806 17450
rect 471474 17382 471674 17426
rect 471689 17416 471713 17426
rect 471689 17392 471723 17416
rect 471734 17392 471806 17426
rect 471689 17382 471806 17392
rect 471461 17358 471806 17382
rect 471474 17314 471674 17358
rect 471689 17348 471713 17358
rect 471689 17324 471723 17348
rect 471734 17324 471806 17358
rect 471689 17314 471806 17324
rect 471461 17290 471806 17314
rect 471474 17278 471674 17290
rect 471485 17266 471509 17278
rect 471689 17266 471713 17290
rect 471734 17278 471806 17290
rect 472036 17278 472092 18278
rect 472108 17278 472164 18278
rect 472466 18198 472666 18278
rect 472681 18208 472715 18232
rect 472726 18208 472798 18278
rect 472681 18198 472798 18208
rect 472453 18174 472798 18198
rect 472466 18130 472666 18174
rect 472681 18164 472705 18174
rect 472681 18140 472715 18164
rect 472726 18140 472798 18174
rect 472681 18130 472798 18140
rect 472453 18106 472798 18130
rect 472466 18062 472666 18106
rect 472681 18096 472705 18106
rect 472681 18072 472715 18096
rect 472726 18072 472798 18106
rect 472681 18062 472798 18072
rect 472453 18038 472798 18062
rect 472466 17994 472666 18038
rect 472681 18028 472705 18038
rect 472681 18004 472715 18028
rect 472726 18004 472798 18038
rect 472681 17994 472798 18004
rect 472453 17970 472798 17994
rect 472466 17926 472666 17970
rect 472681 17960 472705 17970
rect 472681 17936 472715 17960
rect 472726 17936 472798 17970
rect 472681 17926 472798 17936
rect 472453 17902 472798 17926
rect 472466 17858 472666 17902
rect 472681 17892 472705 17902
rect 472681 17868 472715 17892
rect 472726 17868 472798 17902
rect 472681 17858 472798 17868
rect 472453 17834 472798 17858
rect 472466 17790 472666 17834
rect 472681 17824 472705 17834
rect 472681 17800 472715 17824
rect 472726 17800 472798 17834
rect 472681 17790 472798 17800
rect 472453 17766 472798 17790
rect 472466 17722 472666 17766
rect 472681 17756 472705 17766
rect 472681 17732 472715 17756
rect 472726 17732 472798 17766
rect 472681 17722 472798 17732
rect 472453 17698 472798 17722
rect 472466 17654 472666 17698
rect 472681 17688 472705 17698
rect 472681 17664 472715 17688
rect 472726 17664 472798 17698
rect 472681 17654 472798 17664
rect 472453 17630 472798 17654
rect 472466 17586 472666 17630
rect 472681 17620 472705 17630
rect 472681 17596 472715 17620
rect 472726 17596 472798 17630
rect 472681 17586 472798 17596
rect 472453 17562 472798 17586
rect 472466 17518 472666 17562
rect 472681 17552 472705 17562
rect 472681 17528 472715 17552
rect 472726 17528 472798 17562
rect 472681 17518 472798 17528
rect 472453 17494 472798 17518
rect 472466 17450 472666 17494
rect 472681 17484 472705 17494
rect 472681 17460 472715 17484
rect 472726 17460 472798 17494
rect 472681 17450 472798 17460
rect 472453 17426 472798 17450
rect 472466 17382 472666 17426
rect 472681 17416 472705 17426
rect 472681 17392 472715 17416
rect 472726 17392 472798 17426
rect 472681 17382 472798 17392
rect 472453 17358 472798 17382
rect 472466 17314 472666 17358
rect 472681 17348 472705 17358
rect 472681 17324 472715 17348
rect 472726 17324 472798 17358
rect 472681 17314 472798 17324
rect 472453 17290 472798 17314
rect 472466 17278 472666 17290
rect 472477 17266 472501 17278
rect 472681 17266 472705 17290
rect 472726 17278 472798 17290
rect 473028 17278 473084 18278
rect 473100 17278 473156 18278
rect 473458 18198 473658 18278
rect 473673 18208 473707 18232
rect 473718 18208 473790 18278
rect 473673 18198 473790 18208
rect 473445 18174 473790 18198
rect 473458 18130 473658 18174
rect 473673 18164 473697 18174
rect 473673 18140 473707 18164
rect 473718 18140 473790 18174
rect 473673 18130 473790 18140
rect 473445 18106 473790 18130
rect 473458 18062 473658 18106
rect 473673 18096 473697 18106
rect 473673 18072 473707 18096
rect 473718 18072 473790 18106
rect 473673 18062 473790 18072
rect 473445 18038 473790 18062
rect 473458 17994 473658 18038
rect 473673 18028 473697 18038
rect 473673 18004 473707 18028
rect 473718 18004 473790 18038
rect 473673 17994 473790 18004
rect 473445 17970 473790 17994
rect 473458 17926 473658 17970
rect 473673 17960 473697 17970
rect 473673 17936 473707 17960
rect 473718 17936 473790 17970
rect 473673 17926 473790 17936
rect 473445 17902 473790 17926
rect 473458 17858 473658 17902
rect 473673 17892 473697 17902
rect 473673 17868 473707 17892
rect 473718 17868 473790 17902
rect 473673 17858 473790 17868
rect 473445 17834 473790 17858
rect 473458 17790 473658 17834
rect 473673 17824 473697 17834
rect 473673 17800 473707 17824
rect 473718 17800 473790 17834
rect 473673 17790 473790 17800
rect 473445 17766 473790 17790
rect 473458 17722 473658 17766
rect 473673 17756 473697 17766
rect 473673 17732 473707 17756
rect 473718 17732 473790 17766
rect 473673 17722 473790 17732
rect 473445 17698 473790 17722
rect 473458 17654 473658 17698
rect 473673 17688 473697 17698
rect 473673 17664 473707 17688
rect 473718 17664 473790 17698
rect 473673 17654 473790 17664
rect 473445 17630 473790 17654
rect 473458 17586 473658 17630
rect 473673 17620 473697 17630
rect 473673 17596 473707 17620
rect 473718 17596 473790 17630
rect 473673 17586 473790 17596
rect 473445 17562 473790 17586
rect 473458 17518 473658 17562
rect 473673 17552 473697 17562
rect 473673 17528 473707 17552
rect 473718 17528 473790 17562
rect 473673 17518 473790 17528
rect 473445 17494 473790 17518
rect 473458 17450 473658 17494
rect 473673 17484 473697 17494
rect 473673 17460 473707 17484
rect 473718 17460 473790 17494
rect 473673 17450 473790 17460
rect 473445 17426 473790 17450
rect 473458 17382 473658 17426
rect 473673 17416 473697 17426
rect 473673 17392 473707 17416
rect 473718 17392 473790 17426
rect 473673 17382 473790 17392
rect 473445 17358 473790 17382
rect 473458 17314 473658 17358
rect 473673 17348 473697 17358
rect 473673 17324 473707 17348
rect 473718 17324 473790 17358
rect 473673 17314 473790 17324
rect 473445 17290 473790 17314
rect 473458 17278 473658 17290
rect 473469 17266 473493 17278
rect 473673 17266 473697 17290
rect 473718 17278 473790 17290
rect 474020 17278 474076 18278
rect 474092 17278 474148 18278
rect 474450 18198 474650 18278
rect 474665 18208 474699 18232
rect 474710 18208 474782 18278
rect 474665 18198 474782 18208
rect 474437 18174 474782 18198
rect 474450 18130 474650 18174
rect 474665 18164 474689 18174
rect 474665 18140 474699 18164
rect 474710 18140 474782 18174
rect 474665 18130 474782 18140
rect 474437 18106 474782 18130
rect 474450 18062 474650 18106
rect 474665 18096 474689 18106
rect 474665 18072 474699 18096
rect 474710 18072 474782 18106
rect 474665 18062 474782 18072
rect 474437 18038 474782 18062
rect 474450 17994 474650 18038
rect 474665 18028 474689 18038
rect 474665 18004 474699 18028
rect 474710 18004 474782 18038
rect 474665 17994 474782 18004
rect 474437 17970 474782 17994
rect 474450 17926 474650 17970
rect 474665 17960 474689 17970
rect 474665 17936 474699 17960
rect 474710 17936 474782 17970
rect 474665 17926 474782 17936
rect 474437 17902 474782 17926
rect 474450 17858 474650 17902
rect 474665 17892 474689 17902
rect 474665 17868 474699 17892
rect 474710 17868 474782 17902
rect 474665 17858 474782 17868
rect 474437 17834 474782 17858
rect 474450 17790 474650 17834
rect 474665 17824 474689 17834
rect 474665 17800 474699 17824
rect 474710 17800 474782 17834
rect 474665 17790 474782 17800
rect 474437 17766 474782 17790
rect 474450 17722 474650 17766
rect 474665 17756 474689 17766
rect 474665 17732 474699 17756
rect 474710 17732 474782 17766
rect 474665 17722 474782 17732
rect 474437 17698 474782 17722
rect 474450 17654 474650 17698
rect 474665 17688 474689 17698
rect 474665 17664 474699 17688
rect 474710 17664 474782 17698
rect 474665 17654 474782 17664
rect 474437 17630 474782 17654
rect 474450 17586 474650 17630
rect 474665 17620 474689 17630
rect 474665 17596 474699 17620
rect 474710 17596 474782 17630
rect 474665 17586 474782 17596
rect 474437 17562 474782 17586
rect 474450 17518 474650 17562
rect 474665 17552 474689 17562
rect 474665 17528 474699 17552
rect 474710 17528 474782 17562
rect 474665 17518 474782 17528
rect 474437 17494 474782 17518
rect 474450 17450 474650 17494
rect 474665 17484 474689 17494
rect 474665 17460 474699 17484
rect 474710 17460 474782 17494
rect 474665 17450 474782 17460
rect 474437 17426 474782 17450
rect 474450 17382 474650 17426
rect 474665 17416 474689 17426
rect 474665 17392 474699 17416
rect 474710 17392 474782 17426
rect 474665 17382 474782 17392
rect 474437 17358 474782 17382
rect 474450 17314 474650 17358
rect 474665 17348 474689 17358
rect 474665 17324 474699 17348
rect 474710 17324 474782 17358
rect 474665 17314 474782 17324
rect 474437 17290 474782 17314
rect 474450 17278 474650 17290
rect 474461 17266 474485 17278
rect 474665 17266 474689 17290
rect 474710 17278 474782 17290
rect 475012 17278 475068 18278
rect 475084 17278 475140 18278
rect 475442 18198 475642 18278
rect 475657 18208 475691 18232
rect 475702 18208 475774 18278
rect 475657 18198 475774 18208
rect 475429 18174 475774 18198
rect 475442 18130 475642 18174
rect 475657 18164 475681 18174
rect 475657 18140 475691 18164
rect 475702 18140 475774 18174
rect 475657 18130 475774 18140
rect 475429 18106 475774 18130
rect 475442 18062 475642 18106
rect 475657 18096 475681 18106
rect 475657 18072 475691 18096
rect 475702 18072 475774 18106
rect 475657 18062 475774 18072
rect 475429 18038 475774 18062
rect 475442 17994 475642 18038
rect 475657 18028 475681 18038
rect 475657 18004 475691 18028
rect 475702 18004 475774 18038
rect 475657 17994 475774 18004
rect 475429 17970 475774 17994
rect 475442 17926 475642 17970
rect 475657 17960 475681 17970
rect 475657 17936 475691 17960
rect 475702 17936 475774 17970
rect 475657 17926 475774 17936
rect 475429 17902 475774 17926
rect 475442 17858 475642 17902
rect 475657 17892 475681 17902
rect 475657 17868 475691 17892
rect 475702 17868 475774 17902
rect 475657 17858 475774 17868
rect 475429 17834 475774 17858
rect 475442 17790 475642 17834
rect 475657 17824 475681 17834
rect 475657 17800 475691 17824
rect 475702 17800 475774 17834
rect 475657 17790 475774 17800
rect 475429 17766 475774 17790
rect 475442 17722 475642 17766
rect 475657 17756 475681 17766
rect 475657 17732 475691 17756
rect 475702 17732 475774 17766
rect 475657 17722 475774 17732
rect 475429 17698 475774 17722
rect 475442 17654 475642 17698
rect 475657 17688 475681 17698
rect 475657 17664 475691 17688
rect 475702 17664 475774 17698
rect 475657 17654 475774 17664
rect 475429 17630 475774 17654
rect 475442 17586 475642 17630
rect 475657 17620 475681 17630
rect 475657 17596 475691 17620
rect 475702 17596 475774 17630
rect 475657 17586 475774 17596
rect 475429 17562 475774 17586
rect 475442 17518 475642 17562
rect 475657 17552 475681 17562
rect 475657 17528 475691 17552
rect 475702 17528 475774 17562
rect 475657 17518 475774 17528
rect 475429 17494 475774 17518
rect 475442 17450 475642 17494
rect 475657 17484 475681 17494
rect 475657 17460 475691 17484
rect 475702 17460 475774 17494
rect 475657 17450 475774 17460
rect 475429 17426 475774 17450
rect 475442 17382 475642 17426
rect 475657 17416 475681 17426
rect 475657 17392 475691 17416
rect 475702 17392 475774 17426
rect 475657 17382 475774 17392
rect 475429 17358 475774 17382
rect 475442 17314 475642 17358
rect 475657 17348 475681 17358
rect 475657 17324 475691 17348
rect 475702 17324 475774 17358
rect 475657 17314 475774 17324
rect 475429 17290 475774 17314
rect 475442 17278 475642 17290
rect 475453 17266 475477 17278
rect 475657 17266 475681 17290
rect 475702 17278 475774 17290
rect 476004 17278 476060 18278
rect 476076 17278 476132 18278
rect 476434 18198 476634 18278
rect 476649 18208 476683 18232
rect 476694 18208 476766 18278
rect 476649 18198 476766 18208
rect 476421 18174 476766 18198
rect 476434 18130 476634 18174
rect 476649 18164 476673 18174
rect 476649 18140 476683 18164
rect 476694 18140 476766 18174
rect 476649 18130 476766 18140
rect 476421 18106 476766 18130
rect 476434 18062 476634 18106
rect 476649 18096 476673 18106
rect 476649 18072 476683 18096
rect 476694 18072 476766 18106
rect 476649 18062 476766 18072
rect 476421 18038 476766 18062
rect 476434 17994 476634 18038
rect 476649 18028 476673 18038
rect 476649 18004 476683 18028
rect 476694 18004 476766 18038
rect 476649 17994 476766 18004
rect 476421 17970 476766 17994
rect 476434 17926 476634 17970
rect 476649 17960 476673 17970
rect 476649 17936 476683 17960
rect 476694 17936 476766 17970
rect 476649 17926 476766 17936
rect 476421 17902 476766 17926
rect 476434 17858 476634 17902
rect 476649 17892 476673 17902
rect 476649 17868 476683 17892
rect 476694 17868 476766 17902
rect 476649 17858 476766 17868
rect 476421 17834 476766 17858
rect 476434 17790 476634 17834
rect 476649 17824 476673 17834
rect 476649 17800 476683 17824
rect 476694 17800 476766 17834
rect 476649 17790 476766 17800
rect 476421 17766 476766 17790
rect 476434 17722 476634 17766
rect 476649 17756 476673 17766
rect 476649 17732 476683 17756
rect 476694 17732 476766 17766
rect 476649 17722 476766 17732
rect 476421 17698 476766 17722
rect 476434 17654 476634 17698
rect 476649 17688 476673 17698
rect 476649 17664 476683 17688
rect 476694 17664 476766 17698
rect 476649 17654 476766 17664
rect 476421 17630 476766 17654
rect 476434 17586 476634 17630
rect 476649 17620 476673 17630
rect 476649 17596 476683 17620
rect 476694 17596 476766 17630
rect 476649 17586 476766 17596
rect 476421 17562 476766 17586
rect 476434 17518 476634 17562
rect 476649 17552 476673 17562
rect 476649 17528 476683 17552
rect 476694 17528 476766 17562
rect 476649 17518 476766 17528
rect 476421 17494 476766 17518
rect 476434 17450 476634 17494
rect 476649 17484 476673 17494
rect 476649 17460 476683 17484
rect 476694 17460 476766 17494
rect 476649 17450 476766 17460
rect 476421 17426 476766 17450
rect 476434 17382 476634 17426
rect 476649 17416 476673 17426
rect 476649 17392 476683 17416
rect 476694 17392 476766 17426
rect 476649 17382 476766 17392
rect 476421 17358 476766 17382
rect 476434 17314 476634 17358
rect 476649 17348 476673 17358
rect 476649 17324 476683 17348
rect 476694 17324 476766 17358
rect 476649 17314 476766 17324
rect 476421 17290 476766 17314
rect 476434 17278 476634 17290
rect 476445 17266 476469 17278
rect 476649 17266 476673 17290
rect 476694 17278 476766 17290
rect 476996 17278 477052 18278
rect 477068 17278 477124 18278
rect 477426 18198 477626 18278
rect 477641 18208 477675 18232
rect 477686 18208 477758 18278
rect 477641 18198 477758 18208
rect 477413 18174 477758 18198
rect 477426 18130 477626 18174
rect 477641 18164 477665 18174
rect 477641 18140 477675 18164
rect 477686 18140 477758 18174
rect 477641 18130 477758 18140
rect 477413 18106 477758 18130
rect 477426 18062 477626 18106
rect 477641 18096 477665 18106
rect 477641 18072 477675 18096
rect 477686 18072 477758 18106
rect 477641 18062 477758 18072
rect 477413 18038 477758 18062
rect 477426 17994 477626 18038
rect 477641 18028 477665 18038
rect 477641 18004 477675 18028
rect 477686 18004 477758 18038
rect 477641 17994 477758 18004
rect 477413 17970 477758 17994
rect 477426 17926 477626 17970
rect 477641 17960 477665 17970
rect 477641 17936 477675 17960
rect 477686 17936 477758 17970
rect 477641 17926 477758 17936
rect 477413 17902 477758 17926
rect 477426 17858 477626 17902
rect 477641 17892 477665 17902
rect 477641 17868 477675 17892
rect 477686 17868 477758 17902
rect 477641 17858 477758 17868
rect 477413 17834 477758 17858
rect 477426 17790 477626 17834
rect 477641 17824 477665 17834
rect 477641 17800 477675 17824
rect 477686 17800 477758 17834
rect 477641 17790 477758 17800
rect 477413 17766 477758 17790
rect 477426 17722 477626 17766
rect 477641 17756 477665 17766
rect 477641 17732 477675 17756
rect 477686 17732 477758 17766
rect 477641 17722 477758 17732
rect 477413 17698 477758 17722
rect 477426 17654 477626 17698
rect 477641 17688 477665 17698
rect 477641 17664 477675 17688
rect 477686 17664 477758 17698
rect 477641 17654 477758 17664
rect 477413 17630 477758 17654
rect 477426 17586 477626 17630
rect 477641 17620 477665 17630
rect 477641 17596 477675 17620
rect 477686 17596 477758 17630
rect 477641 17586 477758 17596
rect 477413 17562 477758 17586
rect 477426 17518 477626 17562
rect 477641 17552 477665 17562
rect 477641 17528 477675 17552
rect 477686 17528 477758 17562
rect 477641 17518 477758 17528
rect 477413 17494 477758 17518
rect 477426 17450 477626 17494
rect 477641 17484 477665 17494
rect 477641 17460 477675 17484
rect 477686 17460 477758 17494
rect 477641 17450 477758 17460
rect 477413 17426 477758 17450
rect 477426 17382 477626 17426
rect 477641 17416 477665 17426
rect 477641 17392 477675 17416
rect 477686 17392 477758 17426
rect 477641 17382 477758 17392
rect 477413 17358 477758 17382
rect 477426 17314 477626 17358
rect 477641 17348 477665 17358
rect 477641 17324 477675 17348
rect 477686 17324 477758 17358
rect 477641 17314 477758 17324
rect 477413 17290 477758 17314
rect 477426 17278 477626 17290
rect 477437 17266 477461 17278
rect 477641 17266 477665 17290
rect 477686 17278 477758 17290
rect 477988 17278 478044 18278
rect 478060 17278 478116 18278
rect 478327 17278 478377 18278
rect 465533 16678 465567 16690
rect 464746 15878 464780 15908
rect 464708 15840 464780 15870
rect 464903 15678 464936 16678
rect 465106 15678 465123 16678
rect 465261 15678 465333 16678
rect 465522 16656 465722 16678
rect 465737 16666 465771 16690
rect 466525 16678 466559 16690
rect 465782 16666 465854 16678
rect 465737 16656 465854 16666
rect 465509 16632 465854 16656
rect 465522 16588 465722 16632
rect 465737 16622 465761 16632
rect 465737 16598 465771 16622
rect 465782 16598 465854 16632
rect 465737 16588 465854 16598
rect 465509 16564 465854 16588
rect 465522 16520 465722 16564
rect 465737 16554 465761 16564
rect 465737 16530 465771 16554
rect 465782 16530 465854 16564
rect 465737 16520 465854 16530
rect 465509 16496 465854 16520
rect 465522 16452 465722 16496
rect 465737 16486 465761 16496
rect 465737 16462 465771 16486
rect 465782 16462 465854 16496
rect 465737 16452 465854 16462
rect 465509 16428 465854 16452
rect 465522 16384 465722 16428
rect 465737 16418 465761 16428
rect 465737 16394 465771 16418
rect 465782 16394 465854 16428
rect 465737 16384 465854 16394
rect 465509 16360 465854 16384
rect 465522 16316 465722 16360
rect 465737 16350 465761 16360
rect 465737 16326 465771 16350
rect 465782 16326 465854 16360
rect 465737 16316 465854 16326
rect 465509 16292 465854 16316
rect 465522 16248 465722 16292
rect 465737 16282 465761 16292
rect 465737 16258 465771 16282
rect 465782 16258 465854 16292
rect 465737 16248 465854 16258
rect 465509 16224 465854 16248
rect 465522 16180 465722 16224
rect 465737 16214 465761 16224
rect 465737 16190 465771 16214
rect 465782 16190 465854 16224
rect 465737 16180 465854 16190
rect 465509 16156 465854 16180
rect 465522 16112 465722 16156
rect 465737 16146 465761 16156
rect 465737 16122 465771 16146
rect 465782 16122 465854 16156
rect 465737 16112 465854 16122
rect 465509 16088 465854 16112
rect 465522 16044 465722 16088
rect 465737 16078 465761 16088
rect 465737 16054 465771 16078
rect 465782 16054 465854 16088
rect 465737 16044 465854 16054
rect 465509 16020 465854 16044
rect 465522 15976 465722 16020
rect 465737 16010 465761 16020
rect 465737 15986 465771 16010
rect 465782 15986 465854 16020
rect 465737 15976 465854 15986
rect 465509 15952 465854 15976
rect 465522 15908 465722 15952
rect 465737 15942 465761 15952
rect 465737 15918 465771 15942
rect 465782 15918 465854 15952
rect 465737 15908 465854 15918
rect 465509 15884 465854 15908
rect 465522 15840 465722 15884
rect 465737 15874 465761 15884
rect 465737 15850 465771 15874
rect 465782 15850 465854 15884
rect 465737 15840 465854 15850
rect 465509 15816 465854 15840
rect 465522 15772 465722 15816
rect 465737 15806 465761 15816
rect 465737 15782 465771 15806
rect 465782 15782 465854 15816
rect 465737 15772 465854 15782
rect 465509 15748 465854 15772
rect 465522 15678 465722 15748
rect 465737 15724 465761 15748
rect 465782 15678 465854 15748
rect 466084 15678 466140 16678
rect 466156 15678 466212 16678
rect 466514 16656 466714 16678
rect 466729 16666 466763 16690
rect 467517 16678 467551 16690
rect 466774 16666 466846 16678
rect 466729 16656 466846 16666
rect 466501 16632 466846 16656
rect 466514 16588 466714 16632
rect 466729 16622 466753 16632
rect 466729 16598 466763 16622
rect 466774 16598 466846 16632
rect 466729 16588 466846 16598
rect 466501 16564 466846 16588
rect 466514 16520 466714 16564
rect 466729 16554 466753 16564
rect 466729 16530 466763 16554
rect 466774 16530 466846 16564
rect 466729 16520 466846 16530
rect 466501 16496 466846 16520
rect 466514 16452 466714 16496
rect 466729 16486 466753 16496
rect 466729 16462 466763 16486
rect 466774 16462 466846 16496
rect 466729 16452 466846 16462
rect 466501 16428 466846 16452
rect 466514 16384 466714 16428
rect 466729 16418 466753 16428
rect 466729 16394 466763 16418
rect 466774 16394 466846 16428
rect 466729 16384 466846 16394
rect 466501 16360 466846 16384
rect 466514 16316 466714 16360
rect 466729 16350 466753 16360
rect 466729 16326 466763 16350
rect 466774 16326 466846 16360
rect 466729 16316 466846 16326
rect 466501 16292 466846 16316
rect 466514 16248 466714 16292
rect 466729 16282 466753 16292
rect 466729 16258 466763 16282
rect 466774 16258 466846 16292
rect 466729 16248 466846 16258
rect 466501 16224 466846 16248
rect 466514 16180 466714 16224
rect 466729 16214 466753 16224
rect 466729 16190 466763 16214
rect 466774 16190 466846 16224
rect 466729 16180 466846 16190
rect 466501 16156 466846 16180
rect 466514 16112 466714 16156
rect 466729 16146 466753 16156
rect 466729 16122 466763 16146
rect 466774 16122 466846 16156
rect 466729 16112 466846 16122
rect 466501 16088 466846 16112
rect 466514 16044 466714 16088
rect 466729 16078 466753 16088
rect 466729 16054 466763 16078
rect 466774 16054 466846 16088
rect 466729 16044 466846 16054
rect 466501 16020 466846 16044
rect 466514 15976 466714 16020
rect 466729 16010 466753 16020
rect 466729 15986 466763 16010
rect 466774 15986 466846 16020
rect 466729 15976 466846 15986
rect 466501 15952 466846 15976
rect 466514 15908 466714 15952
rect 466729 15942 466753 15952
rect 466729 15918 466763 15942
rect 466774 15918 466846 15952
rect 466729 15908 466846 15918
rect 466501 15884 466846 15908
rect 466514 15840 466714 15884
rect 466729 15874 466753 15884
rect 466729 15850 466763 15874
rect 466774 15850 466846 15884
rect 466729 15840 466846 15850
rect 466501 15816 466846 15840
rect 466514 15772 466714 15816
rect 466729 15806 466753 15816
rect 466729 15782 466763 15806
rect 466774 15782 466846 15816
rect 466729 15772 466846 15782
rect 466501 15748 466846 15772
rect 466514 15678 466714 15748
rect 466729 15724 466753 15748
rect 466774 15678 466846 15748
rect 467076 15678 467132 16678
rect 467148 15678 467204 16678
rect 467506 16656 467706 16678
rect 467721 16666 467755 16690
rect 468509 16678 468543 16690
rect 467766 16666 467838 16678
rect 467721 16656 467838 16666
rect 467493 16632 467838 16656
rect 467506 16588 467706 16632
rect 467721 16622 467745 16632
rect 467721 16598 467755 16622
rect 467766 16598 467838 16632
rect 467721 16588 467838 16598
rect 467493 16564 467838 16588
rect 467506 16520 467706 16564
rect 467721 16554 467745 16564
rect 467721 16530 467755 16554
rect 467766 16530 467838 16564
rect 467721 16520 467838 16530
rect 467493 16496 467838 16520
rect 467506 16452 467706 16496
rect 467721 16486 467745 16496
rect 467721 16462 467755 16486
rect 467766 16462 467838 16496
rect 467721 16452 467838 16462
rect 467493 16428 467838 16452
rect 467506 16384 467706 16428
rect 467721 16418 467745 16428
rect 467721 16394 467755 16418
rect 467766 16394 467838 16428
rect 467721 16384 467838 16394
rect 467493 16360 467838 16384
rect 467506 16316 467706 16360
rect 467721 16350 467745 16360
rect 467721 16326 467755 16350
rect 467766 16326 467838 16360
rect 467721 16316 467838 16326
rect 467493 16292 467838 16316
rect 467506 16248 467706 16292
rect 467721 16282 467745 16292
rect 467721 16258 467755 16282
rect 467766 16258 467838 16292
rect 467721 16248 467838 16258
rect 467493 16224 467838 16248
rect 467506 16180 467706 16224
rect 467721 16214 467745 16224
rect 467721 16190 467755 16214
rect 467766 16190 467838 16224
rect 467721 16180 467838 16190
rect 467493 16156 467838 16180
rect 467506 16112 467706 16156
rect 467721 16146 467745 16156
rect 467721 16122 467755 16146
rect 467766 16122 467838 16156
rect 467721 16112 467838 16122
rect 467493 16088 467838 16112
rect 467506 16044 467706 16088
rect 467721 16078 467745 16088
rect 467721 16054 467755 16078
rect 467766 16054 467838 16088
rect 467721 16044 467838 16054
rect 467493 16020 467838 16044
rect 467506 15976 467706 16020
rect 467721 16010 467745 16020
rect 467721 15986 467755 16010
rect 467766 15986 467838 16020
rect 467721 15976 467838 15986
rect 467493 15952 467838 15976
rect 467506 15908 467706 15952
rect 467721 15942 467745 15952
rect 467721 15918 467755 15942
rect 467766 15918 467838 15952
rect 467721 15908 467838 15918
rect 467493 15884 467838 15908
rect 467506 15840 467706 15884
rect 467721 15874 467745 15884
rect 467721 15850 467755 15874
rect 467766 15850 467838 15884
rect 467721 15840 467838 15850
rect 467493 15816 467838 15840
rect 467506 15772 467706 15816
rect 467721 15806 467745 15816
rect 467721 15782 467755 15806
rect 467766 15782 467838 15816
rect 467721 15772 467838 15782
rect 467493 15748 467838 15772
rect 467506 15678 467706 15748
rect 467721 15724 467745 15748
rect 467766 15678 467838 15748
rect 468068 15678 468124 16678
rect 468140 15678 468196 16678
rect 468498 16656 468698 16678
rect 468713 16666 468747 16690
rect 469501 16678 469535 16690
rect 468758 16666 468830 16678
rect 468713 16656 468830 16666
rect 468485 16632 468830 16656
rect 468498 16588 468698 16632
rect 468713 16622 468737 16632
rect 468713 16598 468747 16622
rect 468758 16598 468830 16632
rect 468713 16588 468830 16598
rect 468485 16564 468830 16588
rect 468498 16520 468698 16564
rect 468713 16554 468737 16564
rect 468713 16530 468747 16554
rect 468758 16530 468830 16564
rect 468713 16520 468830 16530
rect 468485 16496 468830 16520
rect 468498 16452 468698 16496
rect 468713 16486 468737 16496
rect 468713 16462 468747 16486
rect 468758 16462 468830 16496
rect 468713 16452 468830 16462
rect 468485 16428 468830 16452
rect 468498 16384 468698 16428
rect 468713 16418 468737 16428
rect 468713 16394 468747 16418
rect 468758 16394 468830 16428
rect 468713 16384 468830 16394
rect 468485 16360 468830 16384
rect 468498 16316 468698 16360
rect 468713 16350 468737 16360
rect 468713 16326 468747 16350
rect 468758 16326 468830 16360
rect 468713 16316 468830 16326
rect 468485 16292 468830 16316
rect 468498 16248 468698 16292
rect 468713 16282 468737 16292
rect 468713 16258 468747 16282
rect 468758 16258 468830 16292
rect 468713 16248 468830 16258
rect 468485 16224 468830 16248
rect 468498 16180 468698 16224
rect 468713 16214 468737 16224
rect 468713 16190 468747 16214
rect 468758 16190 468830 16224
rect 468713 16180 468830 16190
rect 468485 16156 468830 16180
rect 468498 16112 468698 16156
rect 468713 16146 468737 16156
rect 468713 16122 468747 16146
rect 468758 16122 468830 16156
rect 468713 16112 468830 16122
rect 468485 16088 468830 16112
rect 468498 16044 468698 16088
rect 468713 16078 468737 16088
rect 468713 16054 468747 16078
rect 468758 16054 468830 16088
rect 468713 16044 468830 16054
rect 468485 16020 468830 16044
rect 468498 15976 468698 16020
rect 468713 16010 468737 16020
rect 468713 15986 468747 16010
rect 468758 15986 468830 16020
rect 468713 15976 468830 15986
rect 468485 15952 468830 15976
rect 468498 15908 468698 15952
rect 468713 15942 468737 15952
rect 468713 15918 468747 15942
rect 468758 15918 468830 15952
rect 468713 15908 468830 15918
rect 468485 15884 468830 15908
rect 468498 15840 468698 15884
rect 468713 15874 468737 15884
rect 468713 15850 468747 15874
rect 468758 15850 468830 15884
rect 468713 15840 468830 15850
rect 468485 15816 468830 15840
rect 468498 15772 468698 15816
rect 468713 15806 468737 15816
rect 468713 15782 468747 15806
rect 468758 15782 468830 15816
rect 468713 15772 468830 15782
rect 468485 15748 468830 15772
rect 468498 15678 468698 15748
rect 468713 15724 468737 15748
rect 468758 15678 468830 15748
rect 469060 15678 469116 16678
rect 469132 15678 469188 16678
rect 469490 16656 469690 16678
rect 469705 16666 469739 16690
rect 470493 16678 470527 16690
rect 469750 16666 469822 16678
rect 469705 16656 469822 16666
rect 469477 16632 469822 16656
rect 469490 16588 469690 16632
rect 469705 16622 469729 16632
rect 469705 16598 469739 16622
rect 469750 16598 469822 16632
rect 469705 16588 469822 16598
rect 469477 16564 469822 16588
rect 469490 16520 469690 16564
rect 469705 16554 469729 16564
rect 469705 16530 469739 16554
rect 469750 16530 469822 16564
rect 469705 16520 469822 16530
rect 469477 16496 469822 16520
rect 469490 16452 469690 16496
rect 469705 16486 469729 16496
rect 469705 16462 469739 16486
rect 469750 16462 469822 16496
rect 469705 16452 469822 16462
rect 469477 16428 469822 16452
rect 469490 16384 469690 16428
rect 469705 16418 469729 16428
rect 469705 16394 469739 16418
rect 469750 16394 469822 16428
rect 469705 16384 469822 16394
rect 469477 16360 469822 16384
rect 469490 16316 469690 16360
rect 469705 16350 469729 16360
rect 469705 16326 469739 16350
rect 469750 16326 469822 16360
rect 469705 16316 469822 16326
rect 469477 16292 469822 16316
rect 469490 16248 469690 16292
rect 469705 16282 469729 16292
rect 469705 16258 469739 16282
rect 469750 16258 469822 16292
rect 469705 16248 469822 16258
rect 469477 16224 469822 16248
rect 469490 16180 469690 16224
rect 469705 16214 469729 16224
rect 469705 16190 469739 16214
rect 469750 16190 469822 16224
rect 469705 16180 469822 16190
rect 469477 16156 469822 16180
rect 469490 16112 469690 16156
rect 469705 16146 469729 16156
rect 469705 16122 469739 16146
rect 469750 16122 469822 16156
rect 469705 16112 469822 16122
rect 469477 16088 469822 16112
rect 469490 16044 469690 16088
rect 469705 16078 469729 16088
rect 469705 16054 469739 16078
rect 469750 16054 469822 16088
rect 469705 16044 469822 16054
rect 469477 16020 469822 16044
rect 469490 15976 469690 16020
rect 469705 16010 469729 16020
rect 469705 15986 469739 16010
rect 469750 15986 469822 16020
rect 469705 15976 469822 15986
rect 469477 15952 469822 15976
rect 469490 15908 469690 15952
rect 469705 15942 469729 15952
rect 469705 15918 469739 15942
rect 469750 15918 469822 15952
rect 469705 15908 469822 15918
rect 469477 15884 469822 15908
rect 469490 15840 469690 15884
rect 469705 15874 469729 15884
rect 469705 15850 469739 15874
rect 469750 15850 469822 15884
rect 469705 15840 469822 15850
rect 469477 15816 469822 15840
rect 469490 15772 469690 15816
rect 469705 15806 469729 15816
rect 469705 15782 469739 15806
rect 469750 15782 469822 15816
rect 469705 15772 469822 15782
rect 469477 15748 469822 15772
rect 469490 15678 469690 15748
rect 469705 15724 469729 15748
rect 469750 15678 469822 15748
rect 470052 15678 470108 16678
rect 470124 15678 470180 16678
rect 470482 16656 470682 16678
rect 470697 16666 470731 16690
rect 471485 16678 471519 16690
rect 470742 16666 470814 16678
rect 470697 16656 470814 16666
rect 470469 16632 470814 16656
rect 470482 16588 470682 16632
rect 470697 16622 470721 16632
rect 470697 16598 470731 16622
rect 470742 16598 470814 16632
rect 470697 16588 470814 16598
rect 470469 16564 470814 16588
rect 470482 16520 470682 16564
rect 470697 16554 470721 16564
rect 470697 16530 470731 16554
rect 470742 16530 470814 16564
rect 470697 16520 470814 16530
rect 470469 16496 470814 16520
rect 470482 16452 470682 16496
rect 470697 16486 470721 16496
rect 470697 16462 470731 16486
rect 470742 16462 470814 16496
rect 470697 16452 470814 16462
rect 470469 16428 470814 16452
rect 470482 16384 470682 16428
rect 470697 16418 470721 16428
rect 470697 16394 470731 16418
rect 470742 16394 470814 16428
rect 470697 16384 470814 16394
rect 470469 16360 470814 16384
rect 470482 16316 470682 16360
rect 470697 16350 470721 16360
rect 470697 16326 470731 16350
rect 470742 16326 470814 16360
rect 470697 16316 470814 16326
rect 470469 16292 470814 16316
rect 470482 16248 470682 16292
rect 470697 16282 470721 16292
rect 470697 16258 470731 16282
rect 470742 16258 470814 16292
rect 470697 16248 470814 16258
rect 470469 16224 470814 16248
rect 470482 16180 470682 16224
rect 470697 16214 470721 16224
rect 470697 16190 470731 16214
rect 470742 16190 470814 16224
rect 470697 16180 470814 16190
rect 470469 16156 470814 16180
rect 470482 16112 470682 16156
rect 470697 16146 470721 16156
rect 470697 16122 470731 16146
rect 470742 16122 470814 16156
rect 470697 16112 470814 16122
rect 470469 16088 470814 16112
rect 470482 16044 470682 16088
rect 470697 16078 470721 16088
rect 470697 16054 470731 16078
rect 470742 16054 470814 16088
rect 470697 16044 470814 16054
rect 470469 16020 470814 16044
rect 470482 15976 470682 16020
rect 470697 16010 470721 16020
rect 470697 15986 470731 16010
rect 470742 15986 470814 16020
rect 470697 15976 470814 15986
rect 470469 15952 470814 15976
rect 470482 15908 470682 15952
rect 470697 15942 470721 15952
rect 470697 15918 470731 15942
rect 470742 15918 470814 15952
rect 470697 15908 470814 15918
rect 470469 15884 470814 15908
rect 470482 15840 470682 15884
rect 470697 15874 470721 15884
rect 470697 15850 470731 15874
rect 470742 15850 470814 15884
rect 470697 15840 470814 15850
rect 470469 15816 470814 15840
rect 470482 15772 470682 15816
rect 470697 15806 470721 15816
rect 470697 15782 470731 15806
rect 470742 15782 470814 15816
rect 470697 15772 470814 15782
rect 470469 15748 470814 15772
rect 470482 15678 470682 15748
rect 470697 15724 470721 15748
rect 470742 15678 470814 15748
rect 471044 15678 471100 16678
rect 471116 15678 471172 16678
rect 471474 16656 471674 16678
rect 471689 16666 471723 16690
rect 472477 16678 472511 16690
rect 471734 16666 471806 16678
rect 471689 16656 471806 16666
rect 471461 16632 471806 16656
rect 471474 16588 471674 16632
rect 471689 16622 471713 16632
rect 471689 16598 471723 16622
rect 471734 16598 471806 16632
rect 471689 16588 471806 16598
rect 471461 16564 471806 16588
rect 471474 16520 471674 16564
rect 471689 16554 471713 16564
rect 471689 16530 471723 16554
rect 471734 16530 471806 16564
rect 471689 16520 471806 16530
rect 471461 16496 471806 16520
rect 471474 16452 471674 16496
rect 471689 16486 471713 16496
rect 471689 16462 471723 16486
rect 471734 16462 471806 16496
rect 471689 16452 471806 16462
rect 471461 16428 471806 16452
rect 471474 16384 471674 16428
rect 471689 16418 471713 16428
rect 471689 16394 471723 16418
rect 471734 16394 471806 16428
rect 471689 16384 471806 16394
rect 471461 16360 471806 16384
rect 471474 16316 471674 16360
rect 471689 16350 471713 16360
rect 471689 16326 471723 16350
rect 471734 16326 471806 16360
rect 471689 16316 471806 16326
rect 471461 16292 471806 16316
rect 471474 16248 471674 16292
rect 471689 16282 471713 16292
rect 471689 16258 471723 16282
rect 471734 16258 471806 16292
rect 471689 16248 471806 16258
rect 471461 16224 471806 16248
rect 471474 16180 471674 16224
rect 471689 16214 471713 16224
rect 471689 16190 471723 16214
rect 471734 16190 471806 16224
rect 471689 16180 471806 16190
rect 471461 16156 471806 16180
rect 471474 16112 471674 16156
rect 471689 16146 471713 16156
rect 471689 16122 471723 16146
rect 471734 16122 471806 16156
rect 471689 16112 471806 16122
rect 471461 16088 471806 16112
rect 471474 16044 471674 16088
rect 471689 16078 471713 16088
rect 471689 16054 471723 16078
rect 471734 16054 471806 16088
rect 471689 16044 471806 16054
rect 471461 16020 471806 16044
rect 471474 15976 471674 16020
rect 471689 16010 471713 16020
rect 471689 15986 471723 16010
rect 471734 15986 471806 16020
rect 471689 15976 471806 15986
rect 471461 15952 471806 15976
rect 471474 15908 471674 15952
rect 471689 15942 471713 15952
rect 471689 15918 471723 15942
rect 471734 15918 471806 15952
rect 471689 15908 471806 15918
rect 471461 15884 471806 15908
rect 471474 15840 471674 15884
rect 471689 15874 471713 15884
rect 471689 15850 471723 15874
rect 471734 15850 471806 15884
rect 471689 15840 471806 15850
rect 471461 15816 471806 15840
rect 471474 15772 471674 15816
rect 471689 15806 471713 15816
rect 471689 15782 471723 15806
rect 471734 15782 471806 15816
rect 471689 15772 471806 15782
rect 471461 15748 471806 15772
rect 471474 15678 471674 15748
rect 471689 15724 471713 15748
rect 471734 15678 471806 15748
rect 472036 15678 472092 16678
rect 472108 15678 472164 16678
rect 472466 16656 472666 16678
rect 472681 16666 472715 16690
rect 473469 16678 473503 16690
rect 472726 16666 472798 16678
rect 472681 16656 472798 16666
rect 472453 16632 472798 16656
rect 472466 16588 472666 16632
rect 472681 16622 472705 16632
rect 472681 16598 472715 16622
rect 472726 16598 472798 16632
rect 472681 16588 472798 16598
rect 472453 16564 472798 16588
rect 472466 16520 472666 16564
rect 472681 16554 472705 16564
rect 472681 16530 472715 16554
rect 472726 16530 472798 16564
rect 472681 16520 472798 16530
rect 472453 16496 472798 16520
rect 472466 16452 472666 16496
rect 472681 16486 472705 16496
rect 472681 16462 472715 16486
rect 472726 16462 472798 16496
rect 472681 16452 472798 16462
rect 472453 16428 472798 16452
rect 472466 16384 472666 16428
rect 472681 16418 472705 16428
rect 472681 16394 472715 16418
rect 472726 16394 472798 16428
rect 472681 16384 472798 16394
rect 472453 16360 472798 16384
rect 472466 16316 472666 16360
rect 472681 16350 472705 16360
rect 472681 16326 472715 16350
rect 472726 16326 472798 16360
rect 472681 16316 472798 16326
rect 472453 16292 472798 16316
rect 472466 16248 472666 16292
rect 472681 16282 472705 16292
rect 472681 16258 472715 16282
rect 472726 16258 472798 16292
rect 472681 16248 472798 16258
rect 472453 16224 472798 16248
rect 472466 16180 472666 16224
rect 472681 16214 472705 16224
rect 472681 16190 472715 16214
rect 472726 16190 472798 16224
rect 472681 16180 472798 16190
rect 472453 16156 472798 16180
rect 472466 16112 472666 16156
rect 472681 16146 472705 16156
rect 472681 16122 472715 16146
rect 472726 16122 472798 16156
rect 472681 16112 472798 16122
rect 472453 16088 472798 16112
rect 472466 16044 472666 16088
rect 472681 16078 472705 16088
rect 472681 16054 472715 16078
rect 472726 16054 472798 16088
rect 472681 16044 472798 16054
rect 472453 16020 472798 16044
rect 472466 15976 472666 16020
rect 472681 16010 472705 16020
rect 472681 15986 472715 16010
rect 472726 15986 472798 16020
rect 472681 15976 472798 15986
rect 472453 15952 472798 15976
rect 472466 15908 472666 15952
rect 472681 15942 472705 15952
rect 472681 15918 472715 15942
rect 472726 15918 472798 15952
rect 472681 15908 472798 15918
rect 472453 15884 472798 15908
rect 472466 15840 472666 15884
rect 472681 15874 472705 15884
rect 472681 15850 472715 15874
rect 472726 15850 472798 15884
rect 472681 15840 472798 15850
rect 472453 15816 472798 15840
rect 472466 15772 472666 15816
rect 472681 15806 472705 15816
rect 472681 15782 472715 15806
rect 472726 15782 472798 15816
rect 472681 15772 472798 15782
rect 472453 15748 472798 15772
rect 472466 15678 472666 15748
rect 472681 15724 472705 15748
rect 472726 15678 472798 15748
rect 473028 15678 473084 16678
rect 473100 15678 473156 16678
rect 473458 16656 473658 16678
rect 473673 16666 473707 16690
rect 474461 16678 474495 16690
rect 473718 16666 473790 16678
rect 473673 16656 473790 16666
rect 473445 16632 473790 16656
rect 473458 16588 473658 16632
rect 473673 16622 473697 16632
rect 473673 16598 473707 16622
rect 473718 16598 473790 16632
rect 473673 16588 473790 16598
rect 473445 16564 473790 16588
rect 473458 16520 473658 16564
rect 473673 16554 473697 16564
rect 473673 16530 473707 16554
rect 473718 16530 473790 16564
rect 473673 16520 473790 16530
rect 473445 16496 473790 16520
rect 473458 16452 473658 16496
rect 473673 16486 473697 16496
rect 473673 16462 473707 16486
rect 473718 16462 473790 16496
rect 473673 16452 473790 16462
rect 473445 16428 473790 16452
rect 473458 16384 473658 16428
rect 473673 16418 473697 16428
rect 473673 16394 473707 16418
rect 473718 16394 473790 16428
rect 473673 16384 473790 16394
rect 473445 16360 473790 16384
rect 473458 16316 473658 16360
rect 473673 16350 473697 16360
rect 473673 16326 473707 16350
rect 473718 16326 473790 16360
rect 473673 16316 473790 16326
rect 473445 16292 473790 16316
rect 473458 16248 473658 16292
rect 473673 16282 473697 16292
rect 473673 16258 473707 16282
rect 473718 16258 473790 16292
rect 473673 16248 473790 16258
rect 473445 16224 473790 16248
rect 473458 16180 473658 16224
rect 473673 16214 473697 16224
rect 473673 16190 473707 16214
rect 473718 16190 473790 16224
rect 473673 16180 473790 16190
rect 473445 16156 473790 16180
rect 473458 16112 473658 16156
rect 473673 16146 473697 16156
rect 473673 16122 473707 16146
rect 473718 16122 473790 16156
rect 473673 16112 473790 16122
rect 473445 16088 473790 16112
rect 473458 16044 473658 16088
rect 473673 16078 473697 16088
rect 473673 16054 473707 16078
rect 473718 16054 473790 16088
rect 473673 16044 473790 16054
rect 473445 16020 473790 16044
rect 473458 15976 473658 16020
rect 473673 16010 473697 16020
rect 473673 15986 473707 16010
rect 473718 15986 473790 16020
rect 473673 15976 473790 15986
rect 473445 15952 473790 15976
rect 473458 15908 473658 15952
rect 473673 15942 473697 15952
rect 473673 15918 473707 15942
rect 473718 15918 473790 15952
rect 473673 15908 473790 15918
rect 473445 15884 473790 15908
rect 473458 15840 473658 15884
rect 473673 15874 473697 15884
rect 473673 15850 473707 15874
rect 473718 15850 473790 15884
rect 473673 15840 473790 15850
rect 473445 15816 473790 15840
rect 473458 15772 473658 15816
rect 473673 15806 473697 15816
rect 473673 15782 473707 15806
rect 473718 15782 473790 15816
rect 473673 15772 473790 15782
rect 473445 15748 473790 15772
rect 473458 15678 473658 15748
rect 473673 15724 473697 15748
rect 473718 15678 473790 15748
rect 474020 15678 474076 16678
rect 474092 15678 474148 16678
rect 474450 16656 474650 16678
rect 474665 16666 474699 16690
rect 475453 16678 475487 16690
rect 474710 16666 474782 16678
rect 474665 16656 474782 16666
rect 474437 16632 474782 16656
rect 474450 16588 474650 16632
rect 474665 16622 474689 16632
rect 474665 16598 474699 16622
rect 474710 16598 474782 16632
rect 474665 16588 474782 16598
rect 474437 16564 474782 16588
rect 474450 16520 474650 16564
rect 474665 16554 474689 16564
rect 474665 16530 474699 16554
rect 474710 16530 474782 16564
rect 474665 16520 474782 16530
rect 474437 16496 474782 16520
rect 474450 16452 474650 16496
rect 474665 16486 474689 16496
rect 474665 16462 474699 16486
rect 474710 16462 474782 16496
rect 474665 16452 474782 16462
rect 474437 16428 474782 16452
rect 474450 16384 474650 16428
rect 474665 16418 474689 16428
rect 474665 16394 474699 16418
rect 474710 16394 474782 16428
rect 474665 16384 474782 16394
rect 474437 16360 474782 16384
rect 474450 16316 474650 16360
rect 474665 16350 474689 16360
rect 474665 16326 474699 16350
rect 474710 16326 474782 16360
rect 474665 16316 474782 16326
rect 474437 16292 474782 16316
rect 474450 16248 474650 16292
rect 474665 16282 474689 16292
rect 474665 16258 474699 16282
rect 474710 16258 474782 16292
rect 474665 16248 474782 16258
rect 474437 16224 474782 16248
rect 474450 16180 474650 16224
rect 474665 16214 474689 16224
rect 474665 16190 474699 16214
rect 474710 16190 474782 16224
rect 474665 16180 474782 16190
rect 474437 16156 474782 16180
rect 474450 16112 474650 16156
rect 474665 16146 474689 16156
rect 474665 16122 474699 16146
rect 474710 16122 474782 16156
rect 474665 16112 474782 16122
rect 474437 16088 474782 16112
rect 474450 16044 474650 16088
rect 474665 16078 474689 16088
rect 474665 16054 474699 16078
rect 474710 16054 474782 16088
rect 474665 16044 474782 16054
rect 474437 16020 474782 16044
rect 474450 15976 474650 16020
rect 474665 16010 474689 16020
rect 474665 15986 474699 16010
rect 474710 15986 474782 16020
rect 474665 15976 474782 15986
rect 474437 15952 474782 15976
rect 474450 15908 474650 15952
rect 474665 15942 474689 15952
rect 474665 15918 474699 15942
rect 474710 15918 474782 15952
rect 474665 15908 474782 15918
rect 474437 15884 474782 15908
rect 474450 15840 474650 15884
rect 474665 15874 474689 15884
rect 474665 15850 474699 15874
rect 474710 15850 474782 15884
rect 474665 15840 474782 15850
rect 474437 15816 474782 15840
rect 474450 15772 474650 15816
rect 474665 15806 474689 15816
rect 474665 15782 474699 15806
rect 474710 15782 474782 15816
rect 474665 15772 474782 15782
rect 474437 15748 474782 15772
rect 474450 15678 474650 15748
rect 474665 15724 474689 15748
rect 474710 15678 474782 15748
rect 475012 15678 475068 16678
rect 475084 15678 475140 16678
rect 475442 16656 475642 16678
rect 475657 16666 475691 16690
rect 476445 16678 476479 16690
rect 475702 16666 475774 16678
rect 475657 16656 475774 16666
rect 475429 16632 475774 16656
rect 475442 16588 475642 16632
rect 475657 16622 475681 16632
rect 475657 16598 475691 16622
rect 475702 16598 475774 16632
rect 475657 16588 475774 16598
rect 475429 16564 475774 16588
rect 475442 16520 475642 16564
rect 475657 16554 475681 16564
rect 475657 16530 475691 16554
rect 475702 16530 475774 16564
rect 475657 16520 475774 16530
rect 475429 16496 475774 16520
rect 475442 16452 475642 16496
rect 475657 16486 475681 16496
rect 475657 16462 475691 16486
rect 475702 16462 475774 16496
rect 475657 16452 475774 16462
rect 475429 16428 475774 16452
rect 475442 16384 475642 16428
rect 475657 16418 475681 16428
rect 475657 16394 475691 16418
rect 475702 16394 475774 16428
rect 475657 16384 475774 16394
rect 475429 16360 475774 16384
rect 475442 16316 475642 16360
rect 475657 16350 475681 16360
rect 475657 16326 475691 16350
rect 475702 16326 475774 16360
rect 475657 16316 475774 16326
rect 475429 16292 475774 16316
rect 475442 16248 475642 16292
rect 475657 16282 475681 16292
rect 475657 16258 475691 16282
rect 475702 16258 475774 16292
rect 475657 16248 475774 16258
rect 475429 16224 475774 16248
rect 475442 16180 475642 16224
rect 475657 16214 475681 16224
rect 475657 16190 475691 16214
rect 475702 16190 475774 16224
rect 475657 16180 475774 16190
rect 475429 16156 475774 16180
rect 475442 16112 475642 16156
rect 475657 16146 475681 16156
rect 475657 16122 475691 16146
rect 475702 16122 475774 16156
rect 475657 16112 475774 16122
rect 475429 16088 475774 16112
rect 475442 16044 475642 16088
rect 475657 16078 475681 16088
rect 475657 16054 475691 16078
rect 475702 16054 475774 16088
rect 475657 16044 475774 16054
rect 475429 16020 475774 16044
rect 475442 15976 475642 16020
rect 475657 16010 475681 16020
rect 475657 15986 475691 16010
rect 475702 15986 475774 16020
rect 475657 15976 475774 15986
rect 475429 15952 475774 15976
rect 475442 15908 475642 15952
rect 475657 15942 475681 15952
rect 475657 15918 475691 15942
rect 475702 15918 475774 15952
rect 475657 15908 475774 15918
rect 475429 15884 475774 15908
rect 475442 15840 475642 15884
rect 475657 15874 475681 15884
rect 475657 15850 475691 15874
rect 475702 15850 475774 15884
rect 475657 15840 475774 15850
rect 475429 15816 475774 15840
rect 475442 15772 475642 15816
rect 475657 15806 475681 15816
rect 475657 15782 475691 15806
rect 475702 15782 475774 15816
rect 475657 15772 475774 15782
rect 475429 15748 475774 15772
rect 475442 15678 475642 15748
rect 475657 15724 475681 15748
rect 475702 15678 475774 15748
rect 476004 15678 476060 16678
rect 476076 15678 476132 16678
rect 476434 16656 476634 16678
rect 476649 16666 476683 16690
rect 477437 16678 477471 16690
rect 476694 16666 476766 16678
rect 476649 16656 476766 16666
rect 476421 16632 476766 16656
rect 476434 16588 476634 16632
rect 476649 16622 476673 16632
rect 476649 16598 476683 16622
rect 476694 16598 476766 16632
rect 476649 16588 476766 16598
rect 476421 16564 476766 16588
rect 476434 16520 476634 16564
rect 476649 16554 476673 16564
rect 476649 16530 476683 16554
rect 476694 16530 476766 16564
rect 476649 16520 476766 16530
rect 476421 16496 476766 16520
rect 476434 16452 476634 16496
rect 476649 16486 476673 16496
rect 476649 16462 476683 16486
rect 476694 16462 476766 16496
rect 476649 16452 476766 16462
rect 476421 16428 476766 16452
rect 476434 16384 476634 16428
rect 476649 16418 476673 16428
rect 476649 16394 476683 16418
rect 476694 16394 476766 16428
rect 476649 16384 476766 16394
rect 476421 16360 476766 16384
rect 476434 16316 476634 16360
rect 476649 16350 476673 16360
rect 476649 16326 476683 16350
rect 476694 16326 476766 16360
rect 476649 16316 476766 16326
rect 476421 16292 476766 16316
rect 476434 16248 476634 16292
rect 476649 16282 476673 16292
rect 476649 16258 476683 16282
rect 476694 16258 476766 16292
rect 476649 16248 476766 16258
rect 476421 16224 476766 16248
rect 476434 16180 476634 16224
rect 476649 16214 476673 16224
rect 476649 16190 476683 16214
rect 476694 16190 476766 16224
rect 476649 16180 476766 16190
rect 476421 16156 476766 16180
rect 476434 16112 476634 16156
rect 476649 16146 476673 16156
rect 476649 16122 476683 16146
rect 476694 16122 476766 16156
rect 476649 16112 476766 16122
rect 476421 16088 476766 16112
rect 476434 16044 476634 16088
rect 476649 16078 476673 16088
rect 476649 16054 476683 16078
rect 476694 16054 476766 16088
rect 476649 16044 476766 16054
rect 476421 16020 476766 16044
rect 476434 15976 476634 16020
rect 476649 16010 476673 16020
rect 476649 15986 476683 16010
rect 476694 15986 476766 16020
rect 476649 15976 476766 15986
rect 476421 15952 476766 15976
rect 476434 15908 476634 15952
rect 476649 15942 476673 15952
rect 476649 15918 476683 15942
rect 476694 15918 476766 15952
rect 476649 15908 476766 15918
rect 476421 15884 476766 15908
rect 476434 15840 476634 15884
rect 476649 15874 476673 15884
rect 476649 15850 476683 15874
rect 476694 15850 476766 15884
rect 476649 15840 476766 15850
rect 476421 15816 476766 15840
rect 476434 15772 476634 15816
rect 476649 15806 476673 15816
rect 476649 15782 476683 15806
rect 476694 15782 476766 15816
rect 476649 15772 476766 15782
rect 476421 15748 476766 15772
rect 476434 15678 476634 15748
rect 476649 15724 476673 15748
rect 476694 15678 476766 15748
rect 476996 15678 477052 16678
rect 477068 15678 477124 16678
rect 477426 16656 477626 16678
rect 477641 16666 477675 16690
rect 477686 16666 477758 16678
rect 477641 16656 477758 16666
rect 477413 16632 477758 16656
rect 477426 16588 477626 16632
rect 477641 16622 477665 16632
rect 477641 16598 477675 16622
rect 477686 16598 477758 16632
rect 477641 16588 477758 16598
rect 477413 16564 477758 16588
rect 477426 16520 477626 16564
rect 477641 16554 477665 16564
rect 477641 16530 477675 16554
rect 477686 16530 477758 16564
rect 477641 16520 477758 16530
rect 477413 16496 477758 16520
rect 477426 16452 477626 16496
rect 477641 16486 477665 16496
rect 477641 16462 477675 16486
rect 477686 16462 477758 16496
rect 477641 16452 477758 16462
rect 477413 16428 477758 16452
rect 477426 16384 477626 16428
rect 477641 16418 477665 16428
rect 477641 16394 477675 16418
rect 477686 16394 477758 16428
rect 477641 16384 477758 16394
rect 477413 16360 477758 16384
rect 477426 16316 477626 16360
rect 477641 16350 477665 16360
rect 477641 16326 477675 16350
rect 477686 16326 477758 16360
rect 477641 16316 477758 16326
rect 477413 16292 477758 16316
rect 477426 16248 477626 16292
rect 477641 16282 477665 16292
rect 477641 16258 477675 16282
rect 477686 16258 477758 16292
rect 477641 16248 477758 16258
rect 477413 16224 477758 16248
rect 477426 16180 477626 16224
rect 477641 16214 477665 16224
rect 477641 16190 477675 16214
rect 477686 16190 477758 16224
rect 477641 16180 477758 16190
rect 477413 16156 477758 16180
rect 477426 16112 477626 16156
rect 477641 16146 477665 16156
rect 477641 16122 477675 16146
rect 477686 16122 477758 16156
rect 477641 16112 477758 16122
rect 477413 16088 477758 16112
rect 477426 16044 477626 16088
rect 477641 16078 477665 16088
rect 477641 16054 477675 16078
rect 477686 16054 477758 16088
rect 477641 16044 477758 16054
rect 477413 16020 477758 16044
rect 477426 15976 477626 16020
rect 477641 16010 477665 16020
rect 477641 15986 477675 16010
rect 477686 15986 477758 16020
rect 477641 15976 477758 15986
rect 477413 15952 477758 15976
rect 477426 15908 477626 15952
rect 477641 15942 477665 15952
rect 477641 15918 477675 15942
rect 477686 15918 477758 15952
rect 477641 15908 477758 15918
rect 477413 15884 477758 15908
rect 477426 15840 477626 15884
rect 477641 15874 477665 15884
rect 477641 15850 477675 15874
rect 477686 15850 477758 15884
rect 477641 15840 477758 15850
rect 477413 15816 477758 15840
rect 477426 15772 477626 15816
rect 477641 15806 477665 15816
rect 477641 15782 477675 15806
rect 477686 15782 477758 15816
rect 477641 15772 477758 15782
rect 477413 15748 477758 15772
rect 477426 15678 477626 15748
rect 477641 15724 477665 15748
rect 477686 15678 477758 15748
rect 477988 15678 478044 16678
rect 478060 15678 478116 16678
rect 478327 15678 478377 16678
rect 479065 14844 479172 19390
rect 516903 17278 516936 18278
rect 517106 17278 517123 18278
rect 517582 17278 517722 18278
rect 518084 17278 518140 18278
rect 518156 17278 518212 18278
rect 529486 17278 529626 18278
rect 529988 17278 530044 18278
rect 530060 17278 530116 18278
rect 530327 17278 530377 18278
rect 516746 15878 516780 15908
rect 516708 15840 516780 15870
rect 516903 15678 516936 16678
rect 517106 15678 517123 16678
rect 517582 15678 517722 16678
rect 518084 15678 518140 16678
rect 518156 15678 518212 16678
rect 529486 15678 529626 16678
rect 529988 15678 530044 16678
rect 530060 15678 530116 16678
rect 530327 15678 530377 16678
rect 531065 14844 531172 19390
rect 564903 17278 564936 18278
rect 565106 17278 565123 18278
rect 565261 17278 565333 18278
rect 565522 18198 565722 18278
rect 565737 18208 565771 18232
rect 565782 18208 565854 18278
rect 565737 18198 565854 18208
rect 565509 18174 565854 18198
rect 565522 18130 565722 18174
rect 565737 18164 565761 18174
rect 565737 18140 565771 18164
rect 565782 18140 565854 18174
rect 565737 18130 565854 18140
rect 565509 18106 565854 18130
rect 565522 18062 565722 18106
rect 565737 18096 565761 18106
rect 565737 18072 565771 18096
rect 565782 18072 565854 18106
rect 565737 18062 565854 18072
rect 565509 18038 565854 18062
rect 565522 17994 565722 18038
rect 565737 18028 565761 18038
rect 565737 18004 565771 18028
rect 565782 18004 565854 18038
rect 565737 17994 565854 18004
rect 565509 17970 565854 17994
rect 565522 17926 565722 17970
rect 565737 17960 565761 17970
rect 565737 17936 565771 17960
rect 565782 17936 565854 17970
rect 565737 17926 565854 17936
rect 565509 17902 565854 17926
rect 565522 17858 565722 17902
rect 565737 17892 565761 17902
rect 565737 17868 565771 17892
rect 565782 17868 565854 17902
rect 565737 17858 565854 17868
rect 565509 17834 565854 17858
rect 565522 17790 565722 17834
rect 565737 17824 565761 17834
rect 565737 17800 565771 17824
rect 565782 17800 565854 17834
rect 565737 17790 565854 17800
rect 565509 17766 565854 17790
rect 565522 17722 565722 17766
rect 565737 17756 565761 17766
rect 565737 17732 565771 17756
rect 565782 17732 565854 17766
rect 565737 17722 565854 17732
rect 565509 17698 565854 17722
rect 565522 17654 565722 17698
rect 565737 17688 565761 17698
rect 565737 17664 565771 17688
rect 565782 17664 565854 17698
rect 565737 17654 565854 17664
rect 565509 17630 565854 17654
rect 565522 17586 565722 17630
rect 565737 17620 565761 17630
rect 565737 17596 565771 17620
rect 565782 17596 565854 17630
rect 565737 17586 565854 17596
rect 565509 17562 565854 17586
rect 565522 17518 565722 17562
rect 565737 17552 565761 17562
rect 565737 17528 565771 17552
rect 565782 17528 565854 17562
rect 565737 17518 565854 17528
rect 565509 17494 565854 17518
rect 565522 17450 565722 17494
rect 565737 17484 565761 17494
rect 565737 17460 565771 17484
rect 565782 17460 565854 17494
rect 565737 17450 565854 17460
rect 565509 17426 565854 17450
rect 565522 17382 565722 17426
rect 565737 17416 565761 17426
rect 565737 17392 565771 17416
rect 565782 17392 565854 17426
rect 565737 17382 565854 17392
rect 565509 17358 565854 17382
rect 565522 17314 565722 17358
rect 565737 17348 565761 17358
rect 565737 17324 565771 17348
rect 565782 17324 565854 17358
rect 565737 17314 565854 17324
rect 565509 17290 565854 17314
rect 565522 17278 565722 17290
rect 565533 17266 565557 17278
rect 565737 17266 565761 17290
rect 565782 17278 565854 17290
rect 566084 17278 566140 18278
rect 566156 17278 566212 18278
rect 566514 18198 566714 18278
rect 566729 18208 566763 18232
rect 566774 18208 566846 18278
rect 566729 18198 566846 18208
rect 566501 18174 566846 18198
rect 566514 18130 566714 18174
rect 566729 18164 566753 18174
rect 566729 18140 566763 18164
rect 566774 18140 566846 18174
rect 566729 18130 566846 18140
rect 566501 18106 566846 18130
rect 566514 18062 566714 18106
rect 566729 18096 566753 18106
rect 566729 18072 566763 18096
rect 566774 18072 566846 18106
rect 566729 18062 566846 18072
rect 566501 18038 566846 18062
rect 566514 17994 566714 18038
rect 566729 18028 566753 18038
rect 566729 18004 566763 18028
rect 566774 18004 566846 18038
rect 566729 17994 566846 18004
rect 566501 17970 566846 17994
rect 566514 17926 566714 17970
rect 566729 17960 566753 17970
rect 566729 17936 566763 17960
rect 566774 17936 566846 17970
rect 566729 17926 566846 17936
rect 566501 17902 566846 17926
rect 566514 17858 566714 17902
rect 566729 17892 566753 17902
rect 566729 17868 566763 17892
rect 566774 17868 566846 17902
rect 566729 17858 566846 17868
rect 566501 17834 566846 17858
rect 566514 17790 566714 17834
rect 566729 17824 566753 17834
rect 566729 17800 566763 17824
rect 566774 17800 566846 17834
rect 566729 17790 566846 17800
rect 566501 17766 566846 17790
rect 566514 17722 566714 17766
rect 566729 17756 566753 17766
rect 566729 17732 566763 17756
rect 566774 17732 566846 17766
rect 566729 17722 566846 17732
rect 566501 17698 566846 17722
rect 566514 17654 566714 17698
rect 566729 17688 566753 17698
rect 566729 17664 566763 17688
rect 566774 17664 566846 17698
rect 566729 17654 566846 17664
rect 566501 17630 566846 17654
rect 566514 17586 566714 17630
rect 566729 17620 566753 17630
rect 566729 17596 566763 17620
rect 566774 17596 566846 17630
rect 566729 17586 566846 17596
rect 566501 17562 566846 17586
rect 566514 17518 566714 17562
rect 566729 17552 566753 17562
rect 566729 17528 566763 17552
rect 566774 17528 566846 17562
rect 566729 17518 566846 17528
rect 566501 17494 566846 17518
rect 566514 17450 566714 17494
rect 566729 17484 566753 17494
rect 566729 17460 566763 17484
rect 566774 17460 566846 17494
rect 566729 17450 566846 17460
rect 566501 17426 566846 17450
rect 566514 17382 566714 17426
rect 566729 17416 566753 17426
rect 566729 17392 566763 17416
rect 566774 17392 566846 17426
rect 566729 17382 566846 17392
rect 566501 17358 566846 17382
rect 566514 17314 566714 17358
rect 566729 17348 566753 17358
rect 566729 17324 566763 17348
rect 566774 17324 566846 17358
rect 566729 17314 566846 17324
rect 566501 17290 566846 17314
rect 566514 17278 566714 17290
rect 566525 17266 566549 17278
rect 566729 17266 566753 17290
rect 566774 17278 566846 17290
rect 567076 17278 567132 18278
rect 567148 17278 567204 18278
rect 567506 18198 567706 18278
rect 567721 18208 567755 18232
rect 567766 18208 567838 18278
rect 567721 18198 567838 18208
rect 567493 18174 567838 18198
rect 567506 18130 567706 18174
rect 567721 18164 567745 18174
rect 567721 18140 567755 18164
rect 567766 18140 567838 18174
rect 567721 18130 567838 18140
rect 567493 18106 567838 18130
rect 567506 18062 567706 18106
rect 567721 18096 567745 18106
rect 567721 18072 567755 18096
rect 567766 18072 567838 18106
rect 567721 18062 567838 18072
rect 567493 18038 567838 18062
rect 567506 17994 567706 18038
rect 567721 18028 567745 18038
rect 567721 18004 567755 18028
rect 567766 18004 567838 18038
rect 567721 17994 567838 18004
rect 567493 17970 567838 17994
rect 567506 17926 567706 17970
rect 567721 17960 567745 17970
rect 567721 17936 567755 17960
rect 567766 17936 567838 17970
rect 567721 17926 567838 17936
rect 567493 17902 567838 17926
rect 567506 17858 567706 17902
rect 567721 17892 567745 17902
rect 567721 17868 567755 17892
rect 567766 17868 567838 17902
rect 567721 17858 567838 17868
rect 567493 17834 567838 17858
rect 567506 17790 567706 17834
rect 567721 17824 567745 17834
rect 567721 17800 567755 17824
rect 567766 17800 567838 17834
rect 567721 17790 567838 17800
rect 567493 17766 567838 17790
rect 567506 17722 567706 17766
rect 567721 17756 567745 17766
rect 567721 17732 567755 17756
rect 567766 17732 567838 17766
rect 567721 17722 567838 17732
rect 567493 17698 567838 17722
rect 567506 17654 567706 17698
rect 567721 17688 567745 17698
rect 567721 17664 567755 17688
rect 567766 17664 567838 17698
rect 567721 17654 567838 17664
rect 567493 17630 567838 17654
rect 567506 17586 567706 17630
rect 567721 17620 567745 17630
rect 567721 17596 567755 17620
rect 567766 17596 567838 17630
rect 567721 17586 567838 17596
rect 567493 17562 567838 17586
rect 567506 17518 567706 17562
rect 567721 17552 567745 17562
rect 567721 17528 567755 17552
rect 567766 17528 567838 17562
rect 567721 17518 567838 17528
rect 567493 17494 567838 17518
rect 567506 17450 567706 17494
rect 567721 17484 567745 17494
rect 567721 17460 567755 17484
rect 567766 17460 567838 17494
rect 567721 17450 567838 17460
rect 567493 17426 567838 17450
rect 567506 17382 567706 17426
rect 567721 17416 567745 17426
rect 567721 17392 567755 17416
rect 567766 17392 567838 17426
rect 567721 17382 567838 17392
rect 567493 17358 567838 17382
rect 567506 17314 567706 17358
rect 567721 17348 567745 17358
rect 567721 17324 567755 17348
rect 567766 17324 567838 17358
rect 567721 17314 567838 17324
rect 567493 17290 567838 17314
rect 567506 17278 567706 17290
rect 567517 17266 567541 17278
rect 567721 17266 567745 17290
rect 567766 17278 567838 17290
rect 568068 17278 568124 18278
rect 568140 17278 568196 18278
rect 568498 18198 568698 18278
rect 568713 18208 568747 18232
rect 568758 18208 568830 18278
rect 568713 18198 568830 18208
rect 568485 18174 568830 18198
rect 568498 18130 568698 18174
rect 568713 18164 568737 18174
rect 568713 18140 568747 18164
rect 568758 18140 568830 18174
rect 568713 18130 568830 18140
rect 568485 18106 568830 18130
rect 568498 18062 568698 18106
rect 568713 18096 568737 18106
rect 568713 18072 568747 18096
rect 568758 18072 568830 18106
rect 568713 18062 568830 18072
rect 568485 18038 568830 18062
rect 568498 17994 568698 18038
rect 568713 18028 568737 18038
rect 568713 18004 568747 18028
rect 568758 18004 568830 18038
rect 568713 17994 568830 18004
rect 568485 17970 568830 17994
rect 568498 17926 568698 17970
rect 568713 17960 568737 17970
rect 568713 17936 568747 17960
rect 568758 17936 568830 17970
rect 568713 17926 568830 17936
rect 568485 17902 568830 17926
rect 568498 17858 568698 17902
rect 568713 17892 568737 17902
rect 568713 17868 568747 17892
rect 568758 17868 568830 17902
rect 568713 17858 568830 17868
rect 568485 17834 568830 17858
rect 568498 17790 568698 17834
rect 568713 17824 568737 17834
rect 568713 17800 568747 17824
rect 568758 17800 568830 17834
rect 568713 17790 568830 17800
rect 568485 17766 568830 17790
rect 568498 17722 568698 17766
rect 568713 17756 568737 17766
rect 568713 17732 568747 17756
rect 568758 17732 568830 17766
rect 568713 17722 568830 17732
rect 568485 17698 568830 17722
rect 568498 17654 568698 17698
rect 568713 17688 568737 17698
rect 568713 17664 568747 17688
rect 568758 17664 568830 17698
rect 568713 17654 568830 17664
rect 568485 17630 568830 17654
rect 568498 17586 568698 17630
rect 568713 17620 568737 17630
rect 568713 17596 568747 17620
rect 568758 17596 568830 17630
rect 568713 17586 568830 17596
rect 568485 17562 568830 17586
rect 568498 17518 568698 17562
rect 568713 17552 568737 17562
rect 568713 17528 568747 17552
rect 568758 17528 568830 17562
rect 568713 17518 568830 17528
rect 568485 17494 568830 17518
rect 568498 17450 568698 17494
rect 568713 17484 568737 17494
rect 568713 17460 568747 17484
rect 568758 17460 568830 17494
rect 568713 17450 568830 17460
rect 568485 17426 568830 17450
rect 568498 17382 568698 17426
rect 568713 17416 568737 17426
rect 568713 17392 568747 17416
rect 568758 17392 568830 17426
rect 568713 17382 568830 17392
rect 568485 17358 568830 17382
rect 568498 17314 568698 17358
rect 568713 17348 568737 17358
rect 568713 17324 568747 17348
rect 568758 17324 568830 17358
rect 568713 17314 568830 17324
rect 568485 17290 568830 17314
rect 568498 17278 568698 17290
rect 568509 17266 568533 17278
rect 568713 17266 568737 17290
rect 568758 17278 568830 17290
rect 569060 17278 569116 18278
rect 569132 17278 569188 18278
rect 569490 18198 569690 18278
rect 569705 18208 569739 18232
rect 569750 18208 569822 18278
rect 569705 18198 569822 18208
rect 569477 18174 569822 18198
rect 569490 18130 569690 18174
rect 569705 18164 569729 18174
rect 569705 18140 569739 18164
rect 569750 18140 569822 18174
rect 569705 18130 569822 18140
rect 569477 18106 569822 18130
rect 569490 18062 569690 18106
rect 569705 18096 569729 18106
rect 569705 18072 569739 18096
rect 569750 18072 569822 18106
rect 569705 18062 569822 18072
rect 569477 18038 569822 18062
rect 569490 17994 569690 18038
rect 569705 18028 569729 18038
rect 569705 18004 569739 18028
rect 569750 18004 569822 18038
rect 569705 17994 569822 18004
rect 569477 17970 569822 17994
rect 569490 17926 569690 17970
rect 569705 17960 569729 17970
rect 569705 17936 569739 17960
rect 569750 17936 569822 17970
rect 569705 17926 569822 17936
rect 569477 17902 569822 17926
rect 569490 17858 569690 17902
rect 569705 17892 569729 17902
rect 569705 17868 569739 17892
rect 569750 17868 569822 17902
rect 569705 17858 569822 17868
rect 569477 17834 569822 17858
rect 569490 17790 569690 17834
rect 569705 17824 569729 17834
rect 569705 17800 569739 17824
rect 569750 17800 569822 17834
rect 569705 17790 569822 17800
rect 569477 17766 569822 17790
rect 569490 17722 569690 17766
rect 569705 17756 569729 17766
rect 569705 17732 569739 17756
rect 569750 17732 569822 17766
rect 569705 17722 569822 17732
rect 569477 17698 569822 17722
rect 569490 17654 569690 17698
rect 569705 17688 569729 17698
rect 569705 17664 569739 17688
rect 569750 17664 569822 17698
rect 569705 17654 569822 17664
rect 569477 17630 569822 17654
rect 569490 17586 569690 17630
rect 569705 17620 569729 17630
rect 569705 17596 569739 17620
rect 569750 17596 569822 17630
rect 569705 17586 569822 17596
rect 569477 17562 569822 17586
rect 569490 17518 569690 17562
rect 569705 17552 569729 17562
rect 569705 17528 569739 17552
rect 569750 17528 569822 17562
rect 569705 17518 569822 17528
rect 569477 17494 569822 17518
rect 569490 17450 569690 17494
rect 569705 17484 569729 17494
rect 569705 17460 569739 17484
rect 569750 17460 569822 17494
rect 569705 17450 569822 17460
rect 569477 17426 569822 17450
rect 569490 17382 569690 17426
rect 569705 17416 569729 17426
rect 569705 17392 569739 17416
rect 569750 17392 569822 17426
rect 569705 17382 569822 17392
rect 569477 17358 569822 17382
rect 569490 17314 569690 17358
rect 569705 17348 569729 17358
rect 569705 17324 569739 17348
rect 569750 17324 569822 17358
rect 569705 17314 569822 17324
rect 569477 17290 569822 17314
rect 569490 17278 569690 17290
rect 569501 17266 569525 17278
rect 569705 17266 569729 17290
rect 569750 17278 569822 17290
rect 570052 17278 570108 18278
rect 570124 17278 570180 18278
rect 570482 18198 570682 18278
rect 570697 18208 570731 18232
rect 570742 18208 570814 18278
rect 570697 18198 570814 18208
rect 570469 18174 570814 18198
rect 570482 18130 570682 18174
rect 570697 18164 570721 18174
rect 570697 18140 570731 18164
rect 570742 18140 570814 18174
rect 570697 18130 570814 18140
rect 570469 18106 570814 18130
rect 570482 18062 570682 18106
rect 570697 18096 570721 18106
rect 570697 18072 570731 18096
rect 570742 18072 570814 18106
rect 570697 18062 570814 18072
rect 570469 18038 570814 18062
rect 570482 17994 570682 18038
rect 570697 18028 570721 18038
rect 570697 18004 570731 18028
rect 570742 18004 570814 18038
rect 570697 17994 570814 18004
rect 570469 17970 570814 17994
rect 570482 17926 570682 17970
rect 570697 17960 570721 17970
rect 570697 17936 570731 17960
rect 570742 17936 570814 17970
rect 570697 17926 570814 17936
rect 570469 17902 570814 17926
rect 570482 17858 570682 17902
rect 570697 17892 570721 17902
rect 570697 17868 570731 17892
rect 570742 17868 570814 17902
rect 570697 17858 570814 17868
rect 570469 17834 570814 17858
rect 570482 17790 570682 17834
rect 570697 17824 570721 17834
rect 570697 17800 570731 17824
rect 570742 17800 570814 17834
rect 570697 17790 570814 17800
rect 570469 17766 570814 17790
rect 570482 17722 570682 17766
rect 570697 17756 570721 17766
rect 570697 17732 570731 17756
rect 570742 17732 570814 17766
rect 570697 17722 570814 17732
rect 570469 17698 570814 17722
rect 570482 17654 570682 17698
rect 570697 17688 570721 17698
rect 570697 17664 570731 17688
rect 570742 17664 570814 17698
rect 570697 17654 570814 17664
rect 570469 17630 570814 17654
rect 570482 17586 570682 17630
rect 570697 17620 570721 17630
rect 570697 17596 570731 17620
rect 570742 17596 570814 17630
rect 570697 17586 570814 17596
rect 570469 17562 570814 17586
rect 570482 17518 570682 17562
rect 570697 17552 570721 17562
rect 570697 17528 570731 17552
rect 570742 17528 570814 17562
rect 570697 17518 570814 17528
rect 570469 17494 570814 17518
rect 570482 17450 570682 17494
rect 570697 17484 570721 17494
rect 570697 17460 570731 17484
rect 570742 17460 570814 17494
rect 570697 17450 570814 17460
rect 570469 17426 570814 17450
rect 570482 17382 570682 17426
rect 570697 17416 570721 17426
rect 570697 17392 570731 17416
rect 570742 17392 570814 17426
rect 570697 17382 570814 17392
rect 570469 17358 570814 17382
rect 570482 17314 570682 17358
rect 570697 17348 570721 17358
rect 570697 17324 570731 17348
rect 570742 17324 570814 17358
rect 570697 17314 570814 17324
rect 570469 17290 570814 17314
rect 570482 17278 570682 17290
rect 570493 17266 570517 17278
rect 570697 17266 570721 17290
rect 570742 17278 570814 17290
rect 571044 17278 571100 18278
rect 571116 17278 571172 18278
rect 571474 18198 571674 18278
rect 571689 18208 571723 18232
rect 571734 18208 571806 18278
rect 571689 18198 571806 18208
rect 571461 18174 571806 18198
rect 571474 18130 571674 18174
rect 571689 18164 571713 18174
rect 571689 18140 571723 18164
rect 571734 18140 571806 18174
rect 571689 18130 571806 18140
rect 571461 18106 571806 18130
rect 571474 18062 571674 18106
rect 571689 18096 571713 18106
rect 571689 18072 571723 18096
rect 571734 18072 571806 18106
rect 571689 18062 571806 18072
rect 571461 18038 571806 18062
rect 571474 17994 571674 18038
rect 571689 18028 571713 18038
rect 571689 18004 571723 18028
rect 571734 18004 571806 18038
rect 571689 17994 571806 18004
rect 571461 17970 571806 17994
rect 571474 17926 571674 17970
rect 571689 17960 571713 17970
rect 571689 17936 571723 17960
rect 571734 17936 571806 17970
rect 571689 17926 571806 17936
rect 571461 17902 571806 17926
rect 571474 17858 571674 17902
rect 571689 17892 571713 17902
rect 571689 17868 571723 17892
rect 571734 17868 571806 17902
rect 571689 17858 571806 17868
rect 571461 17834 571806 17858
rect 571474 17790 571674 17834
rect 571689 17824 571713 17834
rect 571689 17800 571723 17824
rect 571734 17800 571806 17834
rect 571689 17790 571806 17800
rect 571461 17766 571806 17790
rect 571474 17722 571674 17766
rect 571689 17756 571713 17766
rect 571689 17732 571723 17756
rect 571734 17732 571806 17766
rect 571689 17722 571806 17732
rect 571461 17698 571806 17722
rect 571474 17654 571674 17698
rect 571689 17688 571713 17698
rect 571689 17664 571723 17688
rect 571734 17664 571806 17698
rect 571689 17654 571806 17664
rect 571461 17630 571806 17654
rect 571474 17586 571674 17630
rect 571689 17620 571713 17630
rect 571689 17596 571723 17620
rect 571734 17596 571806 17630
rect 571689 17586 571806 17596
rect 571461 17562 571806 17586
rect 571474 17518 571674 17562
rect 571689 17552 571713 17562
rect 571689 17528 571723 17552
rect 571734 17528 571806 17562
rect 571689 17518 571806 17528
rect 571461 17494 571806 17518
rect 571474 17450 571674 17494
rect 571689 17484 571713 17494
rect 571689 17460 571723 17484
rect 571734 17460 571806 17494
rect 571689 17450 571806 17460
rect 571461 17426 571806 17450
rect 571474 17382 571674 17426
rect 571689 17416 571713 17426
rect 571689 17392 571723 17416
rect 571734 17392 571806 17426
rect 571689 17382 571806 17392
rect 571461 17358 571806 17382
rect 571474 17314 571674 17358
rect 571689 17348 571713 17358
rect 571689 17324 571723 17348
rect 571734 17324 571806 17358
rect 571689 17314 571806 17324
rect 571461 17290 571806 17314
rect 571474 17278 571674 17290
rect 571485 17266 571509 17278
rect 571689 17266 571713 17290
rect 571734 17278 571806 17290
rect 572036 17278 572092 18278
rect 572108 17278 572164 18278
rect 572466 18198 572666 18278
rect 572681 18208 572715 18232
rect 572726 18208 572798 18278
rect 572681 18198 572798 18208
rect 572453 18174 572798 18198
rect 572466 18130 572666 18174
rect 572681 18164 572705 18174
rect 572681 18140 572715 18164
rect 572726 18140 572798 18174
rect 572681 18130 572798 18140
rect 572453 18106 572798 18130
rect 572466 18062 572666 18106
rect 572681 18096 572705 18106
rect 572681 18072 572715 18096
rect 572726 18072 572798 18106
rect 572681 18062 572798 18072
rect 572453 18038 572798 18062
rect 572466 17994 572666 18038
rect 572681 18028 572705 18038
rect 572681 18004 572715 18028
rect 572726 18004 572798 18038
rect 572681 17994 572798 18004
rect 572453 17970 572798 17994
rect 572466 17926 572666 17970
rect 572681 17960 572705 17970
rect 572681 17936 572715 17960
rect 572726 17936 572798 17970
rect 572681 17926 572798 17936
rect 572453 17902 572798 17926
rect 572466 17858 572666 17902
rect 572681 17892 572705 17902
rect 572681 17868 572715 17892
rect 572726 17868 572798 17902
rect 572681 17858 572798 17868
rect 572453 17834 572798 17858
rect 572466 17790 572666 17834
rect 572681 17824 572705 17834
rect 572681 17800 572715 17824
rect 572726 17800 572798 17834
rect 572681 17790 572798 17800
rect 572453 17766 572798 17790
rect 572466 17722 572666 17766
rect 572681 17756 572705 17766
rect 572681 17732 572715 17756
rect 572726 17732 572798 17766
rect 572681 17722 572798 17732
rect 572453 17698 572798 17722
rect 572466 17654 572666 17698
rect 572681 17688 572705 17698
rect 572681 17664 572715 17688
rect 572726 17664 572798 17698
rect 572681 17654 572798 17664
rect 572453 17630 572798 17654
rect 572466 17586 572666 17630
rect 572681 17620 572705 17630
rect 572681 17596 572715 17620
rect 572726 17596 572798 17630
rect 572681 17586 572798 17596
rect 572453 17562 572798 17586
rect 572466 17518 572666 17562
rect 572681 17552 572705 17562
rect 572681 17528 572715 17552
rect 572726 17528 572798 17562
rect 572681 17518 572798 17528
rect 572453 17494 572798 17518
rect 572466 17450 572666 17494
rect 572681 17484 572705 17494
rect 572681 17460 572715 17484
rect 572726 17460 572798 17494
rect 572681 17450 572798 17460
rect 572453 17426 572798 17450
rect 572466 17382 572666 17426
rect 572681 17416 572705 17426
rect 572681 17392 572715 17416
rect 572726 17392 572798 17426
rect 572681 17382 572798 17392
rect 572453 17358 572798 17382
rect 572466 17314 572666 17358
rect 572681 17348 572705 17358
rect 572681 17324 572715 17348
rect 572726 17324 572798 17358
rect 572681 17314 572798 17324
rect 572453 17290 572798 17314
rect 572466 17278 572666 17290
rect 572477 17266 572501 17278
rect 572681 17266 572705 17290
rect 572726 17278 572798 17290
rect 573028 17278 573084 18278
rect 573100 17278 573156 18278
rect 573458 18198 573658 18278
rect 573673 18208 573707 18232
rect 573718 18208 573790 18278
rect 573673 18198 573790 18208
rect 573445 18174 573790 18198
rect 573458 18130 573658 18174
rect 573673 18164 573697 18174
rect 573673 18140 573707 18164
rect 573718 18140 573790 18174
rect 573673 18130 573790 18140
rect 573445 18106 573790 18130
rect 573458 18062 573658 18106
rect 573673 18096 573697 18106
rect 573673 18072 573707 18096
rect 573718 18072 573790 18106
rect 573673 18062 573790 18072
rect 573445 18038 573790 18062
rect 573458 17994 573658 18038
rect 573673 18028 573697 18038
rect 573673 18004 573707 18028
rect 573718 18004 573790 18038
rect 573673 17994 573790 18004
rect 573445 17970 573790 17994
rect 573458 17926 573658 17970
rect 573673 17960 573697 17970
rect 573673 17936 573707 17960
rect 573718 17936 573790 17970
rect 573673 17926 573790 17936
rect 573445 17902 573790 17926
rect 573458 17858 573658 17902
rect 573673 17892 573697 17902
rect 573673 17868 573707 17892
rect 573718 17868 573790 17902
rect 573673 17858 573790 17868
rect 573445 17834 573790 17858
rect 573458 17790 573658 17834
rect 573673 17824 573697 17834
rect 573673 17800 573707 17824
rect 573718 17800 573790 17834
rect 573673 17790 573790 17800
rect 573445 17766 573790 17790
rect 573458 17722 573658 17766
rect 573673 17756 573697 17766
rect 573673 17732 573707 17756
rect 573718 17732 573790 17766
rect 573673 17722 573790 17732
rect 573445 17698 573790 17722
rect 573458 17654 573658 17698
rect 573673 17688 573697 17698
rect 573673 17664 573707 17688
rect 573718 17664 573790 17698
rect 573673 17654 573790 17664
rect 573445 17630 573790 17654
rect 573458 17586 573658 17630
rect 573673 17620 573697 17630
rect 573673 17596 573707 17620
rect 573718 17596 573790 17630
rect 573673 17586 573790 17596
rect 573445 17562 573790 17586
rect 573458 17518 573658 17562
rect 573673 17552 573697 17562
rect 573673 17528 573707 17552
rect 573718 17528 573790 17562
rect 573673 17518 573790 17528
rect 573445 17494 573790 17518
rect 573458 17450 573658 17494
rect 573673 17484 573697 17494
rect 573673 17460 573707 17484
rect 573718 17460 573790 17494
rect 573673 17450 573790 17460
rect 573445 17426 573790 17450
rect 573458 17382 573658 17426
rect 573673 17416 573697 17426
rect 573673 17392 573707 17416
rect 573718 17392 573790 17426
rect 573673 17382 573790 17392
rect 573445 17358 573790 17382
rect 573458 17314 573658 17358
rect 573673 17348 573697 17358
rect 573673 17324 573707 17348
rect 573718 17324 573790 17358
rect 573673 17314 573790 17324
rect 573445 17290 573790 17314
rect 573458 17278 573658 17290
rect 573469 17266 573493 17278
rect 573673 17266 573697 17290
rect 573718 17278 573790 17290
rect 574020 17278 574076 18278
rect 574092 17278 574148 18278
rect 574450 18198 574650 18278
rect 574665 18208 574699 18232
rect 574710 18208 574782 18278
rect 574665 18198 574782 18208
rect 574437 18174 574782 18198
rect 574450 18130 574650 18174
rect 574665 18164 574689 18174
rect 574665 18140 574699 18164
rect 574710 18140 574782 18174
rect 574665 18130 574782 18140
rect 574437 18106 574782 18130
rect 574450 18062 574650 18106
rect 574665 18096 574689 18106
rect 574665 18072 574699 18096
rect 574710 18072 574782 18106
rect 574665 18062 574782 18072
rect 574437 18038 574782 18062
rect 574450 17994 574650 18038
rect 574665 18028 574689 18038
rect 574665 18004 574699 18028
rect 574710 18004 574782 18038
rect 574665 17994 574782 18004
rect 574437 17970 574782 17994
rect 574450 17926 574650 17970
rect 574665 17960 574689 17970
rect 574665 17936 574699 17960
rect 574710 17936 574782 17970
rect 574665 17926 574782 17936
rect 574437 17902 574782 17926
rect 574450 17858 574650 17902
rect 574665 17892 574689 17902
rect 574665 17868 574699 17892
rect 574710 17868 574782 17902
rect 574665 17858 574782 17868
rect 574437 17834 574782 17858
rect 574450 17790 574650 17834
rect 574665 17824 574689 17834
rect 574665 17800 574699 17824
rect 574710 17800 574782 17834
rect 574665 17790 574782 17800
rect 574437 17766 574782 17790
rect 574450 17722 574650 17766
rect 574665 17756 574689 17766
rect 574665 17732 574699 17756
rect 574710 17732 574782 17766
rect 574665 17722 574782 17732
rect 574437 17698 574782 17722
rect 574450 17654 574650 17698
rect 574665 17688 574689 17698
rect 574665 17664 574699 17688
rect 574710 17664 574782 17698
rect 574665 17654 574782 17664
rect 574437 17630 574782 17654
rect 574450 17586 574650 17630
rect 574665 17620 574689 17630
rect 574665 17596 574699 17620
rect 574710 17596 574782 17630
rect 574665 17586 574782 17596
rect 574437 17562 574782 17586
rect 574450 17518 574650 17562
rect 574665 17552 574689 17562
rect 574665 17528 574699 17552
rect 574710 17528 574782 17562
rect 574665 17518 574782 17528
rect 574437 17494 574782 17518
rect 574450 17450 574650 17494
rect 574665 17484 574689 17494
rect 574665 17460 574699 17484
rect 574710 17460 574782 17494
rect 574665 17450 574782 17460
rect 574437 17426 574782 17450
rect 574450 17382 574650 17426
rect 574665 17416 574689 17426
rect 574665 17392 574699 17416
rect 574710 17392 574782 17426
rect 574665 17382 574782 17392
rect 574437 17358 574782 17382
rect 574450 17314 574650 17358
rect 574665 17348 574689 17358
rect 574665 17324 574699 17348
rect 574710 17324 574782 17358
rect 574665 17314 574782 17324
rect 574437 17290 574782 17314
rect 574450 17278 574650 17290
rect 574461 17266 574485 17278
rect 574665 17266 574689 17290
rect 574710 17278 574782 17290
rect 575012 17278 575068 18278
rect 575084 17278 575140 18278
rect 575442 18198 575642 18278
rect 575657 18208 575691 18232
rect 575702 18208 575774 18278
rect 575657 18198 575774 18208
rect 575429 18174 575774 18198
rect 575442 18130 575642 18174
rect 575657 18164 575681 18174
rect 575657 18140 575691 18164
rect 575702 18140 575774 18174
rect 575657 18130 575774 18140
rect 575429 18106 575774 18130
rect 575442 18062 575642 18106
rect 575657 18096 575681 18106
rect 575657 18072 575691 18096
rect 575702 18072 575774 18106
rect 575657 18062 575774 18072
rect 575429 18038 575774 18062
rect 575442 17994 575642 18038
rect 575657 18028 575681 18038
rect 575657 18004 575691 18028
rect 575702 18004 575774 18038
rect 575657 17994 575774 18004
rect 575429 17970 575774 17994
rect 575442 17926 575642 17970
rect 575657 17960 575681 17970
rect 575657 17936 575691 17960
rect 575702 17936 575774 17970
rect 575657 17926 575774 17936
rect 575429 17902 575774 17926
rect 575442 17858 575642 17902
rect 575657 17892 575681 17902
rect 575657 17868 575691 17892
rect 575702 17868 575774 17902
rect 575657 17858 575774 17868
rect 575429 17834 575774 17858
rect 575442 17790 575642 17834
rect 575657 17824 575681 17834
rect 575657 17800 575691 17824
rect 575702 17800 575774 17834
rect 575657 17790 575774 17800
rect 575429 17766 575774 17790
rect 575442 17722 575642 17766
rect 575657 17756 575681 17766
rect 575657 17732 575691 17756
rect 575702 17732 575774 17766
rect 575657 17722 575774 17732
rect 575429 17698 575774 17722
rect 575442 17654 575642 17698
rect 575657 17688 575681 17698
rect 575657 17664 575691 17688
rect 575702 17664 575774 17698
rect 575657 17654 575774 17664
rect 575429 17630 575774 17654
rect 575442 17586 575642 17630
rect 575657 17620 575681 17630
rect 575657 17596 575691 17620
rect 575702 17596 575774 17630
rect 575657 17586 575774 17596
rect 575429 17562 575774 17586
rect 575442 17518 575642 17562
rect 575657 17552 575681 17562
rect 575657 17528 575691 17552
rect 575702 17528 575774 17562
rect 575657 17518 575774 17528
rect 575429 17494 575774 17518
rect 575442 17450 575642 17494
rect 575657 17484 575681 17494
rect 575657 17460 575691 17484
rect 575702 17460 575774 17494
rect 575657 17450 575774 17460
rect 575429 17426 575774 17450
rect 575442 17382 575642 17426
rect 575657 17416 575681 17426
rect 575657 17392 575691 17416
rect 575702 17392 575774 17426
rect 575657 17382 575774 17392
rect 575429 17358 575774 17382
rect 575442 17314 575642 17358
rect 575657 17348 575681 17358
rect 575657 17324 575691 17348
rect 575702 17324 575774 17358
rect 575657 17314 575774 17324
rect 575429 17290 575774 17314
rect 575442 17278 575642 17290
rect 575453 17266 575477 17278
rect 575657 17266 575681 17290
rect 575702 17278 575774 17290
rect 576004 17278 576060 18278
rect 576076 17278 576132 18278
rect 576434 18198 576634 18278
rect 576649 18208 576683 18232
rect 576694 18208 576766 18278
rect 576649 18198 576766 18208
rect 576421 18174 576766 18198
rect 576434 18130 576634 18174
rect 576649 18164 576673 18174
rect 576649 18140 576683 18164
rect 576694 18140 576766 18174
rect 576649 18130 576766 18140
rect 576421 18106 576766 18130
rect 576434 18062 576634 18106
rect 576649 18096 576673 18106
rect 576649 18072 576683 18096
rect 576694 18072 576766 18106
rect 576649 18062 576766 18072
rect 576421 18038 576766 18062
rect 576434 17994 576634 18038
rect 576649 18028 576673 18038
rect 576649 18004 576683 18028
rect 576694 18004 576766 18038
rect 576649 17994 576766 18004
rect 576421 17970 576766 17994
rect 576434 17926 576634 17970
rect 576649 17960 576673 17970
rect 576649 17936 576683 17960
rect 576694 17936 576766 17970
rect 576649 17926 576766 17936
rect 576421 17902 576766 17926
rect 576434 17858 576634 17902
rect 576649 17892 576673 17902
rect 576649 17868 576683 17892
rect 576694 17868 576766 17902
rect 576649 17858 576766 17868
rect 576421 17834 576766 17858
rect 576434 17790 576634 17834
rect 576649 17824 576673 17834
rect 576649 17800 576683 17824
rect 576694 17800 576766 17834
rect 576649 17790 576766 17800
rect 576421 17766 576766 17790
rect 576434 17722 576634 17766
rect 576649 17756 576673 17766
rect 576649 17732 576683 17756
rect 576694 17732 576766 17766
rect 576649 17722 576766 17732
rect 576421 17698 576766 17722
rect 576434 17654 576634 17698
rect 576649 17688 576673 17698
rect 576649 17664 576683 17688
rect 576694 17664 576766 17698
rect 576649 17654 576766 17664
rect 576421 17630 576766 17654
rect 576434 17586 576634 17630
rect 576649 17620 576673 17630
rect 576649 17596 576683 17620
rect 576694 17596 576766 17630
rect 576649 17586 576766 17596
rect 576421 17562 576766 17586
rect 576434 17518 576634 17562
rect 576649 17552 576673 17562
rect 576649 17528 576683 17552
rect 576694 17528 576766 17562
rect 576649 17518 576766 17528
rect 576421 17494 576766 17518
rect 576434 17450 576634 17494
rect 576649 17484 576673 17494
rect 576649 17460 576683 17484
rect 576694 17460 576766 17494
rect 576649 17450 576766 17460
rect 576421 17426 576766 17450
rect 576434 17382 576634 17426
rect 576649 17416 576673 17426
rect 576649 17392 576683 17416
rect 576694 17392 576766 17426
rect 576649 17382 576766 17392
rect 576421 17358 576766 17382
rect 576434 17314 576634 17358
rect 576649 17348 576673 17358
rect 576649 17324 576683 17348
rect 576694 17324 576766 17358
rect 576649 17314 576766 17324
rect 576421 17290 576766 17314
rect 576434 17278 576634 17290
rect 576445 17266 576469 17278
rect 576649 17266 576673 17290
rect 576694 17278 576766 17290
rect 576996 17278 577052 18278
rect 577068 17278 577124 18278
rect 577426 18198 577626 18278
rect 577641 18208 577675 18232
rect 577686 18208 577758 18278
rect 577641 18198 577758 18208
rect 577413 18174 577758 18198
rect 577426 18130 577626 18174
rect 577641 18164 577665 18174
rect 577641 18140 577675 18164
rect 577686 18140 577758 18174
rect 577641 18130 577758 18140
rect 577413 18106 577758 18130
rect 577426 18062 577626 18106
rect 577641 18096 577665 18106
rect 577641 18072 577675 18096
rect 577686 18072 577758 18106
rect 577641 18062 577758 18072
rect 577413 18038 577758 18062
rect 577426 17994 577626 18038
rect 577641 18028 577665 18038
rect 577641 18004 577675 18028
rect 577686 18004 577758 18038
rect 577641 17994 577758 18004
rect 577413 17970 577758 17994
rect 577426 17926 577626 17970
rect 577641 17960 577665 17970
rect 577641 17936 577675 17960
rect 577686 17936 577758 17970
rect 577641 17926 577758 17936
rect 577413 17902 577758 17926
rect 577426 17858 577626 17902
rect 577641 17892 577665 17902
rect 577641 17868 577675 17892
rect 577686 17868 577758 17902
rect 577641 17858 577758 17868
rect 577413 17834 577758 17858
rect 577426 17790 577626 17834
rect 577641 17824 577665 17834
rect 577641 17800 577675 17824
rect 577686 17800 577758 17834
rect 577641 17790 577758 17800
rect 577413 17766 577758 17790
rect 577426 17722 577626 17766
rect 577641 17756 577665 17766
rect 577641 17732 577675 17756
rect 577686 17732 577758 17766
rect 577641 17722 577758 17732
rect 577413 17698 577758 17722
rect 577426 17654 577626 17698
rect 577641 17688 577665 17698
rect 577641 17664 577675 17688
rect 577686 17664 577758 17698
rect 577641 17654 577758 17664
rect 577413 17630 577758 17654
rect 577426 17586 577626 17630
rect 577641 17620 577665 17630
rect 577641 17596 577675 17620
rect 577686 17596 577758 17630
rect 577641 17586 577758 17596
rect 577413 17562 577758 17586
rect 577426 17518 577626 17562
rect 577641 17552 577665 17562
rect 577641 17528 577675 17552
rect 577686 17528 577758 17562
rect 577641 17518 577758 17528
rect 577413 17494 577758 17518
rect 577426 17450 577626 17494
rect 577641 17484 577665 17494
rect 577641 17460 577675 17484
rect 577686 17460 577758 17494
rect 577641 17450 577758 17460
rect 577413 17426 577758 17450
rect 577426 17382 577626 17426
rect 577641 17416 577665 17426
rect 577641 17392 577675 17416
rect 577686 17392 577758 17426
rect 577641 17382 577758 17392
rect 577413 17358 577758 17382
rect 577426 17314 577626 17358
rect 577641 17348 577665 17358
rect 577641 17324 577675 17348
rect 577686 17324 577758 17358
rect 577641 17314 577758 17324
rect 577413 17290 577758 17314
rect 577426 17278 577626 17290
rect 577437 17266 577461 17278
rect 577641 17266 577665 17290
rect 577686 17278 577758 17290
rect 577988 17278 578044 18278
rect 578060 17278 578116 18278
rect 578327 17278 578377 18278
rect 565533 16678 565567 16690
rect 564746 15878 564780 15908
rect 564708 15840 564780 15870
rect 564903 15678 564936 16678
rect 565106 15678 565123 16678
rect 565261 15678 565333 16678
rect 565522 16656 565722 16678
rect 565737 16666 565771 16690
rect 566525 16678 566559 16690
rect 565782 16666 565854 16678
rect 565737 16656 565854 16666
rect 565509 16632 565854 16656
rect 565522 16588 565722 16632
rect 565737 16622 565761 16632
rect 565737 16598 565771 16622
rect 565782 16598 565854 16632
rect 565737 16588 565854 16598
rect 565509 16564 565854 16588
rect 565522 16520 565722 16564
rect 565737 16554 565761 16564
rect 565737 16530 565771 16554
rect 565782 16530 565854 16564
rect 565737 16520 565854 16530
rect 565509 16496 565854 16520
rect 565522 16452 565722 16496
rect 565737 16486 565761 16496
rect 565737 16462 565771 16486
rect 565782 16462 565854 16496
rect 565737 16452 565854 16462
rect 565509 16428 565854 16452
rect 565522 16384 565722 16428
rect 565737 16418 565761 16428
rect 565737 16394 565771 16418
rect 565782 16394 565854 16428
rect 565737 16384 565854 16394
rect 565509 16360 565854 16384
rect 565522 16316 565722 16360
rect 565737 16350 565761 16360
rect 565737 16326 565771 16350
rect 565782 16326 565854 16360
rect 565737 16316 565854 16326
rect 565509 16292 565854 16316
rect 565522 16248 565722 16292
rect 565737 16282 565761 16292
rect 565737 16258 565771 16282
rect 565782 16258 565854 16292
rect 565737 16248 565854 16258
rect 565509 16224 565854 16248
rect 565522 16180 565722 16224
rect 565737 16214 565761 16224
rect 565737 16190 565771 16214
rect 565782 16190 565854 16224
rect 565737 16180 565854 16190
rect 565509 16156 565854 16180
rect 565522 16112 565722 16156
rect 565737 16146 565761 16156
rect 565737 16122 565771 16146
rect 565782 16122 565854 16156
rect 565737 16112 565854 16122
rect 565509 16088 565854 16112
rect 565522 16044 565722 16088
rect 565737 16078 565761 16088
rect 565737 16054 565771 16078
rect 565782 16054 565854 16088
rect 565737 16044 565854 16054
rect 565509 16020 565854 16044
rect 565522 15976 565722 16020
rect 565737 16010 565761 16020
rect 565737 15986 565771 16010
rect 565782 15986 565854 16020
rect 565737 15976 565854 15986
rect 565509 15952 565854 15976
rect 565522 15908 565722 15952
rect 565737 15942 565761 15952
rect 565737 15918 565771 15942
rect 565782 15918 565854 15952
rect 565737 15908 565854 15918
rect 565509 15884 565854 15908
rect 565522 15840 565722 15884
rect 565737 15874 565761 15884
rect 565737 15850 565771 15874
rect 565782 15850 565854 15884
rect 565737 15840 565854 15850
rect 565509 15816 565854 15840
rect 565522 15772 565722 15816
rect 565737 15806 565761 15816
rect 565737 15782 565771 15806
rect 565782 15782 565854 15816
rect 565737 15772 565854 15782
rect 565509 15748 565854 15772
rect 565522 15678 565722 15748
rect 565737 15724 565761 15748
rect 565782 15678 565854 15748
rect 566084 15678 566140 16678
rect 566156 15678 566212 16678
rect 566514 16656 566714 16678
rect 566729 16666 566763 16690
rect 567517 16678 567551 16690
rect 566774 16666 566846 16678
rect 566729 16656 566846 16666
rect 566501 16632 566846 16656
rect 566514 16588 566714 16632
rect 566729 16622 566753 16632
rect 566729 16598 566763 16622
rect 566774 16598 566846 16632
rect 566729 16588 566846 16598
rect 566501 16564 566846 16588
rect 566514 16520 566714 16564
rect 566729 16554 566753 16564
rect 566729 16530 566763 16554
rect 566774 16530 566846 16564
rect 566729 16520 566846 16530
rect 566501 16496 566846 16520
rect 566514 16452 566714 16496
rect 566729 16486 566753 16496
rect 566729 16462 566763 16486
rect 566774 16462 566846 16496
rect 566729 16452 566846 16462
rect 566501 16428 566846 16452
rect 566514 16384 566714 16428
rect 566729 16418 566753 16428
rect 566729 16394 566763 16418
rect 566774 16394 566846 16428
rect 566729 16384 566846 16394
rect 566501 16360 566846 16384
rect 566514 16316 566714 16360
rect 566729 16350 566753 16360
rect 566729 16326 566763 16350
rect 566774 16326 566846 16360
rect 566729 16316 566846 16326
rect 566501 16292 566846 16316
rect 566514 16248 566714 16292
rect 566729 16282 566753 16292
rect 566729 16258 566763 16282
rect 566774 16258 566846 16292
rect 566729 16248 566846 16258
rect 566501 16224 566846 16248
rect 566514 16180 566714 16224
rect 566729 16214 566753 16224
rect 566729 16190 566763 16214
rect 566774 16190 566846 16224
rect 566729 16180 566846 16190
rect 566501 16156 566846 16180
rect 566514 16112 566714 16156
rect 566729 16146 566753 16156
rect 566729 16122 566763 16146
rect 566774 16122 566846 16156
rect 566729 16112 566846 16122
rect 566501 16088 566846 16112
rect 566514 16044 566714 16088
rect 566729 16078 566753 16088
rect 566729 16054 566763 16078
rect 566774 16054 566846 16088
rect 566729 16044 566846 16054
rect 566501 16020 566846 16044
rect 566514 15976 566714 16020
rect 566729 16010 566753 16020
rect 566729 15986 566763 16010
rect 566774 15986 566846 16020
rect 566729 15976 566846 15986
rect 566501 15952 566846 15976
rect 566514 15908 566714 15952
rect 566729 15942 566753 15952
rect 566729 15918 566763 15942
rect 566774 15918 566846 15952
rect 566729 15908 566846 15918
rect 566501 15884 566846 15908
rect 566514 15840 566714 15884
rect 566729 15874 566753 15884
rect 566729 15850 566763 15874
rect 566774 15850 566846 15884
rect 566729 15840 566846 15850
rect 566501 15816 566846 15840
rect 566514 15772 566714 15816
rect 566729 15806 566753 15816
rect 566729 15782 566763 15806
rect 566774 15782 566846 15816
rect 566729 15772 566846 15782
rect 566501 15748 566846 15772
rect 566514 15678 566714 15748
rect 566729 15724 566753 15748
rect 566774 15678 566846 15748
rect 567076 15678 567132 16678
rect 567148 15678 567204 16678
rect 567506 16656 567706 16678
rect 567721 16666 567755 16690
rect 568509 16678 568543 16690
rect 567766 16666 567838 16678
rect 567721 16656 567838 16666
rect 567493 16632 567838 16656
rect 567506 16588 567706 16632
rect 567721 16622 567745 16632
rect 567721 16598 567755 16622
rect 567766 16598 567838 16632
rect 567721 16588 567838 16598
rect 567493 16564 567838 16588
rect 567506 16520 567706 16564
rect 567721 16554 567745 16564
rect 567721 16530 567755 16554
rect 567766 16530 567838 16564
rect 567721 16520 567838 16530
rect 567493 16496 567838 16520
rect 567506 16452 567706 16496
rect 567721 16486 567745 16496
rect 567721 16462 567755 16486
rect 567766 16462 567838 16496
rect 567721 16452 567838 16462
rect 567493 16428 567838 16452
rect 567506 16384 567706 16428
rect 567721 16418 567745 16428
rect 567721 16394 567755 16418
rect 567766 16394 567838 16428
rect 567721 16384 567838 16394
rect 567493 16360 567838 16384
rect 567506 16316 567706 16360
rect 567721 16350 567745 16360
rect 567721 16326 567755 16350
rect 567766 16326 567838 16360
rect 567721 16316 567838 16326
rect 567493 16292 567838 16316
rect 567506 16248 567706 16292
rect 567721 16282 567745 16292
rect 567721 16258 567755 16282
rect 567766 16258 567838 16292
rect 567721 16248 567838 16258
rect 567493 16224 567838 16248
rect 567506 16180 567706 16224
rect 567721 16214 567745 16224
rect 567721 16190 567755 16214
rect 567766 16190 567838 16224
rect 567721 16180 567838 16190
rect 567493 16156 567838 16180
rect 567506 16112 567706 16156
rect 567721 16146 567745 16156
rect 567721 16122 567755 16146
rect 567766 16122 567838 16156
rect 567721 16112 567838 16122
rect 567493 16088 567838 16112
rect 567506 16044 567706 16088
rect 567721 16078 567745 16088
rect 567721 16054 567755 16078
rect 567766 16054 567838 16088
rect 567721 16044 567838 16054
rect 567493 16020 567838 16044
rect 567506 15976 567706 16020
rect 567721 16010 567745 16020
rect 567721 15986 567755 16010
rect 567766 15986 567838 16020
rect 567721 15976 567838 15986
rect 567493 15952 567838 15976
rect 567506 15908 567706 15952
rect 567721 15942 567745 15952
rect 567721 15918 567755 15942
rect 567766 15918 567838 15952
rect 567721 15908 567838 15918
rect 567493 15884 567838 15908
rect 567506 15840 567706 15884
rect 567721 15874 567745 15884
rect 567721 15850 567755 15874
rect 567766 15850 567838 15884
rect 567721 15840 567838 15850
rect 567493 15816 567838 15840
rect 567506 15772 567706 15816
rect 567721 15806 567745 15816
rect 567721 15782 567755 15806
rect 567766 15782 567838 15816
rect 567721 15772 567838 15782
rect 567493 15748 567838 15772
rect 567506 15678 567706 15748
rect 567721 15724 567745 15748
rect 567766 15678 567838 15748
rect 568068 15678 568124 16678
rect 568140 15678 568196 16678
rect 568498 16656 568698 16678
rect 568713 16666 568747 16690
rect 569501 16678 569535 16690
rect 568758 16666 568830 16678
rect 568713 16656 568830 16666
rect 568485 16632 568830 16656
rect 568498 16588 568698 16632
rect 568713 16622 568737 16632
rect 568713 16598 568747 16622
rect 568758 16598 568830 16632
rect 568713 16588 568830 16598
rect 568485 16564 568830 16588
rect 568498 16520 568698 16564
rect 568713 16554 568737 16564
rect 568713 16530 568747 16554
rect 568758 16530 568830 16564
rect 568713 16520 568830 16530
rect 568485 16496 568830 16520
rect 568498 16452 568698 16496
rect 568713 16486 568737 16496
rect 568713 16462 568747 16486
rect 568758 16462 568830 16496
rect 568713 16452 568830 16462
rect 568485 16428 568830 16452
rect 568498 16384 568698 16428
rect 568713 16418 568737 16428
rect 568713 16394 568747 16418
rect 568758 16394 568830 16428
rect 568713 16384 568830 16394
rect 568485 16360 568830 16384
rect 568498 16316 568698 16360
rect 568713 16350 568737 16360
rect 568713 16326 568747 16350
rect 568758 16326 568830 16360
rect 568713 16316 568830 16326
rect 568485 16292 568830 16316
rect 568498 16248 568698 16292
rect 568713 16282 568737 16292
rect 568713 16258 568747 16282
rect 568758 16258 568830 16292
rect 568713 16248 568830 16258
rect 568485 16224 568830 16248
rect 568498 16180 568698 16224
rect 568713 16214 568737 16224
rect 568713 16190 568747 16214
rect 568758 16190 568830 16224
rect 568713 16180 568830 16190
rect 568485 16156 568830 16180
rect 568498 16112 568698 16156
rect 568713 16146 568737 16156
rect 568713 16122 568747 16146
rect 568758 16122 568830 16156
rect 568713 16112 568830 16122
rect 568485 16088 568830 16112
rect 568498 16044 568698 16088
rect 568713 16078 568737 16088
rect 568713 16054 568747 16078
rect 568758 16054 568830 16088
rect 568713 16044 568830 16054
rect 568485 16020 568830 16044
rect 568498 15976 568698 16020
rect 568713 16010 568737 16020
rect 568713 15986 568747 16010
rect 568758 15986 568830 16020
rect 568713 15976 568830 15986
rect 568485 15952 568830 15976
rect 568498 15908 568698 15952
rect 568713 15942 568737 15952
rect 568713 15918 568747 15942
rect 568758 15918 568830 15952
rect 568713 15908 568830 15918
rect 568485 15884 568830 15908
rect 568498 15840 568698 15884
rect 568713 15874 568737 15884
rect 568713 15850 568747 15874
rect 568758 15850 568830 15884
rect 568713 15840 568830 15850
rect 568485 15816 568830 15840
rect 568498 15772 568698 15816
rect 568713 15806 568737 15816
rect 568713 15782 568747 15806
rect 568758 15782 568830 15816
rect 568713 15772 568830 15782
rect 568485 15748 568830 15772
rect 568498 15678 568698 15748
rect 568713 15724 568737 15748
rect 568758 15678 568830 15748
rect 569060 15678 569116 16678
rect 569132 15678 569188 16678
rect 569490 16656 569690 16678
rect 569705 16666 569739 16690
rect 570493 16678 570527 16690
rect 569750 16666 569822 16678
rect 569705 16656 569822 16666
rect 569477 16632 569822 16656
rect 569490 16588 569690 16632
rect 569705 16622 569729 16632
rect 569705 16598 569739 16622
rect 569750 16598 569822 16632
rect 569705 16588 569822 16598
rect 569477 16564 569822 16588
rect 569490 16520 569690 16564
rect 569705 16554 569729 16564
rect 569705 16530 569739 16554
rect 569750 16530 569822 16564
rect 569705 16520 569822 16530
rect 569477 16496 569822 16520
rect 569490 16452 569690 16496
rect 569705 16486 569729 16496
rect 569705 16462 569739 16486
rect 569750 16462 569822 16496
rect 569705 16452 569822 16462
rect 569477 16428 569822 16452
rect 569490 16384 569690 16428
rect 569705 16418 569729 16428
rect 569705 16394 569739 16418
rect 569750 16394 569822 16428
rect 569705 16384 569822 16394
rect 569477 16360 569822 16384
rect 569490 16316 569690 16360
rect 569705 16350 569729 16360
rect 569705 16326 569739 16350
rect 569750 16326 569822 16360
rect 569705 16316 569822 16326
rect 569477 16292 569822 16316
rect 569490 16248 569690 16292
rect 569705 16282 569729 16292
rect 569705 16258 569739 16282
rect 569750 16258 569822 16292
rect 569705 16248 569822 16258
rect 569477 16224 569822 16248
rect 569490 16180 569690 16224
rect 569705 16214 569729 16224
rect 569705 16190 569739 16214
rect 569750 16190 569822 16224
rect 569705 16180 569822 16190
rect 569477 16156 569822 16180
rect 569490 16112 569690 16156
rect 569705 16146 569729 16156
rect 569705 16122 569739 16146
rect 569750 16122 569822 16156
rect 569705 16112 569822 16122
rect 569477 16088 569822 16112
rect 569490 16044 569690 16088
rect 569705 16078 569729 16088
rect 569705 16054 569739 16078
rect 569750 16054 569822 16088
rect 569705 16044 569822 16054
rect 569477 16020 569822 16044
rect 569490 15976 569690 16020
rect 569705 16010 569729 16020
rect 569705 15986 569739 16010
rect 569750 15986 569822 16020
rect 569705 15976 569822 15986
rect 569477 15952 569822 15976
rect 569490 15908 569690 15952
rect 569705 15942 569729 15952
rect 569705 15918 569739 15942
rect 569750 15918 569822 15952
rect 569705 15908 569822 15918
rect 569477 15884 569822 15908
rect 569490 15840 569690 15884
rect 569705 15874 569729 15884
rect 569705 15850 569739 15874
rect 569750 15850 569822 15884
rect 569705 15840 569822 15850
rect 569477 15816 569822 15840
rect 569490 15772 569690 15816
rect 569705 15806 569729 15816
rect 569705 15782 569739 15806
rect 569750 15782 569822 15816
rect 569705 15772 569822 15782
rect 569477 15748 569822 15772
rect 569490 15678 569690 15748
rect 569705 15724 569729 15748
rect 569750 15678 569822 15748
rect 570052 15678 570108 16678
rect 570124 15678 570180 16678
rect 570482 16656 570682 16678
rect 570697 16666 570731 16690
rect 571485 16678 571519 16690
rect 570742 16666 570814 16678
rect 570697 16656 570814 16666
rect 570469 16632 570814 16656
rect 570482 16588 570682 16632
rect 570697 16622 570721 16632
rect 570697 16598 570731 16622
rect 570742 16598 570814 16632
rect 570697 16588 570814 16598
rect 570469 16564 570814 16588
rect 570482 16520 570682 16564
rect 570697 16554 570721 16564
rect 570697 16530 570731 16554
rect 570742 16530 570814 16564
rect 570697 16520 570814 16530
rect 570469 16496 570814 16520
rect 570482 16452 570682 16496
rect 570697 16486 570721 16496
rect 570697 16462 570731 16486
rect 570742 16462 570814 16496
rect 570697 16452 570814 16462
rect 570469 16428 570814 16452
rect 570482 16384 570682 16428
rect 570697 16418 570721 16428
rect 570697 16394 570731 16418
rect 570742 16394 570814 16428
rect 570697 16384 570814 16394
rect 570469 16360 570814 16384
rect 570482 16316 570682 16360
rect 570697 16350 570721 16360
rect 570697 16326 570731 16350
rect 570742 16326 570814 16360
rect 570697 16316 570814 16326
rect 570469 16292 570814 16316
rect 570482 16248 570682 16292
rect 570697 16282 570721 16292
rect 570697 16258 570731 16282
rect 570742 16258 570814 16292
rect 570697 16248 570814 16258
rect 570469 16224 570814 16248
rect 570482 16180 570682 16224
rect 570697 16214 570721 16224
rect 570697 16190 570731 16214
rect 570742 16190 570814 16224
rect 570697 16180 570814 16190
rect 570469 16156 570814 16180
rect 570482 16112 570682 16156
rect 570697 16146 570721 16156
rect 570697 16122 570731 16146
rect 570742 16122 570814 16156
rect 570697 16112 570814 16122
rect 570469 16088 570814 16112
rect 570482 16044 570682 16088
rect 570697 16078 570721 16088
rect 570697 16054 570731 16078
rect 570742 16054 570814 16088
rect 570697 16044 570814 16054
rect 570469 16020 570814 16044
rect 570482 15976 570682 16020
rect 570697 16010 570721 16020
rect 570697 15986 570731 16010
rect 570742 15986 570814 16020
rect 570697 15976 570814 15986
rect 570469 15952 570814 15976
rect 570482 15908 570682 15952
rect 570697 15942 570721 15952
rect 570697 15918 570731 15942
rect 570742 15918 570814 15952
rect 570697 15908 570814 15918
rect 570469 15884 570814 15908
rect 570482 15840 570682 15884
rect 570697 15874 570721 15884
rect 570697 15850 570731 15874
rect 570742 15850 570814 15884
rect 570697 15840 570814 15850
rect 570469 15816 570814 15840
rect 570482 15772 570682 15816
rect 570697 15806 570721 15816
rect 570697 15782 570731 15806
rect 570742 15782 570814 15816
rect 570697 15772 570814 15782
rect 570469 15748 570814 15772
rect 570482 15678 570682 15748
rect 570697 15724 570721 15748
rect 570742 15678 570814 15748
rect 571044 15678 571100 16678
rect 571116 15678 571172 16678
rect 571474 16656 571674 16678
rect 571689 16666 571723 16690
rect 572477 16678 572511 16690
rect 571734 16666 571806 16678
rect 571689 16656 571806 16666
rect 571461 16632 571806 16656
rect 571474 16588 571674 16632
rect 571689 16622 571713 16632
rect 571689 16598 571723 16622
rect 571734 16598 571806 16632
rect 571689 16588 571806 16598
rect 571461 16564 571806 16588
rect 571474 16520 571674 16564
rect 571689 16554 571713 16564
rect 571689 16530 571723 16554
rect 571734 16530 571806 16564
rect 571689 16520 571806 16530
rect 571461 16496 571806 16520
rect 571474 16452 571674 16496
rect 571689 16486 571713 16496
rect 571689 16462 571723 16486
rect 571734 16462 571806 16496
rect 571689 16452 571806 16462
rect 571461 16428 571806 16452
rect 571474 16384 571674 16428
rect 571689 16418 571713 16428
rect 571689 16394 571723 16418
rect 571734 16394 571806 16428
rect 571689 16384 571806 16394
rect 571461 16360 571806 16384
rect 571474 16316 571674 16360
rect 571689 16350 571713 16360
rect 571689 16326 571723 16350
rect 571734 16326 571806 16360
rect 571689 16316 571806 16326
rect 571461 16292 571806 16316
rect 571474 16248 571674 16292
rect 571689 16282 571713 16292
rect 571689 16258 571723 16282
rect 571734 16258 571806 16292
rect 571689 16248 571806 16258
rect 571461 16224 571806 16248
rect 571474 16180 571674 16224
rect 571689 16214 571713 16224
rect 571689 16190 571723 16214
rect 571734 16190 571806 16224
rect 571689 16180 571806 16190
rect 571461 16156 571806 16180
rect 571474 16112 571674 16156
rect 571689 16146 571713 16156
rect 571689 16122 571723 16146
rect 571734 16122 571806 16156
rect 571689 16112 571806 16122
rect 571461 16088 571806 16112
rect 571474 16044 571674 16088
rect 571689 16078 571713 16088
rect 571689 16054 571723 16078
rect 571734 16054 571806 16088
rect 571689 16044 571806 16054
rect 571461 16020 571806 16044
rect 571474 15976 571674 16020
rect 571689 16010 571713 16020
rect 571689 15986 571723 16010
rect 571734 15986 571806 16020
rect 571689 15976 571806 15986
rect 571461 15952 571806 15976
rect 571474 15908 571674 15952
rect 571689 15942 571713 15952
rect 571689 15918 571723 15942
rect 571734 15918 571806 15952
rect 571689 15908 571806 15918
rect 571461 15884 571806 15908
rect 571474 15840 571674 15884
rect 571689 15874 571713 15884
rect 571689 15850 571723 15874
rect 571734 15850 571806 15884
rect 571689 15840 571806 15850
rect 571461 15816 571806 15840
rect 571474 15772 571674 15816
rect 571689 15806 571713 15816
rect 571689 15782 571723 15806
rect 571734 15782 571806 15816
rect 571689 15772 571806 15782
rect 571461 15748 571806 15772
rect 571474 15678 571674 15748
rect 571689 15724 571713 15748
rect 571734 15678 571806 15748
rect 572036 15678 572092 16678
rect 572108 15678 572164 16678
rect 572466 16656 572666 16678
rect 572681 16666 572715 16690
rect 573469 16678 573503 16690
rect 572726 16666 572798 16678
rect 572681 16656 572798 16666
rect 572453 16632 572798 16656
rect 572466 16588 572666 16632
rect 572681 16622 572705 16632
rect 572681 16598 572715 16622
rect 572726 16598 572798 16632
rect 572681 16588 572798 16598
rect 572453 16564 572798 16588
rect 572466 16520 572666 16564
rect 572681 16554 572705 16564
rect 572681 16530 572715 16554
rect 572726 16530 572798 16564
rect 572681 16520 572798 16530
rect 572453 16496 572798 16520
rect 572466 16452 572666 16496
rect 572681 16486 572705 16496
rect 572681 16462 572715 16486
rect 572726 16462 572798 16496
rect 572681 16452 572798 16462
rect 572453 16428 572798 16452
rect 572466 16384 572666 16428
rect 572681 16418 572705 16428
rect 572681 16394 572715 16418
rect 572726 16394 572798 16428
rect 572681 16384 572798 16394
rect 572453 16360 572798 16384
rect 572466 16316 572666 16360
rect 572681 16350 572705 16360
rect 572681 16326 572715 16350
rect 572726 16326 572798 16360
rect 572681 16316 572798 16326
rect 572453 16292 572798 16316
rect 572466 16248 572666 16292
rect 572681 16282 572705 16292
rect 572681 16258 572715 16282
rect 572726 16258 572798 16292
rect 572681 16248 572798 16258
rect 572453 16224 572798 16248
rect 572466 16180 572666 16224
rect 572681 16214 572705 16224
rect 572681 16190 572715 16214
rect 572726 16190 572798 16224
rect 572681 16180 572798 16190
rect 572453 16156 572798 16180
rect 572466 16112 572666 16156
rect 572681 16146 572705 16156
rect 572681 16122 572715 16146
rect 572726 16122 572798 16156
rect 572681 16112 572798 16122
rect 572453 16088 572798 16112
rect 572466 16044 572666 16088
rect 572681 16078 572705 16088
rect 572681 16054 572715 16078
rect 572726 16054 572798 16088
rect 572681 16044 572798 16054
rect 572453 16020 572798 16044
rect 572466 15976 572666 16020
rect 572681 16010 572705 16020
rect 572681 15986 572715 16010
rect 572726 15986 572798 16020
rect 572681 15976 572798 15986
rect 572453 15952 572798 15976
rect 572466 15908 572666 15952
rect 572681 15942 572705 15952
rect 572681 15918 572715 15942
rect 572726 15918 572798 15952
rect 572681 15908 572798 15918
rect 572453 15884 572798 15908
rect 572466 15840 572666 15884
rect 572681 15874 572705 15884
rect 572681 15850 572715 15874
rect 572726 15850 572798 15884
rect 572681 15840 572798 15850
rect 572453 15816 572798 15840
rect 572466 15772 572666 15816
rect 572681 15806 572705 15816
rect 572681 15782 572715 15806
rect 572726 15782 572798 15816
rect 572681 15772 572798 15782
rect 572453 15748 572798 15772
rect 572466 15678 572666 15748
rect 572681 15724 572705 15748
rect 572726 15678 572798 15748
rect 573028 15678 573084 16678
rect 573100 15678 573156 16678
rect 573458 16656 573658 16678
rect 573673 16666 573707 16690
rect 574461 16678 574495 16690
rect 573718 16666 573790 16678
rect 573673 16656 573790 16666
rect 573445 16632 573790 16656
rect 573458 16588 573658 16632
rect 573673 16622 573697 16632
rect 573673 16598 573707 16622
rect 573718 16598 573790 16632
rect 573673 16588 573790 16598
rect 573445 16564 573790 16588
rect 573458 16520 573658 16564
rect 573673 16554 573697 16564
rect 573673 16530 573707 16554
rect 573718 16530 573790 16564
rect 573673 16520 573790 16530
rect 573445 16496 573790 16520
rect 573458 16452 573658 16496
rect 573673 16486 573697 16496
rect 573673 16462 573707 16486
rect 573718 16462 573790 16496
rect 573673 16452 573790 16462
rect 573445 16428 573790 16452
rect 573458 16384 573658 16428
rect 573673 16418 573697 16428
rect 573673 16394 573707 16418
rect 573718 16394 573790 16428
rect 573673 16384 573790 16394
rect 573445 16360 573790 16384
rect 573458 16316 573658 16360
rect 573673 16350 573697 16360
rect 573673 16326 573707 16350
rect 573718 16326 573790 16360
rect 573673 16316 573790 16326
rect 573445 16292 573790 16316
rect 573458 16248 573658 16292
rect 573673 16282 573697 16292
rect 573673 16258 573707 16282
rect 573718 16258 573790 16292
rect 573673 16248 573790 16258
rect 573445 16224 573790 16248
rect 573458 16180 573658 16224
rect 573673 16214 573697 16224
rect 573673 16190 573707 16214
rect 573718 16190 573790 16224
rect 573673 16180 573790 16190
rect 573445 16156 573790 16180
rect 573458 16112 573658 16156
rect 573673 16146 573697 16156
rect 573673 16122 573707 16146
rect 573718 16122 573790 16156
rect 573673 16112 573790 16122
rect 573445 16088 573790 16112
rect 573458 16044 573658 16088
rect 573673 16078 573697 16088
rect 573673 16054 573707 16078
rect 573718 16054 573790 16088
rect 573673 16044 573790 16054
rect 573445 16020 573790 16044
rect 573458 15976 573658 16020
rect 573673 16010 573697 16020
rect 573673 15986 573707 16010
rect 573718 15986 573790 16020
rect 573673 15976 573790 15986
rect 573445 15952 573790 15976
rect 573458 15908 573658 15952
rect 573673 15942 573697 15952
rect 573673 15918 573707 15942
rect 573718 15918 573790 15952
rect 573673 15908 573790 15918
rect 573445 15884 573790 15908
rect 573458 15840 573658 15884
rect 573673 15874 573697 15884
rect 573673 15850 573707 15874
rect 573718 15850 573790 15884
rect 573673 15840 573790 15850
rect 573445 15816 573790 15840
rect 573458 15772 573658 15816
rect 573673 15806 573697 15816
rect 573673 15782 573707 15806
rect 573718 15782 573790 15816
rect 573673 15772 573790 15782
rect 573445 15748 573790 15772
rect 573458 15678 573658 15748
rect 573673 15724 573697 15748
rect 573718 15678 573790 15748
rect 574020 15678 574076 16678
rect 574092 15678 574148 16678
rect 574450 16656 574650 16678
rect 574665 16666 574699 16690
rect 575453 16678 575487 16690
rect 574710 16666 574782 16678
rect 574665 16656 574782 16666
rect 574437 16632 574782 16656
rect 574450 16588 574650 16632
rect 574665 16622 574689 16632
rect 574665 16598 574699 16622
rect 574710 16598 574782 16632
rect 574665 16588 574782 16598
rect 574437 16564 574782 16588
rect 574450 16520 574650 16564
rect 574665 16554 574689 16564
rect 574665 16530 574699 16554
rect 574710 16530 574782 16564
rect 574665 16520 574782 16530
rect 574437 16496 574782 16520
rect 574450 16452 574650 16496
rect 574665 16486 574689 16496
rect 574665 16462 574699 16486
rect 574710 16462 574782 16496
rect 574665 16452 574782 16462
rect 574437 16428 574782 16452
rect 574450 16384 574650 16428
rect 574665 16418 574689 16428
rect 574665 16394 574699 16418
rect 574710 16394 574782 16428
rect 574665 16384 574782 16394
rect 574437 16360 574782 16384
rect 574450 16316 574650 16360
rect 574665 16350 574689 16360
rect 574665 16326 574699 16350
rect 574710 16326 574782 16360
rect 574665 16316 574782 16326
rect 574437 16292 574782 16316
rect 574450 16248 574650 16292
rect 574665 16282 574689 16292
rect 574665 16258 574699 16282
rect 574710 16258 574782 16292
rect 574665 16248 574782 16258
rect 574437 16224 574782 16248
rect 574450 16180 574650 16224
rect 574665 16214 574689 16224
rect 574665 16190 574699 16214
rect 574710 16190 574782 16224
rect 574665 16180 574782 16190
rect 574437 16156 574782 16180
rect 574450 16112 574650 16156
rect 574665 16146 574689 16156
rect 574665 16122 574699 16146
rect 574710 16122 574782 16156
rect 574665 16112 574782 16122
rect 574437 16088 574782 16112
rect 574450 16044 574650 16088
rect 574665 16078 574689 16088
rect 574665 16054 574699 16078
rect 574710 16054 574782 16088
rect 574665 16044 574782 16054
rect 574437 16020 574782 16044
rect 574450 15976 574650 16020
rect 574665 16010 574689 16020
rect 574665 15986 574699 16010
rect 574710 15986 574782 16020
rect 574665 15976 574782 15986
rect 574437 15952 574782 15976
rect 574450 15908 574650 15952
rect 574665 15942 574689 15952
rect 574665 15918 574699 15942
rect 574710 15918 574782 15952
rect 574665 15908 574782 15918
rect 574437 15884 574782 15908
rect 574450 15840 574650 15884
rect 574665 15874 574689 15884
rect 574665 15850 574699 15874
rect 574710 15850 574782 15884
rect 574665 15840 574782 15850
rect 574437 15816 574782 15840
rect 574450 15772 574650 15816
rect 574665 15806 574689 15816
rect 574665 15782 574699 15806
rect 574710 15782 574782 15816
rect 574665 15772 574782 15782
rect 574437 15748 574782 15772
rect 574450 15678 574650 15748
rect 574665 15724 574689 15748
rect 574710 15678 574782 15748
rect 575012 15678 575068 16678
rect 575084 15678 575140 16678
rect 575442 16656 575642 16678
rect 575657 16666 575691 16690
rect 576445 16678 576479 16690
rect 575702 16666 575774 16678
rect 575657 16656 575774 16666
rect 575429 16632 575774 16656
rect 575442 16588 575642 16632
rect 575657 16622 575681 16632
rect 575657 16598 575691 16622
rect 575702 16598 575774 16632
rect 575657 16588 575774 16598
rect 575429 16564 575774 16588
rect 575442 16520 575642 16564
rect 575657 16554 575681 16564
rect 575657 16530 575691 16554
rect 575702 16530 575774 16564
rect 575657 16520 575774 16530
rect 575429 16496 575774 16520
rect 575442 16452 575642 16496
rect 575657 16486 575681 16496
rect 575657 16462 575691 16486
rect 575702 16462 575774 16496
rect 575657 16452 575774 16462
rect 575429 16428 575774 16452
rect 575442 16384 575642 16428
rect 575657 16418 575681 16428
rect 575657 16394 575691 16418
rect 575702 16394 575774 16428
rect 575657 16384 575774 16394
rect 575429 16360 575774 16384
rect 575442 16316 575642 16360
rect 575657 16350 575681 16360
rect 575657 16326 575691 16350
rect 575702 16326 575774 16360
rect 575657 16316 575774 16326
rect 575429 16292 575774 16316
rect 575442 16248 575642 16292
rect 575657 16282 575681 16292
rect 575657 16258 575691 16282
rect 575702 16258 575774 16292
rect 575657 16248 575774 16258
rect 575429 16224 575774 16248
rect 575442 16180 575642 16224
rect 575657 16214 575681 16224
rect 575657 16190 575691 16214
rect 575702 16190 575774 16224
rect 575657 16180 575774 16190
rect 575429 16156 575774 16180
rect 575442 16112 575642 16156
rect 575657 16146 575681 16156
rect 575657 16122 575691 16146
rect 575702 16122 575774 16156
rect 575657 16112 575774 16122
rect 575429 16088 575774 16112
rect 575442 16044 575642 16088
rect 575657 16078 575681 16088
rect 575657 16054 575691 16078
rect 575702 16054 575774 16088
rect 575657 16044 575774 16054
rect 575429 16020 575774 16044
rect 575442 15976 575642 16020
rect 575657 16010 575681 16020
rect 575657 15986 575691 16010
rect 575702 15986 575774 16020
rect 575657 15976 575774 15986
rect 575429 15952 575774 15976
rect 575442 15908 575642 15952
rect 575657 15942 575681 15952
rect 575657 15918 575691 15942
rect 575702 15918 575774 15952
rect 575657 15908 575774 15918
rect 575429 15884 575774 15908
rect 575442 15840 575642 15884
rect 575657 15874 575681 15884
rect 575657 15850 575691 15874
rect 575702 15850 575774 15884
rect 575657 15840 575774 15850
rect 575429 15816 575774 15840
rect 575442 15772 575642 15816
rect 575657 15806 575681 15816
rect 575657 15782 575691 15806
rect 575702 15782 575774 15816
rect 575657 15772 575774 15782
rect 575429 15748 575774 15772
rect 575442 15678 575642 15748
rect 575657 15724 575681 15748
rect 575702 15678 575774 15748
rect 576004 15678 576060 16678
rect 576076 15678 576132 16678
rect 576434 16656 576634 16678
rect 576649 16666 576683 16690
rect 577437 16678 577471 16690
rect 576694 16666 576766 16678
rect 576649 16656 576766 16666
rect 576421 16632 576766 16656
rect 576434 16588 576634 16632
rect 576649 16622 576673 16632
rect 576649 16598 576683 16622
rect 576694 16598 576766 16632
rect 576649 16588 576766 16598
rect 576421 16564 576766 16588
rect 576434 16520 576634 16564
rect 576649 16554 576673 16564
rect 576649 16530 576683 16554
rect 576694 16530 576766 16564
rect 576649 16520 576766 16530
rect 576421 16496 576766 16520
rect 576434 16452 576634 16496
rect 576649 16486 576673 16496
rect 576649 16462 576683 16486
rect 576694 16462 576766 16496
rect 576649 16452 576766 16462
rect 576421 16428 576766 16452
rect 576434 16384 576634 16428
rect 576649 16418 576673 16428
rect 576649 16394 576683 16418
rect 576694 16394 576766 16428
rect 576649 16384 576766 16394
rect 576421 16360 576766 16384
rect 576434 16316 576634 16360
rect 576649 16350 576673 16360
rect 576649 16326 576683 16350
rect 576694 16326 576766 16360
rect 576649 16316 576766 16326
rect 576421 16292 576766 16316
rect 576434 16248 576634 16292
rect 576649 16282 576673 16292
rect 576649 16258 576683 16282
rect 576694 16258 576766 16292
rect 576649 16248 576766 16258
rect 576421 16224 576766 16248
rect 576434 16180 576634 16224
rect 576649 16214 576673 16224
rect 576649 16190 576683 16214
rect 576694 16190 576766 16224
rect 576649 16180 576766 16190
rect 576421 16156 576766 16180
rect 576434 16112 576634 16156
rect 576649 16146 576673 16156
rect 576649 16122 576683 16146
rect 576694 16122 576766 16156
rect 576649 16112 576766 16122
rect 576421 16088 576766 16112
rect 576434 16044 576634 16088
rect 576649 16078 576673 16088
rect 576649 16054 576683 16078
rect 576694 16054 576766 16088
rect 576649 16044 576766 16054
rect 576421 16020 576766 16044
rect 576434 15976 576634 16020
rect 576649 16010 576673 16020
rect 576649 15986 576683 16010
rect 576694 15986 576766 16020
rect 576649 15976 576766 15986
rect 576421 15952 576766 15976
rect 576434 15908 576634 15952
rect 576649 15942 576673 15952
rect 576649 15918 576683 15942
rect 576694 15918 576766 15952
rect 576649 15908 576766 15918
rect 576421 15884 576766 15908
rect 576434 15840 576634 15884
rect 576649 15874 576673 15884
rect 576649 15850 576683 15874
rect 576694 15850 576766 15884
rect 576649 15840 576766 15850
rect 576421 15816 576766 15840
rect 576434 15772 576634 15816
rect 576649 15806 576673 15816
rect 576649 15782 576683 15806
rect 576694 15782 576766 15816
rect 576649 15772 576766 15782
rect 576421 15748 576766 15772
rect 576434 15678 576634 15748
rect 576649 15724 576673 15748
rect 576694 15678 576766 15748
rect 576996 15678 577052 16678
rect 577068 15678 577124 16678
rect 577426 16656 577626 16678
rect 577641 16666 577675 16690
rect 577686 16666 577758 16678
rect 577641 16656 577758 16666
rect 577413 16632 577758 16656
rect 577426 16588 577626 16632
rect 577641 16622 577665 16632
rect 577641 16598 577675 16622
rect 577686 16598 577758 16632
rect 577641 16588 577758 16598
rect 577413 16564 577758 16588
rect 577426 16520 577626 16564
rect 577641 16554 577665 16564
rect 577641 16530 577675 16554
rect 577686 16530 577758 16564
rect 577641 16520 577758 16530
rect 577413 16496 577758 16520
rect 577426 16452 577626 16496
rect 577641 16486 577665 16496
rect 577641 16462 577675 16486
rect 577686 16462 577758 16496
rect 577641 16452 577758 16462
rect 577413 16428 577758 16452
rect 577426 16384 577626 16428
rect 577641 16418 577665 16428
rect 577641 16394 577675 16418
rect 577686 16394 577758 16428
rect 577641 16384 577758 16394
rect 577413 16360 577758 16384
rect 577426 16316 577626 16360
rect 577641 16350 577665 16360
rect 577641 16326 577675 16350
rect 577686 16326 577758 16360
rect 577641 16316 577758 16326
rect 577413 16292 577758 16316
rect 577426 16248 577626 16292
rect 577641 16282 577665 16292
rect 577641 16258 577675 16282
rect 577686 16258 577758 16292
rect 577641 16248 577758 16258
rect 577413 16224 577758 16248
rect 577426 16180 577626 16224
rect 577641 16214 577665 16224
rect 577641 16190 577675 16214
rect 577686 16190 577758 16224
rect 577641 16180 577758 16190
rect 577413 16156 577758 16180
rect 577426 16112 577626 16156
rect 577641 16146 577665 16156
rect 577641 16122 577675 16146
rect 577686 16122 577758 16156
rect 577641 16112 577758 16122
rect 577413 16088 577758 16112
rect 577426 16044 577626 16088
rect 577641 16078 577665 16088
rect 577641 16054 577675 16078
rect 577686 16054 577758 16088
rect 577641 16044 577758 16054
rect 577413 16020 577758 16044
rect 577426 15976 577626 16020
rect 577641 16010 577665 16020
rect 577641 15986 577675 16010
rect 577686 15986 577758 16020
rect 577641 15976 577758 15986
rect 577413 15952 577758 15976
rect 577426 15908 577626 15952
rect 577641 15942 577665 15952
rect 577641 15918 577675 15942
rect 577686 15918 577758 15952
rect 577641 15908 577758 15918
rect 577413 15884 577758 15908
rect 577426 15840 577626 15884
rect 577641 15874 577665 15884
rect 577641 15850 577675 15874
rect 577686 15850 577758 15884
rect 577641 15840 577758 15850
rect 577413 15816 577758 15840
rect 577426 15772 577626 15816
rect 577641 15806 577665 15816
rect 577641 15782 577675 15806
rect 577686 15782 577758 15816
rect 577641 15772 577758 15782
rect 577413 15748 577758 15772
rect 577426 15678 577626 15748
rect 577641 15724 577665 15748
rect 577686 15678 577758 15748
rect 577988 15678 578044 16678
rect 578060 15678 578116 16678
rect 578327 15678 578377 16678
rect 579065 14844 579172 19390
rect 71017 14747 71172 14844
rect 123017 14747 123172 14844
rect 175017 14747 175172 14844
rect 227017 14747 227172 14844
rect 275017 14747 275172 14844
rect 327017 14747 327172 14844
rect 379017 14747 379172 14844
rect 427017 14747 427172 14844
rect 479017 14747 479172 14844
rect 531017 14747 531172 14844
rect 579017 14747 579172 14844
rect 71017 13955 71041 14747
rect 123017 13955 123041 14747
rect 175017 13955 175041 14747
rect 227017 13955 227041 14747
rect 275017 13955 275041 14747
rect 327017 13955 327041 14747
rect 367710 13901 367714 14061
rect 367856 13899 367860 14059
rect 369052 13899 369056 14059
rect 369198 13899 369202 14059
rect 379017 13955 379041 14747
rect 427017 13955 427041 14747
rect 467710 13901 467714 14061
rect 467856 13899 467860 14059
rect 469052 13899 469056 14059
rect 469198 13899 469202 14059
rect 479017 13955 479041 14747
rect 531017 13955 531041 14747
rect 567710 13901 567714 14061
rect 567856 13899 567860 14059
rect 569052 13899 569056 14059
rect 569198 13899 569202 14059
rect 579017 13955 579041 14747
rect 368269 12865 368285 12881
rect 368167 12559 368285 12865
rect 368269 12543 368285 12559
rect 370457 12865 370473 12881
rect 468269 12865 468285 12881
rect 370457 12559 370575 12865
rect 468167 12559 468285 12865
rect 370457 12543 370473 12559
rect 468269 12543 468285 12559
rect 470457 12865 470473 12881
rect 568269 12865 568285 12881
rect 470457 12559 470575 12865
rect 568167 12559 568285 12865
rect 470457 12543 470473 12559
rect 568269 12543 568285 12559
rect 570457 12865 570473 12881
rect 570457 12559 570575 12865
rect 570457 12543 570473 12559
rect 70648 12427 70664 12493
rect 122648 12427 122664 12493
rect 174648 12427 174664 12493
rect 226648 12427 226664 12493
rect 274648 12427 274664 12493
rect 326648 12427 326664 12493
rect 376624 12427 376640 12493
rect 378648 12427 378664 12493
rect 426648 12427 426664 12493
rect 476624 12427 476640 12493
rect 478648 12427 478664 12493
rect 530648 12427 530664 12493
rect 576624 12427 576640 12493
rect 578648 12427 578664 12493
rect 56970 9990 57252 10026
rect 108970 9990 109252 10026
rect 160970 9990 161252 10026
rect 212970 9990 213252 10026
rect 260970 9990 261252 10026
rect 312970 9990 313252 10026
rect 364970 9990 365252 10026
rect 365701 9990 365814 10026
rect 377866 9990 378076 10026
rect 412970 9990 413252 10026
rect 464970 9990 465252 10026
rect 465701 9990 465814 10026
rect 477866 9990 478076 10026
rect 516970 9990 517252 10026
rect 564970 9990 565252 10026
rect 565701 9990 565814 10026
rect 577866 9990 578076 10026
rect 56559 8990 56663 9990
rect 56759 8990 56831 9990
rect 56970 8990 57010 9990
rect 57047 8990 57103 9990
rect 57119 8990 57175 9990
rect 57216 8990 57252 9990
rect 58039 8990 58095 9990
rect 58111 8990 58167 9990
rect 69901 8990 69902 9990
rect 69943 8990 69999 9990
rect 70040 8990 70041 9990
rect 70383 9976 70487 9990
rect 70383 9942 70477 9976
rect 70383 9905 70487 9942
rect 70383 9871 70477 9905
rect 70383 9831 70487 9871
rect 70383 9797 70477 9831
rect 70383 9760 70487 9797
rect 70383 9726 70477 9760
rect 70383 9686 70487 9726
rect 70383 9652 70477 9686
rect 70383 9615 70487 9652
rect 70383 9581 70477 9615
rect 70383 9541 70487 9581
rect 70383 9507 70477 9541
rect 70383 9470 70487 9507
rect 70383 9436 70477 9470
rect 70383 9396 70487 9436
rect 70383 9362 70477 9396
rect 70383 9325 70487 9362
rect 70383 9291 70477 9325
rect 70383 9231 70487 9291
rect 70383 9197 70477 9231
rect 70383 9154 70487 9197
rect 70383 9120 70477 9154
rect 70383 9078 70487 9120
rect 70383 9044 70477 9078
rect 70383 8996 70487 9044
rect 70383 8990 70477 8996
rect 108559 8990 108663 9990
rect 108759 8990 108831 9990
rect 108970 8990 109010 9990
rect 109047 8990 109103 9990
rect 109119 8990 109175 9990
rect 109216 8990 109252 9990
rect 110039 8990 110095 9990
rect 110111 8990 110167 9990
rect 121901 8990 121902 9990
rect 121943 8990 121999 9990
rect 122040 8990 122041 9990
rect 122383 9976 122487 9990
rect 122383 9942 122477 9976
rect 122383 9905 122487 9942
rect 122383 9871 122477 9905
rect 122383 9831 122487 9871
rect 122383 9797 122477 9831
rect 122383 9760 122487 9797
rect 122383 9726 122477 9760
rect 122383 9686 122487 9726
rect 122383 9652 122477 9686
rect 122383 9615 122487 9652
rect 122383 9581 122477 9615
rect 122383 9541 122487 9581
rect 122383 9507 122477 9541
rect 122383 9470 122487 9507
rect 122383 9436 122477 9470
rect 122383 9396 122487 9436
rect 122383 9362 122477 9396
rect 122383 9325 122487 9362
rect 122383 9291 122477 9325
rect 122383 9231 122487 9291
rect 122383 9197 122477 9231
rect 122383 9154 122487 9197
rect 122383 9120 122477 9154
rect 122383 9078 122487 9120
rect 122383 9044 122477 9078
rect 122383 8996 122487 9044
rect 122383 8990 122477 8996
rect 160559 8990 160663 9990
rect 160759 8990 160831 9990
rect 160970 8990 161010 9990
rect 161047 8990 161103 9990
rect 161119 8990 161175 9990
rect 161216 8990 161252 9990
rect 173901 8990 173902 9990
rect 173943 8990 173999 9990
rect 174040 8990 174041 9990
rect 174383 9976 174487 9990
rect 174383 9942 174477 9976
rect 174383 9905 174487 9942
rect 174383 9871 174477 9905
rect 174383 9831 174487 9871
rect 174383 9797 174477 9831
rect 174383 9760 174487 9797
rect 174383 9726 174477 9760
rect 174383 9686 174487 9726
rect 174383 9652 174477 9686
rect 174383 9615 174487 9652
rect 174383 9581 174477 9615
rect 174383 9541 174487 9581
rect 174383 9507 174477 9541
rect 174383 9470 174487 9507
rect 174383 9436 174477 9470
rect 174383 9396 174487 9436
rect 174383 9362 174477 9396
rect 174383 9325 174487 9362
rect 174383 9291 174477 9325
rect 174383 9231 174487 9291
rect 174383 9197 174477 9231
rect 174383 9154 174487 9197
rect 174383 9120 174477 9154
rect 174383 9078 174487 9120
rect 174383 9044 174477 9078
rect 174383 8996 174487 9044
rect 174383 8990 174477 8996
rect 212559 8990 212663 9990
rect 212759 8990 212831 9990
rect 212970 8990 213010 9990
rect 213047 8990 213103 9990
rect 213119 8990 213175 9990
rect 213216 8990 213252 9990
rect 214039 8990 214095 9990
rect 214111 8990 214167 9990
rect 225901 8990 225902 9990
rect 225943 8990 225999 9990
rect 226040 8990 226041 9990
rect 226383 9976 226487 9990
rect 226383 9942 226477 9976
rect 226383 9905 226487 9942
rect 226383 9871 226477 9905
rect 226383 9831 226487 9871
rect 226383 9797 226477 9831
rect 226383 9760 226487 9797
rect 226383 9726 226477 9760
rect 226383 9686 226487 9726
rect 226383 9652 226477 9686
rect 226383 9615 226487 9652
rect 226383 9581 226477 9615
rect 226383 9541 226487 9581
rect 226383 9507 226477 9541
rect 226383 9470 226487 9507
rect 226383 9436 226477 9470
rect 226383 9396 226487 9436
rect 226383 9362 226477 9396
rect 226383 9325 226487 9362
rect 226383 9291 226477 9325
rect 226383 9231 226487 9291
rect 226383 9197 226477 9231
rect 226383 9154 226487 9197
rect 226383 9120 226477 9154
rect 226383 9078 226487 9120
rect 226383 9044 226477 9078
rect 226383 8996 226487 9044
rect 226383 8990 226477 8996
rect 260559 8990 260663 9990
rect 260759 8990 260831 9990
rect 260970 8990 261010 9990
rect 261047 8990 261103 9990
rect 261119 8990 261175 9990
rect 261216 8990 261252 9990
rect 262039 8990 262080 9990
rect 273901 8990 273902 9990
rect 273943 8990 273999 9990
rect 274040 8990 274041 9990
rect 274383 9976 274487 9990
rect 274383 9942 274477 9976
rect 274383 9905 274487 9942
rect 274383 9871 274477 9905
rect 274383 9831 274487 9871
rect 274383 9797 274477 9831
rect 274383 9760 274487 9797
rect 274383 9726 274477 9760
rect 274383 9686 274487 9726
rect 274383 9652 274477 9686
rect 274383 9615 274487 9652
rect 274383 9581 274477 9615
rect 274383 9541 274487 9581
rect 274383 9507 274477 9541
rect 274383 9470 274487 9507
rect 274383 9436 274477 9470
rect 274383 9396 274487 9436
rect 274383 9362 274477 9396
rect 274383 9325 274487 9362
rect 274383 9291 274477 9325
rect 274383 9231 274487 9291
rect 274383 9197 274477 9231
rect 274383 9154 274487 9197
rect 274383 9120 274477 9154
rect 274383 9078 274487 9120
rect 274383 9044 274477 9078
rect 274383 8996 274487 9044
rect 274383 8990 274477 8996
rect 312559 8990 312663 9990
rect 312759 8990 312831 9990
rect 312970 8990 313010 9990
rect 313047 8990 313103 9990
rect 313119 8990 313175 9990
rect 313216 8990 313252 9990
rect 314039 8990 314095 9990
rect 314111 8990 314167 9990
rect 325901 8990 325902 9990
rect 325943 8990 325999 9990
rect 326040 8990 326041 9990
rect 326383 9976 326487 9990
rect 326383 9942 326477 9976
rect 326383 9905 326487 9942
rect 326383 9871 326477 9905
rect 326383 9831 326487 9871
rect 326383 9797 326477 9831
rect 326383 9760 326487 9797
rect 326383 9726 326477 9760
rect 326383 9686 326487 9726
rect 326383 9652 326477 9686
rect 326383 9615 326487 9652
rect 326383 9581 326477 9615
rect 326383 9541 326487 9581
rect 326383 9507 326477 9541
rect 326383 9470 326487 9507
rect 326383 9436 326477 9470
rect 326383 9396 326487 9436
rect 326383 9362 326477 9396
rect 326383 9325 326487 9362
rect 326383 9291 326477 9325
rect 326383 9231 326487 9291
rect 326383 9197 326477 9231
rect 326383 9154 326487 9197
rect 326383 9120 326477 9154
rect 326383 9078 326487 9120
rect 326383 9044 326477 9078
rect 326383 8996 326487 9044
rect 326383 8990 326477 8996
rect 364559 8990 364663 9990
rect 364759 8990 364831 9990
rect 364970 8990 365010 9990
rect 365047 8990 365103 9990
rect 365119 8990 365175 9990
rect 365216 8990 365252 9990
rect 365266 8990 365270 9990
rect 365477 8990 365537 9990
rect 365701 8990 365737 9990
rect 365778 8990 365814 9990
rect 365828 8990 365832 9990
rect 366039 8990 366095 9990
rect 366111 8990 366167 9990
rect 366469 8990 366529 9990
rect 366729 8990 366801 9990
rect 367031 8990 367087 9990
rect 367103 8990 367159 9990
rect 367461 8990 367521 9990
rect 367721 8990 367793 9990
rect 368023 8990 368079 9990
rect 368095 8990 368151 9990
rect 368453 8990 368513 9990
rect 368713 8990 368785 9990
rect 369015 8990 369071 9990
rect 369087 8990 369143 9990
rect 369445 8990 369505 9990
rect 369705 8990 369777 9990
rect 370007 8990 370063 9990
rect 370079 8990 370135 9990
rect 370437 8990 370497 9990
rect 370697 8990 370769 9990
rect 370999 8990 371055 9990
rect 371071 8990 371127 9990
rect 371429 8990 371489 9990
rect 371689 8990 371761 9990
rect 371991 8990 372047 9990
rect 372063 8990 372119 9990
rect 372421 8990 372481 9990
rect 372681 8990 372753 9990
rect 372983 8990 373039 9990
rect 373055 8990 373111 9990
rect 373413 8990 373473 9990
rect 373673 8990 373745 9990
rect 373975 8990 374031 9990
rect 374047 8990 374103 9990
rect 374405 8990 374465 9990
rect 374665 8990 374737 9990
rect 374967 8990 375023 9990
rect 375039 8990 375095 9990
rect 375397 8990 375457 9990
rect 375657 8990 375729 9990
rect 375959 8990 376015 9990
rect 376031 8990 376087 9990
rect 376389 8990 376449 9990
rect 376649 8990 376721 9990
rect 376951 8990 377007 9990
rect 377023 8990 377079 9990
rect 377381 8990 377441 9990
rect 377641 8990 377713 9990
rect 377901 8990 377906 9990
rect 377943 8990 377999 9990
rect 378040 8990 378041 9990
rect 378287 8990 378347 9990
rect 378383 9976 378487 9990
rect 378383 9942 378477 9976
rect 378487 9942 378521 9976
rect 378383 9905 378487 9942
rect 378383 9871 378477 9905
rect 378487 9871 378521 9905
rect 378383 9831 378487 9871
rect 378383 9797 378477 9831
rect 378487 9797 378521 9831
rect 378383 9760 378487 9797
rect 378383 9726 378477 9760
rect 378487 9726 378521 9760
rect 378383 9686 378487 9726
rect 378383 9652 378477 9686
rect 378487 9652 378521 9686
rect 378383 9615 378487 9652
rect 378383 9581 378477 9615
rect 378487 9581 378521 9615
rect 378383 9541 378487 9581
rect 378383 9507 378477 9541
rect 378487 9507 378521 9541
rect 378383 9470 378487 9507
rect 378383 9436 378477 9470
rect 378487 9436 378521 9470
rect 378383 9396 378487 9436
rect 378383 9362 378477 9396
rect 378487 9362 378521 9396
rect 378383 9325 378487 9362
rect 378383 9291 378477 9325
rect 378487 9291 378521 9325
rect 378383 9231 378487 9291
rect 378383 9197 378477 9231
rect 378487 9197 378521 9231
rect 378383 9154 378487 9197
rect 378383 9120 378477 9154
rect 378487 9120 378521 9154
rect 378383 9078 378487 9120
rect 378383 9044 378477 9078
rect 378487 9044 378521 9078
rect 378383 8996 378487 9044
rect 378383 8990 378521 8996
rect 412559 8990 412663 9990
rect 412759 8990 412831 9990
rect 412970 8990 413010 9990
rect 413047 8990 413103 9990
rect 413119 8990 413175 9990
rect 413216 8990 413252 9990
rect 414039 8990 414095 9990
rect 414111 8990 414167 9990
rect 425901 8990 425902 9990
rect 425943 8990 425999 9990
rect 426040 8990 426041 9990
rect 426383 9976 426487 9990
rect 426383 9942 426477 9976
rect 426383 9905 426487 9942
rect 426383 9871 426477 9905
rect 426383 9831 426487 9871
rect 426383 9797 426477 9831
rect 426383 9760 426487 9797
rect 426383 9726 426477 9760
rect 426383 9686 426487 9726
rect 426383 9652 426477 9686
rect 426383 9615 426487 9652
rect 426383 9581 426477 9615
rect 426383 9541 426487 9581
rect 426383 9507 426477 9541
rect 426383 9470 426487 9507
rect 426383 9436 426477 9470
rect 426383 9396 426487 9436
rect 426383 9362 426477 9396
rect 426383 9325 426487 9362
rect 426383 9291 426477 9325
rect 426383 9231 426487 9291
rect 426383 9197 426477 9231
rect 426383 9154 426487 9197
rect 426383 9120 426477 9154
rect 426383 9078 426487 9120
rect 426383 9044 426477 9078
rect 426383 8996 426487 9044
rect 426383 8990 426477 8996
rect 464559 8990 464663 9990
rect 464759 8990 464831 9990
rect 464970 8990 465010 9990
rect 465047 8990 465103 9990
rect 465119 8990 465175 9990
rect 465216 8990 465252 9990
rect 465266 8990 465270 9990
rect 465477 8990 465537 9990
rect 465701 8990 465737 9990
rect 465778 8990 465814 9990
rect 465828 8990 465832 9990
rect 466039 8990 466095 9990
rect 466111 8990 466167 9990
rect 466469 8990 466529 9990
rect 466729 8990 466801 9990
rect 467031 8990 467087 9990
rect 467103 8990 467159 9990
rect 467461 8990 467521 9990
rect 467721 8990 467793 9990
rect 468023 8990 468079 9990
rect 468095 8990 468151 9990
rect 468453 8990 468513 9990
rect 468713 8990 468785 9990
rect 469015 8990 469071 9990
rect 469087 8990 469143 9990
rect 469445 8990 469505 9990
rect 469705 8990 469777 9990
rect 470007 8990 470063 9990
rect 470079 8990 470135 9990
rect 470437 8990 470497 9990
rect 470697 8990 470769 9990
rect 470999 8990 471055 9990
rect 471071 8990 471127 9990
rect 471429 8990 471489 9990
rect 471689 8990 471761 9990
rect 471991 8990 472047 9990
rect 472063 8990 472119 9990
rect 472421 8990 472481 9990
rect 472681 8990 472753 9990
rect 472983 8990 473039 9990
rect 473055 8990 473111 9990
rect 473413 8990 473473 9990
rect 473673 8990 473745 9990
rect 473975 8990 474031 9990
rect 474047 8990 474103 9990
rect 474405 8990 474465 9990
rect 474665 8990 474737 9990
rect 474967 8990 475023 9990
rect 475039 8990 475095 9990
rect 475397 8990 475457 9990
rect 475657 8990 475729 9990
rect 475959 8990 476015 9990
rect 476031 8990 476087 9990
rect 476389 8990 476449 9990
rect 476649 8990 476721 9990
rect 476951 8990 477007 9990
rect 477023 8990 477079 9990
rect 477381 8990 477441 9990
rect 477641 8990 477713 9990
rect 477901 8990 477906 9990
rect 477943 8990 477999 9990
rect 478040 8990 478041 9990
rect 478287 8990 478347 9990
rect 478383 9976 478487 9990
rect 478383 9942 478477 9976
rect 478487 9942 478521 9976
rect 478383 9905 478487 9942
rect 478383 9871 478477 9905
rect 478487 9871 478521 9905
rect 478383 9831 478487 9871
rect 478383 9797 478477 9831
rect 478487 9797 478521 9831
rect 478383 9760 478487 9797
rect 478383 9726 478477 9760
rect 478487 9726 478521 9760
rect 478383 9686 478487 9726
rect 478383 9652 478477 9686
rect 478487 9652 478521 9686
rect 478383 9615 478487 9652
rect 478383 9581 478477 9615
rect 478487 9581 478521 9615
rect 478383 9541 478487 9581
rect 478383 9507 478477 9541
rect 478487 9507 478521 9541
rect 478383 9470 478487 9507
rect 478383 9436 478477 9470
rect 478487 9436 478521 9470
rect 478383 9396 478487 9436
rect 478383 9362 478477 9396
rect 478487 9362 478521 9396
rect 478383 9325 478487 9362
rect 478383 9291 478477 9325
rect 478487 9291 478521 9325
rect 478383 9231 478487 9291
rect 478383 9197 478477 9231
rect 478487 9197 478521 9231
rect 478383 9154 478487 9197
rect 478383 9120 478477 9154
rect 478487 9120 478521 9154
rect 478383 9078 478487 9120
rect 478383 9044 478477 9078
rect 478487 9044 478521 9078
rect 478383 8996 478487 9044
rect 478383 8990 478521 8996
rect 516559 8990 516663 9990
rect 516759 8990 516831 9990
rect 516970 8990 517010 9990
rect 517047 8990 517103 9990
rect 517119 8990 517175 9990
rect 517216 8990 517252 9990
rect 518039 8990 518095 9990
rect 518111 8990 518167 9990
rect 529901 8990 529902 9990
rect 529943 8990 529999 9990
rect 530040 8990 530041 9990
rect 530383 9976 530487 9990
rect 530383 9942 530477 9976
rect 530383 9905 530487 9942
rect 530383 9871 530477 9905
rect 530383 9831 530487 9871
rect 530383 9797 530477 9831
rect 530383 9760 530487 9797
rect 530383 9726 530477 9760
rect 530383 9686 530487 9726
rect 530383 9652 530477 9686
rect 530383 9615 530487 9652
rect 530383 9581 530477 9615
rect 530383 9541 530487 9581
rect 530383 9507 530477 9541
rect 530383 9470 530487 9507
rect 530383 9436 530477 9470
rect 530383 9396 530487 9436
rect 530383 9362 530477 9396
rect 530383 9325 530487 9362
rect 530383 9291 530477 9325
rect 530383 9231 530487 9291
rect 530383 9197 530477 9231
rect 530383 9154 530487 9197
rect 530383 9120 530477 9154
rect 530383 9078 530487 9120
rect 530383 9044 530477 9078
rect 530383 8996 530487 9044
rect 530383 8990 530477 8996
rect 564559 8990 564663 9990
rect 564759 8990 564831 9990
rect 564970 8990 565010 9990
rect 565047 8990 565103 9990
rect 565119 8990 565175 9990
rect 565216 8990 565252 9990
rect 565266 8990 565270 9990
rect 565477 8990 565537 9990
rect 565701 8990 565737 9990
rect 565778 8990 565814 9990
rect 565828 8990 565832 9990
rect 566039 8990 566095 9990
rect 566111 8990 566167 9990
rect 566469 8990 566529 9990
rect 566729 8990 566801 9990
rect 567031 8990 567087 9990
rect 567103 8990 567159 9990
rect 567461 8990 567521 9990
rect 567721 8990 567793 9990
rect 568023 8990 568079 9990
rect 568095 8990 568151 9990
rect 568453 8990 568513 9990
rect 568713 8990 568785 9990
rect 569015 8990 569071 9990
rect 569087 8990 569143 9990
rect 569445 8990 569505 9990
rect 569705 8990 569777 9990
rect 570007 8990 570063 9990
rect 570079 8990 570135 9990
rect 570437 8990 570497 9990
rect 570697 8990 570769 9990
rect 570999 8990 571055 9990
rect 571071 8990 571127 9990
rect 571429 8990 571489 9990
rect 571689 8990 571761 9990
rect 571991 8990 572047 9990
rect 572063 8990 572119 9990
rect 572421 8990 572481 9990
rect 572681 8990 572753 9990
rect 572983 8990 573039 9990
rect 573055 8990 573111 9990
rect 573413 8990 573473 9990
rect 573673 8990 573745 9990
rect 573975 8990 574031 9990
rect 574047 8990 574103 9990
rect 574405 8990 574465 9990
rect 574665 8990 574737 9990
rect 574967 8990 575023 9990
rect 575039 8990 575095 9990
rect 575397 8990 575457 9990
rect 575657 8990 575729 9990
rect 575959 8990 576015 9990
rect 576031 8990 576087 9990
rect 576389 8990 576449 9990
rect 576649 8990 576721 9990
rect 576951 8990 577007 9990
rect 577023 8990 577079 9990
rect 577381 8990 577441 9990
rect 577641 8990 577713 9990
rect 577901 8990 577906 9990
rect 577943 8990 577999 9990
rect 578040 8990 578041 9990
rect 578287 8990 578347 9990
rect 578383 9976 578487 9990
rect 578383 9942 578477 9976
rect 578487 9942 578521 9976
rect 578383 9905 578487 9942
rect 578383 9871 578477 9905
rect 578487 9871 578521 9905
rect 578383 9831 578487 9871
rect 578383 9797 578477 9831
rect 578487 9797 578521 9831
rect 578383 9760 578487 9797
rect 578383 9726 578477 9760
rect 578487 9726 578521 9760
rect 578383 9686 578487 9726
rect 578383 9652 578477 9686
rect 578487 9652 578521 9686
rect 578383 9615 578487 9652
rect 578383 9581 578477 9615
rect 578487 9581 578521 9615
rect 578383 9541 578487 9581
rect 578383 9507 578477 9541
rect 578487 9507 578521 9541
rect 578383 9470 578487 9507
rect 578383 9436 578477 9470
rect 578487 9436 578521 9470
rect 578383 9396 578487 9436
rect 578383 9362 578477 9396
rect 578487 9362 578521 9396
rect 578383 9325 578487 9362
rect 578383 9291 578477 9325
rect 578487 9291 578521 9325
rect 578383 9231 578487 9291
rect 578383 9197 578477 9231
rect 578487 9197 578521 9231
rect 578383 9154 578487 9197
rect 578383 9120 578477 9154
rect 578487 9120 578521 9154
rect 578383 9078 578487 9120
rect 578383 9044 578477 9078
rect 578487 9044 578521 9078
rect 578383 8996 578487 9044
rect 578383 8990 578521 8996
rect 56970 8954 57252 8990
rect 108970 8954 109252 8990
rect 160970 8954 161252 8990
rect 212970 8954 213252 8990
rect 260970 8954 261252 8990
rect 312970 8954 313252 8990
rect 364970 8954 365252 8990
rect 365701 8954 365814 8990
rect 377866 8954 378076 8990
rect 412970 8954 413252 8990
rect 464970 8954 465252 8990
rect 465701 8954 465814 8990
rect 477866 8954 478076 8990
rect 516970 8954 517252 8990
rect 564970 8954 565252 8990
rect 565701 8954 565814 8990
rect 577866 8954 578076 8990
rect 56559 8389 56569 8413
rect 56970 8389 57252 8425
rect 108559 8389 108569 8413
rect 108970 8389 109252 8425
rect 160559 8389 160569 8413
rect 160970 8389 161252 8425
rect 212559 8389 212569 8413
rect 212970 8389 213252 8425
rect 260559 8389 260569 8413
rect 260970 8389 261252 8425
rect 312559 8389 312569 8413
rect 312970 8389 313252 8425
rect 364559 8389 364569 8413
rect 364970 8389 365252 8425
rect 365701 8389 365814 8425
rect 377866 8389 378076 8425
rect 378477 8415 378521 8423
rect 378477 8389 378487 8415
rect 378511 8389 378521 8415
rect 56559 7389 56663 8389
rect 56759 7389 56831 8389
rect 56970 7389 57010 8389
rect 57047 7389 57103 8389
rect 57119 7389 57175 8389
rect 57216 7389 57252 8389
rect 58039 7389 58095 8389
rect 58111 7389 58167 8389
rect 69943 7389 69999 8389
rect 70040 7389 70064 8389
rect 70409 8381 70477 8389
rect 70409 8330 70487 8381
rect 70409 8296 70477 8330
rect 70409 8236 70487 8296
rect 70409 8202 70477 8236
rect 70409 8165 70487 8202
rect 70409 8131 70477 8165
rect 70409 8091 70487 8131
rect 70409 8057 70477 8091
rect 70409 8020 70487 8057
rect 70409 7986 70477 8020
rect 70409 7946 70487 7986
rect 70409 7912 70477 7946
rect 70409 7875 70487 7912
rect 70409 7841 70477 7875
rect 70409 7801 70487 7841
rect 70409 7767 70477 7801
rect 70409 7730 70487 7767
rect 70409 7696 70477 7730
rect 70409 7656 70487 7696
rect 70409 7622 70477 7656
rect 70409 7585 70487 7622
rect 70409 7551 70477 7585
rect 70409 7511 70487 7551
rect 70409 7477 70477 7511
rect 70409 7440 70487 7477
rect 70409 7406 70477 7440
rect 70409 7389 70487 7406
rect 108559 7389 108663 8389
rect 108759 7389 108831 8389
rect 108970 7389 109010 8389
rect 109047 7389 109103 8389
rect 109119 7389 109175 8389
rect 109216 7389 109252 8389
rect 110039 7389 110095 8389
rect 110111 7389 110167 8389
rect 121943 7389 121999 8389
rect 122040 7389 122064 8389
rect 122409 8381 122477 8389
rect 122409 8330 122487 8381
rect 122409 8296 122477 8330
rect 122409 8236 122487 8296
rect 122409 8202 122477 8236
rect 122409 8165 122487 8202
rect 122409 8131 122477 8165
rect 122409 8091 122487 8131
rect 122409 8057 122477 8091
rect 122409 8020 122487 8057
rect 122409 7986 122477 8020
rect 122409 7946 122487 7986
rect 122409 7912 122477 7946
rect 122409 7875 122487 7912
rect 122409 7841 122477 7875
rect 122409 7801 122487 7841
rect 122409 7767 122477 7801
rect 122409 7730 122487 7767
rect 122409 7696 122477 7730
rect 122409 7656 122487 7696
rect 122409 7622 122477 7656
rect 122409 7585 122487 7622
rect 122409 7551 122477 7585
rect 122409 7511 122487 7551
rect 122409 7477 122477 7511
rect 122409 7440 122487 7477
rect 122409 7406 122477 7440
rect 122409 7389 122487 7406
rect 160559 7389 160663 8389
rect 160759 7389 160831 8389
rect 160970 7389 161010 8389
rect 161047 7389 161103 8389
rect 161119 7389 161175 8389
rect 161216 7389 161252 8389
rect 173943 7389 173999 8389
rect 174040 7389 174064 8389
rect 174409 8381 174477 8389
rect 174409 8330 174487 8381
rect 174409 8296 174477 8330
rect 174409 8236 174487 8296
rect 174409 8202 174477 8236
rect 174409 8165 174487 8202
rect 174409 8131 174477 8165
rect 174409 8091 174487 8131
rect 174409 8057 174477 8091
rect 174409 8020 174487 8057
rect 174409 7986 174477 8020
rect 174409 7946 174487 7986
rect 174409 7912 174477 7946
rect 174409 7875 174487 7912
rect 174409 7841 174477 7875
rect 174409 7801 174487 7841
rect 174409 7767 174477 7801
rect 174409 7730 174487 7767
rect 174409 7696 174477 7730
rect 174409 7656 174487 7696
rect 174409 7622 174477 7656
rect 174409 7585 174487 7622
rect 174409 7551 174477 7585
rect 174409 7511 174487 7551
rect 174409 7477 174477 7511
rect 174409 7440 174487 7477
rect 174409 7406 174477 7440
rect 174409 7389 174487 7406
rect 212559 7389 212663 8389
rect 212759 7389 212831 8389
rect 212970 7389 213010 8389
rect 213047 7389 213103 8389
rect 213119 7389 213175 8389
rect 213216 7389 213252 8389
rect 214039 7389 214095 8389
rect 214111 7389 214167 8389
rect 225943 7389 225999 8389
rect 226040 7389 226064 8389
rect 226409 8381 226477 8389
rect 226409 8330 226487 8381
rect 226409 8296 226477 8330
rect 226409 8236 226487 8296
rect 226409 8202 226477 8236
rect 226409 8165 226487 8202
rect 226409 8131 226477 8165
rect 226409 8091 226487 8131
rect 226409 8057 226477 8091
rect 226409 8020 226487 8057
rect 226409 7986 226477 8020
rect 226409 7946 226487 7986
rect 226409 7912 226477 7946
rect 226409 7875 226487 7912
rect 226409 7841 226477 7875
rect 226409 7801 226487 7841
rect 226409 7767 226477 7801
rect 226409 7730 226487 7767
rect 226409 7696 226477 7730
rect 226409 7656 226487 7696
rect 226409 7622 226477 7656
rect 226409 7585 226487 7622
rect 226409 7551 226477 7585
rect 226409 7511 226487 7551
rect 226409 7477 226477 7511
rect 226409 7440 226487 7477
rect 226409 7406 226477 7440
rect 226409 7389 226487 7406
rect 260559 7389 260663 8389
rect 260759 7389 260831 8389
rect 260970 7389 261010 8389
rect 261047 7389 261103 8389
rect 261119 7389 261175 8389
rect 261216 7389 261252 8389
rect 262039 7389 262080 8389
rect 273943 7389 273999 8389
rect 274040 7389 274064 8389
rect 274409 8381 274477 8389
rect 274409 8330 274487 8381
rect 274409 8296 274477 8330
rect 274409 8236 274487 8296
rect 274409 8202 274477 8236
rect 274409 8165 274487 8202
rect 274409 8131 274477 8165
rect 274409 8091 274487 8131
rect 274409 8057 274477 8091
rect 274409 8020 274487 8057
rect 274409 7986 274477 8020
rect 274409 7946 274487 7986
rect 274409 7912 274477 7946
rect 274409 7875 274487 7912
rect 274409 7841 274477 7875
rect 274409 7801 274487 7841
rect 274409 7767 274477 7801
rect 274409 7730 274487 7767
rect 274409 7696 274477 7730
rect 274409 7656 274487 7696
rect 274409 7622 274477 7656
rect 274409 7585 274487 7622
rect 274409 7551 274477 7585
rect 274409 7511 274487 7551
rect 274409 7477 274477 7511
rect 274409 7440 274487 7477
rect 274409 7406 274477 7440
rect 274409 7389 274487 7406
rect 312559 7389 312663 8389
rect 312759 7389 312831 8389
rect 312970 7389 313010 8389
rect 313047 7389 313103 8389
rect 313119 7389 313175 8389
rect 313216 7389 313252 8389
rect 314039 7389 314095 8389
rect 314111 7389 314167 8389
rect 325943 7389 325999 8389
rect 326040 7389 326064 8389
rect 326409 8381 326477 8389
rect 326409 8330 326487 8381
rect 326409 8296 326477 8330
rect 326409 8236 326487 8296
rect 326409 8202 326477 8236
rect 326409 8165 326487 8202
rect 326409 8131 326477 8165
rect 326409 8091 326487 8131
rect 326409 8057 326477 8091
rect 326409 8020 326487 8057
rect 326409 7986 326477 8020
rect 326409 7946 326487 7986
rect 326409 7912 326477 7946
rect 326409 7875 326487 7912
rect 326409 7841 326477 7875
rect 326409 7801 326487 7841
rect 326409 7767 326477 7801
rect 326409 7730 326487 7767
rect 326409 7696 326477 7730
rect 326409 7656 326487 7696
rect 326409 7622 326477 7656
rect 326409 7585 326487 7622
rect 326409 7551 326477 7585
rect 326409 7511 326487 7551
rect 326409 7477 326477 7511
rect 326409 7440 326487 7477
rect 326409 7406 326477 7440
rect 326409 7389 326487 7406
rect 364559 7389 364663 8389
rect 364759 7389 364831 8389
rect 364970 7389 365010 8389
rect 365047 7389 365103 8389
rect 365119 7389 365175 8389
rect 365216 7389 365252 8389
rect 365266 7389 365270 8389
rect 365477 7389 365537 8389
rect 365701 7389 365737 8389
rect 365778 7389 365814 8389
rect 365828 7389 365832 8389
rect 366039 7389 366095 8389
rect 366111 7389 366167 8389
rect 366469 7389 366529 8389
rect 366729 7389 366801 8389
rect 367031 7389 367087 8389
rect 367103 7389 367159 8389
rect 367461 7389 367521 8389
rect 367721 7389 367793 8389
rect 368023 7389 368079 8389
rect 368095 7389 368151 8389
rect 368453 7389 368513 8389
rect 368713 7389 368785 8389
rect 369015 7389 369071 8389
rect 369087 7389 369143 8389
rect 369445 7389 369505 8389
rect 369705 7389 369777 8389
rect 370007 7389 370063 8389
rect 370079 7389 370135 8389
rect 370437 7389 370497 8389
rect 370697 7389 370769 8389
rect 370999 7389 371055 8389
rect 371071 7389 371127 8389
rect 371429 7389 371489 8389
rect 371689 7389 371761 8389
rect 371991 7389 372047 8389
rect 372063 7389 372119 8389
rect 372421 7389 372481 8389
rect 372681 7389 372753 8389
rect 372983 7389 373039 8389
rect 373055 7389 373111 8389
rect 373413 7389 373473 8389
rect 373673 7389 373745 8389
rect 373975 7389 374031 8389
rect 374047 7389 374103 8389
rect 374405 7389 374465 8389
rect 374665 7389 374737 8389
rect 374967 7389 375023 8389
rect 375039 7389 375095 8389
rect 375397 7389 375457 8389
rect 375657 7389 375729 8389
rect 375959 7389 376015 8389
rect 376031 7389 376087 8389
rect 376389 7389 376449 8389
rect 376649 7389 376721 8389
rect 376951 7389 377007 8389
rect 377023 7389 377079 8389
rect 377381 7389 377441 8389
rect 377641 7389 377713 8389
rect 377866 7389 377906 8389
rect 377943 7389 377999 8389
rect 378040 7389 378064 8389
rect 378287 7389 378347 8389
rect 378409 8381 378477 8389
rect 378487 8381 378521 8389
rect 412559 8389 412569 8413
rect 412970 8389 413252 8425
rect 464559 8389 464569 8413
rect 464970 8389 465252 8425
rect 465701 8389 465814 8425
rect 477866 8389 478076 8425
rect 478477 8415 478521 8423
rect 478477 8389 478487 8415
rect 478511 8389 478521 8415
rect 378409 8330 378487 8381
rect 378409 8296 378477 8330
rect 378487 8296 378521 8330
rect 378409 8236 378487 8296
rect 378409 8202 378477 8236
rect 378487 8202 378521 8236
rect 378409 8165 378487 8202
rect 378409 8131 378477 8165
rect 378487 8131 378521 8165
rect 378409 8091 378487 8131
rect 378409 8057 378477 8091
rect 378487 8057 378521 8091
rect 378409 8020 378487 8057
rect 378409 7986 378477 8020
rect 378487 7986 378521 8020
rect 378409 7946 378487 7986
rect 378409 7912 378477 7946
rect 378487 7912 378521 7946
rect 378409 7875 378487 7912
rect 378409 7841 378477 7875
rect 378487 7841 378521 7875
rect 378409 7801 378487 7841
rect 378409 7767 378477 7801
rect 378487 7767 378521 7801
rect 378409 7730 378487 7767
rect 378409 7696 378477 7730
rect 378487 7696 378521 7730
rect 378409 7656 378487 7696
rect 378409 7622 378477 7656
rect 378487 7622 378521 7656
rect 378409 7585 378487 7622
rect 378409 7551 378477 7585
rect 378487 7551 378521 7585
rect 378409 7511 378487 7551
rect 378409 7477 378477 7511
rect 378487 7477 378521 7511
rect 378409 7440 378487 7477
rect 378409 7406 378477 7440
rect 378487 7406 378521 7440
rect 378409 7389 378487 7406
rect 412559 7389 412663 8389
rect 412759 7389 412831 8389
rect 412970 7389 413010 8389
rect 413047 7389 413103 8389
rect 413119 7389 413175 8389
rect 413216 7389 413252 8389
rect 414039 7389 414095 8389
rect 414111 7389 414167 8389
rect 425943 7389 425999 8389
rect 426040 7389 426064 8389
rect 426409 8381 426477 8389
rect 426409 8330 426487 8381
rect 426409 8296 426477 8330
rect 426409 8236 426487 8296
rect 426409 8202 426477 8236
rect 426409 8165 426487 8202
rect 426409 8131 426477 8165
rect 426409 8091 426487 8131
rect 426409 8057 426477 8091
rect 426409 8020 426487 8057
rect 426409 7986 426477 8020
rect 426409 7946 426487 7986
rect 426409 7912 426477 7946
rect 426409 7875 426487 7912
rect 426409 7841 426477 7875
rect 426409 7801 426487 7841
rect 426409 7767 426477 7801
rect 426409 7730 426487 7767
rect 426409 7696 426477 7730
rect 426409 7656 426487 7696
rect 426409 7622 426477 7656
rect 426409 7585 426487 7622
rect 426409 7551 426477 7585
rect 426409 7511 426487 7551
rect 426409 7477 426477 7511
rect 426409 7440 426487 7477
rect 426409 7406 426477 7440
rect 426409 7389 426487 7406
rect 464559 7389 464663 8389
rect 464759 7389 464831 8389
rect 464970 7389 465010 8389
rect 465047 7389 465103 8389
rect 465119 7389 465175 8389
rect 465216 7389 465252 8389
rect 465266 7389 465270 8389
rect 465477 7389 465537 8389
rect 465701 7389 465737 8389
rect 465778 7389 465814 8389
rect 465828 7389 465832 8389
rect 466039 7389 466095 8389
rect 466111 7389 466167 8389
rect 466469 7389 466529 8389
rect 466729 7389 466801 8389
rect 467031 7389 467087 8389
rect 467103 7389 467159 8389
rect 467461 7389 467521 8389
rect 467721 7389 467793 8389
rect 468023 7389 468079 8389
rect 468095 7389 468151 8389
rect 468453 7389 468513 8389
rect 468713 7389 468785 8389
rect 469015 7389 469071 8389
rect 469087 7389 469143 8389
rect 469445 7389 469505 8389
rect 469705 7389 469777 8389
rect 470007 7389 470063 8389
rect 470079 7389 470135 8389
rect 470437 7389 470497 8389
rect 470697 7389 470769 8389
rect 470999 7389 471055 8389
rect 471071 7389 471127 8389
rect 471429 7389 471489 8389
rect 471689 7389 471761 8389
rect 471991 7389 472047 8389
rect 472063 7389 472119 8389
rect 472421 7389 472481 8389
rect 472681 7389 472753 8389
rect 472983 7389 473039 8389
rect 473055 7389 473111 8389
rect 473413 7389 473473 8389
rect 473673 7389 473745 8389
rect 473975 7389 474031 8389
rect 474047 7389 474103 8389
rect 474405 7389 474465 8389
rect 474665 7389 474737 8389
rect 474967 7389 475023 8389
rect 475039 7389 475095 8389
rect 475397 7389 475457 8389
rect 475657 7389 475729 8389
rect 475959 7389 476015 8389
rect 476031 7389 476087 8389
rect 476389 7389 476449 8389
rect 476649 7389 476721 8389
rect 476951 7389 477007 8389
rect 477023 7389 477079 8389
rect 477381 7389 477441 8389
rect 477641 7389 477713 8389
rect 477866 7389 477906 8389
rect 477943 7389 477999 8389
rect 478040 7389 478064 8389
rect 478287 7389 478347 8389
rect 478409 8381 478477 8389
rect 478487 8381 478521 8389
rect 516559 8389 516569 8413
rect 516970 8389 517252 8425
rect 564559 8389 564569 8413
rect 564970 8389 565252 8425
rect 565701 8389 565814 8425
rect 577866 8389 578076 8425
rect 578477 8415 578521 8423
rect 578477 8389 578487 8415
rect 578511 8389 578521 8415
rect 478409 8330 478487 8381
rect 478409 8296 478477 8330
rect 478487 8296 478521 8330
rect 478409 8236 478487 8296
rect 478409 8202 478477 8236
rect 478487 8202 478521 8236
rect 478409 8165 478487 8202
rect 478409 8131 478477 8165
rect 478487 8131 478521 8165
rect 478409 8091 478487 8131
rect 478409 8057 478477 8091
rect 478487 8057 478521 8091
rect 478409 8020 478487 8057
rect 478409 7986 478477 8020
rect 478487 7986 478521 8020
rect 478409 7946 478487 7986
rect 478409 7912 478477 7946
rect 478487 7912 478521 7946
rect 478409 7875 478487 7912
rect 478409 7841 478477 7875
rect 478487 7841 478521 7875
rect 478409 7801 478487 7841
rect 478409 7767 478477 7801
rect 478487 7767 478521 7801
rect 478409 7730 478487 7767
rect 478409 7696 478477 7730
rect 478487 7696 478521 7730
rect 478409 7656 478487 7696
rect 478409 7622 478477 7656
rect 478487 7622 478521 7656
rect 478409 7585 478487 7622
rect 478409 7551 478477 7585
rect 478487 7551 478521 7585
rect 478409 7511 478487 7551
rect 478409 7477 478477 7511
rect 478487 7477 478521 7511
rect 478409 7440 478487 7477
rect 478409 7406 478477 7440
rect 478487 7406 478521 7440
rect 478409 7389 478487 7406
rect 516559 7389 516663 8389
rect 516759 7389 516831 8389
rect 516970 7389 517010 8389
rect 517047 7389 517103 8389
rect 517119 7389 517175 8389
rect 517216 7389 517252 8389
rect 518039 7389 518095 8389
rect 518111 7389 518167 8389
rect 529943 7389 529999 8389
rect 530040 7389 530064 8389
rect 530409 8381 530477 8389
rect 530409 8330 530487 8381
rect 530409 8296 530477 8330
rect 530409 8236 530487 8296
rect 530409 8202 530477 8236
rect 530409 8165 530487 8202
rect 530409 8131 530477 8165
rect 530409 8091 530487 8131
rect 530409 8057 530477 8091
rect 530409 8020 530487 8057
rect 530409 7986 530477 8020
rect 530409 7946 530487 7986
rect 530409 7912 530477 7946
rect 530409 7875 530487 7912
rect 530409 7841 530477 7875
rect 530409 7801 530487 7841
rect 530409 7767 530477 7801
rect 530409 7730 530487 7767
rect 530409 7696 530477 7730
rect 530409 7656 530487 7696
rect 530409 7622 530477 7656
rect 530409 7585 530487 7622
rect 530409 7551 530477 7585
rect 530409 7511 530487 7551
rect 530409 7477 530477 7511
rect 530409 7440 530487 7477
rect 530409 7406 530477 7440
rect 530409 7389 530487 7406
rect 564559 7389 564663 8389
rect 564759 7389 564831 8389
rect 564970 7389 565010 8389
rect 565047 7389 565103 8389
rect 565119 7389 565175 8389
rect 565216 7389 565252 8389
rect 565266 7389 565270 8389
rect 565477 7389 565537 8389
rect 565701 7389 565737 8389
rect 565778 7389 565814 8389
rect 565828 7389 565832 8389
rect 566039 7389 566095 8389
rect 566111 7389 566167 8389
rect 566469 7389 566529 8389
rect 566729 7389 566801 8389
rect 567031 7389 567087 8389
rect 567103 7389 567159 8389
rect 567461 7389 567521 8389
rect 567721 7389 567793 8389
rect 568023 7389 568079 8389
rect 568095 7389 568151 8389
rect 568453 7389 568513 8389
rect 568713 7389 568785 8389
rect 569015 7389 569071 8389
rect 569087 7389 569143 8389
rect 569445 7389 569505 8389
rect 569705 7389 569777 8389
rect 570007 7389 570063 8389
rect 570079 7389 570135 8389
rect 570437 7389 570497 8389
rect 570697 7389 570769 8389
rect 570999 7389 571055 8389
rect 571071 7389 571127 8389
rect 571429 7389 571489 8389
rect 571689 7389 571761 8389
rect 571991 7389 572047 8389
rect 572063 7389 572119 8389
rect 572421 7389 572481 8389
rect 572681 7389 572753 8389
rect 572983 7389 573039 8389
rect 573055 7389 573111 8389
rect 573413 7389 573473 8389
rect 573673 7389 573745 8389
rect 573975 7389 574031 8389
rect 574047 7389 574103 8389
rect 574405 7389 574465 8389
rect 574665 7389 574737 8389
rect 574967 7389 575023 8389
rect 575039 7389 575095 8389
rect 575397 7389 575457 8389
rect 575657 7389 575729 8389
rect 575959 7389 576015 8389
rect 576031 7389 576087 8389
rect 576389 7389 576449 8389
rect 576649 7389 576721 8389
rect 576951 7389 577007 8389
rect 577023 7389 577079 8389
rect 577381 7389 577441 8389
rect 577641 7389 577713 8389
rect 577866 7389 577906 8389
rect 577943 7389 577999 8389
rect 578040 7389 578064 8389
rect 578287 7389 578347 8389
rect 578409 8381 578477 8389
rect 578487 8381 578521 8389
rect 578409 8330 578487 8381
rect 578409 8296 578477 8330
rect 578487 8296 578521 8330
rect 578409 8236 578487 8296
rect 578409 8202 578477 8236
rect 578487 8202 578521 8236
rect 578409 8165 578487 8202
rect 578409 8131 578477 8165
rect 578487 8131 578521 8165
rect 578409 8091 578487 8131
rect 578409 8057 578477 8091
rect 578487 8057 578521 8091
rect 578409 8020 578487 8057
rect 578409 7986 578477 8020
rect 578487 7986 578521 8020
rect 578409 7946 578487 7986
rect 578409 7912 578477 7946
rect 578487 7912 578521 7946
rect 578409 7875 578487 7912
rect 578409 7841 578477 7875
rect 578487 7841 578521 7875
rect 578409 7801 578487 7841
rect 578409 7767 578477 7801
rect 578487 7767 578521 7801
rect 578409 7730 578487 7767
rect 578409 7696 578477 7730
rect 578487 7696 578521 7730
rect 578409 7656 578487 7696
rect 578409 7622 578477 7656
rect 578487 7622 578521 7656
rect 578409 7585 578487 7622
rect 578409 7551 578477 7585
rect 578487 7551 578521 7585
rect 578409 7511 578487 7551
rect 578409 7477 578477 7511
rect 578487 7477 578521 7511
rect 578409 7440 578487 7477
rect 578409 7406 578477 7440
rect 578487 7406 578521 7440
rect 578409 7389 578487 7406
rect 56970 7353 57252 7389
rect 108970 7353 109252 7389
rect 160970 7353 161252 7389
rect 212970 7353 213252 7389
rect 260970 7353 261252 7389
rect 312970 7353 313252 7389
rect 364970 7353 365252 7389
rect 365701 7353 365814 7389
rect 377866 7353 378076 7389
rect 412970 7353 413252 7389
rect 464970 7353 465252 7389
rect 465701 7353 465814 7389
rect 477866 7353 478076 7389
rect 516970 7353 517252 7389
rect 564970 7353 565252 7389
rect 565701 7353 565814 7389
rect 577866 7353 578076 7389
rect 366447 6059 366586 6089
rect 466447 6059 466586 6089
rect 566447 6059 566586 6089
rect 366447 6021 378698 6059
rect 466447 6021 478698 6059
rect 566447 6021 578698 6059
rect 56669 5995 58475 6021
rect 58505 6005 58520 6021
rect 69480 6005 70699 6021
rect 108669 5995 110475 6021
rect 110505 6005 110520 6021
rect 121480 6005 122699 6021
rect 160669 5995 161280 6021
rect 173480 6005 174699 6021
rect 212669 5995 214475 6021
rect 214505 6005 214520 6021
rect 225480 6005 226699 6021
rect 260669 5995 262080 6021
rect 273480 6005 274699 6021
rect 312669 5995 314475 6021
rect 314505 6005 314520 6021
rect 325480 6005 326699 6021
rect 364669 6005 378699 6021
rect 364669 5995 366475 6005
rect 56669 5981 56693 5995
rect 108669 5981 108693 5995
rect 160669 5981 160693 5995
rect 212669 5981 212693 5995
rect 260669 5981 260693 5995
rect 312669 5981 312693 5995
rect 364669 5981 364693 5995
rect 56669 5137 56683 5981
rect 69480 5658 70303 5708
rect 69480 5488 70303 5538
rect 58515 5169 58520 5191
rect 108669 5137 108683 5981
rect 121480 5658 122303 5708
rect 121480 5488 122303 5538
rect 110515 5169 110520 5191
rect 160669 5137 160683 5981
rect 173480 5658 174303 5708
rect 173480 5488 174303 5538
rect 212669 5137 212683 5981
rect 225480 5658 226303 5708
rect 225480 5488 226303 5538
rect 214515 5169 214520 5191
rect 260669 5137 260683 5981
rect 273480 5658 274303 5708
rect 273480 5488 274303 5538
rect 312669 5137 312683 5981
rect 325480 5658 326303 5708
rect 325480 5488 326303 5538
rect 314515 5169 314520 5191
rect 364669 5137 364683 5981
rect 366505 5967 366515 6005
rect 366518 5971 378698 6005
rect 366518 5967 366539 5971
rect 373655 5967 373689 5971
rect 378563 5967 378698 5971
rect 412669 5995 414475 6021
rect 414505 6005 414520 6021
rect 425480 6005 426699 6021
rect 464669 6005 478699 6021
rect 464669 5995 466475 6005
rect 412669 5981 412693 5995
rect 464669 5981 464693 5995
rect 366800 5658 367800 5708
rect 367921 5658 368921 5708
rect 369042 5658 370042 5708
rect 370152 5658 371152 5708
rect 371273 5658 372273 5708
rect 372394 5658 373394 5708
rect 373951 5658 374951 5708
rect 375072 5658 376072 5708
rect 376193 5658 377193 5708
rect 377303 5658 378303 5708
rect 366800 5488 367800 5538
rect 367921 5488 368921 5538
rect 369042 5488 370042 5538
rect 370152 5488 371152 5538
rect 371273 5488 372273 5538
rect 372394 5488 373394 5538
rect 373951 5488 374951 5538
rect 375072 5488 376072 5538
rect 376193 5488 377193 5538
rect 377303 5488 378303 5538
rect 366515 5169 373629 5191
rect 412669 5137 412683 5981
rect 425480 5658 426303 5708
rect 425480 5488 426303 5538
rect 414515 5169 414520 5191
rect 464669 5137 464683 5981
rect 466505 5967 466515 6005
rect 466518 5971 478698 6005
rect 466518 5967 466539 5971
rect 473655 5967 473689 5971
rect 478563 5967 478698 5971
rect 516669 5995 518475 6021
rect 518505 6005 518520 6021
rect 529480 6005 530699 6021
rect 564669 6005 578699 6021
rect 564669 5995 566475 6005
rect 516669 5981 516693 5995
rect 564669 5981 564693 5995
rect 466800 5658 467800 5708
rect 467921 5658 468921 5708
rect 469042 5658 470042 5708
rect 470152 5658 471152 5708
rect 471273 5658 472273 5708
rect 472394 5658 473394 5708
rect 473951 5658 474951 5708
rect 475072 5658 476072 5708
rect 476193 5658 477193 5708
rect 477303 5658 478303 5708
rect 466800 5488 467800 5538
rect 467921 5488 468921 5538
rect 469042 5488 470042 5538
rect 470152 5488 471152 5538
rect 471273 5488 472273 5538
rect 472394 5488 473394 5538
rect 473951 5488 474951 5538
rect 475072 5488 476072 5538
rect 476193 5488 477193 5538
rect 477303 5488 478303 5538
rect 466515 5169 473629 5191
rect 516669 5137 516683 5981
rect 529480 5658 530303 5708
rect 529480 5488 530303 5538
rect 518515 5169 518520 5191
rect 564669 5137 564683 5981
rect 566505 5967 566515 6005
rect 566518 5971 578698 6005
rect 566518 5967 566539 5971
rect 573655 5967 573689 5971
rect 578563 5967 578698 5971
rect 566800 5658 567800 5708
rect 567921 5658 568921 5708
rect 569042 5658 570042 5708
rect 570152 5658 571152 5708
rect 571273 5658 572273 5708
rect 572394 5658 573394 5708
rect 573951 5658 574951 5708
rect 575072 5658 576072 5708
rect 576193 5658 577193 5708
rect 577303 5658 578303 5708
rect 566800 5488 567800 5538
rect 567921 5488 568921 5538
rect 569042 5488 570042 5538
rect 570152 5488 571152 5538
rect 571273 5488 572273 5538
rect 572394 5488 573394 5538
rect 573951 5488 574951 5538
rect 575072 5488 576072 5538
rect 576193 5488 577193 5538
rect 577303 5488 578303 5538
rect 566515 5169 573629 5191
rect 368539 3967 368655 3989
rect 468539 3967 468655 3989
rect 568539 3967 568655 3989
rect 58215 3959 58520 3960
rect 110215 3959 110520 3960
rect 214215 3959 214520 3960
rect 314215 3959 314520 3960
rect 366215 3926 368539 3960
rect 368655 3926 368691 3960
rect 414215 3959 414520 3960
rect 466215 3926 468539 3960
rect 468655 3926 468691 3960
rect 518215 3959 518520 3960
rect 566215 3926 568539 3960
rect 568655 3926 568691 3960
rect 58178 2850 58228 3850
rect 58388 2850 58438 3850
rect 58504 2850 58520 3850
rect 70002 3375 70602 3425
rect 70002 3125 70602 3175
rect 69643 2848 69677 2955
rect 70877 2914 70911 2955
rect 70877 2874 70979 2914
rect 70877 2848 70911 2874
rect 110178 2850 110228 3850
rect 110388 2850 110438 3850
rect 110504 2850 110520 3850
rect 122002 3375 122602 3425
rect 174002 3375 174602 3425
rect 122002 3125 122602 3175
rect 174002 3125 174602 3175
rect 121643 2848 121677 2955
rect 122877 2914 122911 2955
rect 122877 2874 122979 2914
rect 122877 2848 122911 2874
rect 173643 2848 173677 2955
rect 174877 2914 174911 2955
rect 174877 2874 174979 2914
rect 174877 2848 174911 2874
rect 214178 2850 214228 3850
rect 214388 2850 214438 3850
rect 214504 2850 214520 3850
rect 226002 3375 226602 3425
rect 274002 3375 274602 3425
rect 226002 3125 226602 3175
rect 274002 3125 274602 3175
rect 225643 2848 225677 2955
rect 226877 2914 226911 2955
rect 226877 2874 226979 2914
rect 226877 2848 226911 2874
rect 273643 2848 273677 2955
rect 274877 2914 274911 2955
rect 274877 2874 274979 2914
rect 274877 2848 274911 2874
rect 314178 2850 314228 3850
rect 314388 2850 314438 3850
rect 314504 2850 314520 3850
rect 326002 3375 326602 3425
rect 326002 3125 326602 3175
rect 325643 2848 325677 2955
rect 326877 2914 326911 2955
rect 326877 2874 326979 2914
rect 326877 2848 326911 2874
rect 366178 2850 366228 3850
rect 366388 2850 366438 3850
rect 366504 2850 366554 3850
rect 366714 2850 366842 3850
rect 366930 2850 366986 3850
rect 367146 2850 367274 3850
rect 367362 3122 367412 3850
rect 367362 3050 367415 3122
rect 367362 2850 367412 3050
rect 367475 2850 367487 3050
rect 368636 2850 368686 3850
rect 368786 2850 368842 3850
rect 368942 2850 369070 3850
rect 369098 2850 369226 3850
rect 369254 2850 369310 3850
rect 369410 2850 369538 3850
rect 369566 2850 369694 3850
rect 369722 2850 369850 3850
rect 369878 2850 369928 3850
rect 369994 2850 370044 3850
rect 370144 2850 370272 3850
rect 370300 2850 370428 3850
rect 370456 2850 370584 3850
rect 370612 2850 370668 3850
rect 370768 2850 370896 3850
rect 370924 2850 371052 3850
rect 371080 2850 371130 3850
rect 371208 2850 371258 3850
rect 371358 2850 371414 3850
rect 371514 2850 371564 3850
rect 371630 3250 371680 3850
rect 371780 3250 371908 3850
rect 371936 3250 371992 3850
rect 372092 3250 372220 3850
rect 372248 3250 372304 3850
rect 372504 3250 372554 3850
rect 372620 3107 372670 3850
rect 372617 2850 372670 3107
rect 372830 2850 372880 3850
rect 372946 2850 372996 3850
rect 373156 2850 373206 3850
rect 373272 2850 373322 3850
rect 373482 2850 373532 3850
rect 373598 2850 373648 3850
rect 373808 2850 373936 3850
rect 374024 2850 374152 3850
rect 374240 2850 374368 3850
rect 374456 2850 374512 3850
rect 374672 2850 374800 3850
rect 374888 2850 375016 3850
rect 375104 2850 375232 3850
rect 375320 2850 375448 3850
rect 375536 2850 375592 3850
rect 375752 2850 375808 3850
rect 375968 2850 376096 3850
rect 376184 2850 376312 3850
rect 376400 2850 376528 3850
rect 376616 2850 376744 3850
rect 376832 2850 376882 3850
rect 378002 3375 378602 3425
rect 378002 3125 378602 3175
rect 377643 2914 377677 2955
rect 378877 2914 378911 2955
rect 377643 2874 377745 2914
rect 378877 2874 378979 2914
rect 377643 2848 377677 2874
rect 378877 2848 378911 2874
rect 414178 2850 414228 3850
rect 414388 2850 414438 3850
rect 414504 2850 414520 3850
rect 426002 3375 426602 3425
rect 426002 3125 426602 3175
rect 425643 2848 425677 2955
rect 426877 2914 426911 2955
rect 426877 2874 426979 2914
rect 426877 2848 426911 2874
rect 466178 2850 466228 3850
rect 466388 2850 466438 3850
rect 466504 2850 466554 3850
rect 466714 2850 466842 3850
rect 466930 2850 466986 3850
rect 467146 2850 467274 3850
rect 467362 3122 467412 3850
rect 467362 3050 467415 3122
rect 467362 2850 467412 3050
rect 467475 2850 467487 3050
rect 468636 2850 468686 3850
rect 468786 2850 468842 3850
rect 468942 2850 469070 3850
rect 469098 2850 469226 3850
rect 469254 2850 469310 3850
rect 469410 2850 469538 3850
rect 469566 2850 469694 3850
rect 469722 2850 469850 3850
rect 469878 2850 469928 3850
rect 469994 2850 470044 3850
rect 470144 2850 470272 3850
rect 470300 2850 470428 3850
rect 470456 2850 470584 3850
rect 470612 2850 470668 3850
rect 470768 2850 470896 3850
rect 470924 2850 471052 3850
rect 471080 2850 471130 3850
rect 471208 2850 471258 3850
rect 471358 2850 471414 3850
rect 471514 2850 471564 3850
rect 471630 3250 471680 3850
rect 471780 3250 471908 3850
rect 471936 3250 471992 3850
rect 472092 3250 472220 3850
rect 472248 3250 472304 3850
rect 472504 3250 472554 3850
rect 472620 3107 472670 3850
rect 472617 2850 472670 3107
rect 472830 2850 472880 3850
rect 472946 2850 472996 3850
rect 473156 2850 473206 3850
rect 473272 2850 473322 3850
rect 473482 2850 473532 3850
rect 473598 2850 473648 3850
rect 473808 2850 473936 3850
rect 474024 2850 474152 3850
rect 474240 2850 474368 3850
rect 474456 2850 474512 3850
rect 474672 2850 474800 3850
rect 474888 2850 475016 3850
rect 475104 2850 475232 3850
rect 475320 2850 475448 3850
rect 475536 2850 475592 3850
rect 475752 2850 475808 3850
rect 475968 2850 476096 3850
rect 476184 2850 476312 3850
rect 476400 2850 476528 3850
rect 476616 2850 476744 3850
rect 476832 2850 476882 3850
rect 478002 3375 478602 3425
rect 478002 3125 478602 3175
rect 477643 2914 477677 2955
rect 478877 2914 478911 2955
rect 477643 2874 477745 2914
rect 478877 2874 478979 2914
rect 477643 2848 477677 2874
rect 478877 2848 478911 2874
rect 518178 2850 518228 3850
rect 518388 2850 518438 3850
rect 518504 2850 518520 3850
rect 530002 3375 530602 3425
rect 530002 3125 530602 3175
rect 529643 2848 529677 2955
rect 530877 2914 530911 2955
rect 530877 2874 530979 2914
rect 530877 2848 530911 2874
rect 566178 2850 566228 3850
rect 566388 2850 566438 3850
rect 566504 2850 566554 3850
rect 566714 2850 566842 3850
rect 566930 2850 566986 3850
rect 567146 2850 567274 3850
rect 567362 3122 567412 3850
rect 567362 3050 567415 3122
rect 567362 2850 567412 3050
rect 567475 2850 567487 3050
rect 568636 2850 568686 3850
rect 568786 2850 568842 3850
rect 568942 2850 569070 3850
rect 569098 2850 569226 3850
rect 569254 2850 569310 3850
rect 569410 2850 569538 3850
rect 569566 2850 569694 3850
rect 569722 2850 569850 3850
rect 569878 2850 569928 3850
rect 569994 2850 570044 3850
rect 570144 2850 570272 3850
rect 570300 2850 570428 3850
rect 570456 2850 570584 3850
rect 570612 2850 570668 3850
rect 570768 2850 570896 3850
rect 570924 2850 571052 3850
rect 571080 2850 571130 3850
rect 571208 2850 571258 3850
rect 571358 2850 571414 3850
rect 571514 2850 571564 3850
rect 571630 3250 571680 3850
rect 571780 3250 571908 3850
rect 571936 3250 571992 3850
rect 572092 3250 572220 3850
rect 572248 3250 572304 3850
rect 572504 3250 572554 3850
rect 572620 3107 572670 3850
rect 572617 2850 572670 3107
rect 572830 2850 572880 3850
rect 572946 2850 572996 3850
rect 573156 2850 573206 3850
rect 573272 2850 573322 3850
rect 573482 2850 573532 3850
rect 573598 2850 573648 3850
rect 573808 2850 573936 3850
rect 574024 2850 574152 3850
rect 574240 2850 574368 3850
rect 574456 2850 574512 3850
rect 574672 2850 574800 3850
rect 574888 2850 575016 3850
rect 575104 2850 575232 3850
rect 575320 2850 575448 3850
rect 575536 2850 575592 3850
rect 575752 2850 575808 3850
rect 575968 2850 576096 3850
rect 576184 2850 576312 3850
rect 576400 2850 576528 3850
rect 576616 2850 576744 3850
rect 576832 2850 576882 3850
rect 578002 3375 578602 3425
rect 578002 3125 578602 3175
rect 577643 2914 577677 2955
rect 578877 2914 578911 2955
rect 577643 2874 577745 2914
rect 578877 2874 578979 2914
rect 577643 2848 577677 2874
rect 578877 2848 578911 2874
rect 69774 2737 71692 2819
rect 121774 2737 123692 2819
rect 173774 2737 175692 2819
rect 225774 2737 227692 2819
rect 273774 2737 275692 2819
rect 325774 2737 327692 2819
rect 377774 2737 379692 2819
rect 425774 2737 427692 2819
rect 477774 2737 479692 2819
rect 529774 2737 531692 2819
rect 577774 2737 579692 2819
rect 56703 1594 57703 1644
rect 69671 1602 69753 2636
rect 69963 1772 70045 2466
rect 70085 2455 71391 2537
rect 70281 2261 71223 2311
rect 71328 2218 71368 2258
rect 71244 2178 71338 2218
rect 71244 2018 71338 2058
rect 71328 1978 71368 2018
rect 70281 1917 71223 1967
rect 70085 1703 71391 1785
rect 71531 1772 71613 2466
rect 71823 1602 71905 2636
rect 108703 1594 109703 1644
rect 121671 1602 121753 2636
rect 121963 1772 122045 2466
rect 122085 2455 123391 2537
rect 122281 2261 123223 2311
rect 123328 2218 123368 2258
rect 123244 2178 123338 2218
rect 123244 2018 123338 2058
rect 123328 1978 123368 2018
rect 122281 1917 123223 1967
rect 122085 1703 123391 1785
rect 123531 1772 123613 2466
rect 123823 1602 123905 2636
rect 160703 1594 161280 1644
rect 173671 1602 173753 2636
rect 173963 1772 174045 2466
rect 174085 2455 175391 2537
rect 174281 2261 175223 2311
rect 175328 2218 175368 2258
rect 175244 2178 175338 2218
rect 175244 2018 175338 2058
rect 175328 1978 175368 2018
rect 174281 1917 175223 1967
rect 174085 1703 175391 1785
rect 175531 1772 175613 2466
rect 175823 1602 175905 2636
rect 212703 1594 213703 1644
rect 225671 1602 225753 2636
rect 225963 1772 226045 2466
rect 226085 2455 227391 2537
rect 226281 2261 227223 2311
rect 227328 2218 227368 2258
rect 227244 2178 227338 2218
rect 227244 2018 227338 2058
rect 227328 1978 227368 2018
rect 226281 1917 227223 1967
rect 226085 1703 227391 1785
rect 227531 1772 227613 2466
rect 227823 1602 227905 2636
rect 260703 1594 261703 1644
rect 273671 1602 273753 2636
rect 273963 1772 274045 2466
rect 274085 2455 275391 2537
rect 274281 2261 275223 2311
rect 275328 2218 275368 2258
rect 275244 2178 275338 2218
rect 275244 2018 275338 2058
rect 275328 1978 275368 2018
rect 274281 1917 275223 1967
rect 274085 1703 275391 1785
rect 275531 1772 275613 2466
rect 275823 1602 275905 2636
rect 312703 1594 313703 1644
rect 325671 1602 325753 2636
rect 325963 1772 326045 2466
rect 326085 2455 327391 2537
rect 326281 2261 327223 2311
rect 327328 2218 327368 2258
rect 327244 2178 327338 2218
rect 327244 2018 327338 2058
rect 327328 1978 327368 2018
rect 326281 1917 327223 1967
rect 326085 1703 327391 1785
rect 327531 1772 327613 2466
rect 327823 1602 327905 2636
rect 369813 2196 370413 2246
rect 367069 2064 368069 2114
rect 369813 2040 370413 2096
rect 370809 2040 371809 2090
rect 367069 1848 368069 1976
rect 369813 1884 370413 1940
rect 370809 1884 371809 2012
rect 369813 1728 370413 1784
rect 370809 1728 371809 1856
rect 364703 1594 365703 1644
rect 367069 1638 368069 1688
rect 369813 1578 370413 1628
rect 370809 1578 371809 1628
rect 377671 1602 377753 2636
rect 377963 1772 378045 2466
rect 378085 2455 379391 2537
rect 378281 2261 379223 2311
rect 378208 2249 378217 2258
rect 379359 2249 379368 2258
rect 378217 2218 378248 2249
rect 379328 2218 379359 2249
rect 378238 2196 378332 2218
rect 378238 2178 378248 2196
rect 378270 2178 378332 2196
rect 379244 2196 379338 2218
rect 379244 2178 379306 2196
rect 379328 2178 379338 2196
rect 378238 2040 378248 2058
rect 378270 2040 378332 2058
rect 378238 2018 378332 2040
rect 379244 2040 379306 2058
rect 379328 2040 379338 2058
rect 379244 2018 379338 2040
rect 378208 1978 378248 2018
rect 379328 1978 379368 2018
rect 378281 1917 379223 1967
rect 378085 1703 379391 1785
rect 379531 1772 379613 2466
rect 379823 1602 379905 2636
rect 412703 1594 413703 1644
rect 425671 1602 425753 2636
rect 425963 1772 426045 2466
rect 426085 2455 427391 2537
rect 426281 2261 427223 2311
rect 427328 2218 427368 2258
rect 427244 2178 427338 2218
rect 427244 2018 427338 2058
rect 427328 1978 427368 2018
rect 426281 1917 427223 1967
rect 426085 1703 427391 1785
rect 427531 1772 427613 2466
rect 427823 1602 427905 2636
rect 469813 2196 470413 2246
rect 467069 2064 468069 2114
rect 469813 2040 470413 2096
rect 470809 2040 471809 2090
rect 467069 1848 468069 1976
rect 469813 1884 470413 1940
rect 470809 1884 471809 2012
rect 469813 1728 470413 1784
rect 470809 1728 471809 1856
rect 464703 1594 465703 1644
rect 467069 1638 468069 1688
rect 469813 1578 470413 1628
rect 470809 1578 471809 1628
rect 477671 1602 477753 2636
rect 477963 1772 478045 2466
rect 478085 2455 479391 2537
rect 478281 2261 479223 2311
rect 478208 2249 478217 2258
rect 479359 2249 479368 2258
rect 478217 2218 478248 2249
rect 479328 2218 479359 2249
rect 478238 2196 478332 2218
rect 478238 2178 478248 2196
rect 478270 2178 478332 2196
rect 479244 2196 479338 2218
rect 479244 2178 479306 2196
rect 479328 2178 479338 2196
rect 478238 2040 478248 2058
rect 478270 2040 478332 2058
rect 478238 2018 478332 2040
rect 479244 2040 479306 2058
rect 479328 2040 479338 2058
rect 479244 2018 479338 2040
rect 478208 1978 478248 2018
rect 479328 1978 479368 2018
rect 478281 1917 479223 1967
rect 478085 1703 479391 1785
rect 479531 1772 479613 2466
rect 479823 1602 479905 2636
rect 516703 1594 517703 1644
rect 529671 1602 529753 2636
rect 529963 1772 530045 2466
rect 530085 2455 531391 2537
rect 530281 2261 531223 2311
rect 531328 2218 531368 2258
rect 531244 2178 531338 2218
rect 531244 2018 531338 2058
rect 531328 1978 531368 2018
rect 530281 1917 531223 1967
rect 530085 1703 531391 1785
rect 531531 1772 531613 2466
rect 531823 1602 531905 2636
rect 569813 2196 570413 2246
rect 567069 2064 568069 2114
rect 569813 2040 570413 2096
rect 570809 2040 571809 2090
rect 567069 1848 568069 1976
rect 569813 1884 570413 1940
rect 570809 1884 571809 2012
rect 569813 1728 570413 1784
rect 570809 1728 571809 1856
rect 564703 1594 565703 1644
rect 567069 1638 568069 1688
rect 569813 1578 570413 1628
rect 570809 1578 571809 1628
rect 577671 1602 577753 2636
rect 577963 1772 578045 2466
rect 578085 2455 579391 2537
rect 578281 2261 579223 2311
rect 578208 2249 578217 2258
rect 579359 2249 579368 2258
rect 578217 2218 578248 2249
rect 579328 2218 579359 2249
rect 578238 2196 578332 2218
rect 578238 2178 578248 2196
rect 578270 2178 578332 2196
rect 579244 2196 579338 2218
rect 579244 2178 579306 2196
rect 579328 2178 579338 2196
rect 578238 2040 578248 2058
rect 578270 2040 578332 2058
rect 578238 2018 578332 2040
rect 579244 2040 579306 2058
rect 579328 2040 579338 2058
rect 579244 2018 579338 2040
rect 578208 1978 578248 2018
rect 579328 1978 579368 2018
rect 578281 1917 579223 1967
rect 578085 1703 579391 1785
rect 579531 1772 579613 2466
rect 579823 1602 579905 2636
rect 56703 1438 57260 1566
rect 69642 1528 69645 1529
rect 69642 1527 69643 1528
rect 69644 1527 69645 1528
rect 69642 1526 69645 1527
rect 69774 1418 71692 1500
rect 108703 1438 109260 1566
rect 121642 1528 121645 1529
rect 121642 1527 121643 1528
rect 121644 1527 121645 1528
rect 121642 1526 121645 1527
rect 121774 1418 123692 1500
rect 160703 1438 161260 1566
rect 173642 1528 173645 1529
rect 173642 1527 173643 1528
rect 173644 1527 173645 1528
rect 173642 1526 173645 1527
rect 173774 1418 175692 1500
rect 212703 1438 213260 1566
rect 225642 1528 225645 1529
rect 225642 1527 225643 1528
rect 225644 1527 225645 1528
rect 225642 1526 225645 1527
rect 225774 1418 227692 1500
rect 260703 1438 261260 1566
rect 273642 1528 273645 1529
rect 273642 1527 273643 1528
rect 273644 1527 273645 1528
rect 273642 1526 273645 1527
rect 273774 1418 275692 1500
rect 312703 1438 313260 1566
rect 325642 1528 325645 1529
rect 325642 1527 325643 1528
rect 325644 1527 325645 1528
rect 325642 1526 325645 1527
rect 325774 1418 327692 1500
rect 364703 1438 365703 1566
rect 377642 1528 377645 1529
rect 377642 1527 377643 1528
rect 377644 1527 377645 1528
rect 377642 1526 377645 1527
rect 377774 1418 379692 1500
rect 412703 1438 413260 1566
rect 425642 1528 425645 1529
rect 425642 1527 425643 1528
rect 425644 1527 425645 1528
rect 425642 1526 425645 1527
rect 425774 1418 427692 1500
rect 464703 1438 465703 1566
rect 477642 1528 477645 1529
rect 477642 1527 477643 1528
rect 477644 1527 477645 1528
rect 477642 1526 477645 1527
rect 477774 1418 479692 1500
rect 516703 1438 517260 1566
rect 529642 1528 529645 1529
rect 529642 1527 529643 1528
rect 529644 1527 529645 1528
rect 529642 1526 529645 1527
rect 529774 1418 531692 1500
rect 564703 1438 565703 1566
rect 577642 1528 577645 1529
rect 577642 1527 577643 1528
rect 577644 1527 577645 1528
rect 577642 1526 577645 1527
rect 577774 1418 579692 1500
rect 69642 1391 69645 1392
rect 69642 1390 69643 1391
rect 69644 1390 69645 1391
rect 69642 1389 69645 1390
rect 121642 1391 121645 1392
rect 121642 1390 121643 1391
rect 121644 1390 121645 1391
rect 121642 1389 121645 1390
rect 173642 1391 173645 1392
rect 173642 1390 173643 1391
rect 173644 1390 173645 1391
rect 173642 1389 173645 1390
rect 225642 1391 225645 1392
rect 225642 1390 225643 1391
rect 225644 1390 225645 1391
rect 225642 1389 225645 1390
rect 273642 1391 273645 1392
rect 273642 1390 273643 1391
rect 273644 1390 273645 1391
rect 273642 1389 273645 1390
rect 325642 1391 325645 1392
rect 325642 1390 325643 1391
rect 325644 1390 325645 1391
rect 325642 1389 325645 1390
rect 377642 1391 377645 1392
rect 377642 1390 377643 1391
rect 377644 1390 377645 1391
rect 377642 1389 377645 1390
rect 425642 1391 425645 1392
rect 425642 1390 425643 1391
rect 425644 1390 425645 1391
rect 425642 1389 425645 1390
rect 477642 1391 477645 1392
rect 477642 1390 477643 1391
rect 477644 1390 477645 1391
rect 477642 1389 477645 1390
rect 529642 1391 529645 1392
rect 529642 1390 529643 1391
rect 529644 1390 529645 1391
rect 529642 1389 529645 1390
rect 577642 1391 577645 1392
rect 577642 1390 577643 1391
rect 577644 1390 577645 1391
rect 577642 1389 577645 1390
rect 56703 1288 57703 1338
rect 69671 282 69753 1316
rect 69963 452 70045 1146
rect 70085 1133 71391 1215
rect 70281 951 71223 1001
rect 71328 900 71368 940
rect 71244 860 71338 900
rect 71244 700 71338 740
rect 71328 660 71368 700
rect 70281 607 71223 657
rect 70085 381 71391 463
rect 71531 452 71613 1146
rect 71823 282 71905 1316
rect 108703 1288 109703 1338
rect 121671 282 121753 1316
rect 121963 452 122045 1146
rect 122085 1133 123391 1215
rect 122281 951 123223 1001
rect 123328 900 123368 940
rect 123244 860 123338 900
rect 123244 700 123338 740
rect 123328 660 123368 700
rect 122281 607 123223 657
rect 122085 381 123391 463
rect 123531 452 123613 1146
rect 123823 282 123905 1316
rect 160703 1288 161280 1338
rect 173671 282 173753 1316
rect 173963 452 174045 1146
rect 174085 1133 175391 1215
rect 174281 951 175223 1001
rect 175328 900 175368 940
rect 175244 860 175338 900
rect 175244 700 175338 740
rect 175328 660 175368 700
rect 174281 607 175223 657
rect 174085 381 175391 463
rect 175531 452 175613 1146
rect 175823 282 175905 1316
rect 212703 1288 213703 1338
rect 225671 282 225753 1316
rect 225963 452 226045 1146
rect 226085 1133 227391 1215
rect 226281 951 227223 1001
rect 227328 900 227368 940
rect 227244 860 227338 900
rect 227244 700 227338 740
rect 227328 660 227368 700
rect 226281 607 227223 657
rect 226085 381 227391 463
rect 227531 452 227613 1146
rect 227823 282 227905 1316
rect 260703 1288 261703 1338
rect 273671 282 273753 1316
rect 273963 452 274045 1146
rect 274085 1133 275391 1215
rect 274281 951 275223 1001
rect 275328 900 275368 940
rect 275244 860 275338 900
rect 275244 700 275338 740
rect 275328 660 275368 700
rect 274281 607 275223 657
rect 274085 381 275391 463
rect 275531 452 275613 1146
rect 275823 282 275905 1316
rect 312703 1288 313703 1338
rect 325671 282 325753 1316
rect 325963 452 326045 1146
rect 326085 1133 327391 1215
rect 326281 951 327223 1001
rect 327328 900 327368 940
rect 327244 860 327338 900
rect 327244 700 327338 740
rect 327328 660 327368 700
rect 326281 607 327223 657
rect 326085 381 327391 463
rect 327531 452 327613 1146
rect 327823 282 327905 1316
rect 364703 1288 365703 1338
rect 369351 875 369404 1175
rect 69774 99 71692 181
rect 121774 99 123692 181
rect 173774 99 175692 181
rect 225774 99 227692 181
rect 273774 99 275692 181
rect 325774 99 327692 181
rect 369354 175 369404 875
rect 369504 175 369632 1175
rect 369660 175 369716 1175
rect 369816 175 369944 1175
rect 369972 175 370022 1175
rect 370088 175 370138 1175
rect 370238 175 370366 1175
rect 370394 175 370450 1175
rect 370550 175 370678 1175
rect 370706 175 370756 1175
rect 370822 175 370872 1175
rect 370972 175 371028 1175
rect 371128 175 371178 1175
rect 371244 175 371294 1175
rect 371394 175 371522 1175
rect 371550 175 371678 1175
rect 371706 175 371834 1175
rect 371862 175 371990 1175
rect 372018 175 372068 1175
rect 372860 1153 372918 1187
rect 373798 183 373848 1183
rect 373948 183 374004 1183
rect 374104 183 374154 1183
rect 374220 583 374270 1183
rect 374370 583 374420 1183
rect 374486 183 374536 1183
rect 374636 183 374692 1183
rect 374792 183 374920 1183
rect 374948 183 375004 1183
rect 375104 183 375232 1183
rect 375260 183 375316 1183
rect 375476 183 375526 1183
rect 375642 183 375692 1183
rect 375792 183 375920 1183
rect 375948 183 376004 1183
rect 376164 183 376220 1183
rect 376380 183 376430 1183
rect 376496 183 376546 1183
rect 376646 183 376774 1183
rect 376802 183 376852 1183
rect 377671 282 377753 1316
rect 377963 452 378045 1146
rect 378085 1133 379391 1215
rect 378281 951 379223 1001
rect 378208 900 378248 940
rect 379328 900 379368 940
rect 378238 860 378332 900
rect 379244 860 379338 900
rect 378238 700 378332 740
rect 379244 700 379338 740
rect 378208 660 378248 700
rect 379328 660 379368 700
rect 378281 607 379223 657
rect 378085 381 379391 463
rect 379531 452 379613 1146
rect 379823 282 379905 1316
rect 412703 1288 413703 1338
rect 425671 282 425753 1316
rect 425963 452 426045 1146
rect 426085 1133 427391 1215
rect 426281 951 427223 1001
rect 427328 900 427368 940
rect 427244 860 427338 900
rect 427244 700 427338 740
rect 427328 660 427368 700
rect 426281 607 427223 657
rect 426085 381 427391 463
rect 427531 452 427613 1146
rect 427823 282 427905 1316
rect 464703 1288 465703 1338
rect 469351 875 469404 1175
rect 377774 99 379692 181
rect 425774 99 427692 181
rect 469354 175 469404 875
rect 469504 175 469632 1175
rect 469660 175 469716 1175
rect 469816 175 469944 1175
rect 469972 175 470022 1175
rect 470088 175 470138 1175
rect 470238 175 470366 1175
rect 470394 175 470450 1175
rect 470550 175 470678 1175
rect 470706 175 470756 1175
rect 470822 175 470872 1175
rect 470972 175 471028 1175
rect 471128 175 471178 1175
rect 471244 175 471294 1175
rect 471394 175 471522 1175
rect 471550 175 471678 1175
rect 471706 175 471834 1175
rect 471862 175 471990 1175
rect 472018 175 472068 1175
rect 472860 1153 472918 1187
rect 473798 183 473848 1183
rect 473948 183 474004 1183
rect 474104 183 474154 1183
rect 474220 583 474270 1183
rect 474370 583 474420 1183
rect 474486 183 474536 1183
rect 474636 183 474692 1183
rect 474792 183 474920 1183
rect 474948 183 475004 1183
rect 475104 183 475232 1183
rect 475260 183 475316 1183
rect 475476 183 475526 1183
rect 475642 183 475692 1183
rect 475792 183 475920 1183
rect 475948 183 476004 1183
rect 476164 183 476220 1183
rect 476380 183 476430 1183
rect 476496 183 476546 1183
rect 476646 183 476774 1183
rect 476802 183 476852 1183
rect 477671 282 477753 1316
rect 477963 452 478045 1146
rect 478085 1133 479391 1215
rect 478281 951 479223 1001
rect 478208 900 478248 940
rect 479328 900 479368 940
rect 478238 860 478332 900
rect 479244 860 479338 900
rect 478238 700 478332 740
rect 479244 700 479338 740
rect 478208 660 478248 700
rect 479328 660 479368 700
rect 478281 607 479223 657
rect 478085 381 479391 463
rect 479531 452 479613 1146
rect 479823 282 479905 1316
rect 516703 1288 517703 1338
rect 529671 282 529753 1316
rect 529963 452 530045 1146
rect 530085 1133 531391 1215
rect 530281 951 531223 1001
rect 531328 900 531368 940
rect 531244 860 531338 900
rect 531244 700 531338 740
rect 531328 660 531368 700
rect 530281 607 531223 657
rect 530085 381 531391 463
rect 531531 452 531613 1146
rect 531823 282 531905 1316
rect 564703 1288 565703 1338
rect 569351 875 569404 1175
rect 477774 99 479692 181
rect 529774 99 531692 181
rect 569354 175 569404 875
rect 569504 175 569632 1175
rect 569660 175 569716 1175
rect 569816 175 569944 1175
rect 569972 175 570022 1175
rect 570088 175 570138 1175
rect 570238 175 570366 1175
rect 570394 175 570450 1175
rect 570550 175 570678 1175
rect 570706 175 570756 1175
rect 570822 175 570872 1175
rect 570972 175 571028 1175
rect 571128 175 571178 1175
rect 571244 175 571294 1175
rect 571394 175 571522 1175
rect 571550 175 571678 1175
rect 571706 175 571834 1175
rect 571862 175 571990 1175
rect 572018 175 572068 1175
rect 572860 1153 572918 1187
rect 573798 183 573848 1183
rect 573948 183 574004 1183
rect 574104 183 574154 1183
rect 574220 583 574270 1183
rect 574370 583 574420 1183
rect 574486 183 574536 1183
rect 574636 183 574692 1183
rect 574792 183 574920 1183
rect 574948 183 575004 1183
rect 575104 183 575232 1183
rect 575260 183 575316 1183
rect 575476 183 575526 1183
rect 575642 183 575692 1183
rect 575792 183 575920 1183
rect 575948 183 576004 1183
rect 576164 183 576220 1183
rect 576380 183 576430 1183
rect 576496 183 576546 1183
rect 576646 183 576774 1183
rect 576802 183 576852 1183
rect 577671 282 577753 1316
rect 577963 452 578045 1146
rect 578085 1133 579391 1215
rect 578281 951 579223 1001
rect 578208 900 578248 940
rect 579328 900 579368 940
rect 578238 860 578332 900
rect 579244 860 579338 900
rect 578238 700 578332 740
rect 579244 700 579338 740
rect 578208 660 578248 700
rect 579328 660 579368 700
rect 578281 607 579223 657
rect 578085 381 579391 463
rect 579531 452 579613 1146
rect 579823 282 579905 1316
rect 577774 99 579692 181
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_2 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605576936
transform -1 0 52000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_1
timestamp 1605576936
transform -1 0 48000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_0
timestamp 1605576936
transform -1 0 44000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_521
timestamp 1605576936
transform 0 -1 39593 1 0 40800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_517
timestamp 1605576936
transform 0 -1 39593 1 0 44800
box 0 0 4120 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605576936
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605576936
transform -1 0 72000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_3
timestamp 1605576936
transform -1 0 56000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_4
timestamp 1605576936
transform -1 0 80000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_5
timestamp 1605576936
transform -1 0 76000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_6
timestamp 1605576936
transform -1 0 84000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_7
timestamp 1605576936
transform -1 0 88000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_8
timestamp 1605576936
transform -1 0 92000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_9
timestamp 1605576936
transform -1 0 96000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_10
timestamp 1605576936
transform -1 0 100000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_1
timestamp 1605576936
transform -1 0 124000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_11
timestamp 1605576936
transform -1 0 104000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_12
timestamp 1605576936
transform -1 0 108000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_13
timestamp 1605576936
transform -1 0 128000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_14
timestamp 1605576936
transform -1 0 132000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_16
timestamp 1605576936
transform -1 0 140000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_15
timestamp 1605576936
transform -1 0 136000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_17
timestamp 1605576936
transform -1 0 144000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_19
timestamp 1605576936
transform -1 0 152000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_18
timestamp 1605576936
transform -1 0 148000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_2
timestamp 1605576936
transform -1 0 176000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_20
timestamp 1605576936
transform -1 0 156000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_21
timestamp 1605576936
transform -1 0 160000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_96
timestamp 1605576936
transform -1 0 180000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_22
timestamp 1605576936
transform -1 0 184000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_23
timestamp 1605576936
transform -1 0 188000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_24
timestamp 1605576936
transform -1 0 192000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_61
timestamp 1605576936
transform 0 -1 39593 -1 0 76800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_520
timestamp 1605576936
transform 0 -1 39593 1 0 56800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_518
timestamp 1605576936
transform 0 -1 39593 1 0 48800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_519
timestamp 1605576936
transform 0 -1 39593 1 0 52800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_513
timestamp 1605576936
transform 0 -1 39593 1 0 76800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_514
timestamp 1605576936
transform 0 -1 39593 1 0 80800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_515
timestamp 1605576936
transform 0 -1 39593 1 0 84800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_516
timestamp 1605576936
transform 0 -1 39593 1 0 88800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_512
timestamp 1605576936
transform 0 -1 39593 1 0 92800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_509
timestamp 1605576936
transform 0 -1 39593 1 0 96800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_60
timestamp 1605576936
transform 0 -1 39593 -1 0 124800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_511
timestamp 1605576936
transform 0 -1 39593 1 0 104800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_510
timestamp 1605576936
transform 0 -1 39593 1 0 100800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_505
timestamp 1605576936
transform 0 -1 39593 1 0 136800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_506
timestamp 1605576936
transform 0 -1 39593 1 0 132800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_507
timestamp 1605576936
transform 0 -1 39593 1 0 128800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_508
timestamp 1605576936
transform 0 -1 39593 1 0 124800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_503
timestamp 1605576936
transform 0 -1 39593 1 0 144800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_504
timestamp 1605576936
transform 0 -1 39593 1 0 140800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_59
timestamp 1605576936
transform 0 -1 39593 -1 0 172800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_501
timestamp 1605576936
transform 0 -1 39593 1 0 152800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_502
timestamp 1605576936
transform 0 -1 39593 1 0 148800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_497
timestamp 1605576936
transform 0 -1 39593 1 0 172800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_498
timestamp 1605576936
transform 0 -1 39593 1 0 176800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_499
timestamp 1605576936
transform 0 -1 39593 1 0 180800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_493
timestamp 1605576936
transform 0 -1 39593 1 0 188800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_496
timestamp 1605576936
transform 0 -1 39593 1 0 192800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_500
timestamp 1605576936
transform 0 -1 39593 1 0 184800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_495
timestamp 1605576936
transform 0 -1 39593 1 0 196800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_58
timestamp 1605576936
transform 0 -1 39593 -1 0 220800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_494
timestamp 1605576936
transform 0 -1 39593 1 0 200800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_492
timestamp 1605576936
transform 0 -1 39593 1 0 220800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_490
timestamp 1605576936
transform 0 -1 39593 1 0 228800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_491
timestamp 1605576936
transform 0 -1 39593 1 0 224800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_487
timestamp 1605576936
transform 0 -1 39593 1 0 240800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_488
timestamp 1605576936
transform 0 -1 39593 1 0 236800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_489
timestamp 1605576936
transform 0 -1 39593 1 0 232800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_486
timestamp 1605576936
transform 0 -1 39593 1 0 244800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_485
timestamp 1605576936
transform 0 -1 39593 1 0 248800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_57
timestamp 1605576936
transform 0 -1 39593 -1 0 272800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_484
timestamp 1605576936
transform 0 -1 39593 1 0 252800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_481
timestamp 1605576936
transform 0 -1 39593 1 0 272800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_480
timestamp 1605576936
transform 0 -1 39593 1 0 284800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_479
timestamp 1605576936
transform 0 -1 39593 1 0 288800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_482
timestamp 1605576936
transform 0 -1 39593 1 0 280800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_483
timestamp 1605576936
transform 0 -1 39593 1 0 276800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_477
timestamp 1605576936
transform 0 -1 39593 1 0 296800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_478
timestamp 1605576936
transform 0 -1 39593 1 0 292800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_56
timestamp 1605576936
transform 0 -1 39593 -1 0 320800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_476
timestamp 1605576936
transform 0 -1 39593 1 0 300800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_472
timestamp 1605576936
transform 0 -1 39593 1 0 332800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_473
timestamp 1605576936
transform 0 -1 39593 1 0 328800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_474
timestamp 1605576936
transform 0 -1 39593 1 0 324800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_475
timestamp 1605576936
transform 0 -1 39593 1 0 320800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_469
timestamp 1605576936
transform 0 -1 39593 1 0 348800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_468
timestamp 1605576936
transform 0 -1 39593 1 0 344800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_470
timestamp 1605576936
transform 0 -1 39593 1 0 336800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_471
timestamp 1605576936
transform 0 -1 39593 1 0 340800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_55
timestamp 1605576936
transform 0 -1 39593 -1 0 368800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_464
timestamp 1605576936
transform 0 -1 39593 1 0 380800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_465
timestamp 1605576936
transform 0 -1 39593 1 0 376800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_466
timestamp 1605576936
transform 0 -1 39593 1 0 372800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_467
timestamp 1605576936
transform 0 -1 39593 1 0 368800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_461
timestamp 1605576936
transform 0 -1 39593 1 0 392800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_462
timestamp 1605576936
transform 0 -1 39593 1 0 388800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_463
timestamp 1605576936
transform 0 -1 39593 1 0 384800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_460
timestamp 1605576936
transform 0 -1 39593 1 0 396800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_54
timestamp 1605576936
transform 0 -1 39593 -1 0 416800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_458
timestamp 1605576936
transform 0 -1 39593 1 0 416800
box 0 0 4120 39593
use bump_pad  bump_pad_0
array 0 5 100000 0 9 100000
timestamp 1602626256
transform 1 0 98924 0 1 68694
box -24800 -24800 25000 24800
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_25
timestamp 1605576936
transform -1 0 196000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_26
timestamp 1605576936
transform -1 0 200000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_27
timestamp 1605576936
transform -1 0 204000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_28
timestamp 1605576936
transform -1 0 208000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_3
timestamp 1605576936
transform -1 0 228000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_29
timestamp 1605576936
transform -1 0 212000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_30
timestamp 1605576936
transform -1 0 232000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_33
timestamp 1605576936
transform -1 0 244000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_32
timestamp 1605576936
transform -1 0 240000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_31
timestamp 1605576936
transform -1 0 236000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_34
timestamp 1605576936
transform -1 0 248000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_35
timestamp 1605576936
transform -1 0 252000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_4
timestamp 1605576936
transform -1 0 276000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_37
timestamp 1605576936
transform -1 0 260000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_36
timestamp 1605576936
transform -1 0 256000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_38
timestamp 1605576936
transform -1 0 280000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_39
timestamp 1605576936
transform -1 0 284000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_41
timestamp 1605576936
transform -1 0 292000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_40
timestamp 1605576936
transform -1 0 288000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_42
timestamp 1605576936
transform -1 0 296000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_43
timestamp 1605576936
transform -1 0 300000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_44
timestamp 1605576936
transform -1 0 304000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_45
timestamp 1605576936
transform -1 0 308000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_46
timestamp 1605576936
transform -1 0 312000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_5
timestamp 1605576936
transform -1 0 328000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_50
timestamp 1605576936
transform -1 0 344000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_49
timestamp 1605576936
transform -1 0 340000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_48
timestamp 1605576936
transform -1 0 336000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_47
timestamp 1605576936
transform -1 0 332000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_54
timestamp 1605576936
transform -1 0 360000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_53
timestamp 1605576936
transform -1 0 356000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_52
timestamp 1605576936
transform -1 0 352000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_51
timestamp 1605576936
transform -1 0 348000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_6
timestamp 1605576936
transform -1 0 380000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_55
timestamp 1605576936
transform -1 0 364000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_7
timestamp 1605576936
transform -1 0 428000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_56
timestamp 1605576936
transform -1 0 384000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_58
timestamp 1605576936
transform -1 0 392000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_57
timestamp 1605576936
transform -1 0 388000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_62
timestamp 1605576936
transform -1 0 408000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_61
timestamp 1605576936
transform -1 0 404000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_60
timestamp 1605576936
transform -1 0 400000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_59
timestamp 1605576936
transform -1 0 396000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_63
timestamp 1605576936
transform -1 0 412000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_66
timestamp 1605576936
transform -1 0 440000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_65
timestamp 1605576936
transform -1 0 436000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_64
timestamp 1605576936
transform -1 0 432000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_67
timestamp 1605576936
transform -1 0 444000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_70
timestamp 1605576936
transform -1 0 456000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_68
timestamp 1605576936
transform -1 0 448000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_69
timestamp 1605576936
transform -1 0 452000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_71
timestamp 1605576936
transform -1 0 460000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_72
timestamp 1605576936
transform -1 0 464000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_8
timestamp 1605576936
transform -1 0 480000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_74
timestamp 1605576936
transform -1 0 488000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_73
timestamp 1605576936
transform -1 0 484000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_78
timestamp 1605576936
transform -1 0 504000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_77
timestamp 1605576936
transform -1 0 500000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_76
timestamp 1605576936
transform -1 0 496000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_75
timestamp 1605576936
transform -1 0 492000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_9
timestamp 1605576936
transform -1 0 532000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_81
timestamp 1605576936
transform -1 0 516000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_80
timestamp 1605576936
transform -1 0 512000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_79
timestamp 1605576936
transform -1 0 508000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_82
timestamp 1605576936
transform -1 0 536000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_83
timestamp 1605576936
transform -1 0 540000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_85
timestamp 1605576936
transform -1 0 548000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_84
timestamp 1605576936
transform -1 0 544000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_86
timestamp 1605576936
transform -1 0 552000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_89
timestamp 1605576936
transform -1 0 564000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_88
timestamp 1605576936
transform -1 0 560000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_87
timestamp 1605576936
transform -1 0 556000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_10
timestamp 1605576936
transform -1 0 580000 0 -1 39593
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_92
timestamp 1605576936
transform -1 0 592000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_91
timestamp 1605576936
transform -1 0 588000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_90
timestamp 1605576936
transform -1 0 584000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_93
timestamp 1605576936
transform -1 0 596000 0 -1 39593
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_94
timestamp 1605576936
transform -1 0 600000 0 -1 39593
box 0 0 4120 39593
use sky130_fd_io__corner_bus_overlay  sky130_fd_io__corner_bus_overlay_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1605576936
transform 0 1 676867 -1 0 40000
box 0 0 40000 40733
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_21
timestamp 1605576936
transform 0 1 678007 1 0 56000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_95
timestamp 1605576936
transform 0 1 678007 -1 0 44000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_196
timestamp 1605576936
transform 0 1 678007 -1 0 56000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_195
timestamp 1605576936
transform 0 1 678007 -1 0 52000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_194
timestamp 1605576936
transform 0 1 678007 -1 0 48000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_11
timestamp 1605576936
transform 0 1 678007 1 0 104000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_199
timestamp 1605576936
transform 0 1 678007 -1 0 88000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_198
timestamp 1605576936
transform 0 1 678007 -1 0 84000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_197
timestamp 1605576936
transform 0 1 678007 -1 0 80000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_99
timestamp 1605576936
transform 0 1 678007 -1 0 76000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_203
timestamp 1605576936
transform 0 1 678007 -1 0 104000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_202
timestamp 1605576936
transform 0 1 678007 -1 0 100000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_201
timestamp 1605576936
transform 0 1 678007 -1 0 96000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_200
timestamp 1605576936
transform 0 1 678007 -1 0 92000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_204
timestamp 1605576936
transform 0 1 678007 -1 0 124000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_205
timestamp 1605576936
transform 0 1 678007 -1 0 128000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_206
timestamp 1605576936
transform 0 1 678007 -1 0 132000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_207
timestamp 1605576936
transform 0 1 678007 -1 0 136000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_208
timestamp 1605576936
transform 0 1 678007 -1 0 140000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_209
timestamp 1605576936
transform 0 1 678007 -1 0 144000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_210
timestamp 1605576936
transform 0 1 678007 -1 0 148000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_211
timestamp 1605576936
transform 0 1 678007 -1 0 152000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_12
timestamp 1605576936
transform 0 1 678007 1 0 152000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_214
timestamp 1605576936
transform 0 1 678007 -1 0 180000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_213
timestamp 1605576936
transform 0 1 678007 -1 0 176000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_212
timestamp 1605576936
transform 0 1 678007 -1 0 172000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_215
timestamp 1605576936
transform 0 1 678007 -1 0 184000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_216
timestamp 1605576936
transform 0 1 678007 -1 0 188000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_217
timestamp 1605576936
transform 0 1 678007 -1 0 192000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_218
timestamp 1605576936
transform 0 1 678007 -1 0 196000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_13
timestamp 1605576936
transform 0 1 678007 1 0 200000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_219
timestamp 1605576936
transform 0 1 678007 -1 0 200000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_220
timestamp 1605576936
transform 0 1 678007 -1 0 220000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_221
timestamp 1605576936
transform 0 1 678007 -1 0 224000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_222
timestamp 1605576936
transform 0 1 678007 -1 0 228000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_223
timestamp 1605576936
transform 0 1 678007 -1 0 232000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_225
timestamp 1605576936
transform 0 1 678007 -1 0 240000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_224
timestamp 1605576936
transform 0 1 678007 -1 0 236000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_14
timestamp 1605576936
transform 0 1 678007 1 0 248000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_227
timestamp 1605576936
transform 0 1 678007 -1 0 248000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_226
timestamp 1605576936
transform 0 1 678007 -1 0 244000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_228
timestamp 1605576936
transform 0 1 678007 -1 0 268000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_229
timestamp 1605576936
transform 0 1 678007 -1 0 272000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_230
timestamp 1605576936
transform 0 1 678007 -1 0 276000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_231
timestamp 1605576936
transform 0 1 678007 -1 0 280000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_232
timestamp 1605576936
transform 0 1 678007 -1 0 284000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_233
timestamp 1605576936
transform 0 1 678007 -1 0 288000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_234
timestamp 1605576936
transform 0 1 678007 -1 0 292000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_235
timestamp 1605576936
transform 0 1 678007 -1 0 296000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_15
timestamp 1605576936
transform 0 1 678007 1 0 296000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_239
timestamp 1605576936
transform 0 1 678007 -1 0 328000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_236
timestamp 1605576936
transform 0 1 678007 -1 0 316000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_237
timestamp 1605576936
transform 0 1 678007 -1 0 320000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_238
timestamp 1605576936
transform 0 1 678007 -1 0 324000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_240
timestamp 1605576936
transform 0 1 678007 -1 0 332000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_242
timestamp 1605576936
transform 0 1 678007 -1 0 340000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_241
timestamp 1605576936
transform 0 1 678007 -1 0 336000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_243
timestamp 1605576936
transform 0 1 678007 -1 0 344000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_244
timestamp 1605576936
transform 0 1 678007 -1 0 348000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_16
timestamp 1605576936
transform 0 1 678007 1 0 348000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_245
timestamp 1605576936
transform 0 1 678007 -1 0 368000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_246
timestamp 1605576936
transform 0 1 678007 -1 0 372000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_247
timestamp 1605576936
transform 0 1 678007 -1 0 376000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_248
timestamp 1605576936
transform 0 1 678007 -1 0 380000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_249
timestamp 1605576936
transform 0 1 678007 -1 0 384000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_250
timestamp 1605576936
transform 0 1 678007 -1 0 388000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_17
timestamp 1605576936
transform 0 1 678007 1 0 396000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_251
timestamp 1605576936
transform 0 1 678007 -1 0 392000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_252
timestamp 1605576936
transform 0 1 678007 -1 0 396000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_253
timestamp 1605576936
transform 0 1 678007 -1 0 416000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_254
timestamp 1605576936
transform 0 1 678007 -1 0 420000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_456
timestamp 1605576936
transform 0 -1 39593 1 0 424800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_459
timestamp 1605576936
transform 0 -1 39593 1 0 420800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_455
timestamp 1605576936
transform 0 -1 39593 1 0 432800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_457
timestamp 1605576936
transform 0 -1 39593 1 0 428800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_53
timestamp 1605576936
transform 0 -1 39593 -1 0 464800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_452
timestamp 1605576936
transform 0 -1 39593 1 0 444800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_453
timestamp 1605576936
transform 0 -1 39593 1 0 440800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_454
timestamp 1605576936
transform 0 -1 39593 1 0 436800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_451
timestamp 1605576936
transform 0 -1 39593 1 0 464800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_448
timestamp 1605576936
transform 0 -1 39593 1 0 476800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_449
timestamp 1605576936
transform 0 -1 39593 1 0 472800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_450
timestamp 1605576936
transform 0 -1 39593 1 0 468800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_447
timestamp 1605576936
transform 0 -1 39593 1 0 480800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_443
timestamp 1605576936
transform 0 -1 39593 1 0 488800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_444
timestamp 1605576936
transform 0 -1 39593 1 0 492800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_446
timestamp 1605576936
transform 0 -1 39593 1 0 484800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_52
timestamp 1605576936
transform 0 -1 39593 -1 0 516800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_445
timestamp 1605576936
transform 0 -1 39593 1 0 496800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_440
timestamp 1605576936
transform 0 -1 39593 1 0 524800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_441
timestamp 1605576936
transform 0 -1 39593 1 0 520800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_442
timestamp 1605576936
transform 0 -1 39593 1 0 516800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_439
timestamp 1605576936
transform 0 -1 39593 1 0 528800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_437
timestamp 1605576936
transform 0 -1 39593 1 0 536800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_438
timestamp 1605576936
transform 0 -1 39593 1 0 532800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_51
timestamp 1605576936
transform 0 -1 39593 -1 0 568800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_435
timestamp 1605576936
transform 0 -1 39593 1 0 544800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_436
timestamp 1605576936
transform 0 -1 39593 1 0 540800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_434
timestamp 1605576936
transform 0 -1 39593 1 0 548800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_431
timestamp 1605576936
transform 0 -1 39593 1 0 568800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_433
timestamp 1605576936
transform 0 -1 39593 1 0 576800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_427
timestamp 1605576936
transform 0 -1 39593 1 0 580800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_432
timestamp 1605576936
transform 0 -1 39593 1 0 572800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_428
timestamp 1605576936
transform 0 -1 39593 1 0 584800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_429
timestamp 1605576936
transform 0 -1 39593 1 0 592800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_426
timestamp 1605576936
transform 0 -1 39593 1 0 596800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_430
timestamp 1605576936
transform 0 -1 39593 1 0 588800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_50
timestamp 1605576936
transform 0 -1 39593 -1 0 616800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_425
timestamp 1605576936
transform 0 -1 39593 1 0 616800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_422
timestamp 1605576936
transform 0 -1 39593 1 0 628800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_423
timestamp 1605576936
transform 0 -1 39593 1 0 624800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_424
timestamp 1605576936
transform 0 -1 39593 1 0 620800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_49
timestamp 1605576936
transform 0 -1 39593 -1 0 664800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_421
timestamp 1605576936
transform 0 -1 39593 1 0 632800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_418
timestamp 1605576936
transform 0 -1 39593 1 0 644800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_419
timestamp 1605576936
transform 0 -1 39593 1 0 640800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_420
timestamp 1605576936
transform 0 -1 39593 1 0 636800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_416
timestamp 1605576936
transform 0 -1 39593 1 0 668800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_417
timestamp 1605576936
transform 0 -1 39593 1 0 664800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_415
timestamp 1605576936
transform 0 -1 39593 1 0 672800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_412
timestamp 1605576936
transform 0 -1 39593 1 0 684800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_413
timestamp 1605576936
transform 0 -1 39593 1 0 680800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_414
timestamp 1605576936
transform 0 -1 39593 1 0 676800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_411
timestamp 1605576936
transform 0 -1 39593 1 0 688800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_48
timestamp 1605576936
transform 0 -1 39593 -1 0 712800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_410
timestamp 1605576936
transform 0 -1 39593 1 0 692800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_408
timestamp 1605576936
transform 0 -1 39593 1 0 716800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_409
timestamp 1605576936
transform 0 -1 39593 1 0 712800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_407
timestamp 1605576936
transform 0 -1 39593 1 0 724800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_402
timestamp 1605576936
transform 0 -1 39593 1 0 732800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_405
timestamp 1605576936
transform 0 -1 39593 1 0 728800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_406
timestamp 1605576936
transform 0 -1 39593 1 0 720800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_47
timestamp 1605576936
transform 0 -1 39593 -1 0 764800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_404
timestamp 1605576936
transform 0 -1 39593 1 0 736800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_403
timestamp 1605576936
transform 0 -1 39593 1 0 740800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_401
timestamp 1605576936
transform 0 -1 39593 1 0 744800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_399
timestamp 1605576936
transform 0 -1 39593 1 0 768800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_400
timestamp 1605576936
transform 0 -1 39593 1 0 764800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_398
timestamp 1605576936
transform 0 -1 39593 1 0 772800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_397
timestamp 1605576936
transform 0 -1 39593 1 0 776800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_46
timestamp 1605576936
transform 0 -1 39593 -1 0 812800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_394
timestamp 1605576936
transform 0 -1 39593 1 0 788800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_395
timestamp 1605576936
transform 0 -1 39593 1 0 784800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_396
timestamp 1605576936
transform 0 -1 39593 1 0 780800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_393
timestamp 1605576936
transform 0 -1 39593 1 0 792800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_390
timestamp 1605576936
transform 0 -1 39593 1 0 812800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_392
timestamp 1605576936
transform 0 -1 39593 1 0 820800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_391
timestamp 1605576936
transform 0 -1 39593 1 0 816800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_388
timestamp 1605576936
transform 0 -1 39593 1 0 828800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_389
timestamp 1605576936
transform 0 -1 39593 1 0 824800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_386
timestamp 1605576936
transform 0 -1 39593 1 0 836800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_387
timestamp 1605576936
transform 0 -1 39593 1 0 832800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_45
timestamp 1605576936
transform 0 -1 39593 -1 0 860800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_385
timestamp 1605576936
transform 0 -1 39593 1 0 840800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_381
timestamp 1605576936
transform 0 -1 39593 1 0 872800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_382
timestamp 1605576936
transform 0 -1 39593 1 0 868800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_383
timestamp 1605576936
transform 0 -1 39593 1 0 864800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_384
timestamp 1605576936
transform 0 -1 39593 1 0 860800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_377
timestamp 1605576936
transform 0 -1 39593 1 0 888800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_379
timestamp 1605576936
transform 0 -1 39593 1 0 884800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_378
timestamp 1605576936
transform 0 -1 39593 1 0 880800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_380
timestamp 1605576936
transform 0 -1 39593 1 0 876800
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_44
timestamp 1605576936
transform 0 -1 39593 -1 0 908800
box -143 -515 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_43
timestamp 1605576936
transform 0 -1 39593 -1 0 926800
box -143 -515 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_42
timestamp 1605576936
transform 0 -1 39593 -1 0 981600
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_360
timestamp 1605576936
transform 0 -1 39593 1 0 981600
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_358
timestamp 1605576936
transform 0 -1 39593 1 0 989600
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_359
timestamp 1605576936
transform 0 -1 39593 1 0 985600
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_357
timestamp 1605576936
transform 0 -1 39593 1 0 993600
box 0 0 4120 39593
use sky130_fd_io__corner_bus_overlay  sky130_fd_io__corner_bus_overlay_1
timestamp 1605576936
transform 0 -1 40733 1 0 997600
box 0 0 40000 40733
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_41
timestamp 1605576936
transform 1 0 60733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_193
timestamp 1605576936
transform 1 0 40733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_192
timestamp 1605576936
transform 1 0 44733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_189
timestamp 1605576936
transform 1 0 48733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_190
timestamp 1605576936
transform 1 0 52733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_191
timestamp 1605576936
transform 1 0 56733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_40
timestamp 1605576936
transform 1 0 108733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_182
timestamp 1605576936
transform 1 0 76733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_183
timestamp 1605576936
transform 1 0 80733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_181
timestamp 1605576936
transform 1 0 104733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_186
timestamp 1605576936
transform 1 0 92733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_187
timestamp 1605576936
transform 1 0 96733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_188
timestamp 1605576936
transform 1 0 100733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_184
timestamp 1605576936
transform 1 0 84733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_185
timestamp 1605576936
transform 1 0 88733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_176
timestamp 1605576936
transform 1 0 124733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_179
timestamp 1605576936
transform 1 0 136733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_178
timestamp 1605576936
transform 1 0 132733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_177
timestamp 1605576936
transform 1 0 128733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_180
timestamp 1605576936
transform 1 0 140733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_175
timestamp 1605576936
transform 1 0 144733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_171
timestamp 1605576936
transform 1 0 152733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_170
timestamp 1605576936
transform 1 0 148733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_39
timestamp 1605576936
transform 1 0 160733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_172
timestamp 1605576936
transform 1 0 156733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_173
timestamp 1605576936
transform 1 0 176733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_174
timestamp 1605576936
transform 1 0 180733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_166
timestamp 1605576936
transform 1 0 188733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_169
timestamp 1605576936
transform 1 0 184733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_255
timestamp 1605576936
transform 0 1 678007 -1 0 424000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_256
timestamp 1605576936
transform 0 1 678007 -1 0 428000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_257
timestamp 1605576936
transform 0 1 678007 -1 0 432000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_258
timestamp 1605576936
transform 0 1 678007 -1 0 436000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_18
timestamp 1605576936
transform 0 1 678007 1 0 444000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_259
timestamp 1605576936
transform 0 1 678007 -1 0 440000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_260
timestamp 1605576936
transform 0 1 678007 -1 0 444000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_261
timestamp 1605576936
transform 0 1 678007 -1 0 464000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_262
timestamp 1605576936
transform 0 1 678007 -1 0 468000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_263
timestamp 1605576936
transform 0 1 678007 -1 0 472000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_265
timestamp 1605576936
transform 0 1 678007 -1 0 480000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_264
timestamp 1605576936
transform 0 1 678007 -1 0 476000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_267
timestamp 1605576936
transform 0 1 678007 -1 0 488000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_266
timestamp 1605576936
transform 0 1 678007 -1 0 484000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_19
timestamp 1605576936
transform 0 1 678007 1 0 492000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_268
timestamp 1605576936
transform 0 1 678007 -1 0 492000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_269
timestamp 1605576936
transform 0 1 678007 -1 0 512000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_270
timestamp 1605576936
transform 0 1 678007 -1 0 516000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_271
timestamp 1605576936
transform 0 1 678007 -1 0 520000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_272
timestamp 1605576936
transform 0 1 678007 -1 0 524000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_275
timestamp 1605576936
transform 0 1 678007 -1 0 536000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_273
timestamp 1605576936
transform 0 1 678007 -1 0 528000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_274
timestamp 1605576936
transform 0 1 678007 -1 0 532000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_276
timestamp 1605576936
transform 0 1 678007 -1 0 540000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_20
timestamp 1605576936
transform 0 1 678007 1 0 544000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_277
timestamp 1605576936
transform 0 1 678007 -1 0 544000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_281
timestamp 1605576936
transform 0 1 678007 -1 0 576000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_280
timestamp 1605576936
transform 0 1 678007 -1 0 572000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_279
timestamp 1605576936
transform 0 1 678007 -1 0 568000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_278
timestamp 1605576936
transform 0 1 678007 -1 0 564000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_282
timestamp 1605576936
transform 0 1 678007 -1 0 580000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_283
timestamp 1605576936
transform 0 1 678007 -1 0 584000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_284
timestamp 1605576936
transform 0 1 678007 -1 0 588000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_285
timestamp 1605576936
transform 0 1 678007 -1 0 592000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_22
timestamp 1605576936
transform 0 1 678007 1 0 596000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_286
timestamp 1605576936
transform 0 1 678007 -1 0 596000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_287
timestamp 1605576936
transform 0 1 678007 -1 0 616000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_288
timestamp 1605576936
transform 0 1 678007 -1 0 620000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_289
timestamp 1605576936
transform 0 1 678007 -1 0 624000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_290
timestamp 1605576936
transform 0 1 678007 -1 0 628000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_292
timestamp 1605576936
transform 0 1 678007 -1 0 636000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_291
timestamp 1605576936
transform 0 1 678007 -1 0 632000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_294
timestamp 1605576936
transform 0 1 678007 -1 0 644000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_293
timestamp 1605576936
transform 0 1 678007 -1 0 640000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_23
timestamp 1605576936
transform 0 1 678007 1 0 644000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_295
timestamp 1605576936
transform 0 1 678007 -1 0 664000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_296
timestamp 1605576936
transform 0 1 678007 -1 0 668000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_297
timestamp 1605576936
transform 0 1 678007 -1 0 672000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_298
timestamp 1605576936
transform 0 1 678007 -1 0 676000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_299
timestamp 1605576936
transform 0 1 678007 -1 0 680000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_24
timestamp 1605576936
transform 0 1 678007 1 0 692000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_300
timestamp 1605576936
transform 0 1 678007 -1 0 684000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_301
timestamp 1605576936
transform 0 1 678007 -1 0 688000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_302
timestamp 1605576936
transform 0 1 678007 -1 0 692000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_303
timestamp 1605576936
transform 0 1 678007 -1 0 712000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_304
timestamp 1605576936
transform 0 1 678007 -1 0 716000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_307
timestamp 1605576936
transform 0 1 678007 -1 0 728000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_306
timestamp 1605576936
transform 0 1 678007 -1 0 724000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_305
timestamp 1605576936
transform 0 1 678007 -1 0 720000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_308
timestamp 1605576936
transform 0 1 678007 -1 0 732000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_25
timestamp 1605576936
transform 0 1 678007 1 0 740000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_310
timestamp 1605576936
transform 0 1 678007 -1 0 740000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_309
timestamp 1605576936
transform 0 1 678007 -1 0 736000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_311
timestamp 1605576936
transform 0 1 678007 -1 0 760000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_312
timestamp 1605576936
transform 0 1 678007 -1 0 764000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_313
timestamp 1605576936
transform 0 1 678007 -1 0 768000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_314
timestamp 1605576936
transform 0 1 678007 -1 0 772000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_315
timestamp 1605576936
transform 0 1 678007 -1 0 776000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_316
timestamp 1605576936
transform 0 1 678007 -1 0 780000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_317
timestamp 1605576936
transform 0 1 678007 -1 0 784000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_27
timestamp 1605576936
transform 0 1 678007 1 0 788000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_318
timestamp 1605576936
transform 0 1 678007 -1 0 788000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_319
timestamp 1605576936
transform 0 1 678007 -1 0 808000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_320
timestamp 1605576936
transform 0 1 678007 -1 0 812000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_321
timestamp 1605576936
transform 0 1 678007 -1 0 816000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_323
timestamp 1605576936
transform 0 1 678007 -1 0 824000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_322
timestamp 1605576936
transform 0 1 678007 -1 0 820000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_324
timestamp 1605576936
transform 0 1 678007 -1 0 828000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_325
timestamp 1605576936
transform 0 1 678007 -1 0 832000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_326
timestamp 1605576936
transform 0 1 678007 -1 0 836000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_29
timestamp 1605576936
transform 0 1 678007 1 0 840000
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_327
timestamp 1605576936
transform 0 1 678007 -1 0 840000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_329
timestamp 1605576936
transform 0 1 678007 -1 0 864000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_328
timestamp 1605576936
transform 0 1 678007 -1 0 860000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_330
timestamp 1605576936
transform 0 1 678007 -1 0 868000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_331
timestamp 1605576936
transform 0 1 678007 -1 0 872000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_335
timestamp 1605576936
transform 0 1 678007 -1 0 888000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_334
timestamp 1605576936
transform 0 1 678007 -1 0 884000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_333
timestamp 1605576936
transform 0 1 678007 -1 0 880000
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_332
timestamp 1605576936
transform 0 1 678007 -1 0 876000
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_30
timestamp 1605576936
transform 0 1 678007 1 0 888000
box -143 -515 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_31
timestamp 1605576936
transform 0 1 678007 1 0 906000
box -143 -515 16134 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_32
timestamp 1605576936
transform 0 1 678007 1 0 960800
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_353
timestamp 1605576936
transform 0 1 678007 -1 0 984800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_354
timestamp 1605576936
transform 0 1 678007 -1 0 988800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_352
timestamp 1605576936
transform 0 1 678007 -1 0 980800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_355
timestamp 1605576936
transform 0 1 678007 -1 0 992800
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_165
timestamp 1605576936
transform 1 0 192733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_163
timestamp 1605576936
transform 1 0 196733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_167
timestamp 1605576936
transform 1 0 204733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_164
timestamp 1605576936
transform 1 0 200733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_38
timestamp 1605576936
transform 1 0 212733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_168
timestamp 1605576936
transform 1 0 208733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_162
timestamp 1605576936
transform 1 0 228733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_155
timestamp 1605576936
transform 1 0 232733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_156
timestamp 1605576936
transform 1 0 236733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_157
timestamp 1605576936
transform 1 0 240733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_158
timestamp 1605576936
transform 1 0 244733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_160
timestamp 1605576936
transform 1 0 252733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_161
timestamp 1605576936
transform 1 0 256733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_159
timestamp 1605576936
transform 1 0 248733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_37
timestamp 1605576936
transform 1 0 260733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_154
timestamp 1605576936
transform 1 0 276733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_153
timestamp 1605576936
transform 1 0 280733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_151
timestamp 1605576936
transform 1 0 288733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_152
timestamp 1605576936
transform 1 0 284733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_150
timestamp 1605576936
transform 1 0 292733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_146
timestamp 1605576936
transform 1 0 304733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_147
timestamp 1605576936
transform 1 0 300733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_148
timestamp 1605576936
transform 1 0 296733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_149
timestamp 1605576936
transform 1 0 308733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_36
timestamp 1605576936
transform 1 0 312733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_141
timestamp 1605576936
transform 1 0 328733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_144
timestamp 1605576936
transform 1 0 332733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_143
timestamp 1605576936
transform 1 0 336733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_142
timestamp 1605576936
transform 1 0 340733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_145
timestamp 1605576936
transform 1 0 344733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_140
timestamp 1605576936
transform 1 0 348733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_136
timestamp 1605576936
transform 1 0 356733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_135
timestamp 1605576936
transform 1 0 352733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_137
timestamp 1605576936
transform 1 0 360733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_35
timestamp 1605576936
transform 1 0 364733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_138
timestamp 1605576936
transform 1 0 380733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_139
timestamp 1605576936
transform 1 0 384733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_129
timestamp 1605576936
transform 1 0 392733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_134
timestamp 1605576936
transform 1 0 388733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_130
timestamp 1605576936
transform 1 0 396733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_34
timestamp 1605576936
transform 1 0 412733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_133
timestamp 1605576936
transform 1 0 408733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_131
timestamp 1605576936
transform 1 0 400733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_132
timestamp 1605576936
transform 1 0 404733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_127
timestamp 1605576936
transform 1 0 428733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_128
timestamp 1605576936
transform 1 0 432733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_120
timestamp 1605576936
transform 1 0 436733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_121
timestamp 1605576936
transform 1 0 440733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_122
timestamp 1605576936
transform 1 0 444733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_123
timestamp 1605576936
transform 1 0 448733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_33
timestamp 1605576936
transform 1 0 464733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_124
timestamp 1605576936
transform 1 0 452733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_125
timestamp 1605576936
transform 1 0 456733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_126
timestamp 1605576936
transform 1 0 460733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_119
timestamp 1605576936
transform 1 0 480733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_115
timestamp 1605576936
transform 1 0 496733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_118
timestamp 1605576936
transform 1 0 492733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_116
timestamp 1605576936
transform 1 0 484733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_117
timestamp 1605576936
transform 1 0 488733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_111
timestamp 1605576936
transform 1 0 500733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_28
timestamp 1605576936
transform 1 0 516733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_112
timestamp 1605576936
transform 1 0 508733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_113
timestamp 1605576936
transform 1 0 504733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_114
timestamp 1605576936
transform 1 0 512733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_106
timestamp 1605576936
transform 1 0 532733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_107
timestamp 1605576936
transform 1 0 536733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_108
timestamp 1605576936
transform 1 0 540733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_109
timestamp 1605576936
transform 1 0 544733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_110
timestamp 1605576936
transform 1 0 548733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_105
timestamp 1605576936
transform 1 0 552733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_26
timestamp 1605576936
transform 1 0 568733 0 1 998007
box -143 -515 16134 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_104
timestamp 1605576936
transform 1 0 564733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_101
timestamp 1605576936
transform 1 0 560733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_100
timestamp 1605576936
transform 1 0 556733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_103
timestamp 1605576936
transform 1 0 584733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_102
timestamp 1605576936
transform 1 0 588733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_98
timestamp 1605576936
transform 1 0 592733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_97
timestamp 1605576936
transform 1 0 596733 0 1 998007
box 0 0 4120 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_356
timestamp 1605576936
transform 0 1 678007 -1 0 996800
box 0 0 4120 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_1
timestamp 1605576936
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
<< end >>
