magic
tech sky130A
magscale 12 1
timestamp 1598772956
<< metal5 >>
rect 0 90 45 105
rect 30 70 45 90
rect 25 65 45 70
rect 20 60 45 65
rect 15 55 40 60
rect 10 50 35 55
rect 5 45 30 50
rect 0 40 25 45
rect 0 35 20 40
rect 0 15 15 35
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
