magic
tech sky130A
magscale 12 1
timestamp 1598364576
<< metal5 >>
rect 1680 505 1710 535
rect 1725 505 1755 535
rect 1665 480 1680 490
rect 1755 480 1770 490
rect 1665 475 1685 480
rect 1750 475 1770 480
rect 1665 470 1690 475
rect 1745 470 1770 475
rect 1670 465 1695 470
rect 1740 465 1765 470
rect 1675 460 1760 465
rect 1680 455 1755 460
rect 1685 450 1750 455
<< end >>
